magic
tech sky130A
magscale 1 2
timestamp 1699020319
<< nwell >>
rect 164478 538235 166678 539795
rect 168278 538235 170478 539795
rect 171978 538235 174178 539795
rect 175478 538235 177678 539795
rect 179078 538235 181278 539795
rect 182378 538235 184578 539795
rect 185678 538235 187878 539795
rect 188978 538235 191178 539795
rect 157548 535645 162908 537885
rect 172170 529752 187518 530318
rect 172170 528664 187518 529230
rect 172170 527576 187518 528142
rect 172170 526488 187518 527054
rect 172170 525400 187518 525966
rect 172170 524312 187518 524878
rect 172170 523224 187518 523790
rect 172170 522136 187518 522702
rect 172170 521048 187518 521614
rect 172170 519960 187518 520526
rect 172170 518872 187518 519438
rect 172170 517784 187518 518350
rect 172170 516696 187518 517262
rect 172170 515608 187518 516174
<< pwell >>
rect 164498 539795 166678 541315
rect 168298 539795 170478 541315
rect 171998 539795 174178 541315
rect 175498 539795 177678 541315
rect 179098 539795 181278 541315
rect 182398 539795 184578 541315
rect 185698 539795 187878 541315
rect 188998 539795 191178 541315
rect 157548 537895 162908 538825
rect 164150 535835 166778 538115
rect 167922 535835 169278 538115
rect 171658 535835 172378 538115
rect 175176 535835 175578 538115
rect 178776 536395 179178 538115
rect 182076 536675 182478 538115
rect 185376 536815 185778 538115
rect 188676 536719 189078 538115
rect 164120 533495 166748 535775
rect 172237 530558 172271 530596
rect 172973 530558 173007 530596
rect 173065 530558 173099 530596
rect 174169 530558 174203 530596
rect 174720 530568 174744 530590
rect 175365 530558 175399 530596
rect 175456 530568 175480 530590
rect 177297 530558 177331 530596
rect 177483 530567 177515 530589
rect 178309 530558 178343 530596
rect 178585 530558 178619 530596
rect 179137 530558 179171 530596
rect 179229 530558 179263 530596
rect 179783 530567 179815 530589
rect 180059 530567 180091 530589
rect 180296 530558 180330 530596
rect 181068 530568 181092 530590
rect 181842 530558 181876 530596
rect 181989 530558 182023 530596
rect 182633 530558 182667 530596
rect 183000 530568 183024 530590
rect 183093 530558 183127 530596
rect 183645 530558 183679 530596
rect 184749 530558 184783 530596
rect 185209 530558 185243 530596
rect 185761 530558 185795 530596
rect 186864 530568 186888 530590
rect 186957 530562 186991 530596
rect 187417 530558 187451 530596
rect 172209 530396 172483 530558
rect 172487 530422 173035 530558
rect 173037 530396 174139 530558
rect 174141 530396 174691 530558
rect 174787 530384 174873 530541
rect 174879 530422 175427 530558
rect 175521 530422 177359 530558
rect 175521 530376 175705 530422
rect 176271 530378 176457 530422
rect 177363 530384 177449 530541
rect 177656 530422 178349 530558
rect 177656 530376 177840 530422
rect 178373 530402 178647 530558
rect 178651 530422 179199 530558
rect 179201 530422 179749 530558
rect 179939 530384 180025 530541
rect 180213 530422 180993 530558
rect 181179 530422 181959 530558
rect 181961 530422 182509 530558
rect 180213 530376 180399 530422
rect 181773 530376 181959 530422
rect 182515 530384 182601 530541
rect 182605 530396 182971 530558
rect 183065 530422 183613 530558
rect 183617 530396 184719 530558
rect 184721 530396 185087 530558
rect 185091 530384 185177 530541
rect 185181 530422 185729 530558
rect 185733 530396 186835 530558
rect 187205 530396 187479 530558
rect 172209 529512 172483 529674
rect 172485 529512 173587 529674
rect 173589 529512 174691 529674
rect 175316 529648 175500 529694
rect 176423 529648 176609 529692
rect 177175 529648 177359 529694
rect 174807 529512 175500 529648
rect 175521 529512 177359 529648
rect 177363 529529 177449 529686
rect 178185 529648 178371 529694
rect 177591 529512 178371 529648
rect 178373 529648 178557 529694
rect 179123 529648 179309 529692
rect 181115 529648 181301 529692
rect 181867 529648 182051 529694
rect 178373 529512 180211 529648
rect 180213 529512 182051 529648
rect 182053 529512 182419 529674
rect 182515 529529 182601 529686
rect 182624 529648 182808 529694
rect 182624 529512 183317 529648
rect 183341 529512 184443 529674
rect 184445 529512 185547 529674
rect 185549 529512 186651 529674
rect 186653 529512 187203 529674
rect 187205 529512 187479 529674
rect 172237 529470 172271 529512
rect 172513 529470 172547 529512
rect 173617 529470 173651 529512
rect 174720 529480 174744 529502
rect 174813 529474 174847 529512
rect 174907 529479 174939 529501
rect 175549 529474 175583 529512
rect 175770 529470 175804 529508
rect 177480 529480 177504 529502
rect 177665 529470 177699 529508
rect 177757 529470 177791 529508
rect 178254 529474 178288 529512
rect 179596 529480 179620 529502
rect 179689 529470 179723 529508
rect 180057 529470 180091 529508
rect 180149 529474 180183 529512
rect 180241 529474 180275 529512
rect 180608 529480 180632 529502
rect 180701 529470 180735 529508
rect 182081 529474 182115 529512
rect 182448 529480 182472 529502
rect 182725 529470 182759 529508
rect 182817 529470 182851 529508
rect 183277 529474 183311 529512
rect 183369 529474 183403 529512
rect 183921 529470 183955 529508
rect 184473 529474 184507 529512
rect 185024 529480 185048 529502
rect 185209 529470 185243 529508
rect 185577 529474 185611 529512
rect 186313 529470 186347 529508
rect 186681 529474 186715 529512
rect 187051 529479 187083 529501
rect 187417 529470 187451 529512
rect 172209 529308 172483 529470
rect 172485 529308 173587 529470
rect 173589 529308 174691 529470
rect 174787 529296 174873 529453
rect 175107 529334 175887 529470
rect 175906 529334 177727 529470
rect 177729 529334 179567 529470
rect 175701 529288 175887 529334
rect 178631 529290 178817 529334
rect 179383 529288 179567 529334
rect 179661 529314 179935 529470
rect 179939 529296 180025 529453
rect 180029 529308 180579 529470
rect 180673 529334 182494 529470
rect 182513 529314 182787 529470
rect 182789 529308 183891 529470
rect 183893 529308 184995 529470
rect 185091 529296 185177 529453
rect 185181 529308 186283 529470
rect 186285 529308 187019 529470
rect 187205 529308 187479 529470
rect 172209 528424 172483 528586
rect 172485 528424 173587 528586
rect 173589 528424 174691 528586
rect 174693 528424 175795 528586
rect 175889 528424 176163 528580
rect 176165 528424 176439 528580
rect 177081 528560 177267 528606
rect 176487 528424 177267 528560
rect 177363 528441 177449 528598
rect 177472 528560 177656 528606
rect 177472 528424 178165 528560
rect 178373 528424 180194 528560
rect 180213 528424 180487 528580
rect 181391 528560 181577 528604
rect 182143 528560 182327 528606
rect 180489 528424 182327 528560
rect 182515 528441 182601 528598
rect 182605 528424 183707 528586
rect 183709 528424 184811 528586
rect 184813 528424 185915 528586
rect 185917 528424 187019 528586
rect 187205 528424 187479 528586
rect 172237 528382 172271 528424
rect 172513 528382 172547 528424
rect 173617 528382 173651 528424
rect 174721 528414 174755 528424
rect 174720 528392 174755 528414
rect 174721 528386 174755 528392
rect 174905 528382 174939 528420
rect 175824 528392 175848 528414
rect 175917 528386 175951 528424
rect 176008 528392 176032 528414
rect 176101 528382 176135 528420
rect 176193 528386 176227 528424
rect 177150 528386 177184 528424
rect 177296 528392 177320 528414
rect 178125 528382 178159 528424
rect 178217 528382 178251 528420
rect 178401 528386 178435 528424
rect 179008 528382 179042 528420
rect 179783 528391 179815 528413
rect 180057 528382 180091 528420
rect 180241 528386 180275 528424
rect 180517 528386 180551 528424
rect 180795 528391 180827 528413
rect 181032 528382 181066 528420
rect 181805 528382 181839 528420
rect 182359 528393 182391 528415
rect 182633 528386 182667 528424
rect 182909 528382 182943 528420
rect 183737 528386 183771 528424
rect 184013 528382 184047 528420
rect 184841 528386 184875 528424
rect 185209 528382 185243 528420
rect 185945 528386 185979 528424
rect 186313 528382 186347 528420
rect 187051 528391 187083 528415
rect 187417 528382 187451 528424
rect 172209 528220 172483 528382
rect 172485 528220 173587 528382
rect 173589 528220 174691 528382
rect 174787 528208 174873 528365
rect 174877 528220 175979 528382
rect 176073 528246 177911 528382
rect 176975 528202 177161 528246
rect 177727 528200 177911 528246
rect 177913 528226 178187 528382
rect 178189 528220 178923 528382
rect 178925 528246 179705 528382
rect 178925 528200 179111 528246
rect 179939 528208 180025 528365
rect 180029 528220 180763 528382
rect 180949 528246 181729 528382
rect 180949 528200 181135 528246
rect 181777 528220 182879 528382
rect 182881 528220 183983 528382
rect 183985 528220 185087 528382
rect 185091 528208 185177 528365
rect 185181 528220 186283 528382
rect 186285 528220 187019 528382
rect 187205 528220 187479 528382
rect 172209 527336 172483 527498
rect 172485 527336 173587 527498
rect 173589 527336 174691 527498
rect 174693 527336 175795 527498
rect 175797 527336 176347 527498
rect 176368 527472 176552 527518
rect 176368 527336 177061 527472
rect 177085 527336 177359 527498
rect 177363 527353 177449 527510
rect 177453 527336 178555 527498
rect 178557 527336 178923 527498
rect 178944 527472 179128 527518
rect 178944 527336 179637 527472
rect 179661 527336 180763 527498
rect 180765 527336 181867 527498
rect 181869 527336 182419 527498
rect 182515 527353 182601 527510
rect 182605 527336 183707 527498
rect 183709 527336 184811 527498
rect 184813 527336 185915 527498
rect 185917 527336 187019 527498
rect 187205 527336 187479 527498
rect 172237 527294 172271 527336
rect 172513 527294 172547 527336
rect 173617 527294 173651 527336
rect 174721 527326 174755 527336
rect 174720 527304 174755 527326
rect 174721 527298 174755 527304
rect 174905 527294 174939 527332
rect 175825 527298 175859 527336
rect 176009 527294 176043 527332
rect 177021 527298 177055 527336
rect 177113 527294 177147 527336
rect 177481 527298 177515 527336
rect 178217 527294 178251 527332
rect 178585 527298 178619 527336
rect 179321 527294 179355 527332
rect 179597 527298 179631 527336
rect 179689 527298 179723 527336
rect 179872 527304 179896 527326
rect 180057 527294 180091 527332
rect 180793 527298 180827 527336
rect 181161 527294 181195 527332
rect 181897 527298 181931 527336
rect 182265 527294 182299 527332
rect 182448 527304 182472 527326
rect 182633 527298 182667 527336
rect 183369 527294 183403 527332
rect 183737 527298 183771 527336
rect 184473 527294 184507 527332
rect 184841 527298 184875 527336
rect 185024 527304 185048 527326
rect 185209 527294 185243 527332
rect 185945 527298 185979 527336
rect 186313 527294 186347 527332
rect 187051 527303 187083 527327
rect 187417 527294 187451 527336
rect 172209 527132 172483 527294
rect 172485 527132 173587 527294
rect 173589 527132 174691 527294
rect 174787 527120 174873 527277
rect 174877 527132 175979 527294
rect 175981 527132 177083 527294
rect 177085 527132 178187 527294
rect 178189 527132 179291 527294
rect 179293 527132 179843 527294
rect 179939 527120 180025 527277
rect 180029 527132 181131 527294
rect 181133 527132 182235 527294
rect 182237 527132 183339 527294
rect 183341 527132 184443 527294
rect 184445 527132 184995 527294
rect 185091 527120 185177 527277
rect 185181 527132 186283 527294
rect 186285 527132 187019 527294
rect 187205 527132 187479 527294
rect 172209 526248 172483 526410
rect 172485 526248 173587 526410
rect 173589 526248 174691 526410
rect 174693 526248 175795 526410
rect 175797 526248 176899 526410
rect 176901 526248 177267 526410
rect 177363 526265 177449 526422
rect 177453 526248 178555 526410
rect 178557 526248 179659 526410
rect 179661 526248 180763 526410
rect 180765 526248 181867 526410
rect 181869 526248 182419 526410
rect 182515 526265 182601 526422
rect 182605 526248 183707 526410
rect 183709 526248 184811 526410
rect 184813 526248 185915 526410
rect 185917 526248 187019 526410
rect 187205 526248 187479 526410
rect 172237 526206 172271 526248
rect 172513 526206 172547 526248
rect 173617 526206 173651 526248
rect 174721 526238 174755 526248
rect 174720 526216 174755 526238
rect 174721 526210 174755 526216
rect 174905 526206 174939 526244
rect 175825 526210 175859 526248
rect 176009 526206 176043 526244
rect 176929 526210 176963 526248
rect 177113 526206 177147 526244
rect 177296 526216 177320 526238
rect 177481 526210 177515 526248
rect 178217 526206 178251 526244
rect 178585 526210 178619 526248
rect 179321 526206 179355 526244
rect 179689 526210 179723 526248
rect 179872 526216 179896 526238
rect 180057 526206 180091 526244
rect 180793 526210 180827 526248
rect 181161 526206 181195 526244
rect 181897 526210 181931 526248
rect 182265 526206 182299 526244
rect 182448 526216 182472 526238
rect 182633 526210 182667 526248
rect 183369 526206 183403 526244
rect 183737 526210 183771 526248
rect 184473 526206 184507 526244
rect 184841 526210 184875 526248
rect 185024 526216 185048 526238
rect 185209 526206 185243 526244
rect 185945 526210 185979 526248
rect 186313 526206 186347 526244
rect 187051 526215 187083 526239
rect 187417 526206 187451 526248
rect 172209 526044 172483 526206
rect 172485 526044 173587 526206
rect 173589 526044 174691 526206
rect 174787 526032 174873 526189
rect 174877 526044 175979 526206
rect 175981 526044 177083 526206
rect 177085 526044 178187 526206
rect 178189 526044 179291 526206
rect 179293 526044 179843 526206
rect 179939 526032 180025 526189
rect 180029 526044 181131 526206
rect 181133 526044 182235 526206
rect 182237 526044 183339 526206
rect 183341 526044 184443 526206
rect 184445 526044 184995 526206
rect 185091 526032 185177 526189
rect 185181 526044 186283 526206
rect 186285 526044 187019 526206
rect 187205 526044 187479 526206
rect 172209 525160 172483 525322
rect 172485 525160 173587 525322
rect 173589 525160 174691 525322
rect 174693 525160 175795 525322
rect 175797 525160 176899 525322
rect 176901 525160 177267 525322
rect 177363 525177 177449 525334
rect 177453 525160 178555 525322
rect 178557 525160 179659 525322
rect 179661 525160 180763 525322
rect 180765 525160 181867 525322
rect 181869 525160 182419 525322
rect 182515 525177 182601 525334
rect 182605 525160 183707 525322
rect 183709 525160 184811 525322
rect 184813 525160 185915 525322
rect 185917 525160 187019 525322
rect 187205 525160 187479 525322
rect 172237 525118 172271 525160
rect 172513 525118 172547 525160
rect 173617 525118 173651 525160
rect 174721 525150 174755 525160
rect 174720 525128 174755 525150
rect 174721 525122 174755 525128
rect 174905 525118 174939 525156
rect 175825 525122 175859 525160
rect 176009 525118 176043 525156
rect 176929 525122 176963 525160
rect 177113 525118 177147 525156
rect 177296 525128 177320 525150
rect 177481 525122 177515 525160
rect 178217 525118 178251 525156
rect 178585 525122 178619 525160
rect 179321 525118 179355 525156
rect 179689 525122 179723 525160
rect 179872 525128 179896 525150
rect 180057 525118 180091 525156
rect 180793 525122 180827 525160
rect 181161 525118 181195 525156
rect 181897 525122 181931 525160
rect 182265 525118 182299 525156
rect 182448 525128 182472 525150
rect 182633 525122 182667 525160
rect 183369 525118 183403 525156
rect 183737 525122 183771 525160
rect 184473 525118 184507 525156
rect 184841 525122 184875 525160
rect 185024 525128 185048 525150
rect 185209 525118 185243 525156
rect 185945 525122 185979 525160
rect 186313 525118 186347 525156
rect 187051 525127 187083 525151
rect 187417 525118 187451 525160
rect 172209 524956 172483 525118
rect 172485 524956 173587 525118
rect 173589 524956 174691 525118
rect 174787 524944 174873 525101
rect 174877 524956 175979 525118
rect 175981 524956 177083 525118
rect 177085 524956 178187 525118
rect 178189 524956 179291 525118
rect 179293 524956 179843 525118
rect 179939 524944 180025 525101
rect 180029 524956 181131 525118
rect 181133 524956 182235 525118
rect 182237 524956 183339 525118
rect 183341 524956 184443 525118
rect 184445 524956 184995 525118
rect 185091 524944 185177 525101
rect 185181 524956 186283 525118
rect 186285 524956 187019 525118
rect 187205 524956 187479 525118
rect 172209 524072 172483 524234
rect 172485 524072 173587 524234
rect 173589 524072 174691 524234
rect 174693 524072 175795 524234
rect 175797 524072 176899 524234
rect 176901 524072 177267 524234
rect 177363 524089 177449 524246
rect 177453 524072 178555 524234
rect 178557 524072 179659 524234
rect 179661 524072 180763 524234
rect 180765 524072 181867 524234
rect 181869 524072 182419 524234
rect 182515 524089 182601 524246
rect 182605 524072 183707 524234
rect 183709 524072 184811 524234
rect 184813 524072 185915 524234
rect 185917 524072 187019 524234
rect 187205 524072 187479 524234
rect 172237 524030 172271 524072
rect 172513 524030 172547 524072
rect 173617 524030 173651 524072
rect 174721 524062 174755 524072
rect 174720 524040 174755 524062
rect 174721 524034 174755 524040
rect 174905 524030 174939 524068
rect 175825 524034 175859 524072
rect 176009 524030 176043 524068
rect 176929 524034 176963 524072
rect 177113 524030 177147 524068
rect 177296 524040 177320 524062
rect 177481 524034 177515 524072
rect 178217 524030 178251 524068
rect 178585 524034 178619 524072
rect 179321 524030 179355 524068
rect 179689 524034 179723 524072
rect 179872 524040 179896 524062
rect 180057 524030 180091 524068
rect 180793 524034 180827 524072
rect 181161 524030 181195 524068
rect 181897 524034 181931 524072
rect 182265 524030 182299 524068
rect 182448 524040 182472 524062
rect 182633 524034 182667 524072
rect 183369 524030 183403 524068
rect 183737 524034 183771 524072
rect 184473 524030 184507 524068
rect 184841 524034 184875 524072
rect 185024 524040 185048 524062
rect 185209 524030 185243 524068
rect 185945 524034 185979 524072
rect 186313 524030 186347 524068
rect 187051 524039 187083 524063
rect 187417 524030 187451 524072
rect 172209 523868 172483 524030
rect 172485 523868 173587 524030
rect 173589 523868 174691 524030
rect 174787 523856 174873 524013
rect 174877 523868 175979 524030
rect 175981 523868 177083 524030
rect 177085 523868 178187 524030
rect 178189 523868 179291 524030
rect 179293 523868 179843 524030
rect 179939 523856 180025 524013
rect 180029 523868 181131 524030
rect 181133 523868 182235 524030
rect 182237 523868 183339 524030
rect 183341 523868 184443 524030
rect 184445 523868 184995 524030
rect 185091 523856 185177 524013
rect 185181 523868 186283 524030
rect 186285 523868 187019 524030
rect 187205 523868 187479 524030
rect 172209 522984 172483 523146
rect 172485 522984 173587 523146
rect 173589 522984 174691 523146
rect 174693 522984 175795 523146
rect 175797 522984 176899 523146
rect 176901 522984 177267 523146
rect 177363 523001 177449 523158
rect 177453 522984 178555 523146
rect 178557 522984 179659 523146
rect 179661 522984 180763 523146
rect 180765 522984 181867 523146
rect 181869 522984 182419 523146
rect 182515 523001 182601 523158
rect 182605 522984 183707 523146
rect 183709 522984 184811 523146
rect 184813 522984 185915 523146
rect 185917 522984 187019 523146
rect 187205 522984 187479 523146
rect 172237 522942 172271 522984
rect 172513 522942 172547 522984
rect 173617 522942 173651 522984
rect 174721 522974 174755 522984
rect 174720 522952 174755 522974
rect 174721 522946 174755 522952
rect 174905 522942 174939 522980
rect 175825 522946 175859 522984
rect 176009 522942 176043 522980
rect 176929 522946 176963 522984
rect 177113 522942 177147 522980
rect 177296 522952 177320 522974
rect 177481 522946 177515 522984
rect 178217 522942 178251 522980
rect 178585 522946 178619 522984
rect 179321 522942 179355 522980
rect 179689 522946 179723 522984
rect 179872 522952 179896 522974
rect 180057 522942 180091 522980
rect 180793 522946 180827 522984
rect 181161 522942 181195 522980
rect 181897 522946 181931 522984
rect 182265 522942 182299 522980
rect 182448 522952 182472 522974
rect 182633 522946 182667 522984
rect 183369 522942 183403 522980
rect 183737 522946 183771 522984
rect 184473 522942 184507 522980
rect 184841 522946 184875 522984
rect 185024 522952 185048 522974
rect 185209 522942 185243 522980
rect 185945 522946 185979 522984
rect 186313 522942 186347 522980
rect 187051 522951 187083 522975
rect 187417 522942 187451 522984
rect 172209 522780 172483 522942
rect 172485 522780 173587 522942
rect 173589 522780 174691 522942
rect 174787 522768 174873 522925
rect 174877 522780 175979 522942
rect 175981 522780 177083 522942
rect 177085 522780 178187 522942
rect 178189 522780 179291 522942
rect 179293 522780 179843 522942
rect 179939 522768 180025 522925
rect 180029 522780 181131 522942
rect 181133 522780 182235 522942
rect 182237 522780 183339 522942
rect 183341 522780 184443 522942
rect 184445 522780 184995 522942
rect 185091 522768 185177 522925
rect 185181 522780 186283 522942
rect 186285 522780 187019 522942
rect 187205 522780 187479 522942
rect 172209 521896 172483 522058
rect 172485 521896 173587 522058
rect 173589 521896 174691 522058
rect 174693 521896 175795 522058
rect 175797 521896 176899 522058
rect 176901 521896 177267 522058
rect 177363 521913 177449 522070
rect 177453 521896 178555 522058
rect 178557 521896 179659 522058
rect 179661 521896 180763 522058
rect 180765 521896 181867 522058
rect 181869 521896 182419 522058
rect 182515 521913 182601 522070
rect 182605 521896 183707 522058
rect 183709 521896 184811 522058
rect 184813 521896 185915 522058
rect 185917 521896 187019 522058
rect 187205 521896 187479 522058
rect 172237 521854 172271 521896
rect 172513 521854 172547 521896
rect 173617 521854 173651 521896
rect 174721 521886 174755 521896
rect 174720 521864 174755 521886
rect 174721 521858 174755 521864
rect 174905 521854 174939 521892
rect 175825 521858 175859 521896
rect 176009 521854 176043 521892
rect 176929 521858 176963 521896
rect 177113 521854 177147 521892
rect 177296 521864 177320 521886
rect 177481 521858 177515 521896
rect 178217 521854 178251 521892
rect 178585 521858 178619 521896
rect 179321 521854 179355 521892
rect 179689 521858 179723 521896
rect 179872 521864 179896 521886
rect 180057 521854 180091 521892
rect 180793 521858 180827 521896
rect 181161 521854 181195 521892
rect 181897 521858 181931 521896
rect 182265 521854 182299 521892
rect 182448 521864 182472 521886
rect 182633 521858 182667 521896
rect 183369 521854 183403 521892
rect 183737 521858 183771 521896
rect 184473 521854 184507 521892
rect 184841 521858 184875 521896
rect 185024 521864 185048 521886
rect 185209 521854 185243 521892
rect 185945 521858 185979 521896
rect 186313 521854 186347 521892
rect 187051 521863 187083 521887
rect 187417 521854 187451 521896
rect 172209 521692 172483 521854
rect 172485 521692 173587 521854
rect 173589 521692 174691 521854
rect 174787 521680 174873 521837
rect 174877 521692 175979 521854
rect 175981 521692 177083 521854
rect 177085 521692 178187 521854
rect 178189 521692 179291 521854
rect 179293 521692 179843 521854
rect 179939 521680 180025 521837
rect 180029 521692 181131 521854
rect 181133 521692 182235 521854
rect 182237 521692 183339 521854
rect 183341 521692 184443 521854
rect 184445 521692 184995 521854
rect 185091 521680 185177 521837
rect 185181 521692 186283 521854
rect 186285 521692 187019 521854
rect 187205 521692 187479 521854
rect 172209 520808 172483 520970
rect 172485 520808 173587 520970
rect 173589 520808 174691 520970
rect 174693 520808 175795 520970
rect 175797 520808 176899 520970
rect 176901 520808 177267 520970
rect 177363 520825 177449 520982
rect 177453 520808 178555 520970
rect 178557 520808 179659 520970
rect 179661 520808 180763 520970
rect 180765 520808 181867 520970
rect 181869 520808 182419 520970
rect 182515 520825 182601 520982
rect 182605 520808 183707 520970
rect 183709 520808 184811 520970
rect 184813 520808 185915 520970
rect 185917 520808 187019 520970
rect 187205 520808 187479 520970
rect 172237 520766 172271 520808
rect 172513 520766 172547 520808
rect 173617 520766 173651 520808
rect 174721 520798 174755 520808
rect 174720 520776 174755 520798
rect 174721 520770 174755 520776
rect 174905 520766 174939 520804
rect 175825 520770 175859 520808
rect 176009 520766 176043 520804
rect 176929 520770 176963 520808
rect 177113 520766 177147 520804
rect 177296 520776 177320 520798
rect 177481 520770 177515 520808
rect 178217 520766 178251 520804
rect 178585 520770 178619 520808
rect 179321 520766 179355 520804
rect 179689 520770 179723 520808
rect 179872 520776 179896 520798
rect 180057 520766 180091 520804
rect 180793 520770 180827 520808
rect 181161 520766 181195 520804
rect 181897 520770 181931 520808
rect 182265 520766 182299 520804
rect 182448 520776 182472 520798
rect 182633 520770 182667 520808
rect 183369 520766 183403 520804
rect 183737 520770 183771 520808
rect 184473 520766 184507 520804
rect 184841 520770 184875 520808
rect 185024 520776 185048 520798
rect 185209 520766 185243 520804
rect 185945 520770 185979 520808
rect 186313 520766 186347 520804
rect 187051 520775 187083 520799
rect 187417 520766 187451 520808
rect 172209 520604 172483 520766
rect 172485 520604 173587 520766
rect 173589 520604 174691 520766
rect 174787 520592 174873 520749
rect 174877 520604 175979 520766
rect 175981 520604 177083 520766
rect 177085 520604 178187 520766
rect 178189 520604 179291 520766
rect 179293 520604 179843 520766
rect 179939 520592 180025 520749
rect 180029 520604 181131 520766
rect 181133 520604 182235 520766
rect 182237 520604 183339 520766
rect 183341 520604 184443 520766
rect 184445 520604 184995 520766
rect 185091 520592 185177 520749
rect 185181 520604 186283 520766
rect 186285 520604 187019 520766
rect 187205 520604 187479 520766
rect 172209 519720 172483 519882
rect 172485 519720 173587 519882
rect 173589 519720 174691 519882
rect 174693 519720 175795 519882
rect 175797 519720 176899 519882
rect 176901 519720 177267 519882
rect 177363 519737 177449 519894
rect 177453 519720 178555 519882
rect 178557 519720 179659 519882
rect 179661 519720 180763 519882
rect 180765 519720 181867 519882
rect 181869 519720 182419 519882
rect 182515 519737 182601 519894
rect 182605 519720 183707 519882
rect 183709 519720 184811 519882
rect 184813 519720 185915 519882
rect 185917 519720 187019 519882
rect 187205 519720 187479 519882
rect 172237 519678 172271 519720
rect 172513 519678 172547 519720
rect 173617 519678 173651 519720
rect 174721 519710 174755 519720
rect 174720 519688 174755 519710
rect 174721 519682 174755 519688
rect 174905 519678 174939 519716
rect 175825 519682 175859 519720
rect 176009 519678 176043 519716
rect 176929 519682 176963 519720
rect 177113 519678 177147 519716
rect 177296 519688 177320 519710
rect 177481 519682 177515 519720
rect 178217 519678 178251 519716
rect 178585 519682 178619 519720
rect 179321 519678 179355 519716
rect 179689 519682 179723 519720
rect 179872 519688 179896 519710
rect 180057 519678 180091 519716
rect 180793 519682 180827 519720
rect 181161 519678 181195 519716
rect 181897 519682 181931 519720
rect 182265 519678 182299 519716
rect 182448 519688 182472 519710
rect 182633 519682 182667 519720
rect 183369 519678 183403 519716
rect 183737 519682 183771 519720
rect 184473 519678 184507 519716
rect 184841 519682 184875 519720
rect 185024 519688 185048 519710
rect 185209 519678 185243 519716
rect 185945 519682 185979 519720
rect 186313 519678 186347 519716
rect 187051 519687 187083 519711
rect 187417 519678 187451 519720
rect 172209 519516 172483 519678
rect 172485 519516 173587 519678
rect 173589 519516 174691 519678
rect 174787 519504 174873 519661
rect 174877 519516 175979 519678
rect 175981 519516 177083 519678
rect 177085 519516 178187 519678
rect 178189 519516 179291 519678
rect 179293 519516 179843 519678
rect 179939 519504 180025 519661
rect 180029 519516 181131 519678
rect 181133 519516 182235 519678
rect 182237 519516 183339 519678
rect 183341 519516 184443 519678
rect 184445 519516 184995 519678
rect 185091 519504 185177 519661
rect 185181 519516 186283 519678
rect 186285 519516 187019 519678
rect 187205 519516 187479 519678
rect 172209 518632 172483 518794
rect 172485 518632 173587 518794
rect 173589 518632 174691 518794
rect 174693 518632 175795 518794
rect 175797 518632 176899 518794
rect 176901 518632 177267 518794
rect 177363 518649 177449 518806
rect 177453 518632 178555 518794
rect 178557 518632 179659 518794
rect 179661 518632 180763 518794
rect 180765 518632 181867 518794
rect 181869 518632 182419 518794
rect 182515 518649 182601 518806
rect 182605 518632 183707 518794
rect 183709 518632 184811 518794
rect 184813 518632 185915 518794
rect 185917 518632 187019 518794
rect 187205 518632 187479 518794
rect 172237 518590 172271 518632
rect 172513 518590 172547 518632
rect 173617 518590 173651 518632
rect 174721 518622 174755 518632
rect 174720 518600 174755 518622
rect 174721 518594 174755 518600
rect 174905 518590 174939 518628
rect 175825 518594 175859 518632
rect 176009 518590 176043 518628
rect 176929 518594 176963 518632
rect 177113 518590 177147 518628
rect 177296 518600 177320 518622
rect 177481 518594 177515 518632
rect 178217 518590 178251 518628
rect 178585 518594 178619 518632
rect 179321 518590 179355 518628
rect 179689 518594 179723 518632
rect 179872 518600 179896 518622
rect 180057 518590 180091 518628
rect 180793 518594 180827 518632
rect 181161 518590 181195 518628
rect 181897 518594 181931 518632
rect 182265 518590 182299 518628
rect 182448 518600 182472 518622
rect 182633 518594 182667 518632
rect 183369 518590 183403 518628
rect 183737 518594 183771 518632
rect 184473 518590 184507 518628
rect 184841 518594 184875 518632
rect 185024 518600 185048 518622
rect 185209 518590 185243 518628
rect 185945 518594 185979 518632
rect 186313 518590 186347 518628
rect 187051 518599 187083 518623
rect 187417 518590 187451 518632
rect 172209 518428 172483 518590
rect 172485 518428 173587 518590
rect 173589 518428 174691 518590
rect 174787 518416 174873 518573
rect 174877 518428 175979 518590
rect 175981 518428 177083 518590
rect 177085 518428 178187 518590
rect 178189 518428 179291 518590
rect 179293 518428 179843 518590
rect 179939 518416 180025 518573
rect 180029 518428 181131 518590
rect 181133 518428 182235 518590
rect 182237 518428 183339 518590
rect 183341 518428 184443 518590
rect 184445 518428 184995 518590
rect 185091 518416 185177 518573
rect 185181 518428 186283 518590
rect 186285 518428 187019 518590
rect 187205 518428 187479 518590
rect 172209 517544 172483 517706
rect 172485 517544 173587 517706
rect 173589 517544 174691 517706
rect 174693 517544 175795 517706
rect 175797 517544 176899 517706
rect 176901 517544 177267 517706
rect 177363 517561 177449 517718
rect 177453 517544 178555 517706
rect 178557 517544 179659 517706
rect 179661 517544 180763 517706
rect 180765 517544 181867 517706
rect 181869 517544 182419 517706
rect 182515 517561 182601 517718
rect 182605 517544 183707 517706
rect 183709 517544 184811 517706
rect 184813 517544 185915 517706
rect 185917 517544 187019 517706
rect 187205 517544 187479 517706
rect 172237 517502 172271 517544
rect 172513 517502 172547 517544
rect 173617 517502 173651 517544
rect 174721 517534 174755 517544
rect 174720 517512 174755 517534
rect 174721 517506 174755 517512
rect 174905 517502 174939 517540
rect 175825 517506 175859 517544
rect 176009 517502 176043 517540
rect 176929 517506 176963 517544
rect 177113 517502 177147 517540
rect 177296 517512 177320 517534
rect 177481 517506 177515 517544
rect 178217 517502 178251 517540
rect 178585 517506 178619 517544
rect 179321 517502 179355 517540
rect 179689 517506 179723 517544
rect 179872 517512 179896 517534
rect 180057 517502 180091 517540
rect 180793 517506 180827 517544
rect 181161 517502 181195 517540
rect 181897 517506 181931 517544
rect 182265 517502 182299 517540
rect 182448 517512 182472 517534
rect 182633 517506 182667 517544
rect 183369 517502 183403 517540
rect 183737 517506 183771 517544
rect 184473 517502 184507 517540
rect 184841 517506 184875 517544
rect 185024 517512 185048 517534
rect 185209 517502 185243 517540
rect 185945 517506 185979 517544
rect 186313 517502 186347 517540
rect 187051 517511 187083 517535
rect 187417 517502 187451 517544
rect 172209 517340 172483 517502
rect 172485 517340 173587 517502
rect 173589 517340 174691 517502
rect 174787 517328 174873 517485
rect 174877 517340 175979 517502
rect 175981 517340 177083 517502
rect 177085 517340 178187 517502
rect 178189 517340 179291 517502
rect 179293 517340 179843 517502
rect 179939 517328 180025 517485
rect 180029 517340 181131 517502
rect 181133 517340 182235 517502
rect 182237 517340 183339 517502
rect 183341 517340 184443 517502
rect 184445 517340 184995 517502
rect 185091 517328 185177 517485
rect 185181 517340 186283 517502
rect 186285 517340 187019 517502
rect 187205 517340 187479 517502
rect 172209 516456 172483 516618
rect 172485 516456 173587 516618
rect 173589 516456 174691 516618
rect 174693 516456 175795 516618
rect 175797 516456 176899 516618
rect 176901 516456 177267 516618
rect 177363 516473 177449 516630
rect 177453 516456 178555 516618
rect 178557 516456 179659 516618
rect 179661 516456 180763 516618
rect 180765 516456 181867 516618
rect 181869 516456 182419 516618
rect 182515 516473 182601 516630
rect 182605 516456 183707 516618
rect 183709 516456 184811 516618
rect 184813 516456 185915 516618
rect 185917 516456 187019 516618
rect 187205 516456 187479 516618
rect 172237 516414 172271 516456
rect 172513 516414 172547 516456
rect 173617 516414 173651 516456
rect 174721 516446 174755 516456
rect 174720 516424 174755 516446
rect 174721 516418 174755 516424
rect 174905 516414 174939 516452
rect 175825 516418 175859 516456
rect 176009 516414 176043 516452
rect 176929 516418 176963 516456
rect 177113 516414 177147 516452
rect 177296 516424 177320 516446
rect 177481 516418 177515 516456
rect 178217 516414 178251 516452
rect 178585 516418 178619 516456
rect 179321 516414 179355 516452
rect 179689 516418 179723 516456
rect 179872 516424 179896 516446
rect 180057 516414 180091 516452
rect 180793 516418 180827 516456
rect 181161 516414 181195 516452
rect 181897 516418 181931 516456
rect 182265 516414 182299 516452
rect 182448 516424 182472 516446
rect 182633 516418 182667 516456
rect 183369 516414 183403 516452
rect 183737 516418 183771 516456
rect 184473 516414 184507 516452
rect 184841 516418 184875 516456
rect 185024 516424 185048 516446
rect 185209 516414 185243 516452
rect 185945 516418 185979 516456
rect 186313 516414 186347 516452
rect 187051 516423 187083 516447
rect 187417 516414 187451 516456
rect 172209 516252 172483 516414
rect 172485 516252 173587 516414
rect 173589 516252 174691 516414
rect 174787 516240 174873 516397
rect 174877 516252 175979 516414
rect 175981 516252 177083 516414
rect 177085 516252 178187 516414
rect 178189 516252 179291 516414
rect 179293 516252 179843 516414
rect 179939 516240 180025 516397
rect 180029 516252 181131 516414
rect 181133 516252 182235 516414
rect 182237 516252 183339 516414
rect 183341 516252 184443 516414
rect 184445 516252 184995 516414
rect 185091 516240 185177 516397
rect 185181 516252 186283 516414
rect 186285 516252 187019 516414
rect 187205 516252 187479 516414
rect 172209 515368 172483 515530
rect 172485 515368 173219 515530
rect 173405 515368 173953 515504
rect 173957 515368 174691 515530
rect 174787 515385 174873 515542
rect 174877 515368 175979 515530
rect 175981 515368 177083 515530
rect 177085 515368 177359 515530
rect 177363 515385 177449 515542
rect 177453 515368 178555 515530
rect 178557 515368 179659 515530
rect 179661 515368 179935 515530
rect 179939 515385 180025 515542
rect 180029 515368 181131 515530
rect 181133 515368 181867 515530
rect 182053 515368 182327 515524
rect 182515 515385 182601 515542
rect 182605 515368 183707 515530
rect 183709 515368 184811 515530
rect 184813 515368 185087 515530
rect 185091 515385 185177 515542
rect 185181 515368 186283 515530
rect 186377 515368 186925 515504
rect 186929 515368 187203 515530
rect 187205 515368 187479 515530
rect 172237 515330 172271 515368
rect 172513 515330 172547 515368
rect 173251 515337 173283 515359
rect 173433 515330 173467 515368
rect 173985 515330 174019 515368
rect 174720 515336 174744 515358
rect 174905 515330 174939 515368
rect 176009 515330 176043 515368
rect 177113 515330 177147 515368
rect 177481 515330 177515 515368
rect 178585 515330 178619 515368
rect 179689 515330 179723 515368
rect 180057 515330 180091 515368
rect 181161 515330 181195 515368
rect 181899 515337 181931 515359
rect 182263 515330 182297 515368
rect 182359 515337 182391 515359
rect 182633 515330 182667 515368
rect 183737 515330 183771 515368
rect 184841 515330 184875 515368
rect 185209 515330 185243 515368
rect 186312 515336 186336 515358
rect 186405 515330 186439 515368
rect 186957 515330 186991 515368
rect 187417 515330 187451 515368
<< nmos >>
rect 164730 540047 164760 541047
rect 164937 540054 164967 541054
rect 165033 540054 165063 541054
rect 165129 540054 165159 541054
rect 165225 540054 165255 541054
rect 165321 540054 165351 541054
rect 165417 540054 165447 541054
rect 165513 540054 165543 541054
rect 165609 540054 165639 541054
rect 165705 540054 165735 541054
rect 165801 540054 165831 541054
rect 165897 540054 165927 541054
rect 165993 540054 166023 541054
rect 166210 540047 166240 540247
rect 166410 540047 166440 541047
rect 168530 540047 168560 541047
rect 168737 540054 168767 541054
rect 168833 540054 168863 541054
rect 168929 540054 168959 541054
rect 169025 540054 169055 541054
rect 169121 540054 169151 541054
rect 169217 540054 169247 541054
rect 169313 540054 169343 541054
rect 169409 540054 169439 541054
rect 169505 540054 169535 541054
rect 169601 540054 169631 541054
rect 169697 540054 169727 541054
rect 169793 540054 169823 541054
rect 170010 540047 170040 540247
rect 170210 540047 170240 541047
rect 172230 540047 172260 541047
rect 172437 540054 172467 541054
rect 172533 540054 172563 541054
rect 172629 540054 172659 541054
rect 172725 540054 172755 541054
rect 172821 540054 172851 541054
rect 172917 540054 172947 541054
rect 173013 540054 173043 541054
rect 173109 540054 173139 541054
rect 173205 540054 173235 541054
rect 173301 540054 173331 541054
rect 173397 540054 173427 541054
rect 173493 540054 173523 541054
rect 173710 540047 173740 540247
rect 173910 540047 173940 541047
rect 175730 540047 175760 541047
rect 175937 540054 175967 541054
rect 176033 540054 176063 541054
rect 176129 540054 176159 541054
rect 176225 540054 176255 541054
rect 176321 540054 176351 541054
rect 176417 540054 176447 541054
rect 176513 540054 176543 541054
rect 176609 540054 176639 541054
rect 176705 540054 176735 541054
rect 176801 540054 176831 541054
rect 176897 540054 176927 541054
rect 176993 540054 177023 541054
rect 177210 540047 177240 540247
rect 177410 540047 177440 541047
rect 179330 540047 179360 541047
rect 179537 540054 179567 541054
rect 179633 540054 179663 541054
rect 179729 540054 179759 541054
rect 179825 540054 179855 541054
rect 179921 540054 179951 541054
rect 180017 540054 180047 541054
rect 180113 540054 180143 541054
rect 180209 540054 180239 541054
rect 180305 540054 180335 541054
rect 180401 540054 180431 541054
rect 180497 540054 180527 541054
rect 180593 540054 180623 541054
rect 180810 540047 180840 540247
rect 181010 540047 181040 541047
rect 182630 540047 182660 541047
rect 182837 540054 182867 541054
rect 182933 540054 182963 541054
rect 183029 540054 183059 541054
rect 183125 540054 183155 541054
rect 183221 540054 183251 541054
rect 183317 540054 183347 541054
rect 183413 540054 183443 541054
rect 183509 540054 183539 541054
rect 183605 540054 183635 541054
rect 183701 540054 183731 541054
rect 183797 540054 183827 541054
rect 183893 540054 183923 541054
rect 184110 540047 184140 540247
rect 184310 540047 184340 541047
rect 185930 540047 185960 541047
rect 186137 540054 186167 541054
rect 186233 540054 186263 541054
rect 186329 540054 186359 541054
rect 186425 540054 186455 541054
rect 186521 540054 186551 541054
rect 186617 540054 186647 541054
rect 186713 540054 186743 541054
rect 186809 540054 186839 541054
rect 186905 540054 186935 541054
rect 187001 540054 187031 541054
rect 187097 540054 187127 541054
rect 187193 540054 187223 541054
rect 187410 540047 187440 540247
rect 187610 540047 187640 541047
rect 189230 540047 189260 541047
rect 189437 540054 189467 541054
rect 189533 540054 189563 541054
rect 189629 540054 189659 541054
rect 189725 540054 189755 541054
rect 189821 540054 189851 541054
rect 189917 540054 189947 541054
rect 190013 540054 190043 541054
rect 190109 540054 190139 541054
rect 190205 540054 190235 541054
rect 190301 540054 190331 541054
rect 190397 540054 190427 541054
rect 190493 540054 190523 541054
rect 190710 540047 190740 540247
rect 190910 540047 190940 541047
rect 158710 538197 158910 538397
rect 159086 538197 159286 538397
rect 159344 538197 159544 538397
rect 159602 538197 159802 538397
rect 159860 538197 160060 538397
rect 160118 538197 160318 538397
rect 160376 538197 160576 538397
rect 160634 538197 160834 538397
rect 160892 538197 161092 538397
rect 161150 538197 161350 538397
rect 161530 538197 161730 538397
rect 161930 538197 162130 538397
rect 162310 538197 162510 538397
<< scnmos >>
rect 172287 530422 172405 530532
rect 172571 530448 172601 530532
rect 172657 530448 172687 530532
rect 172743 530448 172773 530532
rect 172829 530448 172859 530532
rect 172926 530448 172956 530532
rect 173115 530422 174061 530532
rect 174219 530422 174613 530532
rect 174963 530448 174993 530532
rect 175049 530448 175079 530532
rect 175135 530448 175165 530532
rect 175221 530448 175251 530532
rect 175318 530448 175348 530532
rect 175599 530402 175629 530532
rect 175807 530448 175837 530532
rect 175898 530448 175928 530532
rect 176047 530448 176077 530532
rect 176143 530460 176173 530532
rect 176252 530460 176282 530532
rect 176351 530404 176381 530532
rect 176483 530448 176513 530532
rect 176555 530448 176585 530532
rect 176721 530460 176751 530532
rect 176817 530460 176847 530532
rect 176912 530448 176942 530532
rect 177167 530448 177197 530532
rect 177251 530448 177281 530532
rect 177734 530402 177764 530532
rect 177829 530448 177929 530532
rect 178087 530448 178187 530532
rect 178241 530448 178271 530532
rect 178451 530428 178481 530532
rect 178539 530428 178569 530532
rect 178735 530448 178765 530532
rect 178821 530448 178851 530532
rect 178907 530448 178937 530532
rect 178993 530448 179023 530532
rect 179090 530448 179120 530532
rect 179280 530448 179310 530532
rect 179377 530448 179407 530532
rect 179463 530448 179493 530532
rect 179549 530448 179579 530532
rect 179635 530448 179665 530532
rect 180291 530402 180321 530532
rect 180400 530448 180430 530532
rect 180496 530448 180526 530532
rect 180621 530448 180651 530532
rect 180717 530448 180747 530532
rect 180885 530448 180915 530532
rect 181257 530448 181287 530532
rect 181425 530448 181455 530532
rect 181521 530448 181551 530532
rect 181646 530448 181676 530532
rect 181742 530448 181772 530532
rect 181851 530402 181881 530532
rect 182040 530448 182070 530532
rect 182137 530448 182167 530532
rect 182223 530448 182253 530532
rect 182309 530448 182339 530532
rect 182395 530448 182425 530532
rect 182683 530422 182893 530532
rect 183144 530448 183174 530532
rect 183241 530448 183271 530532
rect 183327 530448 183357 530532
rect 183413 530448 183443 530532
rect 183499 530448 183529 530532
rect 183695 530422 184641 530532
rect 184799 530422 185009 530532
rect 185260 530448 185290 530532
rect 185357 530448 185387 530532
rect 185443 530448 185473 530532
rect 185529 530448 185559 530532
rect 185615 530448 185645 530532
rect 185811 530422 186757 530532
rect 187283 530422 187401 530532
rect 172287 529538 172405 529648
rect 172563 529538 173509 529648
rect 173667 529538 174613 529648
rect 174885 529538 174915 529622
rect 174969 529538 175069 529622
rect 175227 529538 175327 529622
rect 175392 529538 175422 529668
rect 175599 529538 175629 529622
rect 175683 529538 175713 529622
rect 175938 529538 175968 529622
rect 176033 529538 176063 529610
rect 176129 529538 176159 529610
rect 176295 529538 176325 529622
rect 176367 529538 176397 529622
rect 176499 529538 176529 529666
rect 176598 529538 176628 529610
rect 176707 529538 176737 529610
rect 176803 529538 176833 529622
rect 176952 529538 176982 529622
rect 177043 529538 177073 529622
rect 177251 529538 177281 529668
rect 177669 529538 177699 529622
rect 177837 529538 177867 529622
rect 177933 529538 177963 529622
rect 178058 529538 178088 529622
rect 178154 529538 178184 529622
rect 178263 529538 178293 529668
rect 178451 529538 178481 529668
rect 178659 529538 178689 529622
rect 178750 529538 178780 529622
rect 178899 529538 178929 529622
rect 178995 529538 179025 529610
rect 179104 529538 179134 529610
rect 179203 529538 179233 529666
rect 179335 529538 179365 529622
rect 179407 529538 179437 529622
rect 179573 529538 179603 529610
rect 179669 529538 179699 529610
rect 179764 529538 179794 529622
rect 180019 529538 180049 529622
rect 180103 529538 180133 529622
rect 180291 529538 180321 529622
rect 180375 529538 180405 529622
rect 180630 529538 180660 529622
rect 180725 529538 180755 529610
rect 180821 529538 180851 529610
rect 180987 529538 181017 529622
rect 181059 529538 181089 529622
rect 181191 529538 181221 529666
rect 181290 529538 181320 529610
rect 181399 529538 181429 529610
rect 181495 529538 181525 529622
rect 181644 529538 181674 529622
rect 181735 529538 181765 529622
rect 181943 529538 181973 529668
rect 182131 529538 182341 529648
rect 182702 529538 182732 529668
rect 182797 529538 182897 529622
rect 183055 529538 183155 529622
rect 183209 529538 183239 529622
rect 183419 529538 184365 529648
rect 184523 529538 185469 529648
rect 185627 529538 186573 529648
rect 186731 529538 187125 529648
rect 187283 529538 187401 529648
rect 172287 529334 172405 529444
rect 172563 529334 173509 529444
rect 173667 529334 174613 529444
rect 175185 529360 175215 529444
rect 175353 529360 175383 529444
rect 175449 529360 175479 529444
rect 175574 529360 175604 529444
rect 175670 529360 175700 529444
rect 175779 529314 175809 529444
rect 175985 529360 176015 529444
rect 176071 529360 176101 529444
rect 176157 529360 176187 529444
rect 176243 529360 176273 529444
rect 176329 529360 176359 529444
rect 176415 529360 176445 529444
rect 176501 529360 176531 529444
rect 176587 529360 176617 529444
rect 176672 529360 176702 529444
rect 176758 529360 176788 529444
rect 176844 529360 176874 529444
rect 176930 529360 176960 529444
rect 177016 529360 177046 529444
rect 177102 529360 177132 529444
rect 177188 529360 177218 529444
rect 177274 529360 177304 529444
rect 177360 529360 177390 529444
rect 177446 529360 177476 529444
rect 177532 529360 177562 529444
rect 177618 529360 177648 529444
rect 177807 529360 177837 529444
rect 177891 529360 177921 529444
rect 178146 529360 178176 529444
rect 178241 529372 178271 529444
rect 178337 529372 178367 529444
rect 178503 529360 178533 529444
rect 178575 529360 178605 529444
rect 178707 529316 178737 529444
rect 178806 529372 178836 529444
rect 178915 529372 178945 529444
rect 179011 529360 179041 529444
rect 179160 529360 179190 529444
rect 179251 529360 179281 529444
rect 179459 529314 179489 529444
rect 179739 529340 179769 529444
rect 179827 529340 179857 529444
rect 180107 529334 180501 529444
rect 180752 529360 180782 529444
rect 180838 529360 180868 529444
rect 180924 529360 180954 529444
rect 181010 529360 181040 529444
rect 181096 529360 181126 529444
rect 181182 529360 181212 529444
rect 181268 529360 181298 529444
rect 181354 529360 181384 529444
rect 181440 529360 181470 529444
rect 181526 529360 181556 529444
rect 181612 529360 181642 529444
rect 181698 529360 181728 529444
rect 181783 529360 181813 529444
rect 181869 529360 181899 529444
rect 181955 529360 181985 529444
rect 182041 529360 182071 529444
rect 182127 529360 182157 529444
rect 182213 529360 182243 529444
rect 182299 529360 182329 529444
rect 182385 529360 182415 529444
rect 182591 529340 182621 529444
rect 182679 529340 182709 529444
rect 182867 529334 183813 529444
rect 183971 529334 184917 529444
rect 185259 529334 186205 529444
rect 186363 529334 186941 529444
rect 187283 529334 187401 529444
rect 172287 528450 172405 528560
rect 172563 528450 173509 528560
rect 173667 528450 174613 528560
rect 174771 528450 175717 528560
rect 175967 528450 175997 528554
rect 176055 528450 176085 528554
rect 176243 528450 176273 528554
rect 176331 528450 176361 528554
rect 176565 528450 176595 528534
rect 176733 528450 176763 528534
rect 176829 528450 176859 528534
rect 176954 528450 176984 528534
rect 177050 528450 177080 528534
rect 177159 528450 177189 528580
rect 177550 528450 177580 528580
rect 177645 528450 177745 528534
rect 177903 528450 178003 528534
rect 178057 528450 178087 528534
rect 178452 528450 178482 528534
rect 178538 528450 178568 528534
rect 178624 528450 178654 528534
rect 178710 528450 178740 528534
rect 178796 528450 178826 528534
rect 178882 528450 178912 528534
rect 178968 528450 178998 528534
rect 179054 528450 179084 528534
rect 179140 528450 179170 528534
rect 179226 528450 179256 528534
rect 179312 528450 179342 528534
rect 179398 528450 179428 528534
rect 179483 528450 179513 528534
rect 179569 528450 179599 528534
rect 179655 528450 179685 528534
rect 179741 528450 179771 528534
rect 179827 528450 179857 528534
rect 179913 528450 179943 528534
rect 179999 528450 180029 528534
rect 180085 528450 180115 528534
rect 180291 528450 180321 528554
rect 180379 528450 180409 528554
rect 180567 528450 180597 528534
rect 180651 528450 180681 528534
rect 180906 528450 180936 528534
rect 181001 528450 181031 528522
rect 181097 528450 181127 528522
rect 181263 528450 181293 528534
rect 181335 528450 181365 528534
rect 181467 528450 181497 528578
rect 181566 528450 181596 528522
rect 181675 528450 181705 528522
rect 181771 528450 181801 528534
rect 181920 528450 181950 528534
rect 182011 528450 182041 528534
rect 182219 528450 182249 528580
rect 182683 528450 183629 528560
rect 183787 528450 184733 528560
rect 184891 528450 185837 528560
rect 185995 528450 186941 528560
rect 187283 528450 187401 528560
rect 172287 528246 172405 528356
rect 172563 528246 173509 528356
rect 173667 528246 174613 528356
rect 174955 528246 175901 528356
rect 176151 528272 176181 528356
rect 176235 528272 176265 528356
rect 176490 528272 176520 528356
rect 176585 528284 176615 528356
rect 176681 528284 176711 528356
rect 176847 528272 176877 528356
rect 176919 528272 176949 528356
rect 177051 528228 177081 528356
rect 177150 528284 177180 528356
rect 177259 528284 177289 528356
rect 177355 528272 177385 528356
rect 177504 528272 177534 528356
rect 177595 528272 177625 528356
rect 177803 528226 177833 528356
rect 177991 528252 178021 528356
rect 178079 528252 178109 528356
rect 178267 528246 178845 528356
rect 179003 528226 179033 528356
rect 179112 528272 179142 528356
rect 179208 528272 179238 528356
rect 179333 528272 179363 528356
rect 179429 528272 179459 528356
rect 179597 528272 179627 528356
rect 180107 528246 180685 528356
rect 181027 528226 181057 528356
rect 181136 528272 181166 528356
rect 181232 528272 181262 528356
rect 181357 528272 181387 528356
rect 181453 528272 181483 528356
rect 181621 528272 181651 528356
rect 181855 528246 182801 528356
rect 182959 528246 183905 528356
rect 184063 528246 185009 528356
rect 185259 528246 186205 528356
rect 186363 528246 186941 528356
rect 187283 528246 187401 528356
rect 172287 527362 172405 527472
rect 172563 527362 173509 527472
rect 173667 527362 174613 527472
rect 174771 527362 175717 527472
rect 175875 527362 176269 527472
rect 176446 527362 176476 527492
rect 176541 527362 176641 527446
rect 176799 527362 176899 527446
rect 176953 527362 176983 527446
rect 177163 527362 177281 527472
rect 177531 527362 178477 527472
rect 178635 527362 178845 527472
rect 179022 527362 179052 527492
rect 179117 527362 179217 527446
rect 179375 527362 179475 527446
rect 179529 527362 179559 527446
rect 179739 527362 180685 527472
rect 180843 527362 181789 527472
rect 181947 527362 182341 527472
rect 182683 527362 183629 527472
rect 183787 527362 184733 527472
rect 184891 527362 185837 527472
rect 185995 527362 186941 527472
rect 187283 527362 187401 527472
rect 172287 527158 172405 527268
rect 172563 527158 173509 527268
rect 173667 527158 174613 527268
rect 174955 527158 175901 527268
rect 176059 527158 177005 527268
rect 177163 527158 178109 527268
rect 178267 527158 179213 527268
rect 179371 527158 179765 527268
rect 180107 527158 181053 527268
rect 181211 527158 182157 527268
rect 182315 527158 183261 527268
rect 183419 527158 184365 527268
rect 184523 527158 184917 527268
rect 185259 527158 186205 527268
rect 186363 527158 186941 527268
rect 187283 527158 187401 527268
rect 172287 526274 172405 526384
rect 172563 526274 173509 526384
rect 173667 526274 174613 526384
rect 174771 526274 175717 526384
rect 175875 526274 176821 526384
rect 176979 526274 177189 526384
rect 177531 526274 178477 526384
rect 178635 526274 179581 526384
rect 179739 526274 180685 526384
rect 180843 526274 181789 526384
rect 181947 526274 182341 526384
rect 182683 526274 183629 526384
rect 183787 526274 184733 526384
rect 184891 526274 185837 526384
rect 185995 526274 186941 526384
rect 187283 526274 187401 526384
rect 172287 526070 172405 526180
rect 172563 526070 173509 526180
rect 173667 526070 174613 526180
rect 174955 526070 175901 526180
rect 176059 526070 177005 526180
rect 177163 526070 178109 526180
rect 178267 526070 179213 526180
rect 179371 526070 179765 526180
rect 180107 526070 181053 526180
rect 181211 526070 182157 526180
rect 182315 526070 183261 526180
rect 183419 526070 184365 526180
rect 184523 526070 184917 526180
rect 185259 526070 186205 526180
rect 186363 526070 186941 526180
rect 187283 526070 187401 526180
rect 172287 525186 172405 525296
rect 172563 525186 173509 525296
rect 173667 525186 174613 525296
rect 174771 525186 175717 525296
rect 175875 525186 176821 525296
rect 176979 525186 177189 525296
rect 177531 525186 178477 525296
rect 178635 525186 179581 525296
rect 179739 525186 180685 525296
rect 180843 525186 181789 525296
rect 181947 525186 182341 525296
rect 182683 525186 183629 525296
rect 183787 525186 184733 525296
rect 184891 525186 185837 525296
rect 185995 525186 186941 525296
rect 187283 525186 187401 525296
rect 172287 524982 172405 525092
rect 172563 524982 173509 525092
rect 173667 524982 174613 525092
rect 174955 524982 175901 525092
rect 176059 524982 177005 525092
rect 177163 524982 178109 525092
rect 178267 524982 179213 525092
rect 179371 524982 179765 525092
rect 180107 524982 181053 525092
rect 181211 524982 182157 525092
rect 182315 524982 183261 525092
rect 183419 524982 184365 525092
rect 184523 524982 184917 525092
rect 185259 524982 186205 525092
rect 186363 524982 186941 525092
rect 187283 524982 187401 525092
rect 172287 524098 172405 524208
rect 172563 524098 173509 524208
rect 173667 524098 174613 524208
rect 174771 524098 175717 524208
rect 175875 524098 176821 524208
rect 176979 524098 177189 524208
rect 177531 524098 178477 524208
rect 178635 524098 179581 524208
rect 179739 524098 180685 524208
rect 180843 524098 181789 524208
rect 181947 524098 182341 524208
rect 182683 524098 183629 524208
rect 183787 524098 184733 524208
rect 184891 524098 185837 524208
rect 185995 524098 186941 524208
rect 187283 524098 187401 524208
rect 172287 523894 172405 524004
rect 172563 523894 173509 524004
rect 173667 523894 174613 524004
rect 174955 523894 175901 524004
rect 176059 523894 177005 524004
rect 177163 523894 178109 524004
rect 178267 523894 179213 524004
rect 179371 523894 179765 524004
rect 180107 523894 181053 524004
rect 181211 523894 182157 524004
rect 182315 523894 183261 524004
rect 183419 523894 184365 524004
rect 184523 523894 184917 524004
rect 185259 523894 186205 524004
rect 186363 523894 186941 524004
rect 187283 523894 187401 524004
rect 172287 523010 172405 523120
rect 172563 523010 173509 523120
rect 173667 523010 174613 523120
rect 174771 523010 175717 523120
rect 175875 523010 176821 523120
rect 176979 523010 177189 523120
rect 177531 523010 178477 523120
rect 178635 523010 179581 523120
rect 179739 523010 180685 523120
rect 180843 523010 181789 523120
rect 181947 523010 182341 523120
rect 182683 523010 183629 523120
rect 183787 523010 184733 523120
rect 184891 523010 185837 523120
rect 185995 523010 186941 523120
rect 187283 523010 187401 523120
rect 172287 522806 172405 522916
rect 172563 522806 173509 522916
rect 173667 522806 174613 522916
rect 174955 522806 175901 522916
rect 176059 522806 177005 522916
rect 177163 522806 178109 522916
rect 178267 522806 179213 522916
rect 179371 522806 179765 522916
rect 180107 522806 181053 522916
rect 181211 522806 182157 522916
rect 182315 522806 183261 522916
rect 183419 522806 184365 522916
rect 184523 522806 184917 522916
rect 185259 522806 186205 522916
rect 186363 522806 186941 522916
rect 187283 522806 187401 522916
rect 172287 521922 172405 522032
rect 172563 521922 173509 522032
rect 173667 521922 174613 522032
rect 174771 521922 175717 522032
rect 175875 521922 176821 522032
rect 176979 521922 177189 522032
rect 177531 521922 178477 522032
rect 178635 521922 179581 522032
rect 179739 521922 180685 522032
rect 180843 521922 181789 522032
rect 181947 521922 182341 522032
rect 182683 521922 183629 522032
rect 183787 521922 184733 522032
rect 184891 521922 185837 522032
rect 185995 521922 186941 522032
rect 187283 521922 187401 522032
rect 172287 521718 172405 521828
rect 172563 521718 173509 521828
rect 173667 521718 174613 521828
rect 174955 521718 175901 521828
rect 176059 521718 177005 521828
rect 177163 521718 178109 521828
rect 178267 521718 179213 521828
rect 179371 521718 179765 521828
rect 180107 521718 181053 521828
rect 181211 521718 182157 521828
rect 182315 521718 183261 521828
rect 183419 521718 184365 521828
rect 184523 521718 184917 521828
rect 185259 521718 186205 521828
rect 186363 521718 186941 521828
rect 187283 521718 187401 521828
rect 172287 520834 172405 520944
rect 172563 520834 173509 520944
rect 173667 520834 174613 520944
rect 174771 520834 175717 520944
rect 175875 520834 176821 520944
rect 176979 520834 177189 520944
rect 177531 520834 178477 520944
rect 178635 520834 179581 520944
rect 179739 520834 180685 520944
rect 180843 520834 181789 520944
rect 181947 520834 182341 520944
rect 182683 520834 183629 520944
rect 183787 520834 184733 520944
rect 184891 520834 185837 520944
rect 185995 520834 186941 520944
rect 187283 520834 187401 520944
rect 172287 520630 172405 520740
rect 172563 520630 173509 520740
rect 173667 520630 174613 520740
rect 174955 520630 175901 520740
rect 176059 520630 177005 520740
rect 177163 520630 178109 520740
rect 178267 520630 179213 520740
rect 179371 520630 179765 520740
rect 180107 520630 181053 520740
rect 181211 520630 182157 520740
rect 182315 520630 183261 520740
rect 183419 520630 184365 520740
rect 184523 520630 184917 520740
rect 185259 520630 186205 520740
rect 186363 520630 186941 520740
rect 187283 520630 187401 520740
rect 172287 519746 172405 519856
rect 172563 519746 173509 519856
rect 173667 519746 174613 519856
rect 174771 519746 175717 519856
rect 175875 519746 176821 519856
rect 176979 519746 177189 519856
rect 177531 519746 178477 519856
rect 178635 519746 179581 519856
rect 179739 519746 180685 519856
rect 180843 519746 181789 519856
rect 181947 519746 182341 519856
rect 182683 519746 183629 519856
rect 183787 519746 184733 519856
rect 184891 519746 185837 519856
rect 185995 519746 186941 519856
rect 187283 519746 187401 519856
rect 172287 519542 172405 519652
rect 172563 519542 173509 519652
rect 173667 519542 174613 519652
rect 174955 519542 175901 519652
rect 176059 519542 177005 519652
rect 177163 519542 178109 519652
rect 178267 519542 179213 519652
rect 179371 519542 179765 519652
rect 180107 519542 181053 519652
rect 181211 519542 182157 519652
rect 182315 519542 183261 519652
rect 183419 519542 184365 519652
rect 184523 519542 184917 519652
rect 185259 519542 186205 519652
rect 186363 519542 186941 519652
rect 187283 519542 187401 519652
rect 172287 518658 172405 518768
rect 172563 518658 173509 518768
rect 173667 518658 174613 518768
rect 174771 518658 175717 518768
rect 175875 518658 176821 518768
rect 176979 518658 177189 518768
rect 177531 518658 178477 518768
rect 178635 518658 179581 518768
rect 179739 518658 180685 518768
rect 180843 518658 181789 518768
rect 181947 518658 182341 518768
rect 182683 518658 183629 518768
rect 183787 518658 184733 518768
rect 184891 518658 185837 518768
rect 185995 518658 186941 518768
rect 187283 518658 187401 518768
rect 172287 518454 172405 518564
rect 172563 518454 173509 518564
rect 173667 518454 174613 518564
rect 174955 518454 175901 518564
rect 176059 518454 177005 518564
rect 177163 518454 178109 518564
rect 178267 518454 179213 518564
rect 179371 518454 179765 518564
rect 180107 518454 181053 518564
rect 181211 518454 182157 518564
rect 182315 518454 183261 518564
rect 183419 518454 184365 518564
rect 184523 518454 184917 518564
rect 185259 518454 186205 518564
rect 186363 518454 186941 518564
rect 187283 518454 187401 518564
rect 172287 517570 172405 517680
rect 172563 517570 173509 517680
rect 173667 517570 174613 517680
rect 174771 517570 175717 517680
rect 175875 517570 176821 517680
rect 176979 517570 177189 517680
rect 177531 517570 178477 517680
rect 178635 517570 179581 517680
rect 179739 517570 180685 517680
rect 180843 517570 181789 517680
rect 181947 517570 182341 517680
rect 182683 517570 183629 517680
rect 183787 517570 184733 517680
rect 184891 517570 185837 517680
rect 185995 517570 186941 517680
rect 187283 517570 187401 517680
rect 172287 517366 172405 517476
rect 172563 517366 173509 517476
rect 173667 517366 174613 517476
rect 174955 517366 175901 517476
rect 176059 517366 177005 517476
rect 177163 517366 178109 517476
rect 178267 517366 179213 517476
rect 179371 517366 179765 517476
rect 180107 517366 181053 517476
rect 181211 517366 182157 517476
rect 182315 517366 183261 517476
rect 183419 517366 184365 517476
rect 184523 517366 184917 517476
rect 185259 517366 186205 517476
rect 186363 517366 186941 517476
rect 187283 517366 187401 517476
rect 172287 516482 172405 516592
rect 172563 516482 173509 516592
rect 173667 516482 174613 516592
rect 174771 516482 175717 516592
rect 175875 516482 176821 516592
rect 176979 516482 177189 516592
rect 177531 516482 178477 516592
rect 178635 516482 179581 516592
rect 179739 516482 180685 516592
rect 180843 516482 181789 516592
rect 181947 516482 182341 516592
rect 182683 516482 183629 516592
rect 183787 516482 184733 516592
rect 184891 516482 185837 516592
rect 185995 516482 186941 516592
rect 187283 516482 187401 516592
rect 172287 516278 172405 516388
rect 172563 516278 173509 516388
rect 173667 516278 174613 516388
rect 174955 516278 175901 516388
rect 176059 516278 177005 516388
rect 177163 516278 178109 516388
rect 178267 516278 179213 516388
rect 179371 516278 179765 516388
rect 180107 516278 181053 516388
rect 181211 516278 182157 516388
rect 182315 516278 183261 516388
rect 183419 516278 184365 516388
rect 184523 516278 184917 516388
rect 185259 516278 186205 516388
rect 186363 516278 186941 516388
rect 187283 516278 187401 516388
rect 172287 515394 172405 515504
rect 172563 515394 173141 515504
rect 173484 515394 173514 515478
rect 173581 515394 173611 515478
rect 173667 515394 173697 515478
rect 173753 515394 173783 515478
rect 173839 515394 173869 515478
rect 174035 515394 174613 515504
rect 174955 515394 175901 515504
rect 176059 515394 177005 515504
rect 177163 515394 177281 515504
rect 177531 515394 178477 515504
rect 178635 515394 179581 515504
rect 179739 515394 179857 515504
rect 180107 515394 181053 515504
rect 181211 515394 181789 515504
rect 182131 515394 182161 515498
rect 182219 515394 182249 515498
rect 182683 515394 183629 515504
rect 183787 515394 184733 515504
rect 184891 515394 185009 515504
rect 185259 515394 186205 515504
rect 186456 515394 186486 515478
rect 186553 515394 186583 515478
rect 186639 515394 186669 515478
rect 186725 515394 186755 515478
rect 186811 515394 186841 515478
rect 187007 515394 187125 515504
rect 187283 515394 187401 515504
<< pmos >>
rect 164714 538525 164744 539525
rect 164941 538532 164971 539532
rect 165037 538532 165067 539532
rect 165133 538532 165163 539532
rect 165229 538532 165259 539532
rect 165325 538532 165355 539532
rect 165421 538532 165451 539532
rect 165517 538532 165547 539532
rect 165613 538532 165643 539532
rect 165709 538532 165739 539532
rect 165805 538532 165835 539532
rect 165901 538532 165931 539532
rect 165997 538532 166027 539532
rect 166214 538925 166244 539525
rect 166414 538525 166444 539525
rect 168514 538525 168544 539525
rect 168741 538532 168771 539532
rect 168837 538532 168867 539532
rect 168933 538532 168963 539532
rect 169029 538532 169059 539532
rect 169125 538532 169155 539532
rect 169221 538532 169251 539532
rect 169317 538532 169347 539532
rect 169413 538532 169443 539532
rect 169509 538532 169539 539532
rect 169605 538532 169635 539532
rect 169701 538532 169731 539532
rect 169797 538532 169827 539532
rect 170014 538925 170044 539525
rect 170214 538525 170244 539525
rect 172214 538525 172244 539525
rect 172441 538532 172471 539532
rect 172537 538532 172567 539532
rect 172633 538532 172663 539532
rect 172729 538532 172759 539532
rect 172825 538532 172855 539532
rect 172921 538532 172951 539532
rect 173017 538532 173047 539532
rect 173113 538532 173143 539532
rect 173209 538532 173239 539532
rect 173305 538532 173335 539532
rect 173401 538532 173431 539532
rect 173497 538532 173527 539532
rect 173714 538925 173744 539525
rect 173914 538525 173944 539525
rect 175714 538525 175744 539525
rect 175941 538532 175971 539532
rect 176037 538532 176067 539532
rect 176133 538532 176163 539532
rect 176229 538532 176259 539532
rect 176325 538532 176355 539532
rect 176421 538532 176451 539532
rect 176517 538532 176547 539532
rect 176613 538532 176643 539532
rect 176709 538532 176739 539532
rect 176805 538532 176835 539532
rect 176901 538532 176931 539532
rect 176997 538532 177027 539532
rect 177214 538925 177244 539525
rect 177414 538525 177444 539525
rect 179314 538525 179344 539525
rect 179541 538532 179571 539532
rect 179637 538532 179667 539532
rect 179733 538532 179763 539532
rect 179829 538532 179859 539532
rect 179925 538532 179955 539532
rect 180021 538532 180051 539532
rect 180117 538532 180147 539532
rect 180213 538532 180243 539532
rect 180309 538532 180339 539532
rect 180405 538532 180435 539532
rect 180501 538532 180531 539532
rect 180597 538532 180627 539532
rect 180814 538925 180844 539525
rect 181014 538525 181044 539525
rect 182614 538525 182644 539525
rect 182841 538532 182871 539532
rect 182937 538532 182967 539532
rect 183033 538532 183063 539532
rect 183129 538532 183159 539532
rect 183225 538532 183255 539532
rect 183321 538532 183351 539532
rect 183417 538532 183447 539532
rect 183513 538532 183543 539532
rect 183609 538532 183639 539532
rect 183705 538532 183735 539532
rect 183801 538532 183831 539532
rect 183897 538532 183927 539532
rect 184114 538925 184144 539525
rect 184314 538525 184344 539525
rect 185914 538525 185944 539525
rect 186141 538532 186171 539532
rect 186237 538532 186267 539532
rect 186333 538532 186363 539532
rect 186429 538532 186459 539532
rect 186525 538532 186555 539532
rect 186621 538532 186651 539532
rect 186717 538532 186747 539532
rect 186813 538532 186843 539532
rect 186909 538532 186939 539532
rect 187005 538532 187035 539532
rect 187101 538532 187131 539532
rect 187197 538532 187227 539532
rect 187414 538925 187444 539525
rect 187614 538525 187644 539525
rect 189214 538525 189244 539525
rect 189441 538532 189471 539532
rect 189537 538532 189567 539532
rect 189633 538532 189663 539532
rect 189729 538532 189759 539532
rect 189825 538532 189855 539532
rect 189921 538532 189951 539532
rect 190017 538532 190047 539532
rect 190113 538532 190143 539532
rect 190209 538532 190239 539532
rect 190305 538532 190335 539532
rect 190401 538532 190431 539532
rect 190497 538532 190527 539532
rect 190714 538925 190744 539525
rect 190914 538525 190944 539525
rect 161304 537025 161334 537625
rect 161508 537025 161538 537625
rect 161604 537025 161634 537625
rect 161700 537025 161730 537625
rect 161908 537025 161938 537625
rect 162004 537025 162034 537625
rect 162100 537025 162130 537625
rect 162324 537025 162354 537625
rect 157794 536005 157994 536605
rect 158172 536005 158372 536605
rect 158430 536005 158630 536605
rect 158688 536005 158888 536605
rect 158946 536005 159146 536605
rect 159204 536005 159404 536605
rect 159462 536005 159662 536605
rect 159720 536005 159920 536605
rect 159978 536005 160178 536605
rect 160236 536005 160436 536605
rect 160494 536005 160694 536605
rect 160878 536005 161078 536605
rect 161136 536005 161336 536605
rect 161394 536005 161594 536605
rect 161776 536005 161976 536605
rect 162034 536005 162234 536605
rect 162414 536005 162614 536605
<< scpmoshvt >>
rect 172287 530082 172405 530256
rect 172572 530082 172602 530282
rect 172658 530082 172688 530282
rect 172744 530082 172774 530282
rect 172830 530082 172860 530282
rect 172926 530082 172956 530282
rect 173115 530082 174061 530256
rect 174219 530082 174613 530256
rect 174964 530082 174994 530282
rect 175050 530082 175080 530282
rect 175136 530082 175166 530282
rect 175222 530082 175252 530282
rect 175318 530082 175348 530282
rect 175599 530082 175629 530282
rect 175814 530082 175844 530166
rect 175898 530082 175928 530166
rect 176006 530082 176036 530166
rect 176090 530082 176120 530166
rect 176176 530082 176206 530166
rect 176275 530082 176305 530250
rect 176472 530082 176502 530166
rect 176569 530082 176599 530166
rect 176709 530082 176739 530166
rect 176808 530082 176838 530166
rect 176900 530082 176930 530166
rect 177167 530088 177197 530216
rect 177251 530088 177281 530216
rect 177734 530082 177764 530282
rect 177829 530082 177929 530166
rect 178087 530082 178187 530166
rect 178241 530082 178271 530166
rect 178451 530082 178481 530240
rect 178539 530082 178569 530240
rect 178736 530082 178766 530282
rect 178822 530082 178852 530282
rect 178908 530082 178938 530282
rect 178994 530082 179024 530282
rect 179090 530082 179120 530282
rect 179280 530082 179310 530282
rect 179376 530082 179406 530282
rect 179462 530082 179492 530282
rect 179548 530082 179578 530282
rect 179634 530082 179664 530282
rect 180291 530082 180321 530282
rect 180400 530121 180430 530205
rect 180503 530121 180533 530205
rect 180717 530121 180747 530205
rect 180789 530121 180819 530205
rect 180885 530121 180915 530205
rect 181257 530121 181287 530205
rect 181353 530121 181383 530205
rect 181425 530121 181455 530205
rect 181639 530121 181669 530205
rect 181742 530121 181772 530205
rect 181851 530082 181881 530282
rect 182040 530082 182070 530282
rect 182136 530082 182166 530282
rect 182222 530082 182252 530282
rect 182308 530082 182338 530282
rect 182394 530082 182424 530282
rect 182683 530082 182893 530256
rect 183144 530082 183174 530282
rect 183240 530082 183270 530282
rect 183326 530082 183356 530282
rect 183412 530082 183442 530282
rect 183498 530082 183528 530282
rect 183695 530082 184641 530256
rect 184799 530082 185009 530256
rect 185260 530082 185290 530282
rect 185356 530082 185386 530282
rect 185442 530082 185472 530282
rect 185528 530082 185558 530282
rect 185614 530082 185644 530282
rect 185811 530082 186757 530256
rect 187283 530082 187401 530256
rect 172287 529814 172405 529988
rect 172563 529814 173509 529988
rect 173667 529814 174613 529988
rect 174885 529904 174915 529988
rect 174969 529904 175069 529988
rect 175227 529904 175327 529988
rect 175392 529788 175422 529988
rect 175599 529854 175629 529982
rect 175683 529854 175713 529982
rect 175950 529904 175980 529988
rect 176042 529904 176072 529988
rect 176141 529904 176171 529988
rect 176281 529904 176311 529988
rect 176378 529904 176408 529988
rect 176575 529820 176605 529988
rect 176674 529904 176704 529988
rect 176760 529904 176790 529988
rect 176844 529904 176874 529988
rect 176952 529904 176982 529988
rect 177036 529904 177066 529988
rect 177251 529788 177281 529988
rect 177669 529865 177699 529949
rect 177765 529865 177795 529949
rect 177837 529865 177867 529949
rect 178051 529865 178081 529949
rect 178154 529865 178184 529949
rect 178263 529788 178293 529988
rect 178451 529788 178481 529988
rect 178666 529904 178696 529988
rect 178750 529904 178780 529988
rect 178858 529904 178888 529988
rect 178942 529904 178972 529988
rect 179028 529904 179058 529988
rect 179127 529820 179157 529988
rect 179324 529904 179354 529988
rect 179421 529904 179451 529988
rect 179561 529904 179591 529988
rect 179660 529904 179690 529988
rect 179752 529904 179782 529988
rect 180019 529854 180049 529982
rect 180103 529854 180133 529982
rect 180291 529854 180321 529982
rect 180375 529854 180405 529982
rect 180642 529904 180672 529988
rect 180734 529904 180764 529988
rect 180833 529904 180863 529988
rect 180973 529904 181003 529988
rect 181070 529904 181100 529988
rect 181267 529820 181297 529988
rect 181366 529904 181396 529988
rect 181452 529904 181482 529988
rect 181536 529904 181566 529988
rect 181644 529904 181674 529988
rect 181728 529904 181758 529988
rect 181943 529788 181973 529988
rect 182131 529814 182341 529988
rect 182702 529788 182732 529988
rect 182797 529904 182897 529988
rect 183055 529904 183155 529988
rect 183209 529904 183239 529988
rect 183419 529814 184365 529988
rect 184523 529814 185469 529988
rect 185627 529814 186573 529988
rect 186731 529814 187125 529988
rect 187283 529814 187401 529988
rect 172287 528994 172405 529168
rect 172563 528994 173509 529168
rect 173667 528994 174613 529168
rect 175185 529033 175215 529117
rect 175281 529033 175311 529117
rect 175353 529033 175383 529117
rect 175567 529033 175597 529117
rect 175670 529033 175700 529117
rect 175779 528994 175809 529194
rect 175985 528994 176015 529194
rect 176071 528994 176101 529194
rect 176157 528994 176187 529194
rect 176243 528994 176273 529194
rect 176329 528994 176359 529194
rect 176415 528994 176445 529194
rect 176501 528994 176531 529194
rect 176587 528994 176617 529194
rect 176672 528994 176702 529194
rect 176758 528994 176788 529194
rect 176844 528994 176874 529194
rect 176930 528994 176960 529194
rect 177016 528994 177046 529194
rect 177102 528994 177132 529194
rect 177188 528994 177218 529194
rect 177274 528994 177304 529194
rect 177360 528994 177390 529194
rect 177446 528994 177476 529194
rect 177532 528994 177562 529194
rect 177618 528994 177648 529194
rect 177807 529000 177837 529128
rect 177891 529000 177921 529128
rect 178158 528994 178188 529078
rect 178250 528994 178280 529078
rect 178349 528994 178379 529078
rect 178489 528994 178519 529078
rect 178586 528994 178616 529078
rect 178783 528994 178813 529162
rect 178882 528994 178912 529078
rect 178968 528994 178998 529078
rect 179052 528994 179082 529078
rect 179160 528994 179190 529078
rect 179244 528994 179274 529078
rect 179459 528994 179489 529194
rect 179739 528994 179769 529152
rect 179827 528994 179857 529152
rect 180107 528994 180501 529168
rect 180752 528994 180782 529194
rect 180838 528994 180868 529194
rect 180924 528994 180954 529194
rect 181010 528994 181040 529194
rect 181096 528994 181126 529194
rect 181182 528994 181212 529194
rect 181268 528994 181298 529194
rect 181354 528994 181384 529194
rect 181440 528994 181470 529194
rect 181526 528994 181556 529194
rect 181612 528994 181642 529194
rect 181698 528994 181728 529194
rect 181783 528994 181813 529194
rect 181869 528994 181899 529194
rect 181955 528994 181985 529194
rect 182041 528994 182071 529194
rect 182127 528994 182157 529194
rect 182213 528994 182243 529194
rect 182299 528994 182329 529194
rect 182385 528994 182415 529194
rect 182591 528994 182621 529152
rect 182679 528994 182709 529152
rect 182867 528994 183813 529168
rect 183971 528994 184917 529168
rect 185259 528994 186205 529168
rect 186363 528994 186941 529168
rect 187283 528994 187401 529168
rect 172287 528726 172405 528900
rect 172563 528726 173509 528900
rect 173667 528726 174613 528900
rect 174771 528726 175717 528900
rect 175967 528742 175997 528900
rect 176055 528742 176085 528900
rect 176243 528742 176273 528900
rect 176331 528742 176361 528900
rect 176565 528777 176595 528861
rect 176661 528777 176691 528861
rect 176733 528777 176763 528861
rect 176947 528777 176977 528861
rect 177050 528777 177080 528861
rect 177159 528700 177189 528900
rect 177550 528700 177580 528900
rect 177645 528816 177745 528900
rect 177903 528816 178003 528900
rect 178057 528816 178087 528900
rect 178452 528700 178482 528900
rect 178538 528700 178568 528900
rect 178624 528700 178654 528900
rect 178710 528700 178740 528900
rect 178796 528700 178826 528900
rect 178882 528700 178912 528900
rect 178968 528700 178998 528900
rect 179054 528700 179084 528900
rect 179140 528700 179170 528900
rect 179226 528700 179256 528900
rect 179312 528700 179342 528900
rect 179398 528700 179428 528900
rect 179483 528700 179513 528900
rect 179569 528700 179599 528900
rect 179655 528700 179685 528900
rect 179741 528700 179771 528900
rect 179827 528700 179857 528900
rect 179913 528700 179943 528900
rect 179999 528700 180029 528900
rect 180085 528700 180115 528900
rect 180291 528742 180321 528900
rect 180379 528742 180409 528900
rect 180567 528766 180597 528894
rect 180651 528766 180681 528894
rect 180918 528816 180948 528900
rect 181010 528816 181040 528900
rect 181109 528816 181139 528900
rect 181249 528816 181279 528900
rect 181346 528816 181376 528900
rect 181543 528732 181573 528900
rect 181642 528816 181672 528900
rect 181728 528816 181758 528900
rect 181812 528816 181842 528900
rect 181920 528816 181950 528900
rect 182004 528816 182034 528900
rect 182219 528700 182249 528900
rect 182683 528726 183629 528900
rect 183787 528726 184733 528900
rect 184891 528726 185837 528900
rect 185995 528726 186941 528900
rect 187283 528726 187401 528900
rect 172287 527906 172405 528080
rect 172563 527906 173509 528080
rect 173667 527906 174613 528080
rect 174955 527906 175901 528080
rect 176151 527912 176181 528040
rect 176235 527912 176265 528040
rect 176502 527906 176532 527990
rect 176594 527906 176624 527990
rect 176693 527906 176723 527990
rect 176833 527906 176863 527990
rect 176930 527906 176960 527990
rect 177127 527906 177157 528074
rect 177226 527906 177256 527990
rect 177312 527906 177342 527990
rect 177396 527906 177426 527990
rect 177504 527906 177534 527990
rect 177588 527906 177618 527990
rect 177803 527906 177833 528106
rect 177991 527906 178021 528064
rect 178079 527906 178109 528064
rect 178267 527906 178845 528080
rect 179003 527906 179033 528106
rect 179112 527945 179142 528029
rect 179215 527945 179245 528029
rect 179429 527945 179459 528029
rect 179501 527945 179531 528029
rect 179597 527945 179627 528029
rect 180107 527906 180685 528080
rect 181027 527906 181057 528106
rect 181136 527945 181166 528029
rect 181239 527945 181269 528029
rect 181453 527945 181483 528029
rect 181525 527945 181555 528029
rect 181621 527945 181651 528029
rect 181855 527906 182801 528080
rect 182959 527906 183905 528080
rect 184063 527906 185009 528080
rect 185259 527906 186205 528080
rect 186363 527906 186941 528080
rect 187283 527906 187401 528080
rect 172287 527638 172405 527812
rect 172563 527638 173509 527812
rect 173667 527638 174613 527812
rect 174771 527638 175717 527812
rect 175875 527638 176269 527812
rect 176446 527612 176476 527812
rect 176541 527728 176641 527812
rect 176799 527728 176899 527812
rect 176953 527728 176983 527812
rect 177163 527638 177281 527812
rect 177531 527638 178477 527812
rect 178635 527638 178845 527812
rect 179022 527612 179052 527812
rect 179117 527728 179217 527812
rect 179375 527728 179475 527812
rect 179529 527728 179559 527812
rect 179739 527638 180685 527812
rect 180843 527638 181789 527812
rect 181947 527638 182341 527812
rect 182683 527638 183629 527812
rect 183787 527638 184733 527812
rect 184891 527638 185837 527812
rect 185995 527638 186941 527812
rect 187283 527638 187401 527812
rect 172287 526818 172405 526992
rect 172563 526818 173509 526992
rect 173667 526818 174613 526992
rect 174955 526818 175901 526992
rect 176059 526818 177005 526992
rect 177163 526818 178109 526992
rect 178267 526818 179213 526992
rect 179371 526818 179765 526992
rect 180107 526818 181053 526992
rect 181211 526818 182157 526992
rect 182315 526818 183261 526992
rect 183419 526818 184365 526992
rect 184523 526818 184917 526992
rect 185259 526818 186205 526992
rect 186363 526818 186941 526992
rect 187283 526818 187401 526992
rect 172287 526550 172405 526724
rect 172563 526550 173509 526724
rect 173667 526550 174613 526724
rect 174771 526550 175717 526724
rect 175875 526550 176821 526724
rect 176979 526550 177189 526724
rect 177531 526550 178477 526724
rect 178635 526550 179581 526724
rect 179739 526550 180685 526724
rect 180843 526550 181789 526724
rect 181947 526550 182341 526724
rect 182683 526550 183629 526724
rect 183787 526550 184733 526724
rect 184891 526550 185837 526724
rect 185995 526550 186941 526724
rect 187283 526550 187401 526724
rect 172287 525730 172405 525904
rect 172563 525730 173509 525904
rect 173667 525730 174613 525904
rect 174955 525730 175901 525904
rect 176059 525730 177005 525904
rect 177163 525730 178109 525904
rect 178267 525730 179213 525904
rect 179371 525730 179765 525904
rect 180107 525730 181053 525904
rect 181211 525730 182157 525904
rect 182315 525730 183261 525904
rect 183419 525730 184365 525904
rect 184523 525730 184917 525904
rect 185259 525730 186205 525904
rect 186363 525730 186941 525904
rect 187283 525730 187401 525904
rect 172287 525462 172405 525636
rect 172563 525462 173509 525636
rect 173667 525462 174613 525636
rect 174771 525462 175717 525636
rect 175875 525462 176821 525636
rect 176979 525462 177189 525636
rect 177531 525462 178477 525636
rect 178635 525462 179581 525636
rect 179739 525462 180685 525636
rect 180843 525462 181789 525636
rect 181947 525462 182341 525636
rect 182683 525462 183629 525636
rect 183787 525462 184733 525636
rect 184891 525462 185837 525636
rect 185995 525462 186941 525636
rect 187283 525462 187401 525636
rect 172287 524642 172405 524816
rect 172563 524642 173509 524816
rect 173667 524642 174613 524816
rect 174955 524642 175901 524816
rect 176059 524642 177005 524816
rect 177163 524642 178109 524816
rect 178267 524642 179213 524816
rect 179371 524642 179765 524816
rect 180107 524642 181053 524816
rect 181211 524642 182157 524816
rect 182315 524642 183261 524816
rect 183419 524642 184365 524816
rect 184523 524642 184917 524816
rect 185259 524642 186205 524816
rect 186363 524642 186941 524816
rect 187283 524642 187401 524816
rect 172287 524374 172405 524548
rect 172563 524374 173509 524548
rect 173667 524374 174613 524548
rect 174771 524374 175717 524548
rect 175875 524374 176821 524548
rect 176979 524374 177189 524548
rect 177531 524374 178477 524548
rect 178635 524374 179581 524548
rect 179739 524374 180685 524548
rect 180843 524374 181789 524548
rect 181947 524374 182341 524548
rect 182683 524374 183629 524548
rect 183787 524374 184733 524548
rect 184891 524374 185837 524548
rect 185995 524374 186941 524548
rect 187283 524374 187401 524548
rect 172287 523554 172405 523728
rect 172563 523554 173509 523728
rect 173667 523554 174613 523728
rect 174955 523554 175901 523728
rect 176059 523554 177005 523728
rect 177163 523554 178109 523728
rect 178267 523554 179213 523728
rect 179371 523554 179765 523728
rect 180107 523554 181053 523728
rect 181211 523554 182157 523728
rect 182315 523554 183261 523728
rect 183419 523554 184365 523728
rect 184523 523554 184917 523728
rect 185259 523554 186205 523728
rect 186363 523554 186941 523728
rect 187283 523554 187401 523728
rect 172287 523286 172405 523460
rect 172563 523286 173509 523460
rect 173667 523286 174613 523460
rect 174771 523286 175717 523460
rect 175875 523286 176821 523460
rect 176979 523286 177189 523460
rect 177531 523286 178477 523460
rect 178635 523286 179581 523460
rect 179739 523286 180685 523460
rect 180843 523286 181789 523460
rect 181947 523286 182341 523460
rect 182683 523286 183629 523460
rect 183787 523286 184733 523460
rect 184891 523286 185837 523460
rect 185995 523286 186941 523460
rect 187283 523286 187401 523460
rect 172287 522466 172405 522640
rect 172563 522466 173509 522640
rect 173667 522466 174613 522640
rect 174955 522466 175901 522640
rect 176059 522466 177005 522640
rect 177163 522466 178109 522640
rect 178267 522466 179213 522640
rect 179371 522466 179765 522640
rect 180107 522466 181053 522640
rect 181211 522466 182157 522640
rect 182315 522466 183261 522640
rect 183419 522466 184365 522640
rect 184523 522466 184917 522640
rect 185259 522466 186205 522640
rect 186363 522466 186941 522640
rect 187283 522466 187401 522640
rect 172287 522198 172405 522372
rect 172563 522198 173509 522372
rect 173667 522198 174613 522372
rect 174771 522198 175717 522372
rect 175875 522198 176821 522372
rect 176979 522198 177189 522372
rect 177531 522198 178477 522372
rect 178635 522198 179581 522372
rect 179739 522198 180685 522372
rect 180843 522198 181789 522372
rect 181947 522198 182341 522372
rect 182683 522198 183629 522372
rect 183787 522198 184733 522372
rect 184891 522198 185837 522372
rect 185995 522198 186941 522372
rect 187283 522198 187401 522372
rect 172287 521378 172405 521552
rect 172563 521378 173509 521552
rect 173667 521378 174613 521552
rect 174955 521378 175901 521552
rect 176059 521378 177005 521552
rect 177163 521378 178109 521552
rect 178267 521378 179213 521552
rect 179371 521378 179765 521552
rect 180107 521378 181053 521552
rect 181211 521378 182157 521552
rect 182315 521378 183261 521552
rect 183419 521378 184365 521552
rect 184523 521378 184917 521552
rect 185259 521378 186205 521552
rect 186363 521378 186941 521552
rect 187283 521378 187401 521552
rect 172287 521110 172405 521284
rect 172563 521110 173509 521284
rect 173667 521110 174613 521284
rect 174771 521110 175717 521284
rect 175875 521110 176821 521284
rect 176979 521110 177189 521284
rect 177531 521110 178477 521284
rect 178635 521110 179581 521284
rect 179739 521110 180685 521284
rect 180843 521110 181789 521284
rect 181947 521110 182341 521284
rect 182683 521110 183629 521284
rect 183787 521110 184733 521284
rect 184891 521110 185837 521284
rect 185995 521110 186941 521284
rect 187283 521110 187401 521284
rect 172287 520290 172405 520464
rect 172563 520290 173509 520464
rect 173667 520290 174613 520464
rect 174955 520290 175901 520464
rect 176059 520290 177005 520464
rect 177163 520290 178109 520464
rect 178267 520290 179213 520464
rect 179371 520290 179765 520464
rect 180107 520290 181053 520464
rect 181211 520290 182157 520464
rect 182315 520290 183261 520464
rect 183419 520290 184365 520464
rect 184523 520290 184917 520464
rect 185259 520290 186205 520464
rect 186363 520290 186941 520464
rect 187283 520290 187401 520464
rect 172287 520022 172405 520196
rect 172563 520022 173509 520196
rect 173667 520022 174613 520196
rect 174771 520022 175717 520196
rect 175875 520022 176821 520196
rect 176979 520022 177189 520196
rect 177531 520022 178477 520196
rect 178635 520022 179581 520196
rect 179739 520022 180685 520196
rect 180843 520022 181789 520196
rect 181947 520022 182341 520196
rect 182683 520022 183629 520196
rect 183787 520022 184733 520196
rect 184891 520022 185837 520196
rect 185995 520022 186941 520196
rect 187283 520022 187401 520196
rect 172287 519202 172405 519376
rect 172563 519202 173509 519376
rect 173667 519202 174613 519376
rect 174955 519202 175901 519376
rect 176059 519202 177005 519376
rect 177163 519202 178109 519376
rect 178267 519202 179213 519376
rect 179371 519202 179765 519376
rect 180107 519202 181053 519376
rect 181211 519202 182157 519376
rect 182315 519202 183261 519376
rect 183419 519202 184365 519376
rect 184523 519202 184917 519376
rect 185259 519202 186205 519376
rect 186363 519202 186941 519376
rect 187283 519202 187401 519376
rect 172287 518934 172405 519108
rect 172563 518934 173509 519108
rect 173667 518934 174613 519108
rect 174771 518934 175717 519108
rect 175875 518934 176821 519108
rect 176979 518934 177189 519108
rect 177531 518934 178477 519108
rect 178635 518934 179581 519108
rect 179739 518934 180685 519108
rect 180843 518934 181789 519108
rect 181947 518934 182341 519108
rect 182683 518934 183629 519108
rect 183787 518934 184733 519108
rect 184891 518934 185837 519108
rect 185995 518934 186941 519108
rect 187283 518934 187401 519108
rect 172287 518114 172405 518288
rect 172563 518114 173509 518288
rect 173667 518114 174613 518288
rect 174955 518114 175901 518288
rect 176059 518114 177005 518288
rect 177163 518114 178109 518288
rect 178267 518114 179213 518288
rect 179371 518114 179765 518288
rect 180107 518114 181053 518288
rect 181211 518114 182157 518288
rect 182315 518114 183261 518288
rect 183419 518114 184365 518288
rect 184523 518114 184917 518288
rect 185259 518114 186205 518288
rect 186363 518114 186941 518288
rect 187283 518114 187401 518288
rect 172287 517846 172405 518020
rect 172563 517846 173509 518020
rect 173667 517846 174613 518020
rect 174771 517846 175717 518020
rect 175875 517846 176821 518020
rect 176979 517846 177189 518020
rect 177531 517846 178477 518020
rect 178635 517846 179581 518020
rect 179739 517846 180685 518020
rect 180843 517846 181789 518020
rect 181947 517846 182341 518020
rect 182683 517846 183629 518020
rect 183787 517846 184733 518020
rect 184891 517846 185837 518020
rect 185995 517846 186941 518020
rect 187283 517846 187401 518020
rect 172287 517026 172405 517200
rect 172563 517026 173509 517200
rect 173667 517026 174613 517200
rect 174955 517026 175901 517200
rect 176059 517026 177005 517200
rect 177163 517026 178109 517200
rect 178267 517026 179213 517200
rect 179371 517026 179765 517200
rect 180107 517026 181053 517200
rect 181211 517026 182157 517200
rect 182315 517026 183261 517200
rect 183419 517026 184365 517200
rect 184523 517026 184917 517200
rect 185259 517026 186205 517200
rect 186363 517026 186941 517200
rect 187283 517026 187401 517200
rect 172287 516758 172405 516932
rect 172563 516758 173509 516932
rect 173667 516758 174613 516932
rect 174771 516758 175717 516932
rect 175875 516758 176821 516932
rect 176979 516758 177189 516932
rect 177531 516758 178477 516932
rect 178635 516758 179581 516932
rect 179739 516758 180685 516932
rect 180843 516758 181789 516932
rect 181947 516758 182341 516932
rect 182683 516758 183629 516932
rect 183787 516758 184733 516932
rect 184891 516758 185837 516932
rect 185995 516758 186941 516932
rect 187283 516758 187401 516932
rect 172287 515938 172405 516112
rect 172563 515938 173509 516112
rect 173667 515938 174613 516112
rect 174955 515938 175901 516112
rect 176059 515938 177005 516112
rect 177163 515938 178109 516112
rect 178267 515938 179213 516112
rect 179371 515938 179765 516112
rect 180107 515938 181053 516112
rect 181211 515938 182157 516112
rect 182315 515938 183261 516112
rect 183419 515938 184365 516112
rect 184523 515938 184917 516112
rect 185259 515938 186205 516112
rect 186363 515938 186941 516112
rect 187283 515938 187401 516112
rect 172287 515670 172405 515844
rect 172563 515670 173141 515844
rect 173484 515644 173514 515844
rect 173580 515644 173610 515844
rect 173666 515644 173696 515844
rect 173752 515644 173782 515844
rect 173838 515644 173868 515844
rect 174035 515670 174613 515844
rect 174955 515670 175901 515844
rect 176059 515670 177005 515844
rect 177163 515670 177281 515844
rect 177531 515670 178477 515844
rect 178635 515670 179581 515844
rect 179739 515670 179857 515844
rect 180107 515670 181053 515844
rect 181211 515670 181789 515844
rect 182131 515686 182161 515844
rect 182219 515686 182249 515844
rect 182683 515670 183629 515844
rect 183787 515670 184733 515844
rect 184891 515670 185009 515844
rect 185259 515670 186205 515844
rect 186456 515644 186486 515844
rect 186552 515644 186582 515844
rect 186638 515644 186668 515844
rect 186724 515644 186754 515844
rect 186810 515644 186840 515844
rect 187007 515670 187125 515844
rect 187283 515670 187401 515844
<< ndiff >>
rect 164672 541035 164730 541047
rect 164672 540059 164684 541035
rect 164718 540059 164730 541035
rect 164672 540047 164730 540059
rect 164760 541035 164818 541047
rect 164760 540059 164772 541035
rect 164806 540059 164818 541035
rect 164760 540047 164818 540059
rect 164875 541042 164937 541054
rect 164875 540066 164887 541042
rect 164921 540066 164937 541042
rect 164875 540054 164937 540066
rect 164967 541042 165033 541054
rect 164967 540066 164983 541042
rect 165017 540066 165033 541042
rect 164967 540054 165033 540066
rect 165063 541042 165129 541054
rect 165063 540066 165079 541042
rect 165113 540066 165129 541042
rect 165063 540054 165129 540066
rect 165159 541042 165225 541054
rect 165159 540066 165175 541042
rect 165209 540066 165225 541042
rect 165159 540054 165225 540066
rect 165255 541042 165321 541054
rect 165255 540066 165271 541042
rect 165305 540066 165321 541042
rect 165255 540054 165321 540066
rect 165351 541042 165417 541054
rect 165351 540066 165367 541042
rect 165401 540066 165417 541042
rect 165351 540054 165417 540066
rect 165447 541042 165513 541054
rect 165447 540066 165463 541042
rect 165497 540066 165513 541042
rect 165447 540054 165513 540066
rect 165543 541042 165609 541054
rect 165543 540066 165559 541042
rect 165593 540066 165609 541042
rect 165543 540054 165609 540066
rect 165639 541042 165705 541054
rect 165639 540066 165655 541042
rect 165689 540066 165705 541042
rect 165639 540054 165705 540066
rect 165735 541042 165801 541054
rect 165735 540066 165751 541042
rect 165785 540066 165801 541042
rect 165735 540054 165801 540066
rect 165831 541042 165897 541054
rect 165831 540066 165847 541042
rect 165881 540066 165897 541042
rect 165831 540054 165897 540066
rect 165927 541042 165993 541054
rect 165927 540066 165943 541042
rect 165977 540066 165993 541042
rect 165927 540054 165993 540066
rect 166023 541042 166085 541054
rect 166023 540066 166039 541042
rect 166073 540066 166085 541042
rect 166352 541035 166410 541047
rect 166023 540054 166085 540066
rect 166152 540235 166210 540247
rect 166152 540059 166164 540235
rect 166198 540059 166210 540235
rect 166152 540047 166210 540059
rect 166240 540235 166298 540247
rect 166240 540059 166252 540235
rect 166286 540059 166298 540235
rect 166240 540047 166298 540059
rect 166352 540059 166364 541035
rect 166398 540059 166410 541035
rect 166352 540047 166410 540059
rect 166440 541035 166498 541047
rect 166440 540059 166452 541035
rect 166486 540059 166498 541035
rect 166440 540047 166498 540059
rect 168472 541035 168530 541047
rect 168472 540059 168484 541035
rect 168518 540059 168530 541035
rect 168472 540047 168530 540059
rect 168560 541035 168618 541047
rect 168560 540059 168572 541035
rect 168606 540059 168618 541035
rect 168560 540047 168618 540059
rect 168675 541042 168737 541054
rect 168675 540066 168687 541042
rect 168721 540066 168737 541042
rect 168675 540054 168737 540066
rect 168767 541042 168833 541054
rect 168767 540066 168783 541042
rect 168817 540066 168833 541042
rect 168767 540054 168833 540066
rect 168863 541042 168929 541054
rect 168863 540066 168879 541042
rect 168913 540066 168929 541042
rect 168863 540054 168929 540066
rect 168959 541042 169025 541054
rect 168959 540066 168975 541042
rect 169009 540066 169025 541042
rect 168959 540054 169025 540066
rect 169055 541042 169121 541054
rect 169055 540066 169071 541042
rect 169105 540066 169121 541042
rect 169055 540054 169121 540066
rect 169151 541042 169217 541054
rect 169151 540066 169167 541042
rect 169201 540066 169217 541042
rect 169151 540054 169217 540066
rect 169247 541042 169313 541054
rect 169247 540066 169263 541042
rect 169297 540066 169313 541042
rect 169247 540054 169313 540066
rect 169343 541042 169409 541054
rect 169343 540066 169359 541042
rect 169393 540066 169409 541042
rect 169343 540054 169409 540066
rect 169439 541042 169505 541054
rect 169439 540066 169455 541042
rect 169489 540066 169505 541042
rect 169439 540054 169505 540066
rect 169535 541042 169601 541054
rect 169535 540066 169551 541042
rect 169585 540066 169601 541042
rect 169535 540054 169601 540066
rect 169631 541042 169697 541054
rect 169631 540066 169647 541042
rect 169681 540066 169697 541042
rect 169631 540054 169697 540066
rect 169727 541042 169793 541054
rect 169727 540066 169743 541042
rect 169777 540066 169793 541042
rect 169727 540054 169793 540066
rect 169823 541042 169885 541054
rect 169823 540066 169839 541042
rect 169873 540066 169885 541042
rect 170152 541035 170210 541047
rect 169823 540054 169885 540066
rect 169952 540235 170010 540247
rect 169952 540059 169964 540235
rect 169998 540059 170010 540235
rect 169952 540047 170010 540059
rect 170040 540235 170098 540247
rect 170040 540059 170052 540235
rect 170086 540059 170098 540235
rect 170040 540047 170098 540059
rect 170152 540059 170164 541035
rect 170198 540059 170210 541035
rect 170152 540047 170210 540059
rect 170240 541035 170298 541047
rect 170240 540059 170252 541035
rect 170286 540059 170298 541035
rect 170240 540047 170298 540059
rect 172172 541035 172230 541047
rect 172172 540059 172184 541035
rect 172218 540059 172230 541035
rect 172172 540047 172230 540059
rect 172260 541035 172318 541047
rect 172260 540059 172272 541035
rect 172306 540059 172318 541035
rect 172260 540047 172318 540059
rect 172375 541042 172437 541054
rect 172375 540066 172387 541042
rect 172421 540066 172437 541042
rect 172375 540054 172437 540066
rect 172467 541042 172533 541054
rect 172467 540066 172483 541042
rect 172517 540066 172533 541042
rect 172467 540054 172533 540066
rect 172563 541042 172629 541054
rect 172563 540066 172579 541042
rect 172613 540066 172629 541042
rect 172563 540054 172629 540066
rect 172659 541042 172725 541054
rect 172659 540066 172675 541042
rect 172709 540066 172725 541042
rect 172659 540054 172725 540066
rect 172755 541042 172821 541054
rect 172755 540066 172771 541042
rect 172805 540066 172821 541042
rect 172755 540054 172821 540066
rect 172851 541042 172917 541054
rect 172851 540066 172867 541042
rect 172901 540066 172917 541042
rect 172851 540054 172917 540066
rect 172947 541042 173013 541054
rect 172947 540066 172963 541042
rect 172997 540066 173013 541042
rect 172947 540054 173013 540066
rect 173043 541042 173109 541054
rect 173043 540066 173059 541042
rect 173093 540066 173109 541042
rect 173043 540054 173109 540066
rect 173139 541042 173205 541054
rect 173139 540066 173155 541042
rect 173189 540066 173205 541042
rect 173139 540054 173205 540066
rect 173235 541042 173301 541054
rect 173235 540066 173251 541042
rect 173285 540066 173301 541042
rect 173235 540054 173301 540066
rect 173331 541042 173397 541054
rect 173331 540066 173347 541042
rect 173381 540066 173397 541042
rect 173331 540054 173397 540066
rect 173427 541042 173493 541054
rect 173427 540066 173443 541042
rect 173477 540066 173493 541042
rect 173427 540054 173493 540066
rect 173523 541042 173585 541054
rect 173523 540066 173539 541042
rect 173573 540066 173585 541042
rect 173852 541035 173910 541047
rect 173523 540054 173585 540066
rect 173652 540235 173710 540247
rect 173652 540059 173664 540235
rect 173698 540059 173710 540235
rect 173652 540047 173710 540059
rect 173740 540235 173798 540247
rect 173740 540059 173752 540235
rect 173786 540059 173798 540235
rect 173740 540047 173798 540059
rect 173852 540059 173864 541035
rect 173898 540059 173910 541035
rect 173852 540047 173910 540059
rect 173940 541035 173998 541047
rect 173940 540059 173952 541035
rect 173986 540059 173998 541035
rect 173940 540047 173998 540059
rect 175672 541035 175730 541047
rect 175672 540059 175684 541035
rect 175718 540059 175730 541035
rect 175672 540047 175730 540059
rect 175760 541035 175818 541047
rect 175760 540059 175772 541035
rect 175806 540059 175818 541035
rect 175760 540047 175818 540059
rect 175875 541042 175937 541054
rect 175875 540066 175887 541042
rect 175921 540066 175937 541042
rect 175875 540054 175937 540066
rect 175967 541042 176033 541054
rect 175967 540066 175983 541042
rect 176017 540066 176033 541042
rect 175967 540054 176033 540066
rect 176063 541042 176129 541054
rect 176063 540066 176079 541042
rect 176113 540066 176129 541042
rect 176063 540054 176129 540066
rect 176159 541042 176225 541054
rect 176159 540066 176175 541042
rect 176209 540066 176225 541042
rect 176159 540054 176225 540066
rect 176255 541042 176321 541054
rect 176255 540066 176271 541042
rect 176305 540066 176321 541042
rect 176255 540054 176321 540066
rect 176351 541042 176417 541054
rect 176351 540066 176367 541042
rect 176401 540066 176417 541042
rect 176351 540054 176417 540066
rect 176447 541042 176513 541054
rect 176447 540066 176463 541042
rect 176497 540066 176513 541042
rect 176447 540054 176513 540066
rect 176543 541042 176609 541054
rect 176543 540066 176559 541042
rect 176593 540066 176609 541042
rect 176543 540054 176609 540066
rect 176639 541042 176705 541054
rect 176639 540066 176655 541042
rect 176689 540066 176705 541042
rect 176639 540054 176705 540066
rect 176735 541042 176801 541054
rect 176735 540066 176751 541042
rect 176785 540066 176801 541042
rect 176735 540054 176801 540066
rect 176831 541042 176897 541054
rect 176831 540066 176847 541042
rect 176881 540066 176897 541042
rect 176831 540054 176897 540066
rect 176927 541042 176993 541054
rect 176927 540066 176943 541042
rect 176977 540066 176993 541042
rect 176927 540054 176993 540066
rect 177023 541042 177085 541054
rect 177023 540066 177039 541042
rect 177073 540066 177085 541042
rect 177352 541035 177410 541047
rect 177023 540054 177085 540066
rect 177152 540235 177210 540247
rect 177152 540059 177164 540235
rect 177198 540059 177210 540235
rect 177152 540047 177210 540059
rect 177240 540235 177298 540247
rect 177240 540059 177252 540235
rect 177286 540059 177298 540235
rect 177240 540047 177298 540059
rect 177352 540059 177364 541035
rect 177398 540059 177410 541035
rect 177352 540047 177410 540059
rect 177440 541035 177498 541047
rect 177440 540059 177452 541035
rect 177486 540059 177498 541035
rect 177440 540047 177498 540059
rect 179272 541035 179330 541047
rect 179272 540059 179284 541035
rect 179318 540059 179330 541035
rect 179272 540047 179330 540059
rect 179360 541035 179418 541047
rect 179360 540059 179372 541035
rect 179406 540059 179418 541035
rect 179360 540047 179418 540059
rect 179475 541042 179537 541054
rect 179475 540066 179487 541042
rect 179521 540066 179537 541042
rect 179475 540054 179537 540066
rect 179567 541042 179633 541054
rect 179567 540066 179583 541042
rect 179617 540066 179633 541042
rect 179567 540054 179633 540066
rect 179663 541042 179729 541054
rect 179663 540066 179679 541042
rect 179713 540066 179729 541042
rect 179663 540054 179729 540066
rect 179759 541042 179825 541054
rect 179759 540066 179775 541042
rect 179809 540066 179825 541042
rect 179759 540054 179825 540066
rect 179855 541042 179921 541054
rect 179855 540066 179871 541042
rect 179905 540066 179921 541042
rect 179855 540054 179921 540066
rect 179951 541042 180017 541054
rect 179951 540066 179967 541042
rect 180001 540066 180017 541042
rect 179951 540054 180017 540066
rect 180047 541042 180113 541054
rect 180047 540066 180063 541042
rect 180097 540066 180113 541042
rect 180047 540054 180113 540066
rect 180143 541042 180209 541054
rect 180143 540066 180159 541042
rect 180193 540066 180209 541042
rect 180143 540054 180209 540066
rect 180239 541042 180305 541054
rect 180239 540066 180255 541042
rect 180289 540066 180305 541042
rect 180239 540054 180305 540066
rect 180335 541042 180401 541054
rect 180335 540066 180351 541042
rect 180385 540066 180401 541042
rect 180335 540054 180401 540066
rect 180431 541042 180497 541054
rect 180431 540066 180447 541042
rect 180481 540066 180497 541042
rect 180431 540054 180497 540066
rect 180527 541042 180593 541054
rect 180527 540066 180543 541042
rect 180577 540066 180593 541042
rect 180527 540054 180593 540066
rect 180623 541042 180685 541054
rect 180623 540066 180639 541042
rect 180673 540066 180685 541042
rect 180952 541035 181010 541047
rect 180623 540054 180685 540066
rect 180752 540235 180810 540247
rect 180752 540059 180764 540235
rect 180798 540059 180810 540235
rect 180752 540047 180810 540059
rect 180840 540235 180898 540247
rect 180840 540059 180852 540235
rect 180886 540059 180898 540235
rect 180840 540047 180898 540059
rect 180952 540059 180964 541035
rect 180998 540059 181010 541035
rect 180952 540047 181010 540059
rect 181040 541035 181098 541047
rect 181040 540059 181052 541035
rect 181086 540059 181098 541035
rect 181040 540047 181098 540059
rect 182572 541035 182630 541047
rect 182572 540059 182584 541035
rect 182618 540059 182630 541035
rect 182572 540047 182630 540059
rect 182660 541035 182718 541047
rect 182660 540059 182672 541035
rect 182706 540059 182718 541035
rect 182660 540047 182718 540059
rect 182775 541042 182837 541054
rect 182775 540066 182787 541042
rect 182821 540066 182837 541042
rect 182775 540054 182837 540066
rect 182867 541042 182933 541054
rect 182867 540066 182883 541042
rect 182917 540066 182933 541042
rect 182867 540054 182933 540066
rect 182963 541042 183029 541054
rect 182963 540066 182979 541042
rect 183013 540066 183029 541042
rect 182963 540054 183029 540066
rect 183059 541042 183125 541054
rect 183059 540066 183075 541042
rect 183109 540066 183125 541042
rect 183059 540054 183125 540066
rect 183155 541042 183221 541054
rect 183155 540066 183171 541042
rect 183205 540066 183221 541042
rect 183155 540054 183221 540066
rect 183251 541042 183317 541054
rect 183251 540066 183267 541042
rect 183301 540066 183317 541042
rect 183251 540054 183317 540066
rect 183347 541042 183413 541054
rect 183347 540066 183363 541042
rect 183397 540066 183413 541042
rect 183347 540054 183413 540066
rect 183443 541042 183509 541054
rect 183443 540066 183459 541042
rect 183493 540066 183509 541042
rect 183443 540054 183509 540066
rect 183539 541042 183605 541054
rect 183539 540066 183555 541042
rect 183589 540066 183605 541042
rect 183539 540054 183605 540066
rect 183635 541042 183701 541054
rect 183635 540066 183651 541042
rect 183685 540066 183701 541042
rect 183635 540054 183701 540066
rect 183731 541042 183797 541054
rect 183731 540066 183747 541042
rect 183781 540066 183797 541042
rect 183731 540054 183797 540066
rect 183827 541042 183893 541054
rect 183827 540066 183843 541042
rect 183877 540066 183893 541042
rect 183827 540054 183893 540066
rect 183923 541042 183985 541054
rect 183923 540066 183939 541042
rect 183973 540066 183985 541042
rect 184252 541035 184310 541047
rect 183923 540054 183985 540066
rect 184052 540235 184110 540247
rect 184052 540059 184064 540235
rect 184098 540059 184110 540235
rect 184052 540047 184110 540059
rect 184140 540235 184198 540247
rect 184140 540059 184152 540235
rect 184186 540059 184198 540235
rect 184140 540047 184198 540059
rect 184252 540059 184264 541035
rect 184298 540059 184310 541035
rect 184252 540047 184310 540059
rect 184340 541035 184398 541047
rect 184340 540059 184352 541035
rect 184386 540059 184398 541035
rect 184340 540047 184398 540059
rect 185872 541035 185930 541047
rect 185872 540059 185884 541035
rect 185918 540059 185930 541035
rect 185872 540047 185930 540059
rect 185960 541035 186018 541047
rect 185960 540059 185972 541035
rect 186006 540059 186018 541035
rect 185960 540047 186018 540059
rect 186075 541042 186137 541054
rect 186075 540066 186087 541042
rect 186121 540066 186137 541042
rect 186075 540054 186137 540066
rect 186167 541042 186233 541054
rect 186167 540066 186183 541042
rect 186217 540066 186233 541042
rect 186167 540054 186233 540066
rect 186263 541042 186329 541054
rect 186263 540066 186279 541042
rect 186313 540066 186329 541042
rect 186263 540054 186329 540066
rect 186359 541042 186425 541054
rect 186359 540066 186375 541042
rect 186409 540066 186425 541042
rect 186359 540054 186425 540066
rect 186455 541042 186521 541054
rect 186455 540066 186471 541042
rect 186505 540066 186521 541042
rect 186455 540054 186521 540066
rect 186551 541042 186617 541054
rect 186551 540066 186567 541042
rect 186601 540066 186617 541042
rect 186551 540054 186617 540066
rect 186647 541042 186713 541054
rect 186647 540066 186663 541042
rect 186697 540066 186713 541042
rect 186647 540054 186713 540066
rect 186743 541042 186809 541054
rect 186743 540066 186759 541042
rect 186793 540066 186809 541042
rect 186743 540054 186809 540066
rect 186839 541042 186905 541054
rect 186839 540066 186855 541042
rect 186889 540066 186905 541042
rect 186839 540054 186905 540066
rect 186935 541042 187001 541054
rect 186935 540066 186951 541042
rect 186985 540066 187001 541042
rect 186935 540054 187001 540066
rect 187031 541042 187097 541054
rect 187031 540066 187047 541042
rect 187081 540066 187097 541042
rect 187031 540054 187097 540066
rect 187127 541042 187193 541054
rect 187127 540066 187143 541042
rect 187177 540066 187193 541042
rect 187127 540054 187193 540066
rect 187223 541042 187285 541054
rect 187223 540066 187239 541042
rect 187273 540066 187285 541042
rect 187552 541035 187610 541047
rect 187223 540054 187285 540066
rect 187352 540235 187410 540247
rect 187352 540059 187364 540235
rect 187398 540059 187410 540235
rect 187352 540047 187410 540059
rect 187440 540235 187498 540247
rect 187440 540059 187452 540235
rect 187486 540059 187498 540235
rect 187440 540047 187498 540059
rect 187552 540059 187564 541035
rect 187598 540059 187610 541035
rect 187552 540047 187610 540059
rect 187640 541035 187698 541047
rect 187640 540059 187652 541035
rect 187686 540059 187698 541035
rect 187640 540047 187698 540059
rect 189172 541035 189230 541047
rect 189172 540059 189184 541035
rect 189218 540059 189230 541035
rect 189172 540047 189230 540059
rect 189260 541035 189318 541047
rect 189260 540059 189272 541035
rect 189306 540059 189318 541035
rect 189260 540047 189318 540059
rect 189375 541042 189437 541054
rect 189375 540066 189387 541042
rect 189421 540066 189437 541042
rect 189375 540054 189437 540066
rect 189467 541042 189533 541054
rect 189467 540066 189483 541042
rect 189517 540066 189533 541042
rect 189467 540054 189533 540066
rect 189563 541042 189629 541054
rect 189563 540066 189579 541042
rect 189613 540066 189629 541042
rect 189563 540054 189629 540066
rect 189659 541042 189725 541054
rect 189659 540066 189675 541042
rect 189709 540066 189725 541042
rect 189659 540054 189725 540066
rect 189755 541042 189821 541054
rect 189755 540066 189771 541042
rect 189805 540066 189821 541042
rect 189755 540054 189821 540066
rect 189851 541042 189917 541054
rect 189851 540066 189867 541042
rect 189901 540066 189917 541042
rect 189851 540054 189917 540066
rect 189947 541042 190013 541054
rect 189947 540066 189963 541042
rect 189997 540066 190013 541042
rect 189947 540054 190013 540066
rect 190043 541042 190109 541054
rect 190043 540066 190059 541042
rect 190093 540066 190109 541042
rect 190043 540054 190109 540066
rect 190139 541042 190205 541054
rect 190139 540066 190155 541042
rect 190189 540066 190205 541042
rect 190139 540054 190205 540066
rect 190235 541042 190301 541054
rect 190235 540066 190251 541042
rect 190285 540066 190301 541042
rect 190235 540054 190301 540066
rect 190331 541042 190397 541054
rect 190331 540066 190347 541042
rect 190381 540066 190397 541042
rect 190331 540054 190397 540066
rect 190427 541042 190493 541054
rect 190427 540066 190443 541042
rect 190477 540066 190493 541042
rect 190427 540054 190493 540066
rect 190523 541042 190585 541054
rect 190523 540066 190539 541042
rect 190573 540066 190585 541042
rect 190852 541035 190910 541047
rect 190523 540054 190585 540066
rect 190652 540235 190710 540247
rect 190652 540059 190664 540235
rect 190698 540059 190710 540235
rect 190652 540047 190710 540059
rect 190740 540235 190798 540247
rect 190740 540059 190752 540235
rect 190786 540059 190798 540235
rect 190740 540047 190798 540059
rect 190852 540059 190864 541035
rect 190898 540059 190910 541035
rect 190852 540047 190910 540059
rect 190940 541035 190998 541047
rect 190940 540059 190952 541035
rect 190986 540059 190998 541035
rect 190940 540047 190998 540059
rect 158652 538385 158710 538397
rect 158652 538209 158664 538385
rect 158698 538209 158710 538385
rect 158652 538197 158710 538209
rect 158910 538385 158968 538397
rect 158910 538209 158922 538385
rect 158956 538209 158968 538385
rect 158910 538197 158968 538209
rect 159028 538385 159086 538397
rect 159028 538209 159040 538385
rect 159074 538209 159086 538385
rect 159028 538197 159086 538209
rect 159286 538385 159344 538397
rect 159286 538209 159298 538385
rect 159332 538209 159344 538385
rect 159286 538197 159344 538209
rect 159544 538385 159602 538397
rect 159544 538209 159556 538385
rect 159590 538209 159602 538385
rect 159544 538197 159602 538209
rect 159802 538385 159860 538397
rect 159802 538209 159814 538385
rect 159848 538209 159860 538385
rect 159802 538197 159860 538209
rect 160060 538385 160118 538397
rect 160060 538209 160072 538385
rect 160106 538209 160118 538385
rect 160060 538197 160118 538209
rect 160318 538385 160376 538397
rect 160318 538209 160330 538385
rect 160364 538209 160376 538385
rect 160318 538197 160376 538209
rect 160576 538385 160634 538397
rect 160576 538209 160588 538385
rect 160622 538209 160634 538385
rect 160576 538197 160634 538209
rect 160834 538385 160892 538397
rect 160834 538209 160846 538385
rect 160880 538209 160892 538385
rect 160834 538197 160892 538209
rect 161092 538385 161150 538397
rect 161092 538209 161104 538385
rect 161138 538209 161150 538385
rect 161092 538197 161150 538209
rect 161350 538385 161408 538397
rect 161350 538209 161362 538385
rect 161396 538209 161408 538385
rect 161350 538197 161408 538209
rect 161472 538385 161530 538397
rect 161472 538209 161484 538385
rect 161518 538209 161530 538385
rect 161472 538197 161530 538209
rect 161730 538385 161788 538397
rect 161730 538209 161742 538385
rect 161776 538209 161788 538385
rect 161730 538197 161788 538209
rect 161872 538385 161930 538397
rect 161872 538209 161884 538385
rect 161918 538209 161930 538385
rect 161872 538197 161930 538209
rect 162130 538385 162188 538397
rect 162130 538209 162142 538385
rect 162176 538209 162188 538385
rect 162130 538197 162188 538209
rect 162252 538385 162310 538397
rect 162252 538209 162264 538385
rect 162298 538209 162310 538385
rect 162252 538197 162310 538209
rect 162510 538385 162568 538397
rect 162510 538209 162522 538385
rect 162556 538209 162568 538385
rect 162510 538197 162568 538209
rect 172235 530499 172287 530532
rect 172235 530465 172243 530499
rect 172277 530465 172287 530499
rect 172235 530422 172287 530465
rect 172405 530499 172457 530532
rect 172405 530465 172415 530499
rect 172449 530465 172457 530499
rect 172405 530422 172457 530465
rect 172513 530516 172571 530532
rect 172513 530482 172526 530516
rect 172560 530482 172571 530516
rect 172513 530448 172571 530482
rect 172601 530494 172657 530532
rect 172601 530460 172612 530494
rect 172646 530460 172657 530494
rect 172601 530448 172657 530460
rect 172687 530516 172743 530532
rect 172687 530482 172698 530516
rect 172732 530482 172743 530516
rect 172687 530448 172743 530482
rect 172773 530494 172829 530532
rect 172773 530460 172784 530494
rect 172818 530460 172829 530494
rect 172773 530448 172829 530460
rect 172859 530516 172926 530532
rect 172859 530482 172881 530516
rect 172915 530482 172926 530516
rect 172859 530448 172926 530482
rect 172956 530512 173009 530532
rect 172956 530478 172967 530512
rect 173001 530478 173009 530512
rect 172956 530448 173009 530478
rect 173063 530501 173115 530532
rect 173063 530467 173071 530501
rect 173105 530467 173115 530501
rect 173063 530422 173115 530467
rect 174061 530501 174113 530532
rect 174061 530467 174071 530501
rect 174105 530467 174113 530501
rect 174061 530422 174113 530467
rect 174167 530501 174219 530532
rect 174167 530467 174175 530501
rect 174209 530467 174219 530501
rect 174167 530422 174219 530467
rect 174613 530501 174665 530532
rect 174905 530516 174963 530532
rect 174613 530467 174623 530501
rect 174657 530467 174665 530501
rect 174613 530422 174665 530467
rect 174905 530482 174918 530516
rect 174952 530482 174963 530516
rect 174905 530448 174963 530482
rect 174993 530494 175049 530532
rect 174993 530460 175004 530494
rect 175038 530460 175049 530494
rect 174993 530448 175049 530460
rect 175079 530516 175135 530532
rect 175079 530482 175090 530516
rect 175124 530482 175135 530516
rect 175079 530448 175135 530482
rect 175165 530494 175221 530532
rect 175165 530460 175176 530494
rect 175210 530460 175221 530494
rect 175165 530448 175221 530460
rect 175251 530516 175318 530532
rect 175251 530482 175273 530516
rect 175307 530482 175318 530516
rect 175251 530448 175318 530482
rect 175348 530512 175401 530532
rect 175348 530478 175359 530512
rect 175393 530478 175401 530512
rect 175348 530448 175401 530478
rect 175547 530470 175599 530532
rect 175547 530436 175555 530470
rect 175589 530436 175599 530470
rect 175547 530402 175599 530436
rect 175629 530520 175701 530532
rect 175629 530486 175639 530520
rect 175673 530486 175701 530520
rect 175629 530448 175701 530486
rect 175755 530504 175807 530532
rect 175755 530470 175763 530504
rect 175797 530470 175807 530504
rect 175755 530448 175807 530470
rect 175837 530448 175898 530532
rect 175928 530524 176047 530532
rect 175928 530490 175981 530524
rect 176015 530490 176047 530524
rect 175928 530448 176047 530490
rect 176077 530460 176143 530532
rect 176173 530520 176252 530532
rect 176173 530486 176193 530520
rect 176227 530486 176252 530520
rect 176173 530460 176252 530486
rect 176282 530524 176351 530532
rect 176282 530490 176303 530524
rect 176337 530490 176351 530524
rect 176282 530460 176351 530490
rect 176077 530448 176127 530460
rect 175629 530402 175679 530448
rect 176297 530404 176351 530460
rect 176381 530520 176483 530532
rect 176381 530486 176415 530520
rect 176449 530486 176483 530520
rect 176381 530448 176483 530486
rect 176513 530448 176555 530532
rect 176585 530460 176721 530532
rect 176751 530518 176817 530532
rect 176751 530484 176761 530518
rect 176795 530484 176817 530518
rect 176751 530460 176817 530484
rect 176847 530518 176912 530532
rect 176847 530484 176868 530518
rect 176902 530484 176912 530518
rect 176847 530460 176912 530484
rect 176585 530448 176703 530460
rect 176381 530404 176431 530448
rect 176862 530448 176912 530460
rect 176942 530524 177047 530532
rect 176942 530490 177001 530524
rect 177035 530490 177047 530524
rect 176942 530448 177047 530490
rect 177115 530494 177167 530532
rect 177115 530460 177123 530494
rect 177157 530460 177167 530494
rect 177115 530448 177167 530460
rect 177197 530520 177251 530532
rect 177197 530486 177207 530520
rect 177241 530486 177251 530520
rect 177197 530448 177251 530486
rect 177281 530494 177333 530532
rect 177281 530460 177291 530494
rect 177325 530460 177333 530494
rect 177281 530448 177333 530460
rect 177682 530494 177734 530532
rect 177682 530460 177690 530494
rect 177724 530460 177734 530494
rect 177682 530402 177734 530460
rect 177764 530520 177829 530532
rect 177764 530486 177780 530520
rect 177814 530486 177829 530520
rect 177764 530448 177829 530486
rect 177929 530494 177981 530532
rect 177929 530460 177939 530494
rect 177973 530460 177981 530494
rect 177929 530448 177981 530460
rect 178035 530494 178087 530532
rect 178035 530460 178043 530494
rect 178077 530460 178087 530494
rect 178035 530448 178087 530460
rect 178187 530520 178241 530532
rect 178187 530486 178197 530520
rect 178231 530486 178241 530520
rect 178187 530448 178241 530486
rect 178271 530494 178323 530532
rect 178271 530460 178281 530494
rect 178315 530460 178323 530494
rect 178271 530448 178323 530460
rect 178399 530490 178451 530532
rect 178399 530456 178407 530490
rect 178441 530456 178451 530490
rect 177764 530402 177814 530448
rect 178399 530428 178451 530456
rect 178481 530520 178539 530532
rect 178481 530486 178493 530520
rect 178527 530486 178539 530520
rect 178481 530428 178539 530486
rect 178569 530507 178621 530532
rect 178569 530473 178579 530507
rect 178613 530473 178621 530507
rect 178569 530428 178621 530473
rect 178677 530516 178735 530532
rect 178677 530482 178690 530516
rect 178724 530482 178735 530516
rect 178677 530448 178735 530482
rect 178765 530494 178821 530532
rect 178765 530460 178776 530494
rect 178810 530460 178821 530494
rect 178765 530448 178821 530460
rect 178851 530516 178907 530532
rect 178851 530482 178862 530516
rect 178896 530482 178907 530516
rect 178851 530448 178907 530482
rect 178937 530494 178993 530532
rect 178937 530460 178948 530494
rect 178982 530460 178993 530494
rect 178937 530448 178993 530460
rect 179023 530516 179090 530532
rect 179023 530482 179045 530516
rect 179079 530482 179090 530516
rect 179023 530448 179090 530482
rect 179120 530512 179173 530532
rect 179120 530478 179131 530512
rect 179165 530478 179173 530512
rect 179120 530448 179173 530478
rect 179227 530512 179280 530532
rect 179227 530478 179235 530512
rect 179269 530478 179280 530512
rect 179227 530448 179280 530478
rect 179310 530516 179377 530532
rect 179310 530482 179321 530516
rect 179355 530482 179377 530516
rect 179310 530448 179377 530482
rect 179407 530494 179463 530532
rect 179407 530460 179418 530494
rect 179452 530460 179463 530494
rect 179407 530448 179463 530460
rect 179493 530516 179549 530532
rect 179493 530482 179504 530516
rect 179538 530482 179549 530516
rect 179493 530448 179549 530482
rect 179579 530494 179635 530532
rect 179579 530460 179590 530494
rect 179624 530460 179635 530494
rect 179579 530448 179635 530460
rect 179665 530516 179723 530532
rect 179665 530482 179676 530516
rect 179710 530482 179723 530516
rect 179665 530448 179723 530482
rect 180239 530501 180291 530532
rect 180239 530467 180247 530501
rect 180281 530467 180291 530501
rect 180239 530402 180291 530467
rect 180321 530520 180400 530532
rect 180321 530486 180331 530520
rect 180365 530486 180400 530520
rect 180321 530448 180400 530486
rect 180430 530448 180496 530532
rect 180526 530505 180621 530532
rect 180526 530471 180538 530505
rect 180572 530471 180621 530505
rect 180526 530448 180621 530471
rect 180651 530448 180717 530532
rect 180747 530505 180885 530532
rect 180747 530471 180773 530505
rect 180807 530471 180841 530505
rect 180875 530471 180885 530505
rect 180747 530448 180885 530471
rect 180915 530505 180967 530532
rect 180915 530471 180925 530505
rect 180959 530471 180967 530505
rect 180915 530448 180967 530471
rect 181205 530505 181257 530532
rect 181205 530471 181213 530505
rect 181247 530471 181257 530505
rect 181205 530448 181257 530471
rect 181287 530505 181425 530532
rect 181287 530471 181297 530505
rect 181331 530471 181365 530505
rect 181399 530471 181425 530505
rect 181287 530448 181425 530471
rect 181455 530448 181521 530532
rect 181551 530505 181646 530532
rect 181551 530471 181600 530505
rect 181634 530471 181646 530505
rect 181551 530448 181646 530471
rect 181676 530448 181742 530532
rect 181772 530520 181851 530532
rect 181772 530486 181807 530520
rect 181841 530486 181851 530520
rect 181772 530448 181851 530486
rect 180321 530402 180373 530448
rect 181799 530402 181851 530448
rect 181881 530501 181933 530532
rect 181881 530467 181891 530501
rect 181925 530467 181933 530501
rect 181881 530402 181933 530467
rect 181987 530512 182040 530532
rect 181987 530478 181995 530512
rect 182029 530478 182040 530512
rect 181987 530448 182040 530478
rect 182070 530516 182137 530532
rect 182070 530482 182081 530516
rect 182115 530482 182137 530516
rect 182070 530448 182137 530482
rect 182167 530494 182223 530532
rect 182167 530460 182178 530494
rect 182212 530460 182223 530494
rect 182167 530448 182223 530460
rect 182253 530516 182309 530532
rect 182253 530482 182264 530516
rect 182298 530482 182309 530516
rect 182253 530448 182309 530482
rect 182339 530494 182395 530532
rect 182339 530460 182350 530494
rect 182384 530460 182395 530494
rect 182339 530448 182395 530460
rect 182425 530516 182483 530532
rect 182425 530482 182436 530516
rect 182470 530482 182483 530516
rect 182425 530448 182483 530482
rect 182631 530494 182683 530532
rect 182631 530460 182639 530494
rect 182673 530460 182683 530494
rect 182631 530422 182683 530460
rect 182893 530494 182945 530532
rect 182893 530460 182903 530494
rect 182937 530460 182945 530494
rect 182893 530422 182945 530460
rect 183091 530512 183144 530532
rect 183091 530478 183099 530512
rect 183133 530478 183144 530512
rect 183091 530448 183144 530478
rect 183174 530516 183241 530532
rect 183174 530482 183185 530516
rect 183219 530482 183241 530516
rect 183174 530448 183241 530482
rect 183271 530494 183327 530532
rect 183271 530460 183282 530494
rect 183316 530460 183327 530494
rect 183271 530448 183327 530460
rect 183357 530516 183413 530532
rect 183357 530482 183368 530516
rect 183402 530482 183413 530516
rect 183357 530448 183413 530482
rect 183443 530494 183499 530532
rect 183443 530460 183454 530494
rect 183488 530460 183499 530494
rect 183443 530448 183499 530460
rect 183529 530516 183587 530532
rect 183529 530482 183540 530516
rect 183574 530482 183587 530516
rect 183529 530448 183587 530482
rect 183643 530501 183695 530532
rect 183643 530467 183651 530501
rect 183685 530467 183695 530501
rect 183643 530422 183695 530467
rect 184641 530501 184693 530532
rect 184641 530467 184651 530501
rect 184685 530467 184693 530501
rect 184641 530422 184693 530467
rect 184747 530494 184799 530532
rect 184747 530460 184755 530494
rect 184789 530460 184799 530494
rect 184747 530422 184799 530460
rect 185009 530494 185061 530532
rect 185009 530460 185019 530494
rect 185053 530460 185061 530494
rect 185009 530422 185061 530460
rect 185207 530512 185260 530532
rect 185207 530478 185215 530512
rect 185249 530478 185260 530512
rect 185207 530448 185260 530478
rect 185290 530516 185357 530532
rect 185290 530482 185301 530516
rect 185335 530482 185357 530516
rect 185290 530448 185357 530482
rect 185387 530494 185443 530532
rect 185387 530460 185398 530494
rect 185432 530460 185443 530494
rect 185387 530448 185443 530460
rect 185473 530516 185529 530532
rect 185473 530482 185484 530516
rect 185518 530482 185529 530516
rect 185473 530448 185529 530482
rect 185559 530494 185615 530532
rect 185559 530460 185570 530494
rect 185604 530460 185615 530494
rect 185559 530448 185615 530460
rect 185645 530516 185703 530532
rect 185645 530482 185656 530516
rect 185690 530482 185703 530516
rect 185645 530448 185703 530482
rect 185759 530501 185811 530532
rect 185759 530467 185767 530501
rect 185801 530467 185811 530501
rect 185759 530422 185811 530467
rect 186757 530501 186809 530532
rect 186757 530467 186767 530501
rect 186801 530467 186809 530501
rect 186757 530422 186809 530467
rect 187231 530499 187283 530532
rect 187231 530465 187239 530499
rect 187273 530465 187283 530499
rect 187231 530422 187283 530465
rect 187401 530499 187453 530532
rect 187401 530465 187411 530499
rect 187445 530465 187453 530499
rect 187401 530422 187453 530465
rect 172235 529605 172287 529648
rect 172235 529571 172243 529605
rect 172277 529571 172287 529605
rect 172235 529538 172287 529571
rect 172405 529605 172457 529648
rect 172405 529571 172415 529605
rect 172449 529571 172457 529605
rect 172405 529538 172457 529571
rect 172511 529603 172563 529648
rect 172511 529569 172519 529603
rect 172553 529569 172563 529603
rect 172511 529538 172563 529569
rect 173509 529603 173561 529648
rect 173509 529569 173519 529603
rect 173553 529569 173561 529603
rect 173509 529538 173561 529569
rect 173615 529603 173667 529648
rect 173615 529569 173623 529603
rect 173657 529569 173667 529603
rect 173615 529538 173667 529569
rect 174613 529603 174665 529648
rect 175342 529622 175392 529668
rect 174613 529569 174623 529603
rect 174657 529569 174665 529603
rect 174613 529538 174665 529569
rect 174833 529610 174885 529622
rect 174833 529576 174841 529610
rect 174875 529576 174885 529610
rect 174833 529538 174885 529576
rect 174915 529584 174969 529622
rect 174915 529550 174925 529584
rect 174959 529550 174969 529584
rect 174915 529538 174969 529550
rect 175069 529610 175121 529622
rect 175069 529576 175079 529610
rect 175113 529576 175121 529610
rect 175069 529538 175121 529576
rect 175175 529610 175227 529622
rect 175175 529576 175183 529610
rect 175217 529576 175227 529610
rect 175175 529538 175227 529576
rect 175327 529584 175392 529622
rect 175327 529550 175342 529584
rect 175376 529550 175392 529584
rect 175327 529538 175392 529550
rect 175422 529610 175474 529668
rect 175422 529576 175432 529610
rect 175466 529576 175474 529610
rect 175422 529538 175474 529576
rect 175547 529610 175599 529622
rect 175547 529576 175555 529610
rect 175589 529576 175599 529610
rect 175547 529538 175599 529576
rect 175629 529584 175683 529622
rect 175629 529550 175639 529584
rect 175673 529550 175683 529584
rect 175629 529538 175683 529550
rect 175713 529610 175765 529622
rect 175713 529576 175723 529610
rect 175757 529576 175765 529610
rect 175713 529538 175765 529576
rect 175833 529580 175938 529622
rect 175833 529546 175845 529580
rect 175879 529546 175938 529580
rect 175833 529538 175938 529546
rect 175968 529610 176018 529622
rect 176449 529622 176499 529666
rect 176177 529610 176295 529622
rect 175968 529586 176033 529610
rect 175968 529552 175978 529586
rect 176012 529552 176033 529586
rect 175968 529538 176033 529552
rect 176063 529586 176129 529610
rect 176063 529552 176085 529586
rect 176119 529552 176129 529586
rect 176063 529538 176129 529552
rect 176159 529538 176295 529610
rect 176325 529538 176367 529622
rect 176397 529584 176499 529622
rect 176397 529550 176431 529584
rect 176465 529550 176499 529584
rect 176397 529538 176499 529550
rect 176529 529610 176583 529666
rect 177201 529622 177251 529668
rect 176753 529610 176803 529622
rect 176529 529580 176598 529610
rect 176529 529546 176543 529580
rect 176577 529546 176598 529580
rect 176529 529538 176598 529546
rect 176628 529584 176707 529610
rect 176628 529550 176653 529584
rect 176687 529550 176707 529584
rect 176628 529538 176707 529550
rect 176737 529538 176803 529610
rect 176833 529580 176952 529622
rect 176833 529546 176865 529580
rect 176899 529546 176952 529580
rect 176833 529538 176952 529546
rect 176982 529538 177043 529622
rect 177073 529600 177125 529622
rect 177073 529566 177083 529600
rect 177117 529566 177125 529600
rect 177073 529538 177125 529566
rect 177179 529584 177251 529622
rect 177179 529550 177207 529584
rect 177241 529550 177251 529584
rect 177179 529538 177251 529550
rect 177281 529634 177333 529668
rect 177281 529600 177291 529634
rect 177325 529600 177333 529634
rect 177281 529538 177333 529600
rect 178211 529622 178263 529668
rect 177617 529599 177669 529622
rect 177617 529565 177625 529599
rect 177659 529565 177669 529599
rect 177617 529538 177669 529565
rect 177699 529599 177837 529622
rect 177699 529565 177709 529599
rect 177743 529565 177777 529599
rect 177811 529565 177837 529599
rect 177699 529538 177837 529565
rect 177867 529538 177933 529622
rect 177963 529599 178058 529622
rect 177963 529565 178012 529599
rect 178046 529565 178058 529599
rect 177963 529538 178058 529565
rect 178088 529538 178154 529622
rect 178184 529584 178263 529622
rect 178184 529550 178219 529584
rect 178253 529550 178263 529584
rect 178184 529538 178263 529550
rect 178293 529603 178345 529668
rect 178293 529569 178303 529603
rect 178337 529569 178345 529603
rect 178293 529538 178345 529569
rect 178399 529634 178451 529668
rect 178399 529600 178407 529634
rect 178441 529600 178451 529634
rect 178399 529538 178451 529600
rect 178481 529622 178531 529668
rect 178481 529584 178553 529622
rect 178481 529550 178491 529584
rect 178525 529550 178553 529584
rect 178481 529538 178553 529550
rect 178607 529600 178659 529622
rect 178607 529566 178615 529600
rect 178649 529566 178659 529600
rect 178607 529538 178659 529566
rect 178689 529538 178750 529622
rect 178780 529580 178899 529622
rect 178780 529546 178833 529580
rect 178867 529546 178899 529580
rect 178780 529538 178899 529546
rect 178929 529610 178979 529622
rect 179149 529610 179203 529666
rect 178929 529538 178995 529610
rect 179025 529584 179104 529610
rect 179025 529550 179045 529584
rect 179079 529550 179104 529584
rect 179025 529538 179104 529550
rect 179134 529580 179203 529610
rect 179134 529546 179155 529580
rect 179189 529546 179203 529580
rect 179134 529538 179203 529546
rect 179233 529622 179283 529666
rect 179233 529584 179335 529622
rect 179233 529550 179267 529584
rect 179301 529550 179335 529584
rect 179233 529538 179335 529550
rect 179365 529538 179407 529622
rect 179437 529610 179555 529622
rect 179714 529610 179764 529622
rect 179437 529538 179573 529610
rect 179603 529586 179669 529610
rect 179603 529552 179613 529586
rect 179647 529552 179669 529586
rect 179603 529538 179669 529552
rect 179699 529586 179764 529610
rect 179699 529552 179720 529586
rect 179754 529552 179764 529586
rect 179699 529538 179764 529552
rect 179794 529580 179899 529622
rect 179794 529546 179853 529580
rect 179887 529546 179899 529580
rect 179794 529538 179899 529546
rect 179967 529610 180019 529622
rect 179967 529576 179975 529610
rect 180009 529576 180019 529610
rect 179967 529538 180019 529576
rect 180049 529584 180103 529622
rect 180049 529550 180059 529584
rect 180093 529550 180103 529584
rect 180049 529538 180103 529550
rect 180133 529610 180185 529622
rect 180133 529576 180143 529610
rect 180177 529576 180185 529610
rect 180133 529538 180185 529576
rect 180239 529610 180291 529622
rect 180239 529576 180247 529610
rect 180281 529576 180291 529610
rect 180239 529538 180291 529576
rect 180321 529584 180375 529622
rect 180321 529550 180331 529584
rect 180365 529550 180375 529584
rect 180321 529538 180375 529550
rect 180405 529610 180457 529622
rect 180405 529576 180415 529610
rect 180449 529576 180457 529610
rect 180405 529538 180457 529576
rect 180525 529580 180630 529622
rect 180525 529546 180537 529580
rect 180571 529546 180630 529580
rect 180525 529538 180630 529546
rect 180660 529610 180710 529622
rect 181141 529622 181191 529666
rect 180869 529610 180987 529622
rect 180660 529586 180725 529610
rect 180660 529552 180670 529586
rect 180704 529552 180725 529586
rect 180660 529538 180725 529552
rect 180755 529586 180821 529610
rect 180755 529552 180777 529586
rect 180811 529552 180821 529586
rect 180755 529538 180821 529552
rect 180851 529538 180987 529610
rect 181017 529538 181059 529622
rect 181089 529584 181191 529622
rect 181089 529550 181123 529584
rect 181157 529550 181191 529584
rect 181089 529538 181191 529550
rect 181221 529610 181275 529666
rect 181893 529622 181943 529668
rect 181445 529610 181495 529622
rect 181221 529580 181290 529610
rect 181221 529546 181235 529580
rect 181269 529546 181290 529580
rect 181221 529538 181290 529546
rect 181320 529584 181399 529610
rect 181320 529550 181345 529584
rect 181379 529550 181399 529584
rect 181320 529538 181399 529550
rect 181429 529538 181495 529610
rect 181525 529580 181644 529622
rect 181525 529546 181557 529580
rect 181591 529546 181644 529580
rect 181525 529538 181644 529546
rect 181674 529538 181735 529622
rect 181765 529600 181817 529622
rect 181765 529566 181775 529600
rect 181809 529566 181817 529600
rect 181765 529538 181817 529566
rect 181871 529584 181943 529622
rect 181871 529550 181899 529584
rect 181933 529550 181943 529584
rect 181871 529538 181943 529550
rect 181973 529634 182025 529668
rect 181973 529600 181983 529634
rect 182017 529600 182025 529634
rect 181973 529538 182025 529600
rect 182079 529610 182131 529648
rect 182079 529576 182087 529610
rect 182121 529576 182131 529610
rect 182079 529538 182131 529576
rect 182341 529610 182393 529648
rect 182341 529576 182351 529610
rect 182385 529576 182393 529610
rect 182341 529538 182393 529576
rect 182650 529610 182702 529668
rect 182650 529576 182658 529610
rect 182692 529576 182702 529610
rect 182650 529538 182702 529576
rect 182732 529622 182782 529668
rect 182732 529584 182797 529622
rect 182732 529550 182748 529584
rect 182782 529550 182797 529584
rect 182732 529538 182797 529550
rect 182897 529610 182949 529622
rect 182897 529576 182907 529610
rect 182941 529576 182949 529610
rect 182897 529538 182949 529576
rect 183003 529610 183055 529622
rect 183003 529576 183011 529610
rect 183045 529576 183055 529610
rect 183003 529538 183055 529576
rect 183155 529584 183209 529622
rect 183155 529550 183165 529584
rect 183199 529550 183209 529584
rect 183155 529538 183209 529550
rect 183239 529610 183291 529622
rect 183239 529576 183249 529610
rect 183283 529576 183291 529610
rect 183239 529538 183291 529576
rect 183367 529603 183419 529648
rect 183367 529569 183375 529603
rect 183409 529569 183419 529603
rect 183367 529538 183419 529569
rect 184365 529603 184417 529648
rect 184365 529569 184375 529603
rect 184409 529569 184417 529603
rect 184365 529538 184417 529569
rect 184471 529603 184523 529648
rect 184471 529569 184479 529603
rect 184513 529569 184523 529603
rect 184471 529538 184523 529569
rect 185469 529603 185521 529648
rect 185469 529569 185479 529603
rect 185513 529569 185521 529603
rect 185469 529538 185521 529569
rect 185575 529603 185627 529648
rect 185575 529569 185583 529603
rect 185617 529569 185627 529603
rect 185575 529538 185627 529569
rect 186573 529603 186625 529648
rect 186573 529569 186583 529603
rect 186617 529569 186625 529603
rect 186573 529538 186625 529569
rect 186679 529603 186731 529648
rect 186679 529569 186687 529603
rect 186721 529569 186731 529603
rect 186679 529538 186731 529569
rect 187125 529603 187177 529648
rect 187125 529569 187135 529603
rect 187169 529569 187177 529603
rect 187125 529538 187177 529569
rect 187231 529605 187283 529648
rect 187231 529571 187239 529605
rect 187273 529571 187283 529605
rect 187231 529538 187283 529571
rect 187401 529605 187453 529648
rect 187401 529571 187411 529605
rect 187445 529571 187453 529605
rect 187401 529538 187453 529571
rect 172235 529411 172287 529444
rect 172235 529377 172243 529411
rect 172277 529377 172287 529411
rect 172235 529334 172287 529377
rect 172405 529411 172457 529444
rect 172405 529377 172415 529411
rect 172449 529377 172457 529411
rect 172405 529334 172457 529377
rect 172511 529413 172563 529444
rect 172511 529379 172519 529413
rect 172553 529379 172563 529413
rect 172511 529334 172563 529379
rect 173509 529413 173561 529444
rect 173509 529379 173519 529413
rect 173553 529379 173561 529413
rect 173509 529334 173561 529379
rect 173615 529413 173667 529444
rect 173615 529379 173623 529413
rect 173657 529379 173667 529413
rect 173615 529334 173667 529379
rect 174613 529413 174665 529444
rect 174613 529379 174623 529413
rect 174657 529379 174665 529413
rect 174613 529334 174665 529379
rect 175133 529417 175185 529444
rect 175133 529383 175141 529417
rect 175175 529383 175185 529417
rect 175133 529360 175185 529383
rect 175215 529417 175353 529444
rect 175215 529383 175225 529417
rect 175259 529383 175293 529417
rect 175327 529383 175353 529417
rect 175215 529360 175353 529383
rect 175383 529360 175449 529444
rect 175479 529417 175574 529444
rect 175479 529383 175528 529417
rect 175562 529383 175574 529417
rect 175479 529360 175574 529383
rect 175604 529360 175670 529444
rect 175700 529432 175779 529444
rect 175700 529398 175735 529432
rect 175769 529398 175779 529432
rect 175700 529360 175779 529398
rect 175727 529314 175779 529360
rect 175809 529413 175861 529444
rect 175809 529379 175819 529413
rect 175853 529379 175861 529413
rect 175809 529314 175861 529379
rect 175932 529428 175985 529444
rect 175932 529394 175940 529428
rect 175974 529394 175985 529428
rect 175932 529360 175985 529394
rect 176015 529419 176071 529444
rect 176015 529385 176026 529419
rect 176060 529385 176071 529419
rect 176015 529360 176071 529385
rect 176101 529428 176157 529444
rect 176101 529394 176112 529428
rect 176146 529394 176157 529428
rect 176101 529360 176157 529394
rect 176187 529419 176243 529444
rect 176187 529385 176198 529419
rect 176232 529385 176243 529419
rect 176187 529360 176243 529385
rect 176273 529428 176329 529444
rect 176273 529394 176284 529428
rect 176318 529394 176329 529428
rect 176273 529360 176329 529394
rect 176359 529419 176415 529444
rect 176359 529385 176370 529419
rect 176404 529385 176415 529419
rect 176359 529360 176415 529385
rect 176445 529428 176501 529444
rect 176445 529394 176456 529428
rect 176490 529394 176501 529428
rect 176445 529360 176501 529394
rect 176531 529419 176587 529444
rect 176531 529385 176542 529419
rect 176576 529385 176587 529419
rect 176531 529360 176587 529385
rect 176617 529428 176672 529444
rect 176617 529394 176627 529428
rect 176661 529394 176672 529428
rect 176617 529360 176672 529394
rect 176702 529419 176758 529444
rect 176702 529385 176713 529419
rect 176747 529385 176758 529419
rect 176702 529360 176758 529385
rect 176788 529428 176844 529444
rect 176788 529394 176799 529428
rect 176833 529394 176844 529428
rect 176788 529360 176844 529394
rect 176874 529419 176930 529444
rect 176874 529385 176885 529419
rect 176919 529385 176930 529419
rect 176874 529360 176930 529385
rect 176960 529428 177016 529444
rect 176960 529394 176971 529428
rect 177005 529394 177016 529428
rect 176960 529360 177016 529394
rect 177046 529419 177102 529444
rect 177046 529385 177057 529419
rect 177091 529385 177102 529419
rect 177046 529360 177102 529385
rect 177132 529428 177188 529444
rect 177132 529394 177143 529428
rect 177177 529394 177188 529428
rect 177132 529360 177188 529394
rect 177218 529419 177274 529444
rect 177218 529385 177229 529419
rect 177263 529385 177274 529419
rect 177218 529360 177274 529385
rect 177304 529419 177360 529444
rect 177304 529385 177315 529419
rect 177349 529385 177360 529419
rect 177304 529360 177360 529385
rect 177390 529419 177446 529444
rect 177390 529385 177401 529419
rect 177435 529385 177446 529419
rect 177390 529360 177446 529385
rect 177476 529419 177532 529444
rect 177476 529385 177487 529419
rect 177521 529385 177532 529419
rect 177476 529360 177532 529385
rect 177562 529419 177618 529444
rect 177562 529385 177573 529419
rect 177607 529385 177618 529419
rect 177562 529360 177618 529385
rect 177648 529432 177701 529444
rect 177648 529398 177659 529432
rect 177693 529398 177701 529432
rect 177648 529360 177701 529398
rect 177755 529406 177807 529444
rect 177755 529372 177763 529406
rect 177797 529372 177807 529406
rect 177755 529360 177807 529372
rect 177837 529432 177891 529444
rect 177837 529398 177847 529432
rect 177881 529398 177891 529432
rect 177837 529360 177891 529398
rect 177921 529406 177973 529444
rect 177921 529372 177931 529406
rect 177965 529372 177973 529406
rect 177921 529360 177973 529372
rect 178041 529436 178146 529444
rect 178041 529402 178053 529436
rect 178087 529402 178146 529436
rect 178041 529360 178146 529402
rect 178176 529430 178241 529444
rect 178176 529396 178186 529430
rect 178220 529396 178241 529430
rect 178176 529372 178241 529396
rect 178271 529430 178337 529444
rect 178271 529396 178293 529430
rect 178327 529396 178337 529430
rect 178271 529372 178337 529396
rect 178367 529372 178503 529444
rect 178176 529360 178226 529372
rect 178385 529360 178503 529372
rect 178533 529360 178575 529444
rect 178605 529432 178707 529444
rect 178605 529398 178639 529432
rect 178673 529398 178707 529432
rect 178605 529360 178707 529398
rect 178657 529316 178707 529360
rect 178737 529436 178806 529444
rect 178737 529402 178751 529436
rect 178785 529402 178806 529436
rect 178737 529372 178806 529402
rect 178836 529432 178915 529444
rect 178836 529398 178861 529432
rect 178895 529398 178915 529432
rect 178836 529372 178915 529398
rect 178945 529372 179011 529444
rect 178737 529316 178791 529372
rect 178961 529360 179011 529372
rect 179041 529436 179160 529444
rect 179041 529402 179073 529436
rect 179107 529402 179160 529436
rect 179041 529360 179160 529402
rect 179190 529360 179251 529444
rect 179281 529416 179333 529444
rect 179281 529382 179291 529416
rect 179325 529382 179333 529416
rect 179281 529360 179333 529382
rect 179387 529432 179459 529444
rect 179387 529398 179415 529432
rect 179449 529398 179459 529432
rect 179387 529360 179459 529398
rect 179409 529314 179459 529360
rect 179489 529382 179541 529444
rect 179489 529348 179499 529382
rect 179533 529348 179541 529382
rect 179489 529314 179541 529348
rect 179687 529419 179739 529444
rect 179687 529385 179695 529419
rect 179729 529385 179739 529419
rect 179687 529340 179739 529385
rect 179769 529432 179827 529444
rect 179769 529398 179781 529432
rect 179815 529398 179827 529432
rect 179769 529340 179827 529398
rect 179857 529402 179909 529444
rect 179857 529368 179867 529402
rect 179901 529368 179909 529402
rect 179857 529340 179909 529368
rect 180055 529413 180107 529444
rect 180055 529379 180063 529413
rect 180097 529379 180107 529413
rect 180055 529334 180107 529379
rect 180501 529413 180553 529444
rect 180501 529379 180511 529413
rect 180545 529379 180553 529413
rect 180501 529334 180553 529379
rect 180699 529432 180752 529444
rect 180699 529398 180707 529432
rect 180741 529398 180752 529432
rect 180699 529360 180752 529398
rect 180782 529419 180838 529444
rect 180782 529385 180793 529419
rect 180827 529385 180838 529419
rect 180782 529360 180838 529385
rect 180868 529419 180924 529444
rect 180868 529385 180879 529419
rect 180913 529385 180924 529419
rect 180868 529360 180924 529385
rect 180954 529419 181010 529444
rect 180954 529385 180965 529419
rect 180999 529385 181010 529419
rect 180954 529360 181010 529385
rect 181040 529419 181096 529444
rect 181040 529385 181051 529419
rect 181085 529385 181096 529419
rect 181040 529360 181096 529385
rect 181126 529419 181182 529444
rect 181126 529385 181137 529419
rect 181171 529385 181182 529419
rect 181126 529360 181182 529385
rect 181212 529428 181268 529444
rect 181212 529394 181223 529428
rect 181257 529394 181268 529428
rect 181212 529360 181268 529394
rect 181298 529419 181354 529444
rect 181298 529385 181309 529419
rect 181343 529385 181354 529419
rect 181298 529360 181354 529385
rect 181384 529428 181440 529444
rect 181384 529394 181395 529428
rect 181429 529394 181440 529428
rect 181384 529360 181440 529394
rect 181470 529419 181526 529444
rect 181470 529385 181481 529419
rect 181515 529385 181526 529419
rect 181470 529360 181526 529385
rect 181556 529428 181612 529444
rect 181556 529394 181567 529428
rect 181601 529394 181612 529428
rect 181556 529360 181612 529394
rect 181642 529419 181698 529444
rect 181642 529385 181653 529419
rect 181687 529385 181698 529419
rect 181642 529360 181698 529385
rect 181728 529428 181783 529444
rect 181728 529394 181739 529428
rect 181773 529394 181783 529428
rect 181728 529360 181783 529394
rect 181813 529419 181869 529444
rect 181813 529385 181824 529419
rect 181858 529385 181869 529419
rect 181813 529360 181869 529385
rect 181899 529428 181955 529444
rect 181899 529394 181910 529428
rect 181944 529394 181955 529428
rect 181899 529360 181955 529394
rect 181985 529419 182041 529444
rect 181985 529385 181996 529419
rect 182030 529385 182041 529419
rect 181985 529360 182041 529385
rect 182071 529428 182127 529444
rect 182071 529394 182082 529428
rect 182116 529394 182127 529428
rect 182071 529360 182127 529394
rect 182157 529419 182213 529444
rect 182157 529385 182168 529419
rect 182202 529385 182213 529419
rect 182157 529360 182213 529385
rect 182243 529428 182299 529444
rect 182243 529394 182254 529428
rect 182288 529394 182299 529428
rect 182243 529360 182299 529394
rect 182329 529419 182385 529444
rect 182329 529385 182340 529419
rect 182374 529385 182385 529419
rect 182329 529360 182385 529385
rect 182415 529428 182468 529444
rect 182415 529394 182426 529428
rect 182460 529394 182468 529428
rect 182415 529360 182468 529394
rect 182539 529402 182591 529444
rect 182539 529368 182547 529402
rect 182581 529368 182591 529402
rect 182539 529340 182591 529368
rect 182621 529432 182679 529444
rect 182621 529398 182633 529432
rect 182667 529398 182679 529432
rect 182621 529340 182679 529398
rect 182709 529419 182761 529444
rect 182709 529385 182719 529419
rect 182753 529385 182761 529419
rect 182709 529340 182761 529385
rect 182815 529413 182867 529444
rect 182815 529379 182823 529413
rect 182857 529379 182867 529413
rect 182815 529334 182867 529379
rect 183813 529413 183865 529444
rect 183813 529379 183823 529413
rect 183857 529379 183865 529413
rect 183813 529334 183865 529379
rect 183919 529413 183971 529444
rect 183919 529379 183927 529413
rect 183961 529379 183971 529413
rect 183919 529334 183971 529379
rect 184917 529413 184969 529444
rect 184917 529379 184927 529413
rect 184961 529379 184969 529413
rect 184917 529334 184969 529379
rect 185207 529413 185259 529444
rect 185207 529379 185215 529413
rect 185249 529379 185259 529413
rect 185207 529334 185259 529379
rect 186205 529413 186257 529444
rect 186205 529379 186215 529413
rect 186249 529379 186257 529413
rect 186205 529334 186257 529379
rect 186311 529413 186363 529444
rect 186311 529379 186319 529413
rect 186353 529379 186363 529413
rect 186311 529334 186363 529379
rect 186941 529413 186993 529444
rect 186941 529379 186951 529413
rect 186985 529379 186993 529413
rect 186941 529334 186993 529379
rect 187231 529411 187283 529444
rect 187231 529377 187239 529411
rect 187273 529377 187283 529411
rect 187231 529334 187283 529377
rect 187401 529411 187453 529444
rect 187401 529377 187411 529411
rect 187445 529377 187453 529411
rect 187401 529334 187453 529377
rect 172235 528517 172287 528560
rect 172235 528483 172243 528517
rect 172277 528483 172287 528517
rect 172235 528450 172287 528483
rect 172405 528517 172457 528560
rect 172405 528483 172415 528517
rect 172449 528483 172457 528517
rect 172405 528450 172457 528483
rect 172511 528515 172563 528560
rect 172511 528481 172519 528515
rect 172553 528481 172563 528515
rect 172511 528450 172563 528481
rect 173509 528515 173561 528560
rect 173509 528481 173519 528515
rect 173553 528481 173561 528515
rect 173509 528450 173561 528481
rect 173615 528515 173667 528560
rect 173615 528481 173623 528515
rect 173657 528481 173667 528515
rect 173615 528450 173667 528481
rect 174613 528515 174665 528560
rect 174613 528481 174623 528515
rect 174657 528481 174665 528515
rect 174613 528450 174665 528481
rect 174719 528515 174771 528560
rect 174719 528481 174727 528515
rect 174761 528481 174771 528515
rect 174719 528450 174771 528481
rect 175717 528515 175769 528560
rect 175717 528481 175727 528515
rect 175761 528481 175769 528515
rect 175717 528450 175769 528481
rect 175915 528509 175967 528554
rect 175915 528475 175923 528509
rect 175957 528475 175967 528509
rect 175915 528450 175967 528475
rect 175997 528496 176055 528554
rect 175997 528462 176009 528496
rect 176043 528462 176055 528496
rect 175997 528450 176055 528462
rect 176085 528526 176137 528554
rect 176085 528492 176095 528526
rect 176129 528492 176137 528526
rect 176085 528450 176137 528492
rect 176191 528509 176243 528554
rect 176191 528475 176199 528509
rect 176233 528475 176243 528509
rect 176191 528450 176243 528475
rect 176273 528496 176331 528554
rect 176273 528462 176285 528496
rect 176319 528462 176331 528496
rect 176273 528450 176331 528462
rect 176361 528526 176413 528554
rect 177107 528534 177159 528580
rect 176361 528492 176371 528526
rect 176405 528492 176413 528526
rect 176361 528450 176413 528492
rect 176513 528511 176565 528534
rect 176513 528477 176521 528511
rect 176555 528477 176565 528511
rect 176513 528450 176565 528477
rect 176595 528511 176733 528534
rect 176595 528477 176605 528511
rect 176639 528477 176673 528511
rect 176707 528477 176733 528511
rect 176595 528450 176733 528477
rect 176763 528450 176829 528534
rect 176859 528511 176954 528534
rect 176859 528477 176908 528511
rect 176942 528477 176954 528511
rect 176859 528450 176954 528477
rect 176984 528450 177050 528534
rect 177080 528496 177159 528534
rect 177080 528462 177115 528496
rect 177149 528462 177159 528496
rect 177080 528450 177159 528462
rect 177189 528515 177241 528580
rect 177189 528481 177199 528515
rect 177233 528481 177241 528515
rect 177189 528450 177241 528481
rect 177498 528522 177550 528580
rect 177498 528488 177506 528522
rect 177540 528488 177550 528522
rect 177498 528450 177550 528488
rect 177580 528534 177630 528580
rect 177580 528496 177645 528534
rect 177580 528462 177596 528496
rect 177630 528462 177645 528496
rect 177580 528450 177645 528462
rect 177745 528522 177797 528534
rect 177745 528488 177755 528522
rect 177789 528488 177797 528522
rect 177745 528450 177797 528488
rect 177851 528522 177903 528534
rect 177851 528488 177859 528522
rect 177893 528488 177903 528522
rect 177851 528450 177903 528488
rect 178003 528496 178057 528534
rect 178003 528462 178013 528496
rect 178047 528462 178057 528496
rect 178003 528450 178057 528462
rect 178087 528522 178139 528534
rect 178087 528488 178097 528522
rect 178131 528488 178139 528522
rect 178087 528450 178139 528488
rect 178399 528496 178452 528534
rect 178399 528462 178407 528496
rect 178441 528462 178452 528496
rect 178399 528450 178452 528462
rect 178482 528509 178538 528534
rect 178482 528475 178493 528509
rect 178527 528475 178538 528509
rect 178482 528450 178538 528475
rect 178568 528509 178624 528534
rect 178568 528475 178579 528509
rect 178613 528475 178624 528509
rect 178568 528450 178624 528475
rect 178654 528509 178710 528534
rect 178654 528475 178665 528509
rect 178699 528475 178710 528509
rect 178654 528450 178710 528475
rect 178740 528509 178796 528534
rect 178740 528475 178751 528509
rect 178785 528475 178796 528509
rect 178740 528450 178796 528475
rect 178826 528509 178882 528534
rect 178826 528475 178837 528509
rect 178871 528475 178882 528509
rect 178826 528450 178882 528475
rect 178912 528500 178968 528534
rect 178912 528466 178923 528500
rect 178957 528466 178968 528500
rect 178912 528450 178968 528466
rect 178998 528509 179054 528534
rect 178998 528475 179009 528509
rect 179043 528475 179054 528509
rect 178998 528450 179054 528475
rect 179084 528500 179140 528534
rect 179084 528466 179095 528500
rect 179129 528466 179140 528500
rect 179084 528450 179140 528466
rect 179170 528509 179226 528534
rect 179170 528475 179181 528509
rect 179215 528475 179226 528509
rect 179170 528450 179226 528475
rect 179256 528500 179312 528534
rect 179256 528466 179267 528500
rect 179301 528466 179312 528500
rect 179256 528450 179312 528466
rect 179342 528509 179398 528534
rect 179342 528475 179353 528509
rect 179387 528475 179398 528509
rect 179342 528450 179398 528475
rect 179428 528500 179483 528534
rect 179428 528466 179439 528500
rect 179473 528466 179483 528500
rect 179428 528450 179483 528466
rect 179513 528509 179569 528534
rect 179513 528475 179524 528509
rect 179558 528475 179569 528509
rect 179513 528450 179569 528475
rect 179599 528500 179655 528534
rect 179599 528466 179610 528500
rect 179644 528466 179655 528500
rect 179599 528450 179655 528466
rect 179685 528509 179741 528534
rect 179685 528475 179696 528509
rect 179730 528475 179741 528509
rect 179685 528450 179741 528475
rect 179771 528500 179827 528534
rect 179771 528466 179782 528500
rect 179816 528466 179827 528500
rect 179771 528450 179827 528466
rect 179857 528509 179913 528534
rect 179857 528475 179868 528509
rect 179902 528475 179913 528509
rect 179857 528450 179913 528475
rect 179943 528500 179999 528534
rect 179943 528466 179954 528500
rect 179988 528466 179999 528500
rect 179943 528450 179999 528466
rect 180029 528509 180085 528534
rect 180029 528475 180040 528509
rect 180074 528475 180085 528509
rect 180029 528450 180085 528475
rect 180115 528500 180168 528534
rect 180115 528466 180126 528500
rect 180160 528466 180168 528500
rect 180115 528450 180168 528466
rect 180239 528509 180291 528554
rect 180239 528475 180247 528509
rect 180281 528475 180291 528509
rect 180239 528450 180291 528475
rect 180321 528496 180379 528554
rect 180321 528462 180333 528496
rect 180367 528462 180379 528496
rect 180321 528450 180379 528462
rect 180409 528526 180461 528554
rect 180409 528492 180419 528526
rect 180453 528492 180461 528526
rect 180409 528450 180461 528492
rect 180515 528522 180567 528534
rect 180515 528488 180523 528522
rect 180557 528488 180567 528522
rect 180515 528450 180567 528488
rect 180597 528496 180651 528534
rect 180597 528462 180607 528496
rect 180641 528462 180651 528496
rect 180597 528450 180651 528462
rect 180681 528522 180733 528534
rect 180681 528488 180691 528522
rect 180725 528488 180733 528522
rect 180681 528450 180733 528488
rect 180801 528492 180906 528534
rect 180801 528458 180813 528492
rect 180847 528458 180906 528492
rect 180801 528450 180906 528458
rect 180936 528522 180986 528534
rect 181417 528534 181467 528578
rect 181145 528522 181263 528534
rect 180936 528498 181001 528522
rect 180936 528464 180946 528498
rect 180980 528464 181001 528498
rect 180936 528450 181001 528464
rect 181031 528498 181097 528522
rect 181031 528464 181053 528498
rect 181087 528464 181097 528498
rect 181031 528450 181097 528464
rect 181127 528450 181263 528522
rect 181293 528450 181335 528534
rect 181365 528496 181467 528534
rect 181365 528462 181399 528496
rect 181433 528462 181467 528496
rect 181365 528450 181467 528462
rect 181497 528522 181551 528578
rect 182169 528534 182219 528580
rect 181721 528522 181771 528534
rect 181497 528492 181566 528522
rect 181497 528458 181511 528492
rect 181545 528458 181566 528492
rect 181497 528450 181566 528458
rect 181596 528496 181675 528522
rect 181596 528462 181621 528496
rect 181655 528462 181675 528496
rect 181596 528450 181675 528462
rect 181705 528450 181771 528522
rect 181801 528492 181920 528534
rect 181801 528458 181833 528492
rect 181867 528458 181920 528492
rect 181801 528450 181920 528458
rect 181950 528450 182011 528534
rect 182041 528512 182093 528534
rect 182041 528478 182051 528512
rect 182085 528478 182093 528512
rect 182041 528450 182093 528478
rect 182147 528496 182219 528534
rect 182147 528462 182175 528496
rect 182209 528462 182219 528496
rect 182147 528450 182219 528462
rect 182249 528546 182301 528580
rect 182249 528512 182259 528546
rect 182293 528512 182301 528546
rect 182249 528450 182301 528512
rect 182631 528515 182683 528560
rect 182631 528481 182639 528515
rect 182673 528481 182683 528515
rect 182631 528450 182683 528481
rect 183629 528515 183681 528560
rect 183629 528481 183639 528515
rect 183673 528481 183681 528515
rect 183629 528450 183681 528481
rect 183735 528515 183787 528560
rect 183735 528481 183743 528515
rect 183777 528481 183787 528515
rect 183735 528450 183787 528481
rect 184733 528515 184785 528560
rect 184733 528481 184743 528515
rect 184777 528481 184785 528515
rect 184733 528450 184785 528481
rect 184839 528515 184891 528560
rect 184839 528481 184847 528515
rect 184881 528481 184891 528515
rect 184839 528450 184891 528481
rect 185837 528515 185889 528560
rect 185837 528481 185847 528515
rect 185881 528481 185889 528515
rect 185837 528450 185889 528481
rect 185943 528515 185995 528560
rect 185943 528481 185951 528515
rect 185985 528481 185995 528515
rect 185943 528450 185995 528481
rect 186941 528515 186993 528560
rect 186941 528481 186951 528515
rect 186985 528481 186993 528515
rect 186941 528450 186993 528481
rect 187231 528517 187283 528560
rect 187231 528483 187239 528517
rect 187273 528483 187283 528517
rect 187231 528450 187283 528483
rect 187401 528517 187453 528560
rect 187401 528483 187411 528517
rect 187445 528483 187453 528517
rect 187401 528450 187453 528483
rect 172235 528323 172287 528356
rect 172235 528289 172243 528323
rect 172277 528289 172287 528323
rect 172235 528246 172287 528289
rect 172405 528323 172457 528356
rect 172405 528289 172415 528323
rect 172449 528289 172457 528323
rect 172405 528246 172457 528289
rect 172511 528325 172563 528356
rect 172511 528291 172519 528325
rect 172553 528291 172563 528325
rect 172511 528246 172563 528291
rect 173509 528325 173561 528356
rect 173509 528291 173519 528325
rect 173553 528291 173561 528325
rect 173509 528246 173561 528291
rect 173615 528325 173667 528356
rect 173615 528291 173623 528325
rect 173657 528291 173667 528325
rect 173615 528246 173667 528291
rect 174613 528325 174665 528356
rect 174613 528291 174623 528325
rect 174657 528291 174665 528325
rect 174613 528246 174665 528291
rect 174903 528325 174955 528356
rect 174903 528291 174911 528325
rect 174945 528291 174955 528325
rect 174903 528246 174955 528291
rect 175901 528325 175953 528356
rect 175901 528291 175911 528325
rect 175945 528291 175953 528325
rect 175901 528246 175953 528291
rect 176099 528318 176151 528356
rect 176099 528284 176107 528318
rect 176141 528284 176151 528318
rect 176099 528272 176151 528284
rect 176181 528344 176235 528356
rect 176181 528310 176191 528344
rect 176225 528310 176235 528344
rect 176181 528272 176235 528310
rect 176265 528318 176317 528356
rect 176265 528284 176275 528318
rect 176309 528284 176317 528318
rect 176265 528272 176317 528284
rect 176385 528348 176490 528356
rect 176385 528314 176397 528348
rect 176431 528314 176490 528348
rect 176385 528272 176490 528314
rect 176520 528342 176585 528356
rect 176520 528308 176530 528342
rect 176564 528308 176585 528342
rect 176520 528284 176585 528308
rect 176615 528342 176681 528356
rect 176615 528308 176637 528342
rect 176671 528308 176681 528342
rect 176615 528284 176681 528308
rect 176711 528284 176847 528356
rect 176520 528272 176570 528284
rect 176729 528272 176847 528284
rect 176877 528272 176919 528356
rect 176949 528344 177051 528356
rect 176949 528310 176983 528344
rect 177017 528310 177051 528344
rect 176949 528272 177051 528310
rect 177001 528228 177051 528272
rect 177081 528348 177150 528356
rect 177081 528314 177095 528348
rect 177129 528314 177150 528348
rect 177081 528284 177150 528314
rect 177180 528344 177259 528356
rect 177180 528310 177205 528344
rect 177239 528310 177259 528344
rect 177180 528284 177259 528310
rect 177289 528284 177355 528356
rect 177081 528228 177135 528284
rect 177305 528272 177355 528284
rect 177385 528348 177504 528356
rect 177385 528314 177417 528348
rect 177451 528314 177504 528348
rect 177385 528272 177504 528314
rect 177534 528272 177595 528356
rect 177625 528328 177677 528356
rect 177625 528294 177635 528328
rect 177669 528294 177677 528328
rect 177625 528272 177677 528294
rect 177731 528344 177803 528356
rect 177731 528310 177759 528344
rect 177793 528310 177803 528344
rect 177731 528272 177803 528310
rect 177753 528226 177803 528272
rect 177833 528294 177885 528356
rect 177833 528260 177843 528294
rect 177877 528260 177885 528294
rect 177833 528226 177885 528260
rect 177939 528314 177991 528356
rect 177939 528280 177947 528314
rect 177981 528280 177991 528314
rect 177939 528252 177991 528280
rect 178021 528344 178079 528356
rect 178021 528310 178033 528344
rect 178067 528310 178079 528344
rect 178021 528252 178079 528310
rect 178109 528331 178161 528356
rect 178109 528297 178119 528331
rect 178153 528297 178161 528331
rect 178109 528252 178161 528297
rect 178215 528325 178267 528356
rect 178215 528291 178223 528325
rect 178257 528291 178267 528325
rect 178215 528246 178267 528291
rect 178845 528325 178897 528356
rect 178845 528291 178855 528325
rect 178889 528291 178897 528325
rect 178845 528246 178897 528291
rect 178951 528325 179003 528356
rect 178951 528291 178959 528325
rect 178993 528291 179003 528325
rect 178951 528226 179003 528291
rect 179033 528344 179112 528356
rect 179033 528310 179043 528344
rect 179077 528310 179112 528344
rect 179033 528272 179112 528310
rect 179142 528272 179208 528356
rect 179238 528329 179333 528356
rect 179238 528295 179250 528329
rect 179284 528295 179333 528329
rect 179238 528272 179333 528295
rect 179363 528272 179429 528356
rect 179459 528329 179597 528356
rect 179459 528295 179485 528329
rect 179519 528295 179553 528329
rect 179587 528295 179597 528329
rect 179459 528272 179597 528295
rect 179627 528329 179679 528356
rect 179627 528295 179637 528329
rect 179671 528295 179679 528329
rect 179627 528272 179679 528295
rect 179033 528226 179085 528272
rect 180055 528325 180107 528356
rect 180055 528291 180063 528325
rect 180097 528291 180107 528325
rect 180055 528246 180107 528291
rect 180685 528325 180737 528356
rect 180685 528291 180695 528325
rect 180729 528291 180737 528325
rect 180685 528246 180737 528291
rect 180975 528325 181027 528356
rect 180975 528291 180983 528325
rect 181017 528291 181027 528325
rect 180975 528226 181027 528291
rect 181057 528344 181136 528356
rect 181057 528310 181067 528344
rect 181101 528310 181136 528344
rect 181057 528272 181136 528310
rect 181166 528272 181232 528356
rect 181262 528329 181357 528356
rect 181262 528295 181274 528329
rect 181308 528295 181357 528329
rect 181262 528272 181357 528295
rect 181387 528272 181453 528356
rect 181483 528329 181621 528356
rect 181483 528295 181509 528329
rect 181543 528295 181577 528329
rect 181611 528295 181621 528329
rect 181483 528272 181621 528295
rect 181651 528329 181703 528356
rect 181651 528295 181661 528329
rect 181695 528295 181703 528329
rect 181651 528272 181703 528295
rect 181803 528325 181855 528356
rect 181803 528291 181811 528325
rect 181845 528291 181855 528325
rect 181057 528226 181109 528272
rect 181803 528246 181855 528291
rect 182801 528325 182853 528356
rect 182801 528291 182811 528325
rect 182845 528291 182853 528325
rect 182801 528246 182853 528291
rect 182907 528325 182959 528356
rect 182907 528291 182915 528325
rect 182949 528291 182959 528325
rect 182907 528246 182959 528291
rect 183905 528325 183957 528356
rect 183905 528291 183915 528325
rect 183949 528291 183957 528325
rect 183905 528246 183957 528291
rect 184011 528325 184063 528356
rect 184011 528291 184019 528325
rect 184053 528291 184063 528325
rect 184011 528246 184063 528291
rect 185009 528325 185061 528356
rect 185009 528291 185019 528325
rect 185053 528291 185061 528325
rect 185009 528246 185061 528291
rect 185207 528325 185259 528356
rect 185207 528291 185215 528325
rect 185249 528291 185259 528325
rect 185207 528246 185259 528291
rect 186205 528325 186257 528356
rect 186205 528291 186215 528325
rect 186249 528291 186257 528325
rect 186205 528246 186257 528291
rect 186311 528325 186363 528356
rect 186311 528291 186319 528325
rect 186353 528291 186363 528325
rect 186311 528246 186363 528291
rect 186941 528325 186993 528356
rect 186941 528291 186951 528325
rect 186985 528291 186993 528325
rect 186941 528246 186993 528291
rect 187231 528323 187283 528356
rect 187231 528289 187239 528323
rect 187273 528289 187283 528323
rect 187231 528246 187283 528289
rect 187401 528323 187453 528356
rect 187401 528289 187411 528323
rect 187445 528289 187453 528323
rect 187401 528246 187453 528289
rect 172235 527429 172287 527472
rect 172235 527395 172243 527429
rect 172277 527395 172287 527429
rect 172235 527362 172287 527395
rect 172405 527429 172457 527472
rect 172405 527395 172415 527429
rect 172449 527395 172457 527429
rect 172405 527362 172457 527395
rect 172511 527427 172563 527472
rect 172511 527393 172519 527427
rect 172553 527393 172563 527427
rect 172511 527362 172563 527393
rect 173509 527427 173561 527472
rect 173509 527393 173519 527427
rect 173553 527393 173561 527427
rect 173509 527362 173561 527393
rect 173615 527427 173667 527472
rect 173615 527393 173623 527427
rect 173657 527393 173667 527427
rect 173615 527362 173667 527393
rect 174613 527427 174665 527472
rect 174613 527393 174623 527427
rect 174657 527393 174665 527427
rect 174613 527362 174665 527393
rect 174719 527427 174771 527472
rect 174719 527393 174727 527427
rect 174761 527393 174771 527427
rect 174719 527362 174771 527393
rect 175717 527427 175769 527472
rect 175717 527393 175727 527427
rect 175761 527393 175769 527427
rect 175717 527362 175769 527393
rect 175823 527427 175875 527472
rect 175823 527393 175831 527427
rect 175865 527393 175875 527427
rect 175823 527362 175875 527393
rect 176269 527427 176321 527472
rect 176269 527393 176279 527427
rect 176313 527393 176321 527427
rect 176269 527362 176321 527393
rect 176394 527434 176446 527492
rect 176394 527400 176402 527434
rect 176436 527400 176446 527434
rect 176394 527362 176446 527400
rect 176476 527446 176526 527492
rect 176476 527408 176541 527446
rect 176476 527374 176492 527408
rect 176526 527374 176541 527408
rect 176476 527362 176541 527374
rect 176641 527434 176693 527446
rect 176641 527400 176651 527434
rect 176685 527400 176693 527434
rect 176641 527362 176693 527400
rect 176747 527434 176799 527446
rect 176747 527400 176755 527434
rect 176789 527400 176799 527434
rect 176747 527362 176799 527400
rect 176899 527408 176953 527446
rect 176899 527374 176909 527408
rect 176943 527374 176953 527408
rect 176899 527362 176953 527374
rect 176983 527434 177035 527446
rect 176983 527400 176993 527434
rect 177027 527400 177035 527434
rect 176983 527362 177035 527400
rect 177111 527429 177163 527472
rect 177111 527395 177119 527429
rect 177153 527395 177163 527429
rect 177111 527362 177163 527395
rect 177281 527429 177333 527472
rect 177281 527395 177291 527429
rect 177325 527395 177333 527429
rect 177281 527362 177333 527395
rect 177479 527427 177531 527472
rect 177479 527393 177487 527427
rect 177521 527393 177531 527427
rect 177479 527362 177531 527393
rect 178477 527427 178529 527472
rect 178477 527393 178487 527427
rect 178521 527393 178529 527427
rect 178477 527362 178529 527393
rect 178583 527434 178635 527472
rect 178583 527400 178591 527434
rect 178625 527400 178635 527434
rect 178583 527362 178635 527400
rect 178845 527434 178897 527472
rect 178845 527400 178855 527434
rect 178889 527400 178897 527434
rect 178845 527362 178897 527400
rect 178970 527434 179022 527492
rect 178970 527400 178978 527434
rect 179012 527400 179022 527434
rect 178970 527362 179022 527400
rect 179052 527446 179102 527492
rect 179052 527408 179117 527446
rect 179052 527374 179068 527408
rect 179102 527374 179117 527408
rect 179052 527362 179117 527374
rect 179217 527434 179269 527446
rect 179217 527400 179227 527434
rect 179261 527400 179269 527434
rect 179217 527362 179269 527400
rect 179323 527434 179375 527446
rect 179323 527400 179331 527434
rect 179365 527400 179375 527434
rect 179323 527362 179375 527400
rect 179475 527408 179529 527446
rect 179475 527374 179485 527408
rect 179519 527374 179529 527408
rect 179475 527362 179529 527374
rect 179559 527434 179611 527446
rect 179559 527400 179569 527434
rect 179603 527400 179611 527434
rect 179559 527362 179611 527400
rect 179687 527427 179739 527472
rect 179687 527393 179695 527427
rect 179729 527393 179739 527427
rect 179687 527362 179739 527393
rect 180685 527427 180737 527472
rect 180685 527393 180695 527427
rect 180729 527393 180737 527427
rect 180685 527362 180737 527393
rect 180791 527427 180843 527472
rect 180791 527393 180799 527427
rect 180833 527393 180843 527427
rect 180791 527362 180843 527393
rect 181789 527427 181841 527472
rect 181789 527393 181799 527427
rect 181833 527393 181841 527427
rect 181789 527362 181841 527393
rect 181895 527427 181947 527472
rect 181895 527393 181903 527427
rect 181937 527393 181947 527427
rect 181895 527362 181947 527393
rect 182341 527427 182393 527472
rect 182341 527393 182351 527427
rect 182385 527393 182393 527427
rect 182341 527362 182393 527393
rect 182631 527427 182683 527472
rect 182631 527393 182639 527427
rect 182673 527393 182683 527427
rect 182631 527362 182683 527393
rect 183629 527427 183681 527472
rect 183629 527393 183639 527427
rect 183673 527393 183681 527427
rect 183629 527362 183681 527393
rect 183735 527427 183787 527472
rect 183735 527393 183743 527427
rect 183777 527393 183787 527427
rect 183735 527362 183787 527393
rect 184733 527427 184785 527472
rect 184733 527393 184743 527427
rect 184777 527393 184785 527427
rect 184733 527362 184785 527393
rect 184839 527427 184891 527472
rect 184839 527393 184847 527427
rect 184881 527393 184891 527427
rect 184839 527362 184891 527393
rect 185837 527427 185889 527472
rect 185837 527393 185847 527427
rect 185881 527393 185889 527427
rect 185837 527362 185889 527393
rect 185943 527427 185995 527472
rect 185943 527393 185951 527427
rect 185985 527393 185995 527427
rect 185943 527362 185995 527393
rect 186941 527427 186993 527472
rect 186941 527393 186951 527427
rect 186985 527393 186993 527427
rect 186941 527362 186993 527393
rect 187231 527429 187283 527472
rect 187231 527395 187239 527429
rect 187273 527395 187283 527429
rect 187231 527362 187283 527395
rect 187401 527429 187453 527472
rect 187401 527395 187411 527429
rect 187445 527395 187453 527429
rect 187401 527362 187453 527395
rect 172235 527235 172287 527268
rect 172235 527201 172243 527235
rect 172277 527201 172287 527235
rect 172235 527158 172287 527201
rect 172405 527235 172457 527268
rect 172405 527201 172415 527235
rect 172449 527201 172457 527235
rect 172405 527158 172457 527201
rect 172511 527237 172563 527268
rect 172511 527203 172519 527237
rect 172553 527203 172563 527237
rect 172511 527158 172563 527203
rect 173509 527237 173561 527268
rect 173509 527203 173519 527237
rect 173553 527203 173561 527237
rect 173509 527158 173561 527203
rect 173615 527237 173667 527268
rect 173615 527203 173623 527237
rect 173657 527203 173667 527237
rect 173615 527158 173667 527203
rect 174613 527237 174665 527268
rect 174613 527203 174623 527237
rect 174657 527203 174665 527237
rect 174613 527158 174665 527203
rect 174903 527237 174955 527268
rect 174903 527203 174911 527237
rect 174945 527203 174955 527237
rect 174903 527158 174955 527203
rect 175901 527237 175953 527268
rect 175901 527203 175911 527237
rect 175945 527203 175953 527237
rect 175901 527158 175953 527203
rect 176007 527237 176059 527268
rect 176007 527203 176015 527237
rect 176049 527203 176059 527237
rect 176007 527158 176059 527203
rect 177005 527237 177057 527268
rect 177005 527203 177015 527237
rect 177049 527203 177057 527237
rect 177005 527158 177057 527203
rect 177111 527237 177163 527268
rect 177111 527203 177119 527237
rect 177153 527203 177163 527237
rect 177111 527158 177163 527203
rect 178109 527237 178161 527268
rect 178109 527203 178119 527237
rect 178153 527203 178161 527237
rect 178109 527158 178161 527203
rect 178215 527237 178267 527268
rect 178215 527203 178223 527237
rect 178257 527203 178267 527237
rect 178215 527158 178267 527203
rect 179213 527237 179265 527268
rect 179213 527203 179223 527237
rect 179257 527203 179265 527237
rect 179213 527158 179265 527203
rect 179319 527237 179371 527268
rect 179319 527203 179327 527237
rect 179361 527203 179371 527237
rect 179319 527158 179371 527203
rect 179765 527237 179817 527268
rect 179765 527203 179775 527237
rect 179809 527203 179817 527237
rect 179765 527158 179817 527203
rect 180055 527237 180107 527268
rect 180055 527203 180063 527237
rect 180097 527203 180107 527237
rect 180055 527158 180107 527203
rect 181053 527237 181105 527268
rect 181053 527203 181063 527237
rect 181097 527203 181105 527237
rect 181053 527158 181105 527203
rect 181159 527237 181211 527268
rect 181159 527203 181167 527237
rect 181201 527203 181211 527237
rect 181159 527158 181211 527203
rect 182157 527237 182209 527268
rect 182157 527203 182167 527237
rect 182201 527203 182209 527237
rect 182157 527158 182209 527203
rect 182263 527237 182315 527268
rect 182263 527203 182271 527237
rect 182305 527203 182315 527237
rect 182263 527158 182315 527203
rect 183261 527237 183313 527268
rect 183261 527203 183271 527237
rect 183305 527203 183313 527237
rect 183261 527158 183313 527203
rect 183367 527237 183419 527268
rect 183367 527203 183375 527237
rect 183409 527203 183419 527237
rect 183367 527158 183419 527203
rect 184365 527237 184417 527268
rect 184365 527203 184375 527237
rect 184409 527203 184417 527237
rect 184365 527158 184417 527203
rect 184471 527237 184523 527268
rect 184471 527203 184479 527237
rect 184513 527203 184523 527237
rect 184471 527158 184523 527203
rect 184917 527237 184969 527268
rect 184917 527203 184927 527237
rect 184961 527203 184969 527237
rect 184917 527158 184969 527203
rect 185207 527237 185259 527268
rect 185207 527203 185215 527237
rect 185249 527203 185259 527237
rect 185207 527158 185259 527203
rect 186205 527237 186257 527268
rect 186205 527203 186215 527237
rect 186249 527203 186257 527237
rect 186205 527158 186257 527203
rect 186311 527237 186363 527268
rect 186311 527203 186319 527237
rect 186353 527203 186363 527237
rect 186311 527158 186363 527203
rect 186941 527237 186993 527268
rect 186941 527203 186951 527237
rect 186985 527203 186993 527237
rect 186941 527158 186993 527203
rect 187231 527235 187283 527268
rect 187231 527201 187239 527235
rect 187273 527201 187283 527235
rect 187231 527158 187283 527201
rect 187401 527235 187453 527268
rect 187401 527201 187411 527235
rect 187445 527201 187453 527235
rect 187401 527158 187453 527201
rect 172235 526341 172287 526384
rect 172235 526307 172243 526341
rect 172277 526307 172287 526341
rect 172235 526274 172287 526307
rect 172405 526341 172457 526384
rect 172405 526307 172415 526341
rect 172449 526307 172457 526341
rect 172405 526274 172457 526307
rect 172511 526339 172563 526384
rect 172511 526305 172519 526339
rect 172553 526305 172563 526339
rect 172511 526274 172563 526305
rect 173509 526339 173561 526384
rect 173509 526305 173519 526339
rect 173553 526305 173561 526339
rect 173509 526274 173561 526305
rect 173615 526339 173667 526384
rect 173615 526305 173623 526339
rect 173657 526305 173667 526339
rect 173615 526274 173667 526305
rect 174613 526339 174665 526384
rect 174613 526305 174623 526339
rect 174657 526305 174665 526339
rect 174613 526274 174665 526305
rect 174719 526339 174771 526384
rect 174719 526305 174727 526339
rect 174761 526305 174771 526339
rect 174719 526274 174771 526305
rect 175717 526339 175769 526384
rect 175717 526305 175727 526339
rect 175761 526305 175769 526339
rect 175717 526274 175769 526305
rect 175823 526339 175875 526384
rect 175823 526305 175831 526339
rect 175865 526305 175875 526339
rect 175823 526274 175875 526305
rect 176821 526339 176873 526384
rect 176821 526305 176831 526339
rect 176865 526305 176873 526339
rect 176821 526274 176873 526305
rect 176927 526346 176979 526384
rect 176927 526312 176935 526346
rect 176969 526312 176979 526346
rect 176927 526274 176979 526312
rect 177189 526346 177241 526384
rect 177189 526312 177199 526346
rect 177233 526312 177241 526346
rect 177189 526274 177241 526312
rect 177479 526339 177531 526384
rect 177479 526305 177487 526339
rect 177521 526305 177531 526339
rect 177479 526274 177531 526305
rect 178477 526339 178529 526384
rect 178477 526305 178487 526339
rect 178521 526305 178529 526339
rect 178477 526274 178529 526305
rect 178583 526339 178635 526384
rect 178583 526305 178591 526339
rect 178625 526305 178635 526339
rect 178583 526274 178635 526305
rect 179581 526339 179633 526384
rect 179581 526305 179591 526339
rect 179625 526305 179633 526339
rect 179581 526274 179633 526305
rect 179687 526339 179739 526384
rect 179687 526305 179695 526339
rect 179729 526305 179739 526339
rect 179687 526274 179739 526305
rect 180685 526339 180737 526384
rect 180685 526305 180695 526339
rect 180729 526305 180737 526339
rect 180685 526274 180737 526305
rect 180791 526339 180843 526384
rect 180791 526305 180799 526339
rect 180833 526305 180843 526339
rect 180791 526274 180843 526305
rect 181789 526339 181841 526384
rect 181789 526305 181799 526339
rect 181833 526305 181841 526339
rect 181789 526274 181841 526305
rect 181895 526339 181947 526384
rect 181895 526305 181903 526339
rect 181937 526305 181947 526339
rect 181895 526274 181947 526305
rect 182341 526339 182393 526384
rect 182341 526305 182351 526339
rect 182385 526305 182393 526339
rect 182341 526274 182393 526305
rect 182631 526339 182683 526384
rect 182631 526305 182639 526339
rect 182673 526305 182683 526339
rect 182631 526274 182683 526305
rect 183629 526339 183681 526384
rect 183629 526305 183639 526339
rect 183673 526305 183681 526339
rect 183629 526274 183681 526305
rect 183735 526339 183787 526384
rect 183735 526305 183743 526339
rect 183777 526305 183787 526339
rect 183735 526274 183787 526305
rect 184733 526339 184785 526384
rect 184733 526305 184743 526339
rect 184777 526305 184785 526339
rect 184733 526274 184785 526305
rect 184839 526339 184891 526384
rect 184839 526305 184847 526339
rect 184881 526305 184891 526339
rect 184839 526274 184891 526305
rect 185837 526339 185889 526384
rect 185837 526305 185847 526339
rect 185881 526305 185889 526339
rect 185837 526274 185889 526305
rect 185943 526339 185995 526384
rect 185943 526305 185951 526339
rect 185985 526305 185995 526339
rect 185943 526274 185995 526305
rect 186941 526339 186993 526384
rect 186941 526305 186951 526339
rect 186985 526305 186993 526339
rect 186941 526274 186993 526305
rect 187231 526341 187283 526384
rect 187231 526307 187239 526341
rect 187273 526307 187283 526341
rect 187231 526274 187283 526307
rect 187401 526341 187453 526384
rect 187401 526307 187411 526341
rect 187445 526307 187453 526341
rect 187401 526274 187453 526307
rect 172235 526147 172287 526180
rect 172235 526113 172243 526147
rect 172277 526113 172287 526147
rect 172235 526070 172287 526113
rect 172405 526147 172457 526180
rect 172405 526113 172415 526147
rect 172449 526113 172457 526147
rect 172405 526070 172457 526113
rect 172511 526149 172563 526180
rect 172511 526115 172519 526149
rect 172553 526115 172563 526149
rect 172511 526070 172563 526115
rect 173509 526149 173561 526180
rect 173509 526115 173519 526149
rect 173553 526115 173561 526149
rect 173509 526070 173561 526115
rect 173615 526149 173667 526180
rect 173615 526115 173623 526149
rect 173657 526115 173667 526149
rect 173615 526070 173667 526115
rect 174613 526149 174665 526180
rect 174613 526115 174623 526149
rect 174657 526115 174665 526149
rect 174613 526070 174665 526115
rect 174903 526149 174955 526180
rect 174903 526115 174911 526149
rect 174945 526115 174955 526149
rect 174903 526070 174955 526115
rect 175901 526149 175953 526180
rect 175901 526115 175911 526149
rect 175945 526115 175953 526149
rect 175901 526070 175953 526115
rect 176007 526149 176059 526180
rect 176007 526115 176015 526149
rect 176049 526115 176059 526149
rect 176007 526070 176059 526115
rect 177005 526149 177057 526180
rect 177005 526115 177015 526149
rect 177049 526115 177057 526149
rect 177005 526070 177057 526115
rect 177111 526149 177163 526180
rect 177111 526115 177119 526149
rect 177153 526115 177163 526149
rect 177111 526070 177163 526115
rect 178109 526149 178161 526180
rect 178109 526115 178119 526149
rect 178153 526115 178161 526149
rect 178109 526070 178161 526115
rect 178215 526149 178267 526180
rect 178215 526115 178223 526149
rect 178257 526115 178267 526149
rect 178215 526070 178267 526115
rect 179213 526149 179265 526180
rect 179213 526115 179223 526149
rect 179257 526115 179265 526149
rect 179213 526070 179265 526115
rect 179319 526149 179371 526180
rect 179319 526115 179327 526149
rect 179361 526115 179371 526149
rect 179319 526070 179371 526115
rect 179765 526149 179817 526180
rect 179765 526115 179775 526149
rect 179809 526115 179817 526149
rect 179765 526070 179817 526115
rect 180055 526149 180107 526180
rect 180055 526115 180063 526149
rect 180097 526115 180107 526149
rect 180055 526070 180107 526115
rect 181053 526149 181105 526180
rect 181053 526115 181063 526149
rect 181097 526115 181105 526149
rect 181053 526070 181105 526115
rect 181159 526149 181211 526180
rect 181159 526115 181167 526149
rect 181201 526115 181211 526149
rect 181159 526070 181211 526115
rect 182157 526149 182209 526180
rect 182157 526115 182167 526149
rect 182201 526115 182209 526149
rect 182157 526070 182209 526115
rect 182263 526149 182315 526180
rect 182263 526115 182271 526149
rect 182305 526115 182315 526149
rect 182263 526070 182315 526115
rect 183261 526149 183313 526180
rect 183261 526115 183271 526149
rect 183305 526115 183313 526149
rect 183261 526070 183313 526115
rect 183367 526149 183419 526180
rect 183367 526115 183375 526149
rect 183409 526115 183419 526149
rect 183367 526070 183419 526115
rect 184365 526149 184417 526180
rect 184365 526115 184375 526149
rect 184409 526115 184417 526149
rect 184365 526070 184417 526115
rect 184471 526149 184523 526180
rect 184471 526115 184479 526149
rect 184513 526115 184523 526149
rect 184471 526070 184523 526115
rect 184917 526149 184969 526180
rect 184917 526115 184927 526149
rect 184961 526115 184969 526149
rect 184917 526070 184969 526115
rect 185207 526149 185259 526180
rect 185207 526115 185215 526149
rect 185249 526115 185259 526149
rect 185207 526070 185259 526115
rect 186205 526149 186257 526180
rect 186205 526115 186215 526149
rect 186249 526115 186257 526149
rect 186205 526070 186257 526115
rect 186311 526149 186363 526180
rect 186311 526115 186319 526149
rect 186353 526115 186363 526149
rect 186311 526070 186363 526115
rect 186941 526149 186993 526180
rect 186941 526115 186951 526149
rect 186985 526115 186993 526149
rect 186941 526070 186993 526115
rect 187231 526147 187283 526180
rect 187231 526113 187239 526147
rect 187273 526113 187283 526147
rect 187231 526070 187283 526113
rect 187401 526147 187453 526180
rect 187401 526113 187411 526147
rect 187445 526113 187453 526147
rect 187401 526070 187453 526113
rect 172235 525253 172287 525296
rect 172235 525219 172243 525253
rect 172277 525219 172287 525253
rect 172235 525186 172287 525219
rect 172405 525253 172457 525296
rect 172405 525219 172415 525253
rect 172449 525219 172457 525253
rect 172405 525186 172457 525219
rect 172511 525251 172563 525296
rect 172511 525217 172519 525251
rect 172553 525217 172563 525251
rect 172511 525186 172563 525217
rect 173509 525251 173561 525296
rect 173509 525217 173519 525251
rect 173553 525217 173561 525251
rect 173509 525186 173561 525217
rect 173615 525251 173667 525296
rect 173615 525217 173623 525251
rect 173657 525217 173667 525251
rect 173615 525186 173667 525217
rect 174613 525251 174665 525296
rect 174613 525217 174623 525251
rect 174657 525217 174665 525251
rect 174613 525186 174665 525217
rect 174719 525251 174771 525296
rect 174719 525217 174727 525251
rect 174761 525217 174771 525251
rect 174719 525186 174771 525217
rect 175717 525251 175769 525296
rect 175717 525217 175727 525251
rect 175761 525217 175769 525251
rect 175717 525186 175769 525217
rect 175823 525251 175875 525296
rect 175823 525217 175831 525251
rect 175865 525217 175875 525251
rect 175823 525186 175875 525217
rect 176821 525251 176873 525296
rect 176821 525217 176831 525251
rect 176865 525217 176873 525251
rect 176821 525186 176873 525217
rect 176927 525258 176979 525296
rect 176927 525224 176935 525258
rect 176969 525224 176979 525258
rect 176927 525186 176979 525224
rect 177189 525258 177241 525296
rect 177189 525224 177199 525258
rect 177233 525224 177241 525258
rect 177189 525186 177241 525224
rect 177479 525251 177531 525296
rect 177479 525217 177487 525251
rect 177521 525217 177531 525251
rect 177479 525186 177531 525217
rect 178477 525251 178529 525296
rect 178477 525217 178487 525251
rect 178521 525217 178529 525251
rect 178477 525186 178529 525217
rect 178583 525251 178635 525296
rect 178583 525217 178591 525251
rect 178625 525217 178635 525251
rect 178583 525186 178635 525217
rect 179581 525251 179633 525296
rect 179581 525217 179591 525251
rect 179625 525217 179633 525251
rect 179581 525186 179633 525217
rect 179687 525251 179739 525296
rect 179687 525217 179695 525251
rect 179729 525217 179739 525251
rect 179687 525186 179739 525217
rect 180685 525251 180737 525296
rect 180685 525217 180695 525251
rect 180729 525217 180737 525251
rect 180685 525186 180737 525217
rect 180791 525251 180843 525296
rect 180791 525217 180799 525251
rect 180833 525217 180843 525251
rect 180791 525186 180843 525217
rect 181789 525251 181841 525296
rect 181789 525217 181799 525251
rect 181833 525217 181841 525251
rect 181789 525186 181841 525217
rect 181895 525251 181947 525296
rect 181895 525217 181903 525251
rect 181937 525217 181947 525251
rect 181895 525186 181947 525217
rect 182341 525251 182393 525296
rect 182341 525217 182351 525251
rect 182385 525217 182393 525251
rect 182341 525186 182393 525217
rect 182631 525251 182683 525296
rect 182631 525217 182639 525251
rect 182673 525217 182683 525251
rect 182631 525186 182683 525217
rect 183629 525251 183681 525296
rect 183629 525217 183639 525251
rect 183673 525217 183681 525251
rect 183629 525186 183681 525217
rect 183735 525251 183787 525296
rect 183735 525217 183743 525251
rect 183777 525217 183787 525251
rect 183735 525186 183787 525217
rect 184733 525251 184785 525296
rect 184733 525217 184743 525251
rect 184777 525217 184785 525251
rect 184733 525186 184785 525217
rect 184839 525251 184891 525296
rect 184839 525217 184847 525251
rect 184881 525217 184891 525251
rect 184839 525186 184891 525217
rect 185837 525251 185889 525296
rect 185837 525217 185847 525251
rect 185881 525217 185889 525251
rect 185837 525186 185889 525217
rect 185943 525251 185995 525296
rect 185943 525217 185951 525251
rect 185985 525217 185995 525251
rect 185943 525186 185995 525217
rect 186941 525251 186993 525296
rect 186941 525217 186951 525251
rect 186985 525217 186993 525251
rect 186941 525186 186993 525217
rect 187231 525253 187283 525296
rect 187231 525219 187239 525253
rect 187273 525219 187283 525253
rect 187231 525186 187283 525219
rect 187401 525253 187453 525296
rect 187401 525219 187411 525253
rect 187445 525219 187453 525253
rect 187401 525186 187453 525219
rect 172235 525059 172287 525092
rect 172235 525025 172243 525059
rect 172277 525025 172287 525059
rect 172235 524982 172287 525025
rect 172405 525059 172457 525092
rect 172405 525025 172415 525059
rect 172449 525025 172457 525059
rect 172405 524982 172457 525025
rect 172511 525061 172563 525092
rect 172511 525027 172519 525061
rect 172553 525027 172563 525061
rect 172511 524982 172563 525027
rect 173509 525061 173561 525092
rect 173509 525027 173519 525061
rect 173553 525027 173561 525061
rect 173509 524982 173561 525027
rect 173615 525061 173667 525092
rect 173615 525027 173623 525061
rect 173657 525027 173667 525061
rect 173615 524982 173667 525027
rect 174613 525061 174665 525092
rect 174613 525027 174623 525061
rect 174657 525027 174665 525061
rect 174613 524982 174665 525027
rect 174903 525061 174955 525092
rect 174903 525027 174911 525061
rect 174945 525027 174955 525061
rect 174903 524982 174955 525027
rect 175901 525061 175953 525092
rect 175901 525027 175911 525061
rect 175945 525027 175953 525061
rect 175901 524982 175953 525027
rect 176007 525061 176059 525092
rect 176007 525027 176015 525061
rect 176049 525027 176059 525061
rect 176007 524982 176059 525027
rect 177005 525061 177057 525092
rect 177005 525027 177015 525061
rect 177049 525027 177057 525061
rect 177005 524982 177057 525027
rect 177111 525061 177163 525092
rect 177111 525027 177119 525061
rect 177153 525027 177163 525061
rect 177111 524982 177163 525027
rect 178109 525061 178161 525092
rect 178109 525027 178119 525061
rect 178153 525027 178161 525061
rect 178109 524982 178161 525027
rect 178215 525061 178267 525092
rect 178215 525027 178223 525061
rect 178257 525027 178267 525061
rect 178215 524982 178267 525027
rect 179213 525061 179265 525092
rect 179213 525027 179223 525061
rect 179257 525027 179265 525061
rect 179213 524982 179265 525027
rect 179319 525061 179371 525092
rect 179319 525027 179327 525061
rect 179361 525027 179371 525061
rect 179319 524982 179371 525027
rect 179765 525061 179817 525092
rect 179765 525027 179775 525061
rect 179809 525027 179817 525061
rect 179765 524982 179817 525027
rect 180055 525061 180107 525092
rect 180055 525027 180063 525061
rect 180097 525027 180107 525061
rect 180055 524982 180107 525027
rect 181053 525061 181105 525092
rect 181053 525027 181063 525061
rect 181097 525027 181105 525061
rect 181053 524982 181105 525027
rect 181159 525061 181211 525092
rect 181159 525027 181167 525061
rect 181201 525027 181211 525061
rect 181159 524982 181211 525027
rect 182157 525061 182209 525092
rect 182157 525027 182167 525061
rect 182201 525027 182209 525061
rect 182157 524982 182209 525027
rect 182263 525061 182315 525092
rect 182263 525027 182271 525061
rect 182305 525027 182315 525061
rect 182263 524982 182315 525027
rect 183261 525061 183313 525092
rect 183261 525027 183271 525061
rect 183305 525027 183313 525061
rect 183261 524982 183313 525027
rect 183367 525061 183419 525092
rect 183367 525027 183375 525061
rect 183409 525027 183419 525061
rect 183367 524982 183419 525027
rect 184365 525061 184417 525092
rect 184365 525027 184375 525061
rect 184409 525027 184417 525061
rect 184365 524982 184417 525027
rect 184471 525061 184523 525092
rect 184471 525027 184479 525061
rect 184513 525027 184523 525061
rect 184471 524982 184523 525027
rect 184917 525061 184969 525092
rect 184917 525027 184927 525061
rect 184961 525027 184969 525061
rect 184917 524982 184969 525027
rect 185207 525061 185259 525092
rect 185207 525027 185215 525061
rect 185249 525027 185259 525061
rect 185207 524982 185259 525027
rect 186205 525061 186257 525092
rect 186205 525027 186215 525061
rect 186249 525027 186257 525061
rect 186205 524982 186257 525027
rect 186311 525061 186363 525092
rect 186311 525027 186319 525061
rect 186353 525027 186363 525061
rect 186311 524982 186363 525027
rect 186941 525061 186993 525092
rect 186941 525027 186951 525061
rect 186985 525027 186993 525061
rect 186941 524982 186993 525027
rect 187231 525059 187283 525092
rect 187231 525025 187239 525059
rect 187273 525025 187283 525059
rect 187231 524982 187283 525025
rect 187401 525059 187453 525092
rect 187401 525025 187411 525059
rect 187445 525025 187453 525059
rect 187401 524982 187453 525025
rect 172235 524165 172287 524208
rect 172235 524131 172243 524165
rect 172277 524131 172287 524165
rect 172235 524098 172287 524131
rect 172405 524165 172457 524208
rect 172405 524131 172415 524165
rect 172449 524131 172457 524165
rect 172405 524098 172457 524131
rect 172511 524163 172563 524208
rect 172511 524129 172519 524163
rect 172553 524129 172563 524163
rect 172511 524098 172563 524129
rect 173509 524163 173561 524208
rect 173509 524129 173519 524163
rect 173553 524129 173561 524163
rect 173509 524098 173561 524129
rect 173615 524163 173667 524208
rect 173615 524129 173623 524163
rect 173657 524129 173667 524163
rect 173615 524098 173667 524129
rect 174613 524163 174665 524208
rect 174613 524129 174623 524163
rect 174657 524129 174665 524163
rect 174613 524098 174665 524129
rect 174719 524163 174771 524208
rect 174719 524129 174727 524163
rect 174761 524129 174771 524163
rect 174719 524098 174771 524129
rect 175717 524163 175769 524208
rect 175717 524129 175727 524163
rect 175761 524129 175769 524163
rect 175717 524098 175769 524129
rect 175823 524163 175875 524208
rect 175823 524129 175831 524163
rect 175865 524129 175875 524163
rect 175823 524098 175875 524129
rect 176821 524163 176873 524208
rect 176821 524129 176831 524163
rect 176865 524129 176873 524163
rect 176821 524098 176873 524129
rect 176927 524170 176979 524208
rect 176927 524136 176935 524170
rect 176969 524136 176979 524170
rect 176927 524098 176979 524136
rect 177189 524170 177241 524208
rect 177189 524136 177199 524170
rect 177233 524136 177241 524170
rect 177189 524098 177241 524136
rect 177479 524163 177531 524208
rect 177479 524129 177487 524163
rect 177521 524129 177531 524163
rect 177479 524098 177531 524129
rect 178477 524163 178529 524208
rect 178477 524129 178487 524163
rect 178521 524129 178529 524163
rect 178477 524098 178529 524129
rect 178583 524163 178635 524208
rect 178583 524129 178591 524163
rect 178625 524129 178635 524163
rect 178583 524098 178635 524129
rect 179581 524163 179633 524208
rect 179581 524129 179591 524163
rect 179625 524129 179633 524163
rect 179581 524098 179633 524129
rect 179687 524163 179739 524208
rect 179687 524129 179695 524163
rect 179729 524129 179739 524163
rect 179687 524098 179739 524129
rect 180685 524163 180737 524208
rect 180685 524129 180695 524163
rect 180729 524129 180737 524163
rect 180685 524098 180737 524129
rect 180791 524163 180843 524208
rect 180791 524129 180799 524163
rect 180833 524129 180843 524163
rect 180791 524098 180843 524129
rect 181789 524163 181841 524208
rect 181789 524129 181799 524163
rect 181833 524129 181841 524163
rect 181789 524098 181841 524129
rect 181895 524163 181947 524208
rect 181895 524129 181903 524163
rect 181937 524129 181947 524163
rect 181895 524098 181947 524129
rect 182341 524163 182393 524208
rect 182341 524129 182351 524163
rect 182385 524129 182393 524163
rect 182341 524098 182393 524129
rect 182631 524163 182683 524208
rect 182631 524129 182639 524163
rect 182673 524129 182683 524163
rect 182631 524098 182683 524129
rect 183629 524163 183681 524208
rect 183629 524129 183639 524163
rect 183673 524129 183681 524163
rect 183629 524098 183681 524129
rect 183735 524163 183787 524208
rect 183735 524129 183743 524163
rect 183777 524129 183787 524163
rect 183735 524098 183787 524129
rect 184733 524163 184785 524208
rect 184733 524129 184743 524163
rect 184777 524129 184785 524163
rect 184733 524098 184785 524129
rect 184839 524163 184891 524208
rect 184839 524129 184847 524163
rect 184881 524129 184891 524163
rect 184839 524098 184891 524129
rect 185837 524163 185889 524208
rect 185837 524129 185847 524163
rect 185881 524129 185889 524163
rect 185837 524098 185889 524129
rect 185943 524163 185995 524208
rect 185943 524129 185951 524163
rect 185985 524129 185995 524163
rect 185943 524098 185995 524129
rect 186941 524163 186993 524208
rect 186941 524129 186951 524163
rect 186985 524129 186993 524163
rect 186941 524098 186993 524129
rect 187231 524165 187283 524208
rect 187231 524131 187239 524165
rect 187273 524131 187283 524165
rect 187231 524098 187283 524131
rect 187401 524165 187453 524208
rect 187401 524131 187411 524165
rect 187445 524131 187453 524165
rect 187401 524098 187453 524131
rect 172235 523971 172287 524004
rect 172235 523937 172243 523971
rect 172277 523937 172287 523971
rect 172235 523894 172287 523937
rect 172405 523971 172457 524004
rect 172405 523937 172415 523971
rect 172449 523937 172457 523971
rect 172405 523894 172457 523937
rect 172511 523973 172563 524004
rect 172511 523939 172519 523973
rect 172553 523939 172563 523973
rect 172511 523894 172563 523939
rect 173509 523973 173561 524004
rect 173509 523939 173519 523973
rect 173553 523939 173561 523973
rect 173509 523894 173561 523939
rect 173615 523973 173667 524004
rect 173615 523939 173623 523973
rect 173657 523939 173667 523973
rect 173615 523894 173667 523939
rect 174613 523973 174665 524004
rect 174613 523939 174623 523973
rect 174657 523939 174665 523973
rect 174613 523894 174665 523939
rect 174903 523973 174955 524004
rect 174903 523939 174911 523973
rect 174945 523939 174955 523973
rect 174903 523894 174955 523939
rect 175901 523973 175953 524004
rect 175901 523939 175911 523973
rect 175945 523939 175953 523973
rect 175901 523894 175953 523939
rect 176007 523973 176059 524004
rect 176007 523939 176015 523973
rect 176049 523939 176059 523973
rect 176007 523894 176059 523939
rect 177005 523973 177057 524004
rect 177005 523939 177015 523973
rect 177049 523939 177057 523973
rect 177005 523894 177057 523939
rect 177111 523973 177163 524004
rect 177111 523939 177119 523973
rect 177153 523939 177163 523973
rect 177111 523894 177163 523939
rect 178109 523973 178161 524004
rect 178109 523939 178119 523973
rect 178153 523939 178161 523973
rect 178109 523894 178161 523939
rect 178215 523973 178267 524004
rect 178215 523939 178223 523973
rect 178257 523939 178267 523973
rect 178215 523894 178267 523939
rect 179213 523973 179265 524004
rect 179213 523939 179223 523973
rect 179257 523939 179265 523973
rect 179213 523894 179265 523939
rect 179319 523973 179371 524004
rect 179319 523939 179327 523973
rect 179361 523939 179371 523973
rect 179319 523894 179371 523939
rect 179765 523973 179817 524004
rect 179765 523939 179775 523973
rect 179809 523939 179817 523973
rect 179765 523894 179817 523939
rect 180055 523973 180107 524004
rect 180055 523939 180063 523973
rect 180097 523939 180107 523973
rect 180055 523894 180107 523939
rect 181053 523973 181105 524004
rect 181053 523939 181063 523973
rect 181097 523939 181105 523973
rect 181053 523894 181105 523939
rect 181159 523973 181211 524004
rect 181159 523939 181167 523973
rect 181201 523939 181211 523973
rect 181159 523894 181211 523939
rect 182157 523973 182209 524004
rect 182157 523939 182167 523973
rect 182201 523939 182209 523973
rect 182157 523894 182209 523939
rect 182263 523973 182315 524004
rect 182263 523939 182271 523973
rect 182305 523939 182315 523973
rect 182263 523894 182315 523939
rect 183261 523973 183313 524004
rect 183261 523939 183271 523973
rect 183305 523939 183313 523973
rect 183261 523894 183313 523939
rect 183367 523973 183419 524004
rect 183367 523939 183375 523973
rect 183409 523939 183419 523973
rect 183367 523894 183419 523939
rect 184365 523973 184417 524004
rect 184365 523939 184375 523973
rect 184409 523939 184417 523973
rect 184365 523894 184417 523939
rect 184471 523973 184523 524004
rect 184471 523939 184479 523973
rect 184513 523939 184523 523973
rect 184471 523894 184523 523939
rect 184917 523973 184969 524004
rect 184917 523939 184927 523973
rect 184961 523939 184969 523973
rect 184917 523894 184969 523939
rect 185207 523973 185259 524004
rect 185207 523939 185215 523973
rect 185249 523939 185259 523973
rect 185207 523894 185259 523939
rect 186205 523973 186257 524004
rect 186205 523939 186215 523973
rect 186249 523939 186257 523973
rect 186205 523894 186257 523939
rect 186311 523973 186363 524004
rect 186311 523939 186319 523973
rect 186353 523939 186363 523973
rect 186311 523894 186363 523939
rect 186941 523973 186993 524004
rect 186941 523939 186951 523973
rect 186985 523939 186993 523973
rect 186941 523894 186993 523939
rect 187231 523971 187283 524004
rect 187231 523937 187239 523971
rect 187273 523937 187283 523971
rect 187231 523894 187283 523937
rect 187401 523971 187453 524004
rect 187401 523937 187411 523971
rect 187445 523937 187453 523971
rect 187401 523894 187453 523937
rect 172235 523077 172287 523120
rect 172235 523043 172243 523077
rect 172277 523043 172287 523077
rect 172235 523010 172287 523043
rect 172405 523077 172457 523120
rect 172405 523043 172415 523077
rect 172449 523043 172457 523077
rect 172405 523010 172457 523043
rect 172511 523075 172563 523120
rect 172511 523041 172519 523075
rect 172553 523041 172563 523075
rect 172511 523010 172563 523041
rect 173509 523075 173561 523120
rect 173509 523041 173519 523075
rect 173553 523041 173561 523075
rect 173509 523010 173561 523041
rect 173615 523075 173667 523120
rect 173615 523041 173623 523075
rect 173657 523041 173667 523075
rect 173615 523010 173667 523041
rect 174613 523075 174665 523120
rect 174613 523041 174623 523075
rect 174657 523041 174665 523075
rect 174613 523010 174665 523041
rect 174719 523075 174771 523120
rect 174719 523041 174727 523075
rect 174761 523041 174771 523075
rect 174719 523010 174771 523041
rect 175717 523075 175769 523120
rect 175717 523041 175727 523075
rect 175761 523041 175769 523075
rect 175717 523010 175769 523041
rect 175823 523075 175875 523120
rect 175823 523041 175831 523075
rect 175865 523041 175875 523075
rect 175823 523010 175875 523041
rect 176821 523075 176873 523120
rect 176821 523041 176831 523075
rect 176865 523041 176873 523075
rect 176821 523010 176873 523041
rect 176927 523082 176979 523120
rect 176927 523048 176935 523082
rect 176969 523048 176979 523082
rect 176927 523010 176979 523048
rect 177189 523082 177241 523120
rect 177189 523048 177199 523082
rect 177233 523048 177241 523082
rect 177189 523010 177241 523048
rect 177479 523075 177531 523120
rect 177479 523041 177487 523075
rect 177521 523041 177531 523075
rect 177479 523010 177531 523041
rect 178477 523075 178529 523120
rect 178477 523041 178487 523075
rect 178521 523041 178529 523075
rect 178477 523010 178529 523041
rect 178583 523075 178635 523120
rect 178583 523041 178591 523075
rect 178625 523041 178635 523075
rect 178583 523010 178635 523041
rect 179581 523075 179633 523120
rect 179581 523041 179591 523075
rect 179625 523041 179633 523075
rect 179581 523010 179633 523041
rect 179687 523075 179739 523120
rect 179687 523041 179695 523075
rect 179729 523041 179739 523075
rect 179687 523010 179739 523041
rect 180685 523075 180737 523120
rect 180685 523041 180695 523075
rect 180729 523041 180737 523075
rect 180685 523010 180737 523041
rect 180791 523075 180843 523120
rect 180791 523041 180799 523075
rect 180833 523041 180843 523075
rect 180791 523010 180843 523041
rect 181789 523075 181841 523120
rect 181789 523041 181799 523075
rect 181833 523041 181841 523075
rect 181789 523010 181841 523041
rect 181895 523075 181947 523120
rect 181895 523041 181903 523075
rect 181937 523041 181947 523075
rect 181895 523010 181947 523041
rect 182341 523075 182393 523120
rect 182341 523041 182351 523075
rect 182385 523041 182393 523075
rect 182341 523010 182393 523041
rect 182631 523075 182683 523120
rect 182631 523041 182639 523075
rect 182673 523041 182683 523075
rect 182631 523010 182683 523041
rect 183629 523075 183681 523120
rect 183629 523041 183639 523075
rect 183673 523041 183681 523075
rect 183629 523010 183681 523041
rect 183735 523075 183787 523120
rect 183735 523041 183743 523075
rect 183777 523041 183787 523075
rect 183735 523010 183787 523041
rect 184733 523075 184785 523120
rect 184733 523041 184743 523075
rect 184777 523041 184785 523075
rect 184733 523010 184785 523041
rect 184839 523075 184891 523120
rect 184839 523041 184847 523075
rect 184881 523041 184891 523075
rect 184839 523010 184891 523041
rect 185837 523075 185889 523120
rect 185837 523041 185847 523075
rect 185881 523041 185889 523075
rect 185837 523010 185889 523041
rect 185943 523075 185995 523120
rect 185943 523041 185951 523075
rect 185985 523041 185995 523075
rect 185943 523010 185995 523041
rect 186941 523075 186993 523120
rect 186941 523041 186951 523075
rect 186985 523041 186993 523075
rect 186941 523010 186993 523041
rect 187231 523077 187283 523120
rect 187231 523043 187239 523077
rect 187273 523043 187283 523077
rect 187231 523010 187283 523043
rect 187401 523077 187453 523120
rect 187401 523043 187411 523077
rect 187445 523043 187453 523077
rect 187401 523010 187453 523043
rect 172235 522883 172287 522916
rect 172235 522849 172243 522883
rect 172277 522849 172287 522883
rect 172235 522806 172287 522849
rect 172405 522883 172457 522916
rect 172405 522849 172415 522883
rect 172449 522849 172457 522883
rect 172405 522806 172457 522849
rect 172511 522885 172563 522916
rect 172511 522851 172519 522885
rect 172553 522851 172563 522885
rect 172511 522806 172563 522851
rect 173509 522885 173561 522916
rect 173509 522851 173519 522885
rect 173553 522851 173561 522885
rect 173509 522806 173561 522851
rect 173615 522885 173667 522916
rect 173615 522851 173623 522885
rect 173657 522851 173667 522885
rect 173615 522806 173667 522851
rect 174613 522885 174665 522916
rect 174613 522851 174623 522885
rect 174657 522851 174665 522885
rect 174613 522806 174665 522851
rect 174903 522885 174955 522916
rect 174903 522851 174911 522885
rect 174945 522851 174955 522885
rect 174903 522806 174955 522851
rect 175901 522885 175953 522916
rect 175901 522851 175911 522885
rect 175945 522851 175953 522885
rect 175901 522806 175953 522851
rect 176007 522885 176059 522916
rect 176007 522851 176015 522885
rect 176049 522851 176059 522885
rect 176007 522806 176059 522851
rect 177005 522885 177057 522916
rect 177005 522851 177015 522885
rect 177049 522851 177057 522885
rect 177005 522806 177057 522851
rect 177111 522885 177163 522916
rect 177111 522851 177119 522885
rect 177153 522851 177163 522885
rect 177111 522806 177163 522851
rect 178109 522885 178161 522916
rect 178109 522851 178119 522885
rect 178153 522851 178161 522885
rect 178109 522806 178161 522851
rect 178215 522885 178267 522916
rect 178215 522851 178223 522885
rect 178257 522851 178267 522885
rect 178215 522806 178267 522851
rect 179213 522885 179265 522916
rect 179213 522851 179223 522885
rect 179257 522851 179265 522885
rect 179213 522806 179265 522851
rect 179319 522885 179371 522916
rect 179319 522851 179327 522885
rect 179361 522851 179371 522885
rect 179319 522806 179371 522851
rect 179765 522885 179817 522916
rect 179765 522851 179775 522885
rect 179809 522851 179817 522885
rect 179765 522806 179817 522851
rect 180055 522885 180107 522916
rect 180055 522851 180063 522885
rect 180097 522851 180107 522885
rect 180055 522806 180107 522851
rect 181053 522885 181105 522916
rect 181053 522851 181063 522885
rect 181097 522851 181105 522885
rect 181053 522806 181105 522851
rect 181159 522885 181211 522916
rect 181159 522851 181167 522885
rect 181201 522851 181211 522885
rect 181159 522806 181211 522851
rect 182157 522885 182209 522916
rect 182157 522851 182167 522885
rect 182201 522851 182209 522885
rect 182157 522806 182209 522851
rect 182263 522885 182315 522916
rect 182263 522851 182271 522885
rect 182305 522851 182315 522885
rect 182263 522806 182315 522851
rect 183261 522885 183313 522916
rect 183261 522851 183271 522885
rect 183305 522851 183313 522885
rect 183261 522806 183313 522851
rect 183367 522885 183419 522916
rect 183367 522851 183375 522885
rect 183409 522851 183419 522885
rect 183367 522806 183419 522851
rect 184365 522885 184417 522916
rect 184365 522851 184375 522885
rect 184409 522851 184417 522885
rect 184365 522806 184417 522851
rect 184471 522885 184523 522916
rect 184471 522851 184479 522885
rect 184513 522851 184523 522885
rect 184471 522806 184523 522851
rect 184917 522885 184969 522916
rect 184917 522851 184927 522885
rect 184961 522851 184969 522885
rect 184917 522806 184969 522851
rect 185207 522885 185259 522916
rect 185207 522851 185215 522885
rect 185249 522851 185259 522885
rect 185207 522806 185259 522851
rect 186205 522885 186257 522916
rect 186205 522851 186215 522885
rect 186249 522851 186257 522885
rect 186205 522806 186257 522851
rect 186311 522885 186363 522916
rect 186311 522851 186319 522885
rect 186353 522851 186363 522885
rect 186311 522806 186363 522851
rect 186941 522885 186993 522916
rect 186941 522851 186951 522885
rect 186985 522851 186993 522885
rect 186941 522806 186993 522851
rect 187231 522883 187283 522916
rect 187231 522849 187239 522883
rect 187273 522849 187283 522883
rect 187231 522806 187283 522849
rect 187401 522883 187453 522916
rect 187401 522849 187411 522883
rect 187445 522849 187453 522883
rect 187401 522806 187453 522849
rect 172235 521989 172287 522032
rect 172235 521955 172243 521989
rect 172277 521955 172287 521989
rect 172235 521922 172287 521955
rect 172405 521989 172457 522032
rect 172405 521955 172415 521989
rect 172449 521955 172457 521989
rect 172405 521922 172457 521955
rect 172511 521987 172563 522032
rect 172511 521953 172519 521987
rect 172553 521953 172563 521987
rect 172511 521922 172563 521953
rect 173509 521987 173561 522032
rect 173509 521953 173519 521987
rect 173553 521953 173561 521987
rect 173509 521922 173561 521953
rect 173615 521987 173667 522032
rect 173615 521953 173623 521987
rect 173657 521953 173667 521987
rect 173615 521922 173667 521953
rect 174613 521987 174665 522032
rect 174613 521953 174623 521987
rect 174657 521953 174665 521987
rect 174613 521922 174665 521953
rect 174719 521987 174771 522032
rect 174719 521953 174727 521987
rect 174761 521953 174771 521987
rect 174719 521922 174771 521953
rect 175717 521987 175769 522032
rect 175717 521953 175727 521987
rect 175761 521953 175769 521987
rect 175717 521922 175769 521953
rect 175823 521987 175875 522032
rect 175823 521953 175831 521987
rect 175865 521953 175875 521987
rect 175823 521922 175875 521953
rect 176821 521987 176873 522032
rect 176821 521953 176831 521987
rect 176865 521953 176873 521987
rect 176821 521922 176873 521953
rect 176927 521994 176979 522032
rect 176927 521960 176935 521994
rect 176969 521960 176979 521994
rect 176927 521922 176979 521960
rect 177189 521994 177241 522032
rect 177189 521960 177199 521994
rect 177233 521960 177241 521994
rect 177189 521922 177241 521960
rect 177479 521987 177531 522032
rect 177479 521953 177487 521987
rect 177521 521953 177531 521987
rect 177479 521922 177531 521953
rect 178477 521987 178529 522032
rect 178477 521953 178487 521987
rect 178521 521953 178529 521987
rect 178477 521922 178529 521953
rect 178583 521987 178635 522032
rect 178583 521953 178591 521987
rect 178625 521953 178635 521987
rect 178583 521922 178635 521953
rect 179581 521987 179633 522032
rect 179581 521953 179591 521987
rect 179625 521953 179633 521987
rect 179581 521922 179633 521953
rect 179687 521987 179739 522032
rect 179687 521953 179695 521987
rect 179729 521953 179739 521987
rect 179687 521922 179739 521953
rect 180685 521987 180737 522032
rect 180685 521953 180695 521987
rect 180729 521953 180737 521987
rect 180685 521922 180737 521953
rect 180791 521987 180843 522032
rect 180791 521953 180799 521987
rect 180833 521953 180843 521987
rect 180791 521922 180843 521953
rect 181789 521987 181841 522032
rect 181789 521953 181799 521987
rect 181833 521953 181841 521987
rect 181789 521922 181841 521953
rect 181895 521987 181947 522032
rect 181895 521953 181903 521987
rect 181937 521953 181947 521987
rect 181895 521922 181947 521953
rect 182341 521987 182393 522032
rect 182341 521953 182351 521987
rect 182385 521953 182393 521987
rect 182341 521922 182393 521953
rect 182631 521987 182683 522032
rect 182631 521953 182639 521987
rect 182673 521953 182683 521987
rect 182631 521922 182683 521953
rect 183629 521987 183681 522032
rect 183629 521953 183639 521987
rect 183673 521953 183681 521987
rect 183629 521922 183681 521953
rect 183735 521987 183787 522032
rect 183735 521953 183743 521987
rect 183777 521953 183787 521987
rect 183735 521922 183787 521953
rect 184733 521987 184785 522032
rect 184733 521953 184743 521987
rect 184777 521953 184785 521987
rect 184733 521922 184785 521953
rect 184839 521987 184891 522032
rect 184839 521953 184847 521987
rect 184881 521953 184891 521987
rect 184839 521922 184891 521953
rect 185837 521987 185889 522032
rect 185837 521953 185847 521987
rect 185881 521953 185889 521987
rect 185837 521922 185889 521953
rect 185943 521987 185995 522032
rect 185943 521953 185951 521987
rect 185985 521953 185995 521987
rect 185943 521922 185995 521953
rect 186941 521987 186993 522032
rect 186941 521953 186951 521987
rect 186985 521953 186993 521987
rect 186941 521922 186993 521953
rect 187231 521989 187283 522032
rect 187231 521955 187239 521989
rect 187273 521955 187283 521989
rect 187231 521922 187283 521955
rect 187401 521989 187453 522032
rect 187401 521955 187411 521989
rect 187445 521955 187453 521989
rect 187401 521922 187453 521955
rect 172235 521795 172287 521828
rect 172235 521761 172243 521795
rect 172277 521761 172287 521795
rect 172235 521718 172287 521761
rect 172405 521795 172457 521828
rect 172405 521761 172415 521795
rect 172449 521761 172457 521795
rect 172405 521718 172457 521761
rect 172511 521797 172563 521828
rect 172511 521763 172519 521797
rect 172553 521763 172563 521797
rect 172511 521718 172563 521763
rect 173509 521797 173561 521828
rect 173509 521763 173519 521797
rect 173553 521763 173561 521797
rect 173509 521718 173561 521763
rect 173615 521797 173667 521828
rect 173615 521763 173623 521797
rect 173657 521763 173667 521797
rect 173615 521718 173667 521763
rect 174613 521797 174665 521828
rect 174613 521763 174623 521797
rect 174657 521763 174665 521797
rect 174613 521718 174665 521763
rect 174903 521797 174955 521828
rect 174903 521763 174911 521797
rect 174945 521763 174955 521797
rect 174903 521718 174955 521763
rect 175901 521797 175953 521828
rect 175901 521763 175911 521797
rect 175945 521763 175953 521797
rect 175901 521718 175953 521763
rect 176007 521797 176059 521828
rect 176007 521763 176015 521797
rect 176049 521763 176059 521797
rect 176007 521718 176059 521763
rect 177005 521797 177057 521828
rect 177005 521763 177015 521797
rect 177049 521763 177057 521797
rect 177005 521718 177057 521763
rect 177111 521797 177163 521828
rect 177111 521763 177119 521797
rect 177153 521763 177163 521797
rect 177111 521718 177163 521763
rect 178109 521797 178161 521828
rect 178109 521763 178119 521797
rect 178153 521763 178161 521797
rect 178109 521718 178161 521763
rect 178215 521797 178267 521828
rect 178215 521763 178223 521797
rect 178257 521763 178267 521797
rect 178215 521718 178267 521763
rect 179213 521797 179265 521828
rect 179213 521763 179223 521797
rect 179257 521763 179265 521797
rect 179213 521718 179265 521763
rect 179319 521797 179371 521828
rect 179319 521763 179327 521797
rect 179361 521763 179371 521797
rect 179319 521718 179371 521763
rect 179765 521797 179817 521828
rect 179765 521763 179775 521797
rect 179809 521763 179817 521797
rect 179765 521718 179817 521763
rect 180055 521797 180107 521828
rect 180055 521763 180063 521797
rect 180097 521763 180107 521797
rect 180055 521718 180107 521763
rect 181053 521797 181105 521828
rect 181053 521763 181063 521797
rect 181097 521763 181105 521797
rect 181053 521718 181105 521763
rect 181159 521797 181211 521828
rect 181159 521763 181167 521797
rect 181201 521763 181211 521797
rect 181159 521718 181211 521763
rect 182157 521797 182209 521828
rect 182157 521763 182167 521797
rect 182201 521763 182209 521797
rect 182157 521718 182209 521763
rect 182263 521797 182315 521828
rect 182263 521763 182271 521797
rect 182305 521763 182315 521797
rect 182263 521718 182315 521763
rect 183261 521797 183313 521828
rect 183261 521763 183271 521797
rect 183305 521763 183313 521797
rect 183261 521718 183313 521763
rect 183367 521797 183419 521828
rect 183367 521763 183375 521797
rect 183409 521763 183419 521797
rect 183367 521718 183419 521763
rect 184365 521797 184417 521828
rect 184365 521763 184375 521797
rect 184409 521763 184417 521797
rect 184365 521718 184417 521763
rect 184471 521797 184523 521828
rect 184471 521763 184479 521797
rect 184513 521763 184523 521797
rect 184471 521718 184523 521763
rect 184917 521797 184969 521828
rect 184917 521763 184927 521797
rect 184961 521763 184969 521797
rect 184917 521718 184969 521763
rect 185207 521797 185259 521828
rect 185207 521763 185215 521797
rect 185249 521763 185259 521797
rect 185207 521718 185259 521763
rect 186205 521797 186257 521828
rect 186205 521763 186215 521797
rect 186249 521763 186257 521797
rect 186205 521718 186257 521763
rect 186311 521797 186363 521828
rect 186311 521763 186319 521797
rect 186353 521763 186363 521797
rect 186311 521718 186363 521763
rect 186941 521797 186993 521828
rect 186941 521763 186951 521797
rect 186985 521763 186993 521797
rect 186941 521718 186993 521763
rect 187231 521795 187283 521828
rect 187231 521761 187239 521795
rect 187273 521761 187283 521795
rect 187231 521718 187283 521761
rect 187401 521795 187453 521828
rect 187401 521761 187411 521795
rect 187445 521761 187453 521795
rect 187401 521718 187453 521761
rect 172235 520901 172287 520944
rect 172235 520867 172243 520901
rect 172277 520867 172287 520901
rect 172235 520834 172287 520867
rect 172405 520901 172457 520944
rect 172405 520867 172415 520901
rect 172449 520867 172457 520901
rect 172405 520834 172457 520867
rect 172511 520899 172563 520944
rect 172511 520865 172519 520899
rect 172553 520865 172563 520899
rect 172511 520834 172563 520865
rect 173509 520899 173561 520944
rect 173509 520865 173519 520899
rect 173553 520865 173561 520899
rect 173509 520834 173561 520865
rect 173615 520899 173667 520944
rect 173615 520865 173623 520899
rect 173657 520865 173667 520899
rect 173615 520834 173667 520865
rect 174613 520899 174665 520944
rect 174613 520865 174623 520899
rect 174657 520865 174665 520899
rect 174613 520834 174665 520865
rect 174719 520899 174771 520944
rect 174719 520865 174727 520899
rect 174761 520865 174771 520899
rect 174719 520834 174771 520865
rect 175717 520899 175769 520944
rect 175717 520865 175727 520899
rect 175761 520865 175769 520899
rect 175717 520834 175769 520865
rect 175823 520899 175875 520944
rect 175823 520865 175831 520899
rect 175865 520865 175875 520899
rect 175823 520834 175875 520865
rect 176821 520899 176873 520944
rect 176821 520865 176831 520899
rect 176865 520865 176873 520899
rect 176821 520834 176873 520865
rect 176927 520906 176979 520944
rect 176927 520872 176935 520906
rect 176969 520872 176979 520906
rect 176927 520834 176979 520872
rect 177189 520906 177241 520944
rect 177189 520872 177199 520906
rect 177233 520872 177241 520906
rect 177189 520834 177241 520872
rect 177479 520899 177531 520944
rect 177479 520865 177487 520899
rect 177521 520865 177531 520899
rect 177479 520834 177531 520865
rect 178477 520899 178529 520944
rect 178477 520865 178487 520899
rect 178521 520865 178529 520899
rect 178477 520834 178529 520865
rect 178583 520899 178635 520944
rect 178583 520865 178591 520899
rect 178625 520865 178635 520899
rect 178583 520834 178635 520865
rect 179581 520899 179633 520944
rect 179581 520865 179591 520899
rect 179625 520865 179633 520899
rect 179581 520834 179633 520865
rect 179687 520899 179739 520944
rect 179687 520865 179695 520899
rect 179729 520865 179739 520899
rect 179687 520834 179739 520865
rect 180685 520899 180737 520944
rect 180685 520865 180695 520899
rect 180729 520865 180737 520899
rect 180685 520834 180737 520865
rect 180791 520899 180843 520944
rect 180791 520865 180799 520899
rect 180833 520865 180843 520899
rect 180791 520834 180843 520865
rect 181789 520899 181841 520944
rect 181789 520865 181799 520899
rect 181833 520865 181841 520899
rect 181789 520834 181841 520865
rect 181895 520899 181947 520944
rect 181895 520865 181903 520899
rect 181937 520865 181947 520899
rect 181895 520834 181947 520865
rect 182341 520899 182393 520944
rect 182341 520865 182351 520899
rect 182385 520865 182393 520899
rect 182341 520834 182393 520865
rect 182631 520899 182683 520944
rect 182631 520865 182639 520899
rect 182673 520865 182683 520899
rect 182631 520834 182683 520865
rect 183629 520899 183681 520944
rect 183629 520865 183639 520899
rect 183673 520865 183681 520899
rect 183629 520834 183681 520865
rect 183735 520899 183787 520944
rect 183735 520865 183743 520899
rect 183777 520865 183787 520899
rect 183735 520834 183787 520865
rect 184733 520899 184785 520944
rect 184733 520865 184743 520899
rect 184777 520865 184785 520899
rect 184733 520834 184785 520865
rect 184839 520899 184891 520944
rect 184839 520865 184847 520899
rect 184881 520865 184891 520899
rect 184839 520834 184891 520865
rect 185837 520899 185889 520944
rect 185837 520865 185847 520899
rect 185881 520865 185889 520899
rect 185837 520834 185889 520865
rect 185943 520899 185995 520944
rect 185943 520865 185951 520899
rect 185985 520865 185995 520899
rect 185943 520834 185995 520865
rect 186941 520899 186993 520944
rect 186941 520865 186951 520899
rect 186985 520865 186993 520899
rect 186941 520834 186993 520865
rect 187231 520901 187283 520944
rect 187231 520867 187239 520901
rect 187273 520867 187283 520901
rect 187231 520834 187283 520867
rect 187401 520901 187453 520944
rect 187401 520867 187411 520901
rect 187445 520867 187453 520901
rect 187401 520834 187453 520867
rect 172235 520707 172287 520740
rect 172235 520673 172243 520707
rect 172277 520673 172287 520707
rect 172235 520630 172287 520673
rect 172405 520707 172457 520740
rect 172405 520673 172415 520707
rect 172449 520673 172457 520707
rect 172405 520630 172457 520673
rect 172511 520709 172563 520740
rect 172511 520675 172519 520709
rect 172553 520675 172563 520709
rect 172511 520630 172563 520675
rect 173509 520709 173561 520740
rect 173509 520675 173519 520709
rect 173553 520675 173561 520709
rect 173509 520630 173561 520675
rect 173615 520709 173667 520740
rect 173615 520675 173623 520709
rect 173657 520675 173667 520709
rect 173615 520630 173667 520675
rect 174613 520709 174665 520740
rect 174613 520675 174623 520709
rect 174657 520675 174665 520709
rect 174613 520630 174665 520675
rect 174903 520709 174955 520740
rect 174903 520675 174911 520709
rect 174945 520675 174955 520709
rect 174903 520630 174955 520675
rect 175901 520709 175953 520740
rect 175901 520675 175911 520709
rect 175945 520675 175953 520709
rect 175901 520630 175953 520675
rect 176007 520709 176059 520740
rect 176007 520675 176015 520709
rect 176049 520675 176059 520709
rect 176007 520630 176059 520675
rect 177005 520709 177057 520740
rect 177005 520675 177015 520709
rect 177049 520675 177057 520709
rect 177005 520630 177057 520675
rect 177111 520709 177163 520740
rect 177111 520675 177119 520709
rect 177153 520675 177163 520709
rect 177111 520630 177163 520675
rect 178109 520709 178161 520740
rect 178109 520675 178119 520709
rect 178153 520675 178161 520709
rect 178109 520630 178161 520675
rect 178215 520709 178267 520740
rect 178215 520675 178223 520709
rect 178257 520675 178267 520709
rect 178215 520630 178267 520675
rect 179213 520709 179265 520740
rect 179213 520675 179223 520709
rect 179257 520675 179265 520709
rect 179213 520630 179265 520675
rect 179319 520709 179371 520740
rect 179319 520675 179327 520709
rect 179361 520675 179371 520709
rect 179319 520630 179371 520675
rect 179765 520709 179817 520740
rect 179765 520675 179775 520709
rect 179809 520675 179817 520709
rect 179765 520630 179817 520675
rect 180055 520709 180107 520740
rect 180055 520675 180063 520709
rect 180097 520675 180107 520709
rect 180055 520630 180107 520675
rect 181053 520709 181105 520740
rect 181053 520675 181063 520709
rect 181097 520675 181105 520709
rect 181053 520630 181105 520675
rect 181159 520709 181211 520740
rect 181159 520675 181167 520709
rect 181201 520675 181211 520709
rect 181159 520630 181211 520675
rect 182157 520709 182209 520740
rect 182157 520675 182167 520709
rect 182201 520675 182209 520709
rect 182157 520630 182209 520675
rect 182263 520709 182315 520740
rect 182263 520675 182271 520709
rect 182305 520675 182315 520709
rect 182263 520630 182315 520675
rect 183261 520709 183313 520740
rect 183261 520675 183271 520709
rect 183305 520675 183313 520709
rect 183261 520630 183313 520675
rect 183367 520709 183419 520740
rect 183367 520675 183375 520709
rect 183409 520675 183419 520709
rect 183367 520630 183419 520675
rect 184365 520709 184417 520740
rect 184365 520675 184375 520709
rect 184409 520675 184417 520709
rect 184365 520630 184417 520675
rect 184471 520709 184523 520740
rect 184471 520675 184479 520709
rect 184513 520675 184523 520709
rect 184471 520630 184523 520675
rect 184917 520709 184969 520740
rect 184917 520675 184927 520709
rect 184961 520675 184969 520709
rect 184917 520630 184969 520675
rect 185207 520709 185259 520740
rect 185207 520675 185215 520709
rect 185249 520675 185259 520709
rect 185207 520630 185259 520675
rect 186205 520709 186257 520740
rect 186205 520675 186215 520709
rect 186249 520675 186257 520709
rect 186205 520630 186257 520675
rect 186311 520709 186363 520740
rect 186311 520675 186319 520709
rect 186353 520675 186363 520709
rect 186311 520630 186363 520675
rect 186941 520709 186993 520740
rect 186941 520675 186951 520709
rect 186985 520675 186993 520709
rect 186941 520630 186993 520675
rect 187231 520707 187283 520740
rect 187231 520673 187239 520707
rect 187273 520673 187283 520707
rect 187231 520630 187283 520673
rect 187401 520707 187453 520740
rect 187401 520673 187411 520707
rect 187445 520673 187453 520707
rect 187401 520630 187453 520673
rect 172235 519813 172287 519856
rect 172235 519779 172243 519813
rect 172277 519779 172287 519813
rect 172235 519746 172287 519779
rect 172405 519813 172457 519856
rect 172405 519779 172415 519813
rect 172449 519779 172457 519813
rect 172405 519746 172457 519779
rect 172511 519811 172563 519856
rect 172511 519777 172519 519811
rect 172553 519777 172563 519811
rect 172511 519746 172563 519777
rect 173509 519811 173561 519856
rect 173509 519777 173519 519811
rect 173553 519777 173561 519811
rect 173509 519746 173561 519777
rect 173615 519811 173667 519856
rect 173615 519777 173623 519811
rect 173657 519777 173667 519811
rect 173615 519746 173667 519777
rect 174613 519811 174665 519856
rect 174613 519777 174623 519811
rect 174657 519777 174665 519811
rect 174613 519746 174665 519777
rect 174719 519811 174771 519856
rect 174719 519777 174727 519811
rect 174761 519777 174771 519811
rect 174719 519746 174771 519777
rect 175717 519811 175769 519856
rect 175717 519777 175727 519811
rect 175761 519777 175769 519811
rect 175717 519746 175769 519777
rect 175823 519811 175875 519856
rect 175823 519777 175831 519811
rect 175865 519777 175875 519811
rect 175823 519746 175875 519777
rect 176821 519811 176873 519856
rect 176821 519777 176831 519811
rect 176865 519777 176873 519811
rect 176821 519746 176873 519777
rect 176927 519818 176979 519856
rect 176927 519784 176935 519818
rect 176969 519784 176979 519818
rect 176927 519746 176979 519784
rect 177189 519818 177241 519856
rect 177189 519784 177199 519818
rect 177233 519784 177241 519818
rect 177189 519746 177241 519784
rect 177479 519811 177531 519856
rect 177479 519777 177487 519811
rect 177521 519777 177531 519811
rect 177479 519746 177531 519777
rect 178477 519811 178529 519856
rect 178477 519777 178487 519811
rect 178521 519777 178529 519811
rect 178477 519746 178529 519777
rect 178583 519811 178635 519856
rect 178583 519777 178591 519811
rect 178625 519777 178635 519811
rect 178583 519746 178635 519777
rect 179581 519811 179633 519856
rect 179581 519777 179591 519811
rect 179625 519777 179633 519811
rect 179581 519746 179633 519777
rect 179687 519811 179739 519856
rect 179687 519777 179695 519811
rect 179729 519777 179739 519811
rect 179687 519746 179739 519777
rect 180685 519811 180737 519856
rect 180685 519777 180695 519811
rect 180729 519777 180737 519811
rect 180685 519746 180737 519777
rect 180791 519811 180843 519856
rect 180791 519777 180799 519811
rect 180833 519777 180843 519811
rect 180791 519746 180843 519777
rect 181789 519811 181841 519856
rect 181789 519777 181799 519811
rect 181833 519777 181841 519811
rect 181789 519746 181841 519777
rect 181895 519811 181947 519856
rect 181895 519777 181903 519811
rect 181937 519777 181947 519811
rect 181895 519746 181947 519777
rect 182341 519811 182393 519856
rect 182341 519777 182351 519811
rect 182385 519777 182393 519811
rect 182341 519746 182393 519777
rect 182631 519811 182683 519856
rect 182631 519777 182639 519811
rect 182673 519777 182683 519811
rect 182631 519746 182683 519777
rect 183629 519811 183681 519856
rect 183629 519777 183639 519811
rect 183673 519777 183681 519811
rect 183629 519746 183681 519777
rect 183735 519811 183787 519856
rect 183735 519777 183743 519811
rect 183777 519777 183787 519811
rect 183735 519746 183787 519777
rect 184733 519811 184785 519856
rect 184733 519777 184743 519811
rect 184777 519777 184785 519811
rect 184733 519746 184785 519777
rect 184839 519811 184891 519856
rect 184839 519777 184847 519811
rect 184881 519777 184891 519811
rect 184839 519746 184891 519777
rect 185837 519811 185889 519856
rect 185837 519777 185847 519811
rect 185881 519777 185889 519811
rect 185837 519746 185889 519777
rect 185943 519811 185995 519856
rect 185943 519777 185951 519811
rect 185985 519777 185995 519811
rect 185943 519746 185995 519777
rect 186941 519811 186993 519856
rect 186941 519777 186951 519811
rect 186985 519777 186993 519811
rect 186941 519746 186993 519777
rect 187231 519813 187283 519856
rect 187231 519779 187239 519813
rect 187273 519779 187283 519813
rect 187231 519746 187283 519779
rect 187401 519813 187453 519856
rect 187401 519779 187411 519813
rect 187445 519779 187453 519813
rect 187401 519746 187453 519779
rect 172235 519619 172287 519652
rect 172235 519585 172243 519619
rect 172277 519585 172287 519619
rect 172235 519542 172287 519585
rect 172405 519619 172457 519652
rect 172405 519585 172415 519619
rect 172449 519585 172457 519619
rect 172405 519542 172457 519585
rect 172511 519621 172563 519652
rect 172511 519587 172519 519621
rect 172553 519587 172563 519621
rect 172511 519542 172563 519587
rect 173509 519621 173561 519652
rect 173509 519587 173519 519621
rect 173553 519587 173561 519621
rect 173509 519542 173561 519587
rect 173615 519621 173667 519652
rect 173615 519587 173623 519621
rect 173657 519587 173667 519621
rect 173615 519542 173667 519587
rect 174613 519621 174665 519652
rect 174613 519587 174623 519621
rect 174657 519587 174665 519621
rect 174613 519542 174665 519587
rect 174903 519621 174955 519652
rect 174903 519587 174911 519621
rect 174945 519587 174955 519621
rect 174903 519542 174955 519587
rect 175901 519621 175953 519652
rect 175901 519587 175911 519621
rect 175945 519587 175953 519621
rect 175901 519542 175953 519587
rect 176007 519621 176059 519652
rect 176007 519587 176015 519621
rect 176049 519587 176059 519621
rect 176007 519542 176059 519587
rect 177005 519621 177057 519652
rect 177005 519587 177015 519621
rect 177049 519587 177057 519621
rect 177005 519542 177057 519587
rect 177111 519621 177163 519652
rect 177111 519587 177119 519621
rect 177153 519587 177163 519621
rect 177111 519542 177163 519587
rect 178109 519621 178161 519652
rect 178109 519587 178119 519621
rect 178153 519587 178161 519621
rect 178109 519542 178161 519587
rect 178215 519621 178267 519652
rect 178215 519587 178223 519621
rect 178257 519587 178267 519621
rect 178215 519542 178267 519587
rect 179213 519621 179265 519652
rect 179213 519587 179223 519621
rect 179257 519587 179265 519621
rect 179213 519542 179265 519587
rect 179319 519621 179371 519652
rect 179319 519587 179327 519621
rect 179361 519587 179371 519621
rect 179319 519542 179371 519587
rect 179765 519621 179817 519652
rect 179765 519587 179775 519621
rect 179809 519587 179817 519621
rect 179765 519542 179817 519587
rect 180055 519621 180107 519652
rect 180055 519587 180063 519621
rect 180097 519587 180107 519621
rect 180055 519542 180107 519587
rect 181053 519621 181105 519652
rect 181053 519587 181063 519621
rect 181097 519587 181105 519621
rect 181053 519542 181105 519587
rect 181159 519621 181211 519652
rect 181159 519587 181167 519621
rect 181201 519587 181211 519621
rect 181159 519542 181211 519587
rect 182157 519621 182209 519652
rect 182157 519587 182167 519621
rect 182201 519587 182209 519621
rect 182157 519542 182209 519587
rect 182263 519621 182315 519652
rect 182263 519587 182271 519621
rect 182305 519587 182315 519621
rect 182263 519542 182315 519587
rect 183261 519621 183313 519652
rect 183261 519587 183271 519621
rect 183305 519587 183313 519621
rect 183261 519542 183313 519587
rect 183367 519621 183419 519652
rect 183367 519587 183375 519621
rect 183409 519587 183419 519621
rect 183367 519542 183419 519587
rect 184365 519621 184417 519652
rect 184365 519587 184375 519621
rect 184409 519587 184417 519621
rect 184365 519542 184417 519587
rect 184471 519621 184523 519652
rect 184471 519587 184479 519621
rect 184513 519587 184523 519621
rect 184471 519542 184523 519587
rect 184917 519621 184969 519652
rect 184917 519587 184927 519621
rect 184961 519587 184969 519621
rect 184917 519542 184969 519587
rect 185207 519621 185259 519652
rect 185207 519587 185215 519621
rect 185249 519587 185259 519621
rect 185207 519542 185259 519587
rect 186205 519621 186257 519652
rect 186205 519587 186215 519621
rect 186249 519587 186257 519621
rect 186205 519542 186257 519587
rect 186311 519621 186363 519652
rect 186311 519587 186319 519621
rect 186353 519587 186363 519621
rect 186311 519542 186363 519587
rect 186941 519621 186993 519652
rect 186941 519587 186951 519621
rect 186985 519587 186993 519621
rect 186941 519542 186993 519587
rect 187231 519619 187283 519652
rect 187231 519585 187239 519619
rect 187273 519585 187283 519619
rect 187231 519542 187283 519585
rect 187401 519619 187453 519652
rect 187401 519585 187411 519619
rect 187445 519585 187453 519619
rect 187401 519542 187453 519585
rect 172235 518725 172287 518768
rect 172235 518691 172243 518725
rect 172277 518691 172287 518725
rect 172235 518658 172287 518691
rect 172405 518725 172457 518768
rect 172405 518691 172415 518725
rect 172449 518691 172457 518725
rect 172405 518658 172457 518691
rect 172511 518723 172563 518768
rect 172511 518689 172519 518723
rect 172553 518689 172563 518723
rect 172511 518658 172563 518689
rect 173509 518723 173561 518768
rect 173509 518689 173519 518723
rect 173553 518689 173561 518723
rect 173509 518658 173561 518689
rect 173615 518723 173667 518768
rect 173615 518689 173623 518723
rect 173657 518689 173667 518723
rect 173615 518658 173667 518689
rect 174613 518723 174665 518768
rect 174613 518689 174623 518723
rect 174657 518689 174665 518723
rect 174613 518658 174665 518689
rect 174719 518723 174771 518768
rect 174719 518689 174727 518723
rect 174761 518689 174771 518723
rect 174719 518658 174771 518689
rect 175717 518723 175769 518768
rect 175717 518689 175727 518723
rect 175761 518689 175769 518723
rect 175717 518658 175769 518689
rect 175823 518723 175875 518768
rect 175823 518689 175831 518723
rect 175865 518689 175875 518723
rect 175823 518658 175875 518689
rect 176821 518723 176873 518768
rect 176821 518689 176831 518723
rect 176865 518689 176873 518723
rect 176821 518658 176873 518689
rect 176927 518730 176979 518768
rect 176927 518696 176935 518730
rect 176969 518696 176979 518730
rect 176927 518658 176979 518696
rect 177189 518730 177241 518768
rect 177189 518696 177199 518730
rect 177233 518696 177241 518730
rect 177189 518658 177241 518696
rect 177479 518723 177531 518768
rect 177479 518689 177487 518723
rect 177521 518689 177531 518723
rect 177479 518658 177531 518689
rect 178477 518723 178529 518768
rect 178477 518689 178487 518723
rect 178521 518689 178529 518723
rect 178477 518658 178529 518689
rect 178583 518723 178635 518768
rect 178583 518689 178591 518723
rect 178625 518689 178635 518723
rect 178583 518658 178635 518689
rect 179581 518723 179633 518768
rect 179581 518689 179591 518723
rect 179625 518689 179633 518723
rect 179581 518658 179633 518689
rect 179687 518723 179739 518768
rect 179687 518689 179695 518723
rect 179729 518689 179739 518723
rect 179687 518658 179739 518689
rect 180685 518723 180737 518768
rect 180685 518689 180695 518723
rect 180729 518689 180737 518723
rect 180685 518658 180737 518689
rect 180791 518723 180843 518768
rect 180791 518689 180799 518723
rect 180833 518689 180843 518723
rect 180791 518658 180843 518689
rect 181789 518723 181841 518768
rect 181789 518689 181799 518723
rect 181833 518689 181841 518723
rect 181789 518658 181841 518689
rect 181895 518723 181947 518768
rect 181895 518689 181903 518723
rect 181937 518689 181947 518723
rect 181895 518658 181947 518689
rect 182341 518723 182393 518768
rect 182341 518689 182351 518723
rect 182385 518689 182393 518723
rect 182341 518658 182393 518689
rect 182631 518723 182683 518768
rect 182631 518689 182639 518723
rect 182673 518689 182683 518723
rect 182631 518658 182683 518689
rect 183629 518723 183681 518768
rect 183629 518689 183639 518723
rect 183673 518689 183681 518723
rect 183629 518658 183681 518689
rect 183735 518723 183787 518768
rect 183735 518689 183743 518723
rect 183777 518689 183787 518723
rect 183735 518658 183787 518689
rect 184733 518723 184785 518768
rect 184733 518689 184743 518723
rect 184777 518689 184785 518723
rect 184733 518658 184785 518689
rect 184839 518723 184891 518768
rect 184839 518689 184847 518723
rect 184881 518689 184891 518723
rect 184839 518658 184891 518689
rect 185837 518723 185889 518768
rect 185837 518689 185847 518723
rect 185881 518689 185889 518723
rect 185837 518658 185889 518689
rect 185943 518723 185995 518768
rect 185943 518689 185951 518723
rect 185985 518689 185995 518723
rect 185943 518658 185995 518689
rect 186941 518723 186993 518768
rect 186941 518689 186951 518723
rect 186985 518689 186993 518723
rect 186941 518658 186993 518689
rect 187231 518725 187283 518768
rect 187231 518691 187239 518725
rect 187273 518691 187283 518725
rect 187231 518658 187283 518691
rect 187401 518725 187453 518768
rect 187401 518691 187411 518725
rect 187445 518691 187453 518725
rect 187401 518658 187453 518691
rect 172235 518531 172287 518564
rect 172235 518497 172243 518531
rect 172277 518497 172287 518531
rect 172235 518454 172287 518497
rect 172405 518531 172457 518564
rect 172405 518497 172415 518531
rect 172449 518497 172457 518531
rect 172405 518454 172457 518497
rect 172511 518533 172563 518564
rect 172511 518499 172519 518533
rect 172553 518499 172563 518533
rect 172511 518454 172563 518499
rect 173509 518533 173561 518564
rect 173509 518499 173519 518533
rect 173553 518499 173561 518533
rect 173509 518454 173561 518499
rect 173615 518533 173667 518564
rect 173615 518499 173623 518533
rect 173657 518499 173667 518533
rect 173615 518454 173667 518499
rect 174613 518533 174665 518564
rect 174613 518499 174623 518533
rect 174657 518499 174665 518533
rect 174613 518454 174665 518499
rect 174903 518533 174955 518564
rect 174903 518499 174911 518533
rect 174945 518499 174955 518533
rect 174903 518454 174955 518499
rect 175901 518533 175953 518564
rect 175901 518499 175911 518533
rect 175945 518499 175953 518533
rect 175901 518454 175953 518499
rect 176007 518533 176059 518564
rect 176007 518499 176015 518533
rect 176049 518499 176059 518533
rect 176007 518454 176059 518499
rect 177005 518533 177057 518564
rect 177005 518499 177015 518533
rect 177049 518499 177057 518533
rect 177005 518454 177057 518499
rect 177111 518533 177163 518564
rect 177111 518499 177119 518533
rect 177153 518499 177163 518533
rect 177111 518454 177163 518499
rect 178109 518533 178161 518564
rect 178109 518499 178119 518533
rect 178153 518499 178161 518533
rect 178109 518454 178161 518499
rect 178215 518533 178267 518564
rect 178215 518499 178223 518533
rect 178257 518499 178267 518533
rect 178215 518454 178267 518499
rect 179213 518533 179265 518564
rect 179213 518499 179223 518533
rect 179257 518499 179265 518533
rect 179213 518454 179265 518499
rect 179319 518533 179371 518564
rect 179319 518499 179327 518533
rect 179361 518499 179371 518533
rect 179319 518454 179371 518499
rect 179765 518533 179817 518564
rect 179765 518499 179775 518533
rect 179809 518499 179817 518533
rect 179765 518454 179817 518499
rect 180055 518533 180107 518564
rect 180055 518499 180063 518533
rect 180097 518499 180107 518533
rect 180055 518454 180107 518499
rect 181053 518533 181105 518564
rect 181053 518499 181063 518533
rect 181097 518499 181105 518533
rect 181053 518454 181105 518499
rect 181159 518533 181211 518564
rect 181159 518499 181167 518533
rect 181201 518499 181211 518533
rect 181159 518454 181211 518499
rect 182157 518533 182209 518564
rect 182157 518499 182167 518533
rect 182201 518499 182209 518533
rect 182157 518454 182209 518499
rect 182263 518533 182315 518564
rect 182263 518499 182271 518533
rect 182305 518499 182315 518533
rect 182263 518454 182315 518499
rect 183261 518533 183313 518564
rect 183261 518499 183271 518533
rect 183305 518499 183313 518533
rect 183261 518454 183313 518499
rect 183367 518533 183419 518564
rect 183367 518499 183375 518533
rect 183409 518499 183419 518533
rect 183367 518454 183419 518499
rect 184365 518533 184417 518564
rect 184365 518499 184375 518533
rect 184409 518499 184417 518533
rect 184365 518454 184417 518499
rect 184471 518533 184523 518564
rect 184471 518499 184479 518533
rect 184513 518499 184523 518533
rect 184471 518454 184523 518499
rect 184917 518533 184969 518564
rect 184917 518499 184927 518533
rect 184961 518499 184969 518533
rect 184917 518454 184969 518499
rect 185207 518533 185259 518564
rect 185207 518499 185215 518533
rect 185249 518499 185259 518533
rect 185207 518454 185259 518499
rect 186205 518533 186257 518564
rect 186205 518499 186215 518533
rect 186249 518499 186257 518533
rect 186205 518454 186257 518499
rect 186311 518533 186363 518564
rect 186311 518499 186319 518533
rect 186353 518499 186363 518533
rect 186311 518454 186363 518499
rect 186941 518533 186993 518564
rect 186941 518499 186951 518533
rect 186985 518499 186993 518533
rect 186941 518454 186993 518499
rect 187231 518531 187283 518564
rect 187231 518497 187239 518531
rect 187273 518497 187283 518531
rect 187231 518454 187283 518497
rect 187401 518531 187453 518564
rect 187401 518497 187411 518531
rect 187445 518497 187453 518531
rect 187401 518454 187453 518497
rect 172235 517637 172287 517680
rect 172235 517603 172243 517637
rect 172277 517603 172287 517637
rect 172235 517570 172287 517603
rect 172405 517637 172457 517680
rect 172405 517603 172415 517637
rect 172449 517603 172457 517637
rect 172405 517570 172457 517603
rect 172511 517635 172563 517680
rect 172511 517601 172519 517635
rect 172553 517601 172563 517635
rect 172511 517570 172563 517601
rect 173509 517635 173561 517680
rect 173509 517601 173519 517635
rect 173553 517601 173561 517635
rect 173509 517570 173561 517601
rect 173615 517635 173667 517680
rect 173615 517601 173623 517635
rect 173657 517601 173667 517635
rect 173615 517570 173667 517601
rect 174613 517635 174665 517680
rect 174613 517601 174623 517635
rect 174657 517601 174665 517635
rect 174613 517570 174665 517601
rect 174719 517635 174771 517680
rect 174719 517601 174727 517635
rect 174761 517601 174771 517635
rect 174719 517570 174771 517601
rect 175717 517635 175769 517680
rect 175717 517601 175727 517635
rect 175761 517601 175769 517635
rect 175717 517570 175769 517601
rect 175823 517635 175875 517680
rect 175823 517601 175831 517635
rect 175865 517601 175875 517635
rect 175823 517570 175875 517601
rect 176821 517635 176873 517680
rect 176821 517601 176831 517635
rect 176865 517601 176873 517635
rect 176821 517570 176873 517601
rect 176927 517642 176979 517680
rect 176927 517608 176935 517642
rect 176969 517608 176979 517642
rect 176927 517570 176979 517608
rect 177189 517642 177241 517680
rect 177189 517608 177199 517642
rect 177233 517608 177241 517642
rect 177189 517570 177241 517608
rect 177479 517635 177531 517680
rect 177479 517601 177487 517635
rect 177521 517601 177531 517635
rect 177479 517570 177531 517601
rect 178477 517635 178529 517680
rect 178477 517601 178487 517635
rect 178521 517601 178529 517635
rect 178477 517570 178529 517601
rect 178583 517635 178635 517680
rect 178583 517601 178591 517635
rect 178625 517601 178635 517635
rect 178583 517570 178635 517601
rect 179581 517635 179633 517680
rect 179581 517601 179591 517635
rect 179625 517601 179633 517635
rect 179581 517570 179633 517601
rect 179687 517635 179739 517680
rect 179687 517601 179695 517635
rect 179729 517601 179739 517635
rect 179687 517570 179739 517601
rect 180685 517635 180737 517680
rect 180685 517601 180695 517635
rect 180729 517601 180737 517635
rect 180685 517570 180737 517601
rect 180791 517635 180843 517680
rect 180791 517601 180799 517635
rect 180833 517601 180843 517635
rect 180791 517570 180843 517601
rect 181789 517635 181841 517680
rect 181789 517601 181799 517635
rect 181833 517601 181841 517635
rect 181789 517570 181841 517601
rect 181895 517635 181947 517680
rect 181895 517601 181903 517635
rect 181937 517601 181947 517635
rect 181895 517570 181947 517601
rect 182341 517635 182393 517680
rect 182341 517601 182351 517635
rect 182385 517601 182393 517635
rect 182341 517570 182393 517601
rect 182631 517635 182683 517680
rect 182631 517601 182639 517635
rect 182673 517601 182683 517635
rect 182631 517570 182683 517601
rect 183629 517635 183681 517680
rect 183629 517601 183639 517635
rect 183673 517601 183681 517635
rect 183629 517570 183681 517601
rect 183735 517635 183787 517680
rect 183735 517601 183743 517635
rect 183777 517601 183787 517635
rect 183735 517570 183787 517601
rect 184733 517635 184785 517680
rect 184733 517601 184743 517635
rect 184777 517601 184785 517635
rect 184733 517570 184785 517601
rect 184839 517635 184891 517680
rect 184839 517601 184847 517635
rect 184881 517601 184891 517635
rect 184839 517570 184891 517601
rect 185837 517635 185889 517680
rect 185837 517601 185847 517635
rect 185881 517601 185889 517635
rect 185837 517570 185889 517601
rect 185943 517635 185995 517680
rect 185943 517601 185951 517635
rect 185985 517601 185995 517635
rect 185943 517570 185995 517601
rect 186941 517635 186993 517680
rect 186941 517601 186951 517635
rect 186985 517601 186993 517635
rect 186941 517570 186993 517601
rect 187231 517637 187283 517680
rect 187231 517603 187239 517637
rect 187273 517603 187283 517637
rect 187231 517570 187283 517603
rect 187401 517637 187453 517680
rect 187401 517603 187411 517637
rect 187445 517603 187453 517637
rect 187401 517570 187453 517603
rect 172235 517443 172287 517476
rect 172235 517409 172243 517443
rect 172277 517409 172287 517443
rect 172235 517366 172287 517409
rect 172405 517443 172457 517476
rect 172405 517409 172415 517443
rect 172449 517409 172457 517443
rect 172405 517366 172457 517409
rect 172511 517445 172563 517476
rect 172511 517411 172519 517445
rect 172553 517411 172563 517445
rect 172511 517366 172563 517411
rect 173509 517445 173561 517476
rect 173509 517411 173519 517445
rect 173553 517411 173561 517445
rect 173509 517366 173561 517411
rect 173615 517445 173667 517476
rect 173615 517411 173623 517445
rect 173657 517411 173667 517445
rect 173615 517366 173667 517411
rect 174613 517445 174665 517476
rect 174613 517411 174623 517445
rect 174657 517411 174665 517445
rect 174613 517366 174665 517411
rect 174903 517445 174955 517476
rect 174903 517411 174911 517445
rect 174945 517411 174955 517445
rect 174903 517366 174955 517411
rect 175901 517445 175953 517476
rect 175901 517411 175911 517445
rect 175945 517411 175953 517445
rect 175901 517366 175953 517411
rect 176007 517445 176059 517476
rect 176007 517411 176015 517445
rect 176049 517411 176059 517445
rect 176007 517366 176059 517411
rect 177005 517445 177057 517476
rect 177005 517411 177015 517445
rect 177049 517411 177057 517445
rect 177005 517366 177057 517411
rect 177111 517445 177163 517476
rect 177111 517411 177119 517445
rect 177153 517411 177163 517445
rect 177111 517366 177163 517411
rect 178109 517445 178161 517476
rect 178109 517411 178119 517445
rect 178153 517411 178161 517445
rect 178109 517366 178161 517411
rect 178215 517445 178267 517476
rect 178215 517411 178223 517445
rect 178257 517411 178267 517445
rect 178215 517366 178267 517411
rect 179213 517445 179265 517476
rect 179213 517411 179223 517445
rect 179257 517411 179265 517445
rect 179213 517366 179265 517411
rect 179319 517445 179371 517476
rect 179319 517411 179327 517445
rect 179361 517411 179371 517445
rect 179319 517366 179371 517411
rect 179765 517445 179817 517476
rect 179765 517411 179775 517445
rect 179809 517411 179817 517445
rect 179765 517366 179817 517411
rect 180055 517445 180107 517476
rect 180055 517411 180063 517445
rect 180097 517411 180107 517445
rect 180055 517366 180107 517411
rect 181053 517445 181105 517476
rect 181053 517411 181063 517445
rect 181097 517411 181105 517445
rect 181053 517366 181105 517411
rect 181159 517445 181211 517476
rect 181159 517411 181167 517445
rect 181201 517411 181211 517445
rect 181159 517366 181211 517411
rect 182157 517445 182209 517476
rect 182157 517411 182167 517445
rect 182201 517411 182209 517445
rect 182157 517366 182209 517411
rect 182263 517445 182315 517476
rect 182263 517411 182271 517445
rect 182305 517411 182315 517445
rect 182263 517366 182315 517411
rect 183261 517445 183313 517476
rect 183261 517411 183271 517445
rect 183305 517411 183313 517445
rect 183261 517366 183313 517411
rect 183367 517445 183419 517476
rect 183367 517411 183375 517445
rect 183409 517411 183419 517445
rect 183367 517366 183419 517411
rect 184365 517445 184417 517476
rect 184365 517411 184375 517445
rect 184409 517411 184417 517445
rect 184365 517366 184417 517411
rect 184471 517445 184523 517476
rect 184471 517411 184479 517445
rect 184513 517411 184523 517445
rect 184471 517366 184523 517411
rect 184917 517445 184969 517476
rect 184917 517411 184927 517445
rect 184961 517411 184969 517445
rect 184917 517366 184969 517411
rect 185207 517445 185259 517476
rect 185207 517411 185215 517445
rect 185249 517411 185259 517445
rect 185207 517366 185259 517411
rect 186205 517445 186257 517476
rect 186205 517411 186215 517445
rect 186249 517411 186257 517445
rect 186205 517366 186257 517411
rect 186311 517445 186363 517476
rect 186311 517411 186319 517445
rect 186353 517411 186363 517445
rect 186311 517366 186363 517411
rect 186941 517445 186993 517476
rect 186941 517411 186951 517445
rect 186985 517411 186993 517445
rect 186941 517366 186993 517411
rect 187231 517443 187283 517476
rect 187231 517409 187239 517443
rect 187273 517409 187283 517443
rect 187231 517366 187283 517409
rect 187401 517443 187453 517476
rect 187401 517409 187411 517443
rect 187445 517409 187453 517443
rect 187401 517366 187453 517409
rect 172235 516549 172287 516592
rect 172235 516515 172243 516549
rect 172277 516515 172287 516549
rect 172235 516482 172287 516515
rect 172405 516549 172457 516592
rect 172405 516515 172415 516549
rect 172449 516515 172457 516549
rect 172405 516482 172457 516515
rect 172511 516547 172563 516592
rect 172511 516513 172519 516547
rect 172553 516513 172563 516547
rect 172511 516482 172563 516513
rect 173509 516547 173561 516592
rect 173509 516513 173519 516547
rect 173553 516513 173561 516547
rect 173509 516482 173561 516513
rect 173615 516547 173667 516592
rect 173615 516513 173623 516547
rect 173657 516513 173667 516547
rect 173615 516482 173667 516513
rect 174613 516547 174665 516592
rect 174613 516513 174623 516547
rect 174657 516513 174665 516547
rect 174613 516482 174665 516513
rect 174719 516547 174771 516592
rect 174719 516513 174727 516547
rect 174761 516513 174771 516547
rect 174719 516482 174771 516513
rect 175717 516547 175769 516592
rect 175717 516513 175727 516547
rect 175761 516513 175769 516547
rect 175717 516482 175769 516513
rect 175823 516547 175875 516592
rect 175823 516513 175831 516547
rect 175865 516513 175875 516547
rect 175823 516482 175875 516513
rect 176821 516547 176873 516592
rect 176821 516513 176831 516547
rect 176865 516513 176873 516547
rect 176821 516482 176873 516513
rect 176927 516554 176979 516592
rect 176927 516520 176935 516554
rect 176969 516520 176979 516554
rect 176927 516482 176979 516520
rect 177189 516554 177241 516592
rect 177189 516520 177199 516554
rect 177233 516520 177241 516554
rect 177189 516482 177241 516520
rect 177479 516547 177531 516592
rect 177479 516513 177487 516547
rect 177521 516513 177531 516547
rect 177479 516482 177531 516513
rect 178477 516547 178529 516592
rect 178477 516513 178487 516547
rect 178521 516513 178529 516547
rect 178477 516482 178529 516513
rect 178583 516547 178635 516592
rect 178583 516513 178591 516547
rect 178625 516513 178635 516547
rect 178583 516482 178635 516513
rect 179581 516547 179633 516592
rect 179581 516513 179591 516547
rect 179625 516513 179633 516547
rect 179581 516482 179633 516513
rect 179687 516547 179739 516592
rect 179687 516513 179695 516547
rect 179729 516513 179739 516547
rect 179687 516482 179739 516513
rect 180685 516547 180737 516592
rect 180685 516513 180695 516547
rect 180729 516513 180737 516547
rect 180685 516482 180737 516513
rect 180791 516547 180843 516592
rect 180791 516513 180799 516547
rect 180833 516513 180843 516547
rect 180791 516482 180843 516513
rect 181789 516547 181841 516592
rect 181789 516513 181799 516547
rect 181833 516513 181841 516547
rect 181789 516482 181841 516513
rect 181895 516547 181947 516592
rect 181895 516513 181903 516547
rect 181937 516513 181947 516547
rect 181895 516482 181947 516513
rect 182341 516547 182393 516592
rect 182341 516513 182351 516547
rect 182385 516513 182393 516547
rect 182341 516482 182393 516513
rect 182631 516547 182683 516592
rect 182631 516513 182639 516547
rect 182673 516513 182683 516547
rect 182631 516482 182683 516513
rect 183629 516547 183681 516592
rect 183629 516513 183639 516547
rect 183673 516513 183681 516547
rect 183629 516482 183681 516513
rect 183735 516547 183787 516592
rect 183735 516513 183743 516547
rect 183777 516513 183787 516547
rect 183735 516482 183787 516513
rect 184733 516547 184785 516592
rect 184733 516513 184743 516547
rect 184777 516513 184785 516547
rect 184733 516482 184785 516513
rect 184839 516547 184891 516592
rect 184839 516513 184847 516547
rect 184881 516513 184891 516547
rect 184839 516482 184891 516513
rect 185837 516547 185889 516592
rect 185837 516513 185847 516547
rect 185881 516513 185889 516547
rect 185837 516482 185889 516513
rect 185943 516547 185995 516592
rect 185943 516513 185951 516547
rect 185985 516513 185995 516547
rect 185943 516482 185995 516513
rect 186941 516547 186993 516592
rect 186941 516513 186951 516547
rect 186985 516513 186993 516547
rect 186941 516482 186993 516513
rect 187231 516549 187283 516592
rect 187231 516515 187239 516549
rect 187273 516515 187283 516549
rect 187231 516482 187283 516515
rect 187401 516549 187453 516592
rect 187401 516515 187411 516549
rect 187445 516515 187453 516549
rect 187401 516482 187453 516515
rect 172235 516355 172287 516388
rect 172235 516321 172243 516355
rect 172277 516321 172287 516355
rect 172235 516278 172287 516321
rect 172405 516355 172457 516388
rect 172405 516321 172415 516355
rect 172449 516321 172457 516355
rect 172405 516278 172457 516321
rect 172511 516357 172563 516388
rect 172511 516323 172519 516357
rect 172553 516323 172563 516357
rect 172511 516278 172563 516323
rect 173509 516357 173561 516388
rect 173509 516323 173519 516357
rect 173553 516323 173561 516357
rect 173509 516278 173561 516323
rect 173615 516357 173667 516388
rect 173615 516323 173623 516357
rect 173657 516323 173667 516357
rect 173615 516278 173667 516323
rect 174613 516357 174665 516388
rect 174613 516323 174623 516357
rect 174657 516323 174665 516357
rect 174613 516278 174665 516323
rect 174903 516357 174955 516388
rect 174903 516323 174911 516357
rect 174945 516323 174955 516357
rect 174903 516278 174955 516323
rect 175901 516357 175953 516388
rect 175901 516323 175911 516357
rect 175945 516323 175953 516357
rect 175901 516278 175953 516323
rect 176007 516357 176059 516388
rect 176007 516323 176015 516357
rect 176049 516323 176059 516357
rect 176007 516278 176059 516323
rect 177005 516357 177057 516388
rect 177005 516323 177015 516357
rect 177049 516323 177057 516357
rect 177005 516278 177057 516323
rect 177111 516357 177163 516388
rect 177111 516323 177119 516357
rect 177153 516323 177163 516357
rect 177111 516278 177163 516323
rect 178109 516357 178161 516388
rect 178109 516323 178119 516357
rect 178153 516323 178161 516357
rect 178109 516278 178161 516323
rect 178215 516357 178267 516388
rect 178215 516323 178223 516357
rect 178257 516323 178267 516357
rect 178215 516278 178267 516323
rect 179213 516357 179265 516388
rect 179213 516323 179223 516357
rect 179257 516323 179265 516357
rect 179213 516278 179265 516323
rect 179319 516357 179371 516388
rect 179319 516323 179327 516357
rect 179361 516323 179371 516357
rect 179319 516278 179371 516323
rect 179765 516357 179817 516388
rect 179765 516323 179775 516357
rect 179809 516323 179817 516357
rect 179765 516278 179817 516323
rect 180055 516357 180107 516388
rect 180055 516323 180063 516357
rect 180097 516323 180107 516357
rect 180055 516278 180107 516323
rect 181053 516357 181105 516388
rect 181053 516323 181063 516357
rect 181097 516323 181105 516357
rect 181053 516278 181105 516323
rect 181159 516357 181211 516388
rect 181159 516323 181167 516357
rect 181201 516323 181211 516357
rect 181159 516278 181211 516323
rect 182157 516357 182209 516388
rect 182157 516323 182167 516357
rect 182201 516323 182209 516357
rect 182157 516278 182209 516323
rect 182263 516357 182315 516388
rect 182263 516323 182271 516357
rect 182305 516323 182315 516357
rect 182263 516278 182315 516323
rect 183261 516357 183313 516388
rect 183261 516323 183271 516357
rect 183305 516323 183313 516357
rect 183261 516278 183313 516323
rect 183367 516357 183419 516388
rect 183367 516323 183375 516357
rect 183409 516323 183419 516357
rect 183367 516278 183419 516323
rect 184365 516357 184417 516388
rect 184365 516323 184375 516357
rect 184409 516323 184417 516357
rect 184365 516278 184417 516323
rect 184471 516357 184523 516388
rect 184471 516323 184479 516357
rect 184513 516323 184523 516357
rect 184471 516278 184523 516323
rect 184917 516357 184969 516388
rect 184917 516323 184927 516357
rect 184961 516323 184969 516357
rect 184917 516278 184969 516323
rect 185207 516357 185259 516388
rect 185207 516323 185215 516357
rect 185249 516323 185259 516357
rect 185207 516278 185259 516323
rect 186205 516357 186257 516388
rect 186205 516323 186215 516357
rect 186249 516323 186257 516357
rect 186205 516278 186257 516323
rect 186311 516357 186363 516388
rect 186311 516323 186319 516357
rect 186353 516323 186363 516357
rect 186311 516278 186363 516323
rect 186941 516357 186993 516388
rect 186941 516323 186951 516357
rect 186985 516323 186993 516357
rect 186941 516278 186993 516323
rect 187231 516355 187283 516388
rect 187231 516321 187239 516355
rect 187273 516321 187283 516355
rect 187231 516278 187283 516321
rect 187401 516355 187453 516388
rect 187401 516321 187411 516355
rect 187445 516321 187453 516355
rect 187401 516278 187453 516321
rect 172235 515461 172287 515504
rect 172235 515427 172243 515461
rect 172277 515427 172287 515461
rect 172235 515394 172287 515427
rect 172405 515461 172457 515504
rect 172405 515427 172415 515461
rect 172449 515427 172457 515461
rect 172405 515394 172457 515427
rect 172511 515459 172563 515504
rect 172511 515425 172519 515459
rect 172553 515425 172563 515459
rect 172511 515394 172563 515425
rect 173141 515459 173193 515504
rect 173141 515425 173151 515459
rect 173185 515425 173193 515459
rect 173141 515394 173193 515425
rect 173431 515448 173484 515478
rect 173431 515414 173439 515448
rect 173473 515414 173484 515448
rect 173431 515394 173484 515414
rect 173514 515444 173581 515478
rect 173514 515410 173525 515444
rect 173559 515410 173581 515444
rect 173514 515394 173581 515410
rect 173611 515466 173667 515478
rect 173611 515432 173622 515466
rect 173656 515432 173667 515466
rect 173611 515394 173667 515432
rect 173697 515444 173753 515478
rect 173697 515410 173708 515444
rect 173742 515410 173753 515444
rect 173697 515394 173753 515410
rect 173783 515466 173839 515478
rect 173783 515432 173794 515466
rect 173828 515432 173839 515466
rect 173783 515394 173839 515432
rect 173869 515444 173927 515478
rect 173869 515410 173880 515444
rect 173914 515410 173927 515444
rect 173869 515394 173927 515410
rect 173983 515459 174035 515504
rect 173983 515425 173991 515459
rect 174025 515425 174035 515459
rect 173983 515394 174035 515425
rect 174613 515459 174665 515504
rect 174613 515425 174623 515459
rect 174657 515425 174665 515459
rect 174613 515394 174665 515425
rect 174903 515459 174955 515504
rect 174903 515425 174911 515459
rect 174945 515425 174955 515459
rect 174903 515394 174955 515425
rect 175901 515459 175953 515504
rect 175901 515425 175911 515459
rect 175945 515425 175953 515459
rect 175901 515394 175953 515425
rect 176007 515459 176059 515504
rect 176007 515425 176015 515459
rect 176049 515425 176059 515459
rect 176007 515394 176059 515425
rect 177005 515459 177057 515504
rect 177005 515425 177015 515459
rect 177049 515425 177057 515459
rect 177005 515394 177057 515425
rect 177111 515461 177163 515504
rect 177111 515427 177119 515461
rect 177153 515427 177163 515461
rect 177111 515394 177163 515427
rect 177281 515461 177333 515504
rect 177281 515427 177291 515461
rect 177325 515427 177333 515461
rect 177281 515394 177333 515427
rect 177479 515459 177531 515504
rect 177479 515425 177487 515459
rect 177521 515425 177531 515459
rect 177479 515394 177531 515425
rect 178477 515459 178529 515504
rect 178477 515425 178487 515459
rect 178521 515425 178529 515459
rect 178477 515394 178529 515425
rect 178583 515459 178635 515504
rect 178583 515425 178591 515459
rect 178625 515425 178635 515459
rect 178583 515394 178635 515425
rect 179581 515459 179633 515504
rect 179581 515425 179591 515459
rect 179625 515425 179633 515459
rect 179581 515394 179633 515425
rect 179687 515461 179739 515504
rect 179687 515427 179695 515461
rect 179729 515427 179739 515461
rect 179687 515394 179739 515427
rect 179857 515461 179909 515504
rect 179857 515427 179867 515461
rect 179901 515427 179909 515461
rect 179857 515394 179909 515427
rect 180055 515459 180107 515504
rect 180055 515425 180063 515459
rect 180097 515425 180107 515459
rect 180055 515394 180107 515425
rect 181053 515459 181105 515504
rect 181053 515425 181063 515459
rect 181097 515425 181105 515459
rect 181053 515394 181105 515425
rect 181159 515459 181211 515504
rect 181159 515425 181167 515459
rect 181201 515425 181211 515459
rect 181159 515394 181211 515425
rect 181789 515459 181841 515504
rect 181789 515425 181799 515459
rect 181833 515425 181841 515459
rect 181789 515394 181841 515425
rect 182079 515470 182131 515498
rect 182079 515436 182087 515470
rect 182121 515436 182131 515470
rect 182079 515394 182131 515436
rect 182161 515440 182219 515498
rect 182161 515406 182173 515440
rect 182207 515406 182219 515440
rect 182161 515394 182219 515406
rect 182249 515453 182301 515498
rect 182249 515419 182259 515453
rect 182293 515419 182301 515453
rect 182249 515394 182301 515419
rect 182631 515459 182683 515504
rect 182631 515425 182639 515459
rect 182673 515425 182683 515459
rect 182631 515394 182683 515425
rect 183629 515459 183681 515504
rect 183629 515425 183639 515459
rect 183673 515425 183681 515459
rect 183629 515394 183681 515425
rect 183735 515459 183787 515504
rect 183735 515425 183743 515459
rect 183777 515425 183787 515459
rect 183735 515394 183787 515425
rect 184733 515459 184785 515504
rect 184733 515425 184743 515459
rect 184777 515425 184785 515459
rect 184733 515394 184785 515425
rect 184839 515461 184891 515504
rect 184839 515427 184847 515461
rect 184881 515427 184891 515461
rect 184839 515394 184891 515427
rect 185009 515461 185061 515504
rect 185009 515427 185019 515461
rect 185053 515427 185061 515461
rect 185009 515394 185061 515427
rect 185207 515459 185259 515504
rect 185207 515425 185215 515459
rect 185249 515425 185259 515459
rect 185207 515394 185259 515425
rect 186205 515459 186257 515504
rect 186205 515425 186215 515459
rect 186249 515425 186257 515459
rect 186205 515394 186257 515425
rect 186403 515448 186456 515478
rect 186403 515414 186411 515448
rect 186445 515414 186456 515448
rect 186403 515394 186456 515414
rect 186486 515444 186553 515478
rect 186486 515410 186497 515444
rect 186531 515410 186553 515444
rect 186486 515394 186553 515410
rect 186583 515466 186639 515478
rect 186583 515432 186594 515466
rect 186628 515432 186639 515466
rect 186583 515394 186639 515432
rect 186669 515444 186725 515478
rect 186669 515410 186680 515444
rect 186714 515410 186725 515444
rect 186669 515394 186725 515410
rect 186755 515466 186811 515478
rect 186755 515432 186766 515466
rect 186800 515432 186811 515466
rect 186755 515394 186811 515432
rect 186841 515444 186899 515478
rect 186841 515410 186852 515444
rect 186886 515410 186899 515444
rect 186841 515394 186899 515410
rect 186955 515461 187007 515504
rect 186955 515427 186963 515461
rect 186997 515427 187007 515461
rect 186955 515394 187007 515427
rect 187125 515461 187177 515504
rect 187125 515427 187135 515461
rect 187169 515427 187177 515461
rect 187125 515394 187177 515427
rect 187231 515461 187283 515504
rect 187231 515427 187239 515461
rect 187273 515427 187283 515461
rect 187231 515394 187283 515427
rect 187401 515461 187453 515504
rect 187401 515427 187411 515461
rect 187445 515427 187453 515461
rect 187401 515394 187453 515427
<< pdiff >>
rect 164656 539513 164714 539525
rect 164656 538537 164668 539513
rect 164702 538537 164714 539513
rect 164656 538525 164714 538537
rect 164744 539513 164802 539525
rect 164744 538537 164756 539513
rect 164790 538537 164802 539513
rect 164744 538525 164802 538537
rect 164879 539520 164941 539532
rect 164879 538544 164891 539520
rect 164925 538544 164941 539520
rect 164879 538532 164941 538544
rect 164971 539520 165037 539532
rect 164971 538544 164987 539520
rect 165021 538544 165037 539520
rect 164971 538532 165037 538544
rect 165067 539520 165133 539532
rect 165067 538544 165083 539520
rect 165117 538544 165133 539520
rect 165067 538532 165133 538544
rect 165163 539520 165229 539532
rect 165163 538544 165179 539520
rect 165213 538544 165229 539520
rect 165163 538532 165229 538544
rect 165259 539520 165325 539532
rect 165259 538544 165275 539520
rect 165309 538544 165325 539520
rect 165259 538532 165325 538544
rect 165355 539520 165421 539532
rect 165355 538544 165371 539520
rect 165405 538544 165421 539520
rect 165355 538532 165421 538544
rect 165451 539520 165517 539532
rect 165451 538544 165467 539520
rect 165501 538544 165517 539520
rect 165451 538532 165517 538544
rect 165547 539520 165613 539532
rect 165547 538544 165563 539520
rect 165597 538544 165613 539520
rect 165547 538532 165613 538544
rect 165643 539520 165709 539532
rect 165643 538544 165659 539520
rect 165693 538544 165709 539520
rect 165643 538532 165709 538544
rect 165739 539520 165805 539532
rect 165739 538544 165755 539520
rect 165789 538544 165805 539520
rect 165739 538532 165805 538544
rect 165835 539520 165901 539532
rect 165835 538544 165851 539520
rect 165885 538544 165901 539520
rect 165835 538532 165901 538544
rect 165931 539520 165997 539532
rect 165931 538544 165947 539520
rect 165981 538544 165997 539520
rect 165931 538532 165997 538544
rect 166027 539520 166089 539532
rect 166027 538544 166043 539520
rect 166077 538544 166089 539520
rect 166156 539513 166214 539525
rect 166156 538937 166168 539513
rect 166202 538937 166214 539513
rect 166156 538925 166214 538937
rect 166244 539513 166302 539525
rect 166244 538937 166256 539513
rect 166290 538937 166302 539513
rect 166244 538925 166302 538937
rect 166356 539513 166414 539525
rect 166027 538532 166089 538544
rect 166356 538537 166368 539513
rect 166402 538537 166414 539513
rect 166356 538525 166414 538537
rect 166444 539513 166502 539525
rect 166444 538537 166456 539513
rect 166490 538537 166502 539513
rect 166444 538525 166502 538537
rect 168456 539513 168514 539525
rect 168456 538537 168468 539513
rect 168502 538537 168514 539513
rect 168456 538525 168514 538537
rect 168544 539513 168602 539525
rect 168544 538537 168556 539513
rect 168590 538537 168602 539513
rect 168544 538525 168602 538537
rect 168679 539520 168741 539532
rect 168679 538544 168691 539520
rect 168725 538544 168741 539520
rect 168679 538532 168741 538544
rect 168771 539520 168837 539532
rect 168771 538544 168787 539520
rect 168821 538544 168837 539520
rect 168771 538532 168837 538544
rect 168867 539520 168933 539532
rect 168867 538544 168883 539520
rect 168917 538544 168933 539520
rect 168867 538532 168933 538544
rect 168963 539520 169029 539532
rect 168963 538544 168979 539520
rect 169013 538544 169029 539520
rect 168963 538532 169029 538544
rect 169059 539520 169125 539532
rect 169059 538544 169075 539520
rect 169109 538544 169125 539520
rect 169059 538532 169125 538544
rect 169155 539520 169221 539532
rect 169155 538544 169171 539520
rect 169205 538544 169221 539520
rect 169155 538532 169221 538544
rect 169251 539520 169317 539532
rect 169251 538544 169267 539520
rect 169301 538544 169317 539520
rect 169251 538532 169317 538544
rect 169347 539520 169413 539532
rect 169347 538544 169363 539520
rect 169397 538544 169413 539520
rect 169347 538532 169413 538544
rect 169443 539520 169509 539532
rect 169443 538544 169459 539520
rect 169493 538544 169509 539520
rect 169443 538532 169509 538544
rect 169539 539520 169605 539532
rect 169539 538544 169555 539520
rect 169589 538544 169605 539520
rect 169539 538532 169605 538544
rect 169635 539520 169701 539532
rect 169635 538544 169651 539520
rect 169685 538544 169701 539520
rect 169635 538532 169701 538544
rect 169731 539520 169797 539532
rect 169731 538544 169747 539520
rect 169781 538544 169797 539520
rect 169731 538532 169797 538544
rect 169827 539520 169889 539532
rect 169827 538544 169843 539520
rect 169877 538544 169889 539520
rect 169956 539513 170014 539525
rect 169956 538937 169968 539513
rect 170002 538937 170014 539513
rect 169956 538925 170014 538937
rect 170044 539513 170102 539525
rect 170044 538937 170056 539513
rect 170090 538937 170102 539513
rect 170044 538925 170102 538937
rect 170156 539513 170214 539525
rect 169827 538532 169889 538544
rect 170156 538537 170168 539513
rect 170202 538537 170214 539513
rect 170156 538525 170214 538537
rect 170244 539513 170302 539525
rect 170244 538537 170256 539513
rect 170290 538537 170302 539513
rect 170244 538525 170302 538537
rect 172156 539513 172214 539525
rect 172156 538537 172168 539513
rect 172202 538537 172214 539513
rect 172156 538525 172214 538537
rect 172244 539513 172302 539525
rect 172244 538537 172256 539513
rect 172290 538537 172302 539513
rect 172244 538525 172302 538537
rect 172379 539520 172441 539532
rect 172379 538544 172391 539520
rect 172425 538544 172441 539520
rect 172379 538532 172441 538544
rect 172471 539520 172537 539532
rect 172471 538544 172487 539520
rect 172521 538544 172537 539520
rect 172471 538532 172537 538544
rect 172567 539520 172633 539532
rect 172567 538544 172583 539520
rect 172617 538544 172633 539520
rect 172567 538532 172633 538544
rect 172663 539520 172729 539532
rect 172663 538544 172679 539520
rect 172713 538544 172729 539520
rect 172663 538532 172729 538544
rect 172759 539520 172825 539532
rect 172759 538544 172775 539520
rect 172809 538544 172825 539520
rect 172759 538532 172825 538544
rect 172855 539520 172921 539532
rect 172855 538544 172871 539520
rect 172905 538544 172921 539520
rect 172855 538532 172921 538544
rect 172951 539520 173017 539532
rect 172951 538544 172967 539520
rect 173001 538544 173017 539520
rect 172951 538532 173017 538544
rect 173047 539520 173113 539532
rect 173047 538544 173063 539520
rect 173097 538544 173113 539520
rect 173047 538532 173113 538544
rect 173143 539520 173209 539532
rect 173143 538544 173159 539520
rect 173193 538544 173209 539520
rect 173143 538532 173209 538544
rect 173239 539520 173305 539532
rect 173239 538544 173255 539520
rect 173289 538544 173305 539520
rect 173239 538532 173305 538544
rect 173335 539520 173401 539532
rect 173335 538544 173351 539520
rect 173385 538544 173401 539520
rect 173335 538532 173401 538544
rect 173431 539520 173497 539532
rect 173431 538544 173447 539520
rect 173481 538544 173497 539520
rect 173431 538532 173497 538544
rect 173527 539520 173589 539532
rect 173527 538544 173543 539520
rect 173577 538544 173589 539520
rect 173656 539513 173714 539525
rect 173656 538937 173668 539513
rect 173702 538937 173714 539513
rect 173656 538925 173714 538937
rect 173744 539513 173802 539525
rect 173744 538937 173756 539513
rect 173790 538937 173802 539513
rect 173744 538925 173802 538937
rect 173856 539513 173914 539525
rect 173527 538532 173589 538544
rect 173856 538537 173868 539513
rect 173902 538537 173914 539513
rect 173856 538525 173914 538537
rect 173944 539513 174002 539525
rect 173944 538537 173956 539513
rect 173990 538537 174002 539513
rect 173944 538525 174002 538537
rect 175656 539513 175714 539525
rect 175656 538537 175668 539513
rect 175702 538537 175714 539513
rect 175656 538525 175714 538537
rect 175744 539513 175802 539525
rect 175744 538537 175756 539513
rect 175790 538537 175802 539513
rect 175744 538525 175802 538537
rect 175879 539520 175941 539532
rect 175879 538544 175891 539520
rect 175925 538544 175941 539520
rect 175879 538532 175941 538544
rect 175971 539520 176037 539532
rect 175971 538544 175987 539520
rect 176021 538544 176037 539520
rect 175971 538532 176037 538544
rect 176067 539520 176133 539532
rect 176067 538544 176083 539520
rect 176117 538544 176133 539520
rect 176067 538532 176133 538544
rect 176163 539520 176229 539532
rect 176163 538544 176179 539520
rect 176213 538544 176229 539520
rect 176163 538532 176229 538544
rect 176259 539520 176325 539532
rect 176259 538544 176275 539520
rect 176309 538544 176325 539520
rect 176259 538532 176325 538544
rect 176355 539520 176421 539532
rect 176355 538544 176371 539520
rect 176405 538544 176421 539520
rect 176355 538532 176421 538544
rect 176451 539520 176517 539532
rect 176451 538544 176467 539520
rect 176501 538544 176517 539520
rect 176451 538532 176517 538544
rect 176547 539520 176613 539532
rect 176547 538544 176563 539520
rect 176597 538544 176613 539520
rect 176547 538532 176613 538544
rect 176643 539520 176709 539532
rect 176643 538544 176659 539520
rect 176693 538544 176709 539520
rect 176643 538532 176709 538544
rect 176739 539520 176805 539532
rect 176739 538544 176755 539520
rect 176789 538544 176805 539520
rect 176739 538532 176805 538544
rect 176835 539520 176901 539532
rect 176835 538544 176851 539520
rect 176885 538544 176901 539520
rect 176835 538532 176901 538544
rect 176931 539520 176997 539532
rect 176931 538544 176947 539520
rect 176981 538544 176997 539520
rect 176931 538532 176997 538544
rect 177027 539520 177089 539532
rect 177027 538544 177043 539520
rect 177077 538544 177089 539520
rect 177156 539513 177214 539525
rect 177156 538937 177168 539513
rect 177202 538937 177214 539513
rect 177156 538925 177214 538937
rect 177244 539513 177302 539525
rect 177244 538937 177256 539513
rect 177290 538937 177302 539513
rect 177244 538925 177302 538937
rect 177356 539513 177414 539525
rect 177027 538532 177089 538544
rect 177356 538537 177368 539513
rect 177402 538537 177414 539513
rect 177356 538525 177414 538537
rect 177444 539513 177502 539525
rect 177444 538537 177456 539513
rect 177490 538537 177502 539513
rect 177444 538525 177502 538537
rect 179256 539513 179314 539525
rect 179256 538537 179268 539513
rect 179302 538537 179314 539513
rect 179256 538525 179314 538537
rect 179344 539513 179402 539525
rect 179344 538537 179356 539513
rect 179390 538537 179402 539513
rect 179344 538525 179402 538537
rect 179479 539520 179541 539532
rect 179479 538544 179491 539520
rect 179525 538544 179541 539520
rect 179479 538532 179541 538544
rect 179571 539520 179637 539532
rect 179571 538544 179587 539520
rect 179621 538544 179637 539520
rect 179571 538532 179637 538544
rect 179667 539520 179733 539532
rect 179667 538544 179683 539520
rect 179717 538544 179733 539520
rect 179667 538532 179733 538544
rect 179763 539520 179829 539532
rect 179763 538544 179779 539520
rect 179813 538544 179829 539520
rect 179763 538532 179829 538544
rect 179859 539520 179925 539532
rect 179859 538544 179875 539520
rect 179909 538544 179925 539520
rect 179859 538532 179925 538544
rect 179955 539520 180021 539532
rect 179955 538544 179971 539520
rect 180005 538544 180021 539520
rect 179955 538532 180021 538544
rect 180051 539520 180117 539532
rect 180051 538544 180067 539520
rect 180101 538544 180117 539520
rect 180051 538532 180117 538544
rect 180147 539520 180213 539532
rect 180147 538544 180163 539520
rect 180197 538544 180213 539520
rect 180147 538532 180213 538544
rect 180243 539520 180309 539532
rect 180243 538544 180259 539520
rect 180293 538544 180309 539520
rect 180243 538532 180309 538544
rect 180339 539520 180405 539532
rect 180339 538544 180355 539520
rect 180389 538544 180405 539520
rect 180339 538532 180405 538544
rect 180435 539520 180501 539532
rect 180435 538544 180451 539520
rect 180485 538544 180501 539520
rect 180435 538532 180501 538544
rect 180531 539520 180597 539532
rect 180531 538544 180547 539520
rect 180581 538544 180597 539520
rect 180531 538532 180597 538544
rect 180627 539520 180689 539532
rect 180627 538544 180643 539520
rect 180677 538544 180689 539520
rect 180756 539513 180814 539525
rect 180756 538937 180768 539513
rect 180802 538937 180814 539513
rect 180756 538925 180814 538937
rect 180844 539513 180902 539525
rect 180844 538937 180856 539513
rect 180890 538937 180902 539513
rect 180844 538925 180902 538937
rect 180956 539513 181014 539525
rect 180627 538532 180689 538544
rect 180956 538537 180968 539513
rect 181002 538537 181014 539513
rect 180956 538525 181014 538537
rect 181044 539513 181102 539525
rect 181044 538537 181056 539513
rect 181090 538537 181102 539513
rect 181044 538525 181102 538537
rect 182556 539513 182614 539525
rect 182556 538537 182568 539513
rect 182602 538537 182614 539513
rect 182556 538525 182614 538537
rect 182644 539513 182702 539525
rect 182644 538537 182656 539513
rect 182690 538537 182702 539513
rect 182644 538525 182702 538537
rect 182779 539520 182841 539532
rect 182779 538544 182791 539520
rect 182825 538544 182841 539520
rect 182779 538532 182841 538544
rect 182871 539520 182937 539532
rect 182871 538544 182887 539520
rect 182921 538544 182937 539520
rect 182871 538532 182937 538544
rect 182967 539520 183033 539532
rect 182967 538544 182983 539520
rect 183017 538544 183033 539520
rect 182967 538532 183033 538544
rect 183063 539520 183129 539532
rect 183063 538544 183079 539520
rect 183113 538544 183129 539520
rect 183063 538532 183129 538544
rect 183159 539520 183225 539532
rect 183159 538544 183175 539520
rect 183209 538544 183225 539520
rect 183159 538532 183225 538544
rect 183255 539520 183321 539532
rect 183255 538544 183271 539520
rect 183305 538544 183321 539520
rect 183255 538532 183321 538544
rect 183351 539520 183417 539532
rect 183351 538544 183367 539520
rect 183401 538544 183417 539520
rect 183351 538532 183417 538544
rect 183447 539520 183513 539532
rect 183447 538544 183463 539520
rect 183497 538544 183513 539520
rect 183447 538532 183513 538544
rect 183543 539520 183609 539532
rect 183543 538544 183559 539520
rect 183593 538544 183609 539520
rect 183543 538532 183609 538544
rect 183639 539520 183705 539532
rect 183639 538544 183655 539520
rect 183689 538544 183705 539520
rect 183639 538532 183705 538544
rect 183735 539520 183801 539532
rect 183735 538544 183751 539520
rect 183785 538544 183801 539520
rect 183735 538532 183801 538544
rect 183831 539520 183897 539532
rect 183831 538544 183847 539520
rect 183881 538544 183897 539520
rect 183831 538532 183897 538544
rect 183927 539520 183989 539532
rect 183927 538544 183943 539520
rect 183977 538544 183989 539520
rect 184056 539513 184114 539525
rect 184056 538937 184068 539513
rect 184102 538937 184114 539513
rect 184056 538925 184114 538937
rect 184144 539513 184202 539525
rect 184144 538937 184156 539513
rect 184190 538937 184202 539513
rect 184144 538925 184202 538937
rect 184256 539513 184314 539525
rect 183927 538532 183989 538544
rect 184256 538537 184268 539513
rect 184302 538537 184314 539513
rect 184256 538525 184314 538537
rect 184344 539513 184402 539525
rect 184344 538537 184356 539513
rect 184390 538537 184402 539513
rect 184344 538525 184402 538537
rect 185856 539513 185914 539525
rect 185856 538537 185868 539513
rect 185902 538537 185914 539513
rect 185856 538525 185914 538537
rect 185944 539513 186002 539525
rect 185944 538537 185956 539513
rect 185990 538537 186002 539513
rect 185944 538525 186002 538537
rect 186079 539520 186141 539532
rect 186079 538544 186091 539520
rect 186125 538544 186141 539520
rect 186079 538532 186141 538544
rect 186171 539520 186237 539532
rect 186171 538544 186187 539520
rect 186221 538544 186237 539520
rect 186171 538532 186237 538544
rect 186267 539520 186333 539532
rect 186267 538544 186283 539520
rect 186317 538544 186333 539520
rect 186267 538532 186333 538544
rect 186363 539520 186429 539532
rect 186363 538544 186379 539520
rect 186413 538544 186429 539520
rect 186363 538532 186429 538544
rect 186459 539520 186525 539532
rect 186459 538544 186475 539520
rect 186509 538544 186525 539520
rect 186459 538532 186525 538544
rect 186555 539520 186621 539532
rect 186555 538544 186571 539520
rect 186605 538544 186621 539520
rect 186555 538532 186621 538544
rect 186651 539520 186717 539532
rect 186651 538544 186667 539520
rect 186701 538544 186717 539520
rect 186651 538532 186717 538544
rect 186747 539520 186813 539532
rect 186747 538544 186763 539520
rect 186797 538544 186813 539520
rect 186747 538532 186813 538544
rect 186843 539520 186909 539532
rect 186843 538544 186859 539520
rect 186893 538544 186909 539520
rect 186843 538532 186909 538544
rect 186939 539520 187005 539532
rect 186939 538544 186955 539520
rect 186989 538544 187005 539520
rect 186939 538532 187005 538544
rect 187035 539520 187101 539532
rect 187035 538544 187051 539520
rect 187085 538544 187101 539520
rect 187035 538532 187101 538544
rect 187131 539520 187197 539532
rect 187131 538544 187147 539520
rect 187181 538544 187197 539520
rect 187131 538532 187197 538544
rect 187227 539520 187289 539532
rect 187227 538544 187243 539520
rect 187277 538544 187289 539520
rect 187356 539513 187414 539525
rect 187356 538937 187368 539513
rect 187402 538937 187414 539513
rect 187356 538925 187414 538937
rect 187444 539513 187502 539525
rect 187444 538937 187456 539513
rect 187490 538937 187502 539513
rect 187444 538925 187502 538937
rect 187556 539513 187614 539525
rect 187227 538532 187289 538544
rect 187556 538537 187568 539513
rect 187602 538537 187614 539513
rect 187556 538525 187614 538537
rect 187644 539513 187702 539525
rect 187644 538537 187656 539513
rect 187690 538537 187702 539513
rect 187644 538525 187702 538537
rect 189156 539513 189214 539525
rect 189156 538537 189168 539513
rect 189202 538537 189214 539513
rect 189156 538525 189214 538537
rect 189244 539513 189302 539525
rect 189244 538537 189256 539513
rect 189290 538537 189302 539513
rect 189244 538525 189302 538537
rect 189379 539520 189441 539532
rect 189379 538544 189391 539520
rect 189425 538544 189441 539520
rect 189379 538532 189441 538544
rect 189471 539520 189537 539532
rect 189471 538544 189487 539520
rect 189521 538544 189537 539520
rect 189471 538532 189537 538544
rect 189567 539520 189633 539532
rect 189567 538544 189583 539520
rect 189617 538544 189633 539520
rect 189567 538532 189633 538544
rect 189663 539520 189729 539532
rect 189663 538544 189679 539520
rect 189713 538544 189729 539520
rect 189663 538532 189729 538544
rect 189759 539520 189825 539532
rect 189759 538544 189775 539520
rect 189809 538544 189825 539520
rect 189759 538532 189825 538544
rect 189855 539520 189921 539532
rect 189855 538544 189871 539520
rect 189905 538544 189921 539520
rect 189855 538532 189921 538544
rect 189951 539520 190017 539532
rect 189951 538544 189967 539520
rect 190001 538544 190017 539520
rect 189951 538532 190017 538544
rect 190047 539520 190113 539532
rect 190047 538544 190063 539520
rect 190097 538544 190113 539520
rect 190047 538532 190113 538544
rect 190143 539520 190209 539532
rect 190143 538544 190159 539520
rect 190193 538544 190209 539520
rect 190143 538532 190209 538544
rect 190239 539520 190305 539532
rect 190239 538544 190255 539520
rect 190289 538544 190305 539520
rect 190239 538532 190305 538544
rect 190335 539520 190401 539532
rect 190335 538544 190351 539520
rect 190385 538544 190401 539520
rect 190335 538532 190401 538544
rect 190431 539520 190497 539532
rect 190431 538544 190447 539520
rect 190481 538544 190497 539520
rect 190431 538532 190497 538544
rect 190527 539520 190589 539532
rect 190527 538544 190543 539520
rect 190577 538544 190589 539520
rect 190656 539513 190714 539525
rect 190656 538937 190668 539513
rect 190702 538937 190714 539513
rect 190656 538925 190714 538937
rect 190744 539513 190802 539525
rect 190744 538937 190756 539513
rect 190790 538937 190802 539513
rect 190744 538925 190802 538937
rect 190856 539513 190914 539525
rect 190527 538532 190589 538544
rect 190856 538537 190868 539513
rect 190902 538537 190914 539513
rect 190856 538525 190914 538537
rect 190944 539513 191002 539525
rect 190944 538537 190956 539513
rect 190990 538537 191002 539513
rect 190944 538525 191002 538537
rect 161246 537613 161304 537625
rect 161246 537037 161258 537613
rect 161292 537037 161304 537613
rect 161246 537025 161304 537037
rect 161334 537613 161392 537625
rect 161334 537037 161346 537613
rect 161380 537037 161392 537613
rect 161334 537025 161392 537037
rect 161446 537613 161508 537625
rect 161446 537037 161458 537613
rect 161492 537037 161508 537613
rect 161446 537025 161508 537037
rect 161538 537613 161604 537625
rect 161538 537037 161554 537613
rect 161588 537037 161604 537613
rect 161538 537025 161604 537037
rect 161634 537613 161700 537625
rect 161634 537037 161650 537613
rect 161684 537037 161700 537613
rect 161634 537025 161700 537037
rect 161730 537613 161792 537625
rect 161730 537037 161746 537613
rect 161780 537037 161792 537613
rect 161730 537025 161792 537037
rect 161846 537613 161908 537625
rect 161846 537037 161858 537613
rect 161892 537037 161908 537613
rect 161846 537025 161908 537037
rect 161938 537613 162004 537625
rect 161938 537037 161954 537613
rect 161988 537037 162004 537613
rect 161938 537025 162004 537037
rect 162034 537613 162100 537625
rect 162034 537037 162050 537613
rect 162084 537037 162100 537613
rect 162034 537025 162100 537037
rect 162130 537613 162192 537625
rect 162130 537037 162146 537613
rect 162180 537037 162192 537613
rect 162130 537025 162192 537037
rect 162266 537613 162324 537625
rect 162266 537037 162278 537613
rect 162312 537037 162324 537613
rect 162266 537025 162324 537037
rect 162354 537613 162412 537625
rect 162354 537037 162366 537613
rect 162400 537037 162412 537613
rect 162354 537025 162412 537037
rect 157736 536593 157794 536605
rect 157736 536017 157748 536593
rect 157782 536017 157794 536593
rect 157736 536005 157794 536017
rect 157994 536593 158052 536605
rect 157994 536017 158006 536593
rect 158040 536017 158052 536593
rect 157994 536005 158052 536017
rect 158114 536593 158172 536605
rect 158114 536017 158126 536593
rect 158160 536017 158172 536593
rect 158114 536005 158172 536017
rect 158372 536593 158430 536605
rect 158372 536017 158384 536593
rect 158418 536017 158430 536593
rect 158372 536005 158430 536017
rect 158630 536593 158688 536605
rect 158630 536017 158642 536593
rect 158676 536017 158688 536593
rect 158630 536005 158688 536017
rect 158888 536593 158946 536605
rect 158888 536017 158900 536593
rect 158934 536017 158946 536593
rect 158888 536005 158946 536017
rect 159146 536593 159204 536605
rect 159146 536017 159158 536593
rect 159192 536017 159204 536593
rect 159146 536005 159204 536017
rect 159404 536593 159462 536605
rect 159404 536017 159416 536593
rect 159450 536017 159462 536593
rect 159404 536005 159462 536017
rect 159662 536593 159720 536605
rect 159662 536017 159674 536593
rect 159708 536017 159720 536593
rect 159662 536005 159720 536017
rect 159920 536593 159978 536605
rect 159920 536017 159932 536593
rect 159966 536017 159978 536593
rect 159920 536005 159978 536017
rect 160178 536593 160236 536605
rect 160178 536017 160190 536593
rect 160224 536017 160236 536593
rect 160178 536005 160236 536017
rect 160436 536593 160494 536605
rect 160436 536017 160448 536593
rect 160482 536017 160494 536593
rect 160436 536005 160494 536017
rect 160694 536593 160752 536605
rect 160694 536017 160706 536593
rect 160740 536017 160752 536593
rect 160694 536005 160752 536017
rect 160820 536593 160878 536605
rect 160820 536017 160832 536593
rect 160866 536017 160878 536593
rect 160820 536005 160878 536017
rect 161078 536593 161136 536605
rect 161078 536017 161090 536593
rect 161124 536017 161136 536593
rect 161078 536005 161136 536017
rect 161336 536593 161394 536605
rect 161336 536017 161348 536593
rect 161382 536017 161394 536593
rect 161336 536005 161394 536017
rect 161594 536593 161652 536605
rect 161594 536017 161606 536593
rect 161640 536017 161652 536593
rect 161594 536005 161652 536017
rect 161718 536593 161776 536605
rect 161718 536017 161730 536593
rect 161764 536017 161776 536593
rect 161718 536005 161776 536017
rect 161976 536593 162034 536605
rect 161976 536017 161988 536593
rect 162022 536017 162034 536593
rect 161976 536005 162034 536017
rect 162234 536593 162292 536605
rect 162234 536017 162246 536593
rect 162280 536017 162292 536593
rect 162234 536005 162292 536017
rect 162356 536593 162414 536605
rect 162356 536017 162368 536593
rect 162402 536017 162414 536593
rect 162356 536005 162414 536017
rect 162614 536593 162672 536605
rect 162614 536017 162626 536593
rect 162660 536017 162672 536593
rect 162614 536005 162672 536017
rect 172235 530223 172287 530256
rect 172235 530189 172243 530223
rect 172277 530189 172287 530223
rect 172235 530128 172287 530189
rect 172235 530094 172243 530128
rect 172277 530094 172287 530128
rect 172235 530082 172287 530094
rect 172405 530223 172457 530256
rect 172405 530189 172415 530223
rect 172449 530189 172457 530223
rect 172405 530128 172457 530189
rect 172405 530094 172415 530128
rect 172449 530094 172457 530128
rect 172405 530082 172457 530094
rect 172512 530210 172572 530282
rect 172512 530176 172527 530210
rect 172561 530176 172572 530210
rect 172512 530142 172572 530176
rect 172512 530108 172527 530142
rect 172561 530108 172572 530142
rect 172512 530082 172572 530108
rect 172602 530272 172658 530282
rect 172602 530238 172613 530272
rect 172647 530238 172658 530272
rect 172602 530204 172658 530238
rect 172602 530170 172613 530204
rect 172647 530170 172658 530204
rect 172602 530136 172658 530170
rect 172602 530102 172613 530136
rect 172647 530102 172658 530136
rect 172602 530082 172658 530102
rect 172688 530128 172744 530282
rect 172688 530094 172699 530128
rect 172733 530094 172744 530128
rect 172688 530082 172744 530094
rect 172774 530163 172830 530282
rect 172774 530129 172785 530163
rect 172819 530129 172830 530163
rect 172774 530082 172830 530129
rect 172860 530196 172926 530282
rect 172860 530162 172881 530196
rect 172915 530162 172926 530196
rect 172860 530128 172926 530162
rect 172860 530094 172881 530128
rect 172915 530094 172926 530128
rect 172860 530082 172926 530094
rect 172956 530258 173009 530282
rect 172956 530224 172967 530258
rect 173001 530224 173009 530258
rect 172956 530136 173009 530224
rect 172956 530102 172967 530136
rect 173001 530102 173009 530136
rect 172956 530082 173009 530102
rect 173063 530128 173115 530256
rect 173063 530094 173071 530128
rect 173105 530094 173115 530128
rect 173063 530082 173115 530094
rect 174061 530128 174113 530256
rect 174061 530094 174071 530128
rect 174105 530094 174113 530128
rect 174061 530082 174113 530094
rect 174167 530230 174219 530256
rect 174167 530196 174175 530230
rect 174209 530196 174219 530230
rect 174167 530128 174219 530196
rect 174167 530094 174175 530128
rect 174209 530094 174219 530128
rect 174167 530082 174219 530094
rect 174613 530230 174665 530256
rect 174613 530196 174623 530230
rect 174657 530196 174665 530230
rect 174613 530128 174665 530196
rect 174613 530094 174623 530128
rect 174657 530094 174665 530128
rect 174904 530210 174964 530282
rect 174904 530176 174919 530210
rect 174953 530176 174964 530210
rect 174904 530142 174964 530176
rect 174904 530108 174919 530142
rect 174953 530108 174964 530142
rect 174613 530082 174665 530094
rect 174904 530082 174964 530108
rect 174994 530272 175050 530282
rect 174994 530238 175005 530272
rect 175039 530238 175050 530272
rect 174994 530204 175050 530238
rect 174994 530170 175005 530204
rect 175039 530170 175050 530204
rect 174994 530136 175050 530170
rect 174994 530102 175005 530136
rect 175039 530102 175050 530136
rect 174994 530082 175050 530102
rect 175080 530128 175136 530282
rect 175080 530094 175091 530128
rect 175125 530094 175136 530128
rect 175080 530082 175136 530094
rect 175166 530163 175222 530282
rect 175166 530129 175177 530163
rect 175211 530129 175222 530163
rect 175166 530082 175222 530129
rect 175252 530196 175318 530282
rect 175252 530162 175273 530196
rect 175307 530162 175318 530196
rect 175252 530128 175318 530162
rect 175252 530094 175273 530128
rect 175307 530094 175318 530128
rect 175252 530082 175318 530094
rect 175348 530258 175401 530282
rect 175348 530224 175359 530258
rect 175393 530224 175401 530258
rect 175348 530136 175401 530224
rect 175348 530102 175359 530136
rect 175393 530102 175401 530136
rect 175348 530082 175401 530102
rect 175547 530232 175599 530282
rect 175547 530198 175555 530232
rect 175589 530198 175599 530232
rect 175547 530164 175599 530198
rect 175547 530130 175555 530164
rect 175589 530130 175599 530164
rect 175547 530082 175599 530130
rect 175629 530210 175679 530282
rect 175629 530196 175695 530210
rect 175629 530162 175639 530196
rect 175673 530162 175695 530196
rect 176221 530166 176275 530250
rect 175629 530128 175695 530162
rect 175629 530094 175639 530128
rect 175673 530094 175695 530128
rect 175629 530082 175695 530094
rect 175760 530128 175814 530166
rect 175760 530094 175768 530128
rect 175802 530094 175814 530128
rect 175760 530082 175814 530094
rect 175844 530154 175898 530166
rect 175844 530120 175854 530154
rect 175888 530120 175898 530154
rect 175844 530082 175898 530120
rect 175928 530128 176006 530166
rect 175928 530094 175938 530128
rect 175972 530094 176006 530128
rect 175928 530082 176006 530094
rect 176036 530082 176090 530166
rect 176120 530129 176176 530166
rect 176120 530095 176130 530129
rect 176164 530095 176176 530129
rect 176120 530082 176176 530095
rect 176206 530136 176275 530166
rect 176206 530102 176227 530136
rect 176261 530102 176275 530136
rect 176206 530082 176275 530102
rect 176305 530128 176357 530250
rect 177115 530204 177167 530216
rect 177115 530170 177123 530204
rect 177157 530170 177167 530204
rect 176305 530094 176315 530128
rect 176349 530094 176357 530128
rect 176305 530082 176357 530094
rect 176420 530154 176472 530166
rect 176420 530120 176428 530154
rect 176462 530120 176472 530154
rect 176420 530082 176472 530120
rect 176502 530138 176569 530166
rect 176502 530104 176512 530138
rect 176546 530104 176569 530138
rect 176502 530082 176569 530104
rect 176599 530154 176709 530166
rect 176599 530120 176609 530154
rect 176643 530120 176709 530154
rect 176599 530082 176709 530120
rect 176739 530130 176808 530166
rect 176739 530096 176763 530130
rect 176797 530096 176808 530130
rect 176739 530082 176808 530096
rect 176838 530136 176900 530166
rect 176838 530102 176856 530136
rect 176890 530102 176900 530136
rect 176838 530082 176900 530102
rect 176930 530128 176982 530166
rect 176930 530094 176940 530128
rect 176974 530094 176982 530128
rect 176930 530082 176982 530094
rect 177115 530136 177167 530170
rect 177115 530102 177123 530136
rect 177157 530102 177167 530136
rect 177115 530088 177167 530102
rect 177197 530152 177251 530216
rect 177197 530118 177207 530152
rect 177241 530118 177251 530152
rect 177197 530088 177251 530118
rect 177281 530204 177333 530216
rect 177281 530170 177291 530204
rect 177325 530170 177333 530204
rect 177281 530136 177333 530170
rect 177281 530102 177291 530136
rect 177325 530102 177333 530136
rect 177281 530088 177333 530102
rect 177682 530154 177734 530282
rect 177682 530120 177690 530154
rect 177724 530120 177734 530154
rect 177682 530082 177734 530120
rect 177764 530166 177814 530282
rect 178399 530217 178451 530240
rect 178399 530183 178407 530217
rect 178441 530183 178451 530217
rect 177764 530128 177829 530166
rect 177764 530094 177780 530128
rect 177814 530094 177829 530128
rect 177764 530082 177829 530094
rect 177929 530154 177981 530166
rect 177929 530120 177939 530154
rect 177973 530120 177981 530154
rect 177929 530082 177981 530120
rect 178035 530154 178087 530166
rect 178035 530120 178043 530154
rect 178077 530120 178087 530154
rect 178035 530082 178087 530120
rect 178187 530128 178241 530166
rect 178187 530094 178197 530128
rect 178231 530094 178241 530128
rect 178187 530082 178241 530094
rect 178271 530154 178323 530166
rect 178271 530120 178281 530154
rect 178315 530120 178323 530154
rect 178271 530082 178323 530120
rect 178399 530136 178451 530183
rect 178399 530102 178407 530136
rect 178441 530102 178451 530136
rect 178399 530082 178451 530102
rect 178481 530204 178539 530240
rect 178481 530170 178493 530204
rect 178527 530170 178539 530204
rect 178481 530136 178539 530170
rect 178481 530102 178493 530136
rect 178527 530102 178539 530136
rect 178481 530082 178539 530102
rect 178569 530204 178621 530240
rect 178569 530170 178579 530204
rect 178613 530170 178621 530204
rect 178569 530136 178621 530170
rect 178569 530102 178579 530136
rect 178613 530102 178621 530136
rect 178569 530082 178621 530102
rect 178676 530210 178736 530282
rect 178676 530176 178691 530210
rect 178725 530176 178736 530210
rect 178676 530142 178736 530176
rect 178676 530108 178691 530142
rect 178725 530108 178736 530142
rect 178676 530082 178736 530108
rect 178766 530272 178822 530282
rect 178766 530238 178777 530272
rect 178811 530238 178822 530272
rect 178766 530204 178822 530238
rect 178766 530170 178777 530204
rect 178811 530170 178822 530204
rect 178766 530136 178822 530170
rect 178766 530102 178777 530136
rect 178811 530102 178822 530136
rect 178766 530082 178822 530102
rect 178852 530128 178908 530282
rect 178852 530094 178863 530128
rect 178897 530094 178908 530128
rect 178852 530082 178908 530094
rect 178938 530163 178994 530282
rect 178938 530129 178949 530163
rect 178983 530129 178994 530163
rect 178938 530082 178994 530129
rect 179024 530196 179090 530282
rect 179024 530162 179045 530196
rect 179079 530162 179090 530196
rect 179024 530128 179090 530162
rect 179024 530094 179045 530128
rect 179079 530094 179090 530128
rect 179024 530082 179090 530094
rect 179120 530258 179173 530282
rect 179120 530224 179131 530258
rect 179165 530224 179173 530258
rect 179120 530136 179173 530224
rect 179120 530102 179131 530136
rect 179165 530102 179173 530136
rect 179120 530082 179173 530102
rect 179227 530258 179280 530282
rect 179227 530224 179235 530258
rect 179269 530224 179280 530258
rect 179227 530136 179280 530224
rect 179227 530102 179235 530136
rect 179269 530102 179280 530136
rect 179227 530082 179280 530102
rect 179310 530196 179376 530282
rect 179310 530162 179321 530196
rect 179355 530162 179376 530196
rect 179310 530128 179376 530162
rect 179310 530094 179321 530128
rect 179355 530094 179376 530128
rect 179310 530082 179376 530094
rect 179406 530163 179462 530282
rect 179406 530129 179417 530163
rect 179451 530129 179462 530163
rect 179406 530082 179462 530129
rect 179492 530128 179548 530282
rect 179492 530094 179503 530128
rect 179537 530094 179548 530128
rect 179492 530082 179548 530094
rect 179578 530272 179634 530282
rect 179578 530238 179589 530272
rect 179623 530238 179634 530272
rect 179578 530204 179634 530238
rect 179578 530170 179589 530204
rect 179623 530170 179634 530204
rect 179578 530136 179634 530170
rect 179578 530102 179589 530136
rect 179623 530102 179634 530136
rect 179578 530082 179634 530102
rect 179664 530210 179724 530282
rect 179664 530176 179675 530210
rect 179709 530176 179724 530210
rect 179664 530142 179724 530176
rect 179664 530108 179675 530142
rect 179709 530108 179724 530142
rect 179664 530082 179724 530108
rect 180239 530264 180291 530282
rect 180239 530230 180247 530264
rect 180281 530230 180291 530264
rect 180239 530196 180291 530230
rect 180239 530162 180247 530196
rect 180281 530162 180291 530196
rect 180239 530128 180291 530162
rect 180239 530094 180247 530128
rect 180281 530094 180291 530128
rect 180239 530082 180291 530094
rect 180321 530264 180373 530282
rect 180321 530230 180331 530264
rect 180365 530230 180373 530264
rect 180321 530205 180373 530230
rect 181799 530264 181851 530282
rect 181799 530230 181807 530264
rect 181841 530230 181851 530264
rect 181799 530205 181851 530230
rect 180321 530196 180400 530205
rect 180321 530162 180331 530196
rect 180365 530162 180400 530196
rect 180321 530128 180400 530162
rect 180321 530094 180331 530128
rect 180365 530121 180400 530128
rect 180430 530121 180503 530205
rect 180533 530188 180717 530205
rect 180533 530154 180567 530188
rect 180601 530154 180642 530188
rect 180676 530154 180717 530188
rect 180533 530121 180717 530154
rect 180747 530121 180789 530205
rect 180819 530188 180885 530205
rect 180819 530154 180839 530188
rect 180873 530154 180885 530188
rect 180819 530121 180885 530154
rect 180915 530188 180971 530205
rect 180915 530154 180925 530188
rect 180959 530154 180971 530188
rect 180915 530121 180971 530154
rect 181201 530188 181257 530205
rect 181201 530154 181213 530188
rect 181247 530154 181257 530188
rect 181201 530121 181257 530154
rect 181287 530188 181353 530205
rect 181287 530154 181299 530188
rect 181333 530154 181353 530188
rect 181287 530121 181353 530154
rect 181383 530121 181425 530205
rect 181455 530188 181639 530205
rect 181455 530154 181496 530188
rect 181530 530154 181571 530188
rect 181605 530154 181639 530188
rect 181455 530121 181639 530154
rect 181669 530121 181742 530205
rect 181772 530196 181851 530205
rect 181772 530162 181807 530196
rect 181841 530162 181851 530196
rect 181772 530128 181851 530162
rect 181772 530121 181807 530128
rect 180365 530094 180373 530121
rect 180321 530082 180373 530094
rect 181799 530094 181807 530121
rect 181841 530094 181851 530128
rect 181799 530082 181851 530094
rect 181881 530264 181933 530282
rect 181881 530230 181891 530264
rect 181925 530230 181933 530264
rect 181881 530196 181933 530230
rect 181881 530162 181891 530196
rect 181925 530162 181933 530196
rect 181881 530128 181933 530162
rect 181881 530094 181891 530128
rect 181925 530094 181933 530128
rect 181881 530082 181933 530094
rect 181987 530258 182040 530282
rect 181987 530224 181995 530258
rect 182029 530224 182040 530258
rect 181987 530136 182040 530224
rect 181987 530102 181995 530136
rect 182029 530102 182040 530136
rect 181987 530082 182040 530102
rect 182070 530196 182136 530282
rect 182070 530162 182081 530196
rect 182115 530162 182136 530196
rect 182070 530128 182136 530162
rect 182070 530094 182081 530128
rect 182115 530094 182136 530128
rect 182070 530082 182136 530094
rect 182166 530163 182222 530282
rect 182166 530129 182177 530163
rect 182211 530129 182222 530163
rect 182166 530082 182222 530129
rect 182252 530128 182308 530282
rect 182252 530094 182263 530128
rect 182297 530094 182308 530128
rect 182252 530082 182308 530094
rect 182338 530272 182394 530282
rect 182338 530238 182349 530272
rect 182383 530238 182394 530272
rect 182338 530204 182394 530238
rect 182338 530170 182349 530204
rect 182383 530170 182394 530204
rect 182338 530136 182394 530170
rect 182338 530102 182349 530136
rect 182383 530102 182394 530136
rect 182338 530082 182394 530102
rect 182424 530210 182484 530282
rect 182424 530176 182435 530210
rect 182469 530176 182484 530210
rect 182424 530142 182484 530176
rect 182424 530108 182435 530142
rect 182469 530108 182484 530142
rect 182424 530082 182484 530108
rect 183091 530258 183144 530282
rect 182631 530230 182683 530256
rect 182631 530196 182639 530230
rect 182673 530196 182683 530230
rect 182631 530128 182683 530196
rect 182631 530094 182639 530128
rect 182673 530094 182683 530128
rect 182631 530082 182683 530094
rect 182893 530230 182945 530256
rect 182893 530196 182903 530230
rect 182937 530196 182945 530230
rect 182893 530128 182945 530196
rect 182893 530094 182903 530128
rect 182937 530094 182945 530128
rect 182893 530082 182945 530094
rect 183091 530224 183099 530258
rect 183133 530224 183144 530258
rect 183091 530136 183144 530224
rect 183091 530102 183099 530136
rect 183133 530102 183144 530136
rect 183091 530082 183144 530102
rect 183174 530196 183240 530282
rect 183174 530162 183185 530196
rect 183219 530162 183240 530196
rect 183174 530128 183240 530162
rect 183174 530094 183185 530128
rect 183219 530094 183240 530128
rect 183174 530082 183240 530094
rect 183270 530163 183326 530282
rect 183270 530129 183281 530163
rect 183315 530129 183326 530163
rect 183270 530082 183326 530129
rect 183356 530128 183412 530282
rect 183356 530094 183367 530128
rect 183401 530094 183412 530128
rect 183356 530082 183412 530094
rect 183442 530272 183498 530282
rect 183442 530238 183453 530272
rect 183487 530238 183498 530272
rect 183442 530204 183498 530238
rect 183442 530170 183453 530204
rect 183487 530170 183498 530204
rect 183442 530136 183498 530170
rect 183442 530102 183453 530136
rect 183487 530102 183498 530136
rect 183442 530082 183498 530102
rect 183528 530210 183588 530282
rect 183528 530176 183539 530210
rect 183573 530176 183588 530210
rect 183528 530142 183588 530176
rect 183528 530108 183539 530142
rect 183573 530108 183588 530142
rect 183528 530082 183588 530108
rect 183643 530128 183695 530256
rect 183643 530094 183651 530128
rect 183685 530094 183695 530128
rect 183643 530082 183695 530094
rect 184641 530128 184693 530256
rect 184641 530094 184651 530128
rect 184685 530094 184693 530128
rect 184641 530082 184693 530094
rect 184747 530230 184799 530256
rect 184747 530196 184755 530230
rect 184789 530196 184799 530230
rect 184747 530128 184799 530196
rect 184747 530094 184755 530128
rect 184789 530094 184799 530128
rect 184747 530082 184799 530094
rect 185009 530230 185061 530256
rect 185009 530196 185019 530230
rect 185053 530196 185061 530230
rect 185009 530128 185061 530196
rect 185009 530094 185019 530128
rect 185053 530094 185061 530128
rect 185207 530258 185260 530282
rect 185207 530224 185215 530258
rect 185249 530224 185260 530258
rect 185207 530136 185260 530224
rect 185207 530102 185215 530136
rect 185249 530102 185260 530136
rect 185009 530082 185061 530094
rect 185207 530082 185260 530102
rect 185290 530196 185356 530282
rect 185290 530162 185301 530196
rect 185335 530162 185356 530196
rect 185290 530128 185356 530162
rect 185290 530094 185301 530128
rect 185335 530094 185356 530128
rect 185290 530082 185356 530094
rect 185386 530163 185442 530282
rect 185386 530129 185397 530163
rect 185431 530129 185442 530163
rect 185386 530082 185442 530129
rect 185472 530128 185528 530282
rect 185472 530094 185483 530128
rect 185517 530094 185528 530128
rect 185472 530082 185528 530094
rect 185558 530272 185614 530282
rect 185558 530238 185569 530272
rect 185603 530238 185614 530272
rect 185558 530204 185614 530238
rect 185558 530170 185569 530204
rect 185603 530170 185614 530204
rect 185558 530136 185614 530170
rect 185558 530102 185569 530136
rect 185603 530102 185614 530136
rect 185558 530082 185614 530102
rect 185644 530210 185704 530282
rect 185644 530176 185655 530210
rect 185689 530176 185704 530210
rect 185644 530142 185704 530176
rect 185644 530108 185655 530142
rect 185689 530108 185704 530142
rect 185644 530082 185704 530108
rect 185759 530128 185811 530256
rect 185759 530094 185767 530128
rect 185801 530094 185811 530128
rect 185759 530082 185811 530094
rect 186757 530128 186809 530256
rect 186757 530094 186767 530128
rect 186801 530094 186809 530128
rect 186757 530082 186809 530094
rect 187231 530223 187283 530256
rect 187231 530189 187239 530223
rect 187273 530189 187283 530223
rect 187231 530128 187283 530189
rect 187231 530094 187239 530128
rect 187273 530094 187283 530128
rect 187231 530082 187283 530094
rect 187401 530223 187453 530256
rect 187401 530189 187411 530223
rect 187445 530189 187453 530223
rect 187401 530128 187453 530189
rect 187401 530094 187411 530128
rect 187445 530094 187453 530128
rect 187401 530082 187453 530094
rect 172235 529976 172287 529988
rect 172235 529942 172243 529976
rect 172277 529942 172287 529976
rect 172235 529881 172287 529942
rect 172235 529847 172243 529881
rect 172277 529847 172287 529881
rect 172235 529814 172287 529847
rect 172405 529976 172457 529988
rect 172405 529942 172415 529976
rect 172449 529942 172457 529976
rect 172405 529881 172457 529942
rect 172405 529847 172415 529881
rect 172449 529847 172457 529881
rect 172405 529814 172457 529847
rect 172511 529976 172563 529988
rect 172511 529942 172519 529976
rect 172553 529942 172563 529976
rect 172511 529814 172563 529942
rect 173509 529976 173561 529988
rect 173509 529942 173519 529976
rect 173553 529942 173561 529976
rect 173509 529814 173561 529942
rect 173615 529976 173667 529988
rect 173615 529942 173623 529976
rect 173657 529942 173667 529976
rect 173615 529814 173667 529942
rect 174613 529976 174665 529988
rect 174613 529942 174623 529976
rect 174657 529942 174665 529976
rect 174613 529814 174665 529942
rect 174833 529950 174885 529988
rect 174833 529916 174841 529950
rect 174875 529916 174885 529950
rect 174833 529904 174885 529916
rect 174915 529976 174969 529988
rect 174915 529942 174925 529976
rect 174959 529942 174969 529976
rect 174915 529904 174969 529942
rect 175069 529950 175121 529988
rect 175069 529916 175079 529950
rect 175113 529916 175121 529950
rect 175069 529904 175121 529916
rect 175175 529950 175227 529988
rect 175175 529916 175183 529950
rect 175217 529916 175227 529950
rect 175175 529904 175227 529916
rect 175327 529976 175392 529988
rect 175327 529942 175342 529976
rect 175376 529942 175392 529976
rect 175327 529904 175392 529942
rect 175342 529788 175392 529904
rect 175422 529950 175474 529988
rect 175422 529916 175432 529950
rect 175466 529916 175474 529950
rect 175422 529788 175474 529916
rect 175547 529968 175599 529982
rect 175547 529934 175555 529968
rect 175589 529934 175599 529968
rect 175547 529900 175599 529934
rect 175547 529866 175555 529900
rect 175589 529866 175599 529900
rect 175547 529854 175599 529866
rect 175629 529952 175683 529982
rect 175629 529918 175639 529952
rect 175673 529918 175683 529952
rect 175629 529854 175683 529918
rect 175713 529968 175765 529982
rect 175713 529934 175723 529968
rect 175757 529934 175765 529968
rect 175713 529900 175765 529934
rect 175898 529976 175950 529988
rect 175898 529942 175906 529976
rect 175940 529942 175950 529976
rect 175898 529904 175950 529942
rect 175980 529968 176042 529988
rect 175980 529934 175990 529968
rect 176024 529934 176042 529968
rect 175980 529904 176042 529934
rect 176072 529974 176141 529988
rect 176072 529940 176083 529974
rect 176117 529940 176141 529974
rect 176072 529904 176141 529940
rect 176171 529950 176281 529988
rect 176171 529916 176237 529950
rect 176271 529916 176281 529950
rect 176171 529904 176281 529916
rect 176311 529966 176378 529988
rect 176311 529932 176334 529966
rect 176368 529932 176378 529966
rect 176311 529904 176378 529932
rect 176408 529950 176460 529988
rect 176408 529916 176418 529950
rect 176452 529916 176460 529950
rect 176408 529904 176460 529916
rect 176523 529976 176575 529988
rect 176523 529942 176531 529976
rect 176565 529942 176575 529976
rect 175713 529866 175723 529900
rect 175757 529866 175765 529900
rect 175713 529854 175765 529866
rect 176523 529820 176575 529942
rect 176605 529968 176674 529988
rect 176605 529934 176619 529968
rect 176653 529934 176674 529968
rect 176605 529904 176674 529934
rect 176704 529975 176760 529988
rect 176704 529941 176716 529975
rect 176750 529941 176760 529975
rect 176704 529904 176760 529941
rect 176790 529904 176844 529988
rect 176874 529976 176952 529988
rect 176874 529942 176908 529976
rect 176942 529942 176952 529976
rect 176874 529904 176952 529942
rect 176982 529950 177036 529988
rect 176982 529916 176992 529950
rect 177026 529916 177036 529950
rect 176982 529904 177036 529916
rect 177066 529976 177120 529988
rect 177066 529942 177078 529976
rect 177112 529942 177120 529976
rect 177066 529904 177120 529942
rect 177185 529976 177251 529988
rect 177185 529942 177207 529976
rect 177241 529942 177251 529976
rect 177185 529908 177251 529942
rect 176605 529820 176659 529904
rect 177185 529874 177207 529908
rect 177241 529874 177251 529908
rect 177185 529860 177251 529874
rect 177201 529788 177251 529860
rect 177281 529940 177333 529988
rect 178211 529976 178263 529988
rect 177281 529906 177291 529940
rect 177325 529906 177333 529940
rect 177281 529872 177333 529906
rect 177281 529838 177291 529872
rect 177325 529838 177333 529872
rect 177281 529788 177333 529838
rect 178211 529949 178219 529976
rect 177613 529916 177669 529949
rect 177613 529882 177625 529916
rect 177659 529882 177669 529916
rect 177613 529865 177669 529882
rect 177699 529916 177765 529949
rect 177699 529882 177711 529916
rect 177745 529882 177765 529916
rect 177699 529865 177765 529882
rect 177795 529865 177837 529949
rect 177867 529916 178051 529949
rect 177867 529882 177908 529916
rect 177942 529882 177983 529916
rect 178017 529882 178051 529916
rect 177867 529865 178051 529882
rect 178081 529865 178154 529949
rect 178184 529942 178219 529949
rect 178253 529942 178263 529976
rect 178184 529908 178263 529942
rect 178184 529874 178219 529908
rect 178253 529874 178263 529908
rect 178184 529865 178263 529874
rect 178211 529840 178263 529865
rect 178211 529806 178219 529840
rect 178253 529806 178263 529840
rect 178211 529788 178263 529806
rect 178293 529976 178345 529988
rect 178293 529942 178303 529976
rect 178337 529942 178345 529976
rect 178293 529908 178345 529942
rect 178293 529874 178303 529908
rect 178337 529874 178345 529908
rect 178293 529840 178345 529874
rect 178293 529806 178303 529840
rect 178337 529806 178345 529840
rect 178293 529788 178345 529806
rect 178399 529940 178451 529988
rect 178399 529906 178407 529940
rect 178441 529906 178451 529940
rect 178399 529872 178451 529906
rect 178399 529838 178407 529872
rect 178441 529838 178451 529872
rect 178399 529788 178451 529838
rect 178481 529976 178547 529988
rect 178481 529942 178491 529976
rect 178525 529942 178547 529976
rect 178481 529908 178547 529942
rect 178481 529874 178491 529908
rect 178525 529874 178547 529908
rect 178612 529976 178666 529988
rect 178612 529942 178620 529976
rect 178654 529942 178666 529976
rect 178612 529904 178666 529942
rect 178696 529950 178750 529988
rect 178696 529916 178706 529950
rect 178740 529916 178750 529950
rect 178696 529904 178750 529916
rect 178780 529976 178858 529988
rect 178780 529942 178790 529976
rect 178824 529942 178858 529976
rect 178780 529904 178858 529942
rect 178888 529904 178942 529988
rect 178972 529975 179028 529988
rect 178972 529941 178982 529975
rect 179016 529941 179028 529975
rect 178972 529904 179028 529941
rect 179058 529968 179127 529988
rect 179058 529934 179079 529968
rect 179113 529934 179127 529968
rect 179058 529904 179127 529934
rect 178481 529860 178547 529874
rect 178481 529788 178531 529860
rect 179073 529820 179127 529904
rect 179157 529976 179209 529988
rect 179157 529942 179167 529976
rect 179201 529942 179209 529976
rect 179157 529820 179209 529942
rect 179272 529950 179324 529988
rect 179272 529916 179280 529950
rect 179314 529916 179324 529950
rect 179272 529904 179324 529916
rect 179354 529966 179421 529988
rect 179354 529932 179364 529966
rect 179398 529932 179421 529966
rect 179354 529904 179421 529932
rect 179451 529950 179561 529988
rect 179451 529916 179461 529950
rect 179495 529916 179561 529950
rect 179451 529904 179561 529916
rect 179591 529974 179660 529988
rect 179591 529940 179615 529974
rect 179649 529940 179660 529974
rect 179591 529904 179660 529940
rect 179690 529968 179752 529988
rect 179690 529934 179708 529968
rect 179742 529934 179752 529968
rect 179690 529904 179752 529934
rect 179782 529976 179834 529988
rect 179782 529942 179792 529976
rect 179826 529942 179834 529976
rect 179782 529904 179834 529942
rect 179967 529968 180019 529982
rect 179967 529934 179975 529968
rect 180009 529934 180019 529968
rect 179967 529900 180019 529934
rect 179967 529866 179975 529900
rect 180009 529866 180019 529900
rect 179967 529854 180019 529866
rect 180049 529952 180103 529982
rect 180049 529918 180059 529952
rect 180093 529918 180103 529952
rect 180049 529854 180103 529918
rect 180133 529968 180185 529982
rect 180133 529934 180143 529968
rect 180177 529934 180185 529968
rect 180133 529900 180185 529934
rect 180133 529866 180143 529900
rect 180177 529866 180185 529900
rect 180133 529854 180185 529866
rect 180239 529968 180291 529982
rect 180239 529934 180247 529968
rect 180281 529934 180291 529968
rect 180239 529900 180291 529934
rect 180239 529866 180247 529900
rect 180281 529866 180291 529900
rect 180239 529854 180291 529866
rect 180321 529952 180375 529982
rect 180321 529918 180331 529952
rect 180365 529918 180375 529952
rect 180321 529854 180375 529918
rect 180405 529968 180457 529982
rect 180405 529934 180415 529968
rect 180449 529934 180457 529968
rect 180405 529900 180457 529934
rect 180590 529976 180642 529988
rect 180590 529942 180598 529976
rect 180632 529942 180642 529976
rect 180590 529904 180642 529942
rect 180672 529968 180734 529988
rect 180672 529934 180682 529968
rect 180716 529934 180734 529968
rect 180672 529904 180734 529934
rect 180764 529974 180833 529988
rect 180764 529940 180775 529974
rect 180809 529940 180833 529974
rect 180764 529904 180833 529940
rect 180863 529950 180973 529988
rect 180863 529916 180929 529950
rect 180963 529916 180973 529950
rect 180863 529904 180973 529916
rect 181003 529966 181070 529988
rect 181003 529932 181026 529966
rect 181060 529932 181070 529966
rect 181003 529904 181070 529932
rect 181100 529950 181152 529988
rect 181100 529916 181110 529950
rect 181144 529916 181152 529950
rect 181100 529904 181152 529916
rect 181215 529976 181267 529988
rect 181215 529942 181223 529976
rect 181257 529942 181267 529976
rect 180405 529866 180415 529900
rect 180449 529866 180457 529900
rect 180405 529854 180457 529866
rect 181215 529820 181267 529942
rect 181297 529968 181366 529988
rect 181297 529934 181311 529968
rect 181345 529934 181366 529968
rect 181297 529904 181366 529934
rect 181396 529975 181452 529988
rect 181396 529941 181408 529975
rect 181442 529941 181452 529975
rect 181396 529904 181452 529941
rect 181482 529904 181536 529988
rect 181566 529976 181644 529988
rect 181566 529942 181600 529976
rect 181634 529942 181644 529976
rect 181566 529904 181644 529942
rect 181674 529950 181728 529988
rect 181674 529916 181684 529950
rect 181718 529916 181728 529950
rect 181674 529904 181728 529916
rect 181758 529976 181812 529988
rect 181758 529942 181770 529976
rect 181804 529942 181812 529976
rect 181758 529904 181812 529942
rect 181877 529976 181943 529988
rect 181877 529942 181899 529976
rect 181933 529942 181943 529976
rect 181877 529908 181943 529942
rect 181297 529820 181351 529904
rect 181877 529874 181899 529908
rect 181933 529874 181943 529908
rect 181877 529860 181943 529874
rect 181893 529788 181943 529860
rect 181973 529940 182025 529988
rect 181973 529906 181983 529940
rect 182017 529906 182025 529940
rect 181973 529872 182025 529906
rect 181973 529838 181983 529872
rect 182017 529838 182025 529872
rect 181973 529788 182025 529838
rect 182079 529976 182131 529988
rect 182079 529942 182087 529976
rect 182121 529942 182131 529976
rect 182079 529874 182131 529942
rect 182079 529840 182087 529874
rect 182121 529840 182131 529874
rect 182079 529814 182131 529840
rect 182341 529976 182393 529988
rect 182341 529942 182351 529976
rect 182385 529942 182393 529976
rect 182341 529874 182393 529942
rect 182341 529840 182351 529874
rect 182385 529840 182393 529874
rect 182341 529814 182393 529840
rect 182650 529950 182702 529988
rect 182650 529916 182658 529950
rect 182692 529916 182702 529950
rect 182650 529788 182702 529916
rect 182732 529976 182797 529988
rect 182732 529942 182748 529976
rect 182782 529942 182797 529976
rect 182732 529904 182797 529942
rect 182897 529950 182949 529988
rect 182897 529916 182907 529950
rect 182941 529916 182949 529950
rect 182897 529904 182949 529916
rect 183003 529950 183055 529988
rect 183003 529916 183011 529950
rect 183045 529916 183055 529950
rect 183003 529904 183055 529916
rect 183155 529976 183209 529988
rect 183155 529942 183165 529976
rect 183199 529942 183209 529976
rect 183155 529904 183209 529942
rect 183239 529950 183291 529988
rect 183239 529916 183249 529950
rect 183283 529916 183291 529950
rect 183239 529904 183291 529916
rect 183367 529976 183419 529988
rect 183367 529942 183375 529976
rect 183409 529942 183419 529976
rect 182732 529788 182782 529904
rect 183367 529814 183419 529942
rect 184365 529976 184417 529988
rect 184365 529942 184375 529976
rect 184409 529942 184417 529976
rect 184365 529814 184417 529942
rect 184471 529976 184523 529988
rect 184471 529942 184479 529976
rect 184513 529942 184523 529976
rect 184471 529814 184523 529942
rect 185469 529976 185521 529988
rect 185469 529942 185479 529976
rect 185513 529942 185521 529976
rect 185469 529814 185521 529942
rect 185575 529976 185627 529988
rect 185575 529942 185583 529976
rect 185617 529942 185627 529976
rect 185575 529814 185627 529942
rect 186573 529976 186625 529988
rect 186573 529942 186583 529976
rect 186617 529942 186625 529976
rect 186573 529814 186625 529942
rect 186679 529976 186731 529988
rect 186679 529942 186687 529976
rect 186721 529942 186731 529976
rect 186679 529874 186731 529942
rect 186679 529840 186687 529874
rect 186721 529840 186731 529874
rect 186679 529814 186731 529840
rect 187125 529976 187177 529988
rect 187125 529942 187135 529976
rect 187169 529942 187177 529976
rect 187125 529874 187177 529942
rect 187125 529840 187135 529874
rect 187169 529840 187177 529874
rect 187125 529814 187177 529840
rect 187231 529976 187283 529988
rect 187231 529942 187239 529976
rect 187273 529942 187283 529976
rect 187231 529881 187283 529942
rect 187231 529847 187239 529881
rect 187273 529847 187283 529881
rect 187231 529814 187283 529847
rect 187401 529976 187453 529988
rect 187401 529942 187411 529976
rect 187445 529942 187453 529976
rect 187401 529881 187453 529942
rect 187401 529847 187411 529881
rect 187445 529847 187453 529881
rect 187401 529814 187453 529847
rect 172235 529135 172287 529168
rect 172235 529101 172243 529135
rect 172277 529101 172287 529135
rect 172235 529040 172287 529101
rect 172235 529006 172243 529040
rect 172277 529006 172287 529040
rect 172235 528994 172287 529006
rect 172405 529135 172457 529168
rect 172405 529101 172415 529135
rect 172449 529101 172457 529135
rect 172405 529040 172457 529101
rect 172405 529006 172415 529040
rect 172449 529006 172457 529040
rect 172405 528994 172457 529006
rect 172511 529040 172563 529168
rect 172511 529006 172519 529040
rect 172553 529006 172563 529040
rect 172511 528994 172563 529006
rect 173509 529040 173561 529168
rect 173509 529006 173519 529040
rect 173553 529006 173561 529040
rect 173509 528994 173561 529006
rect 173615 529040 173667 529168
rect 173615 529006 173623 529040
rect 173657 529006 173667 529040
rect 173615 528994 173667 529006
rect 174613 529040 174665 529168
rect 174613 529006 174623 529040
rect 174657 529006 174665 529040
rect 175727 529176 175779 529194
rect 175727 529142 175735 529176
rect 175769 529142 175779 529176
rect 175727 529117 175779 529142
rect 175129 529100 175185 529117
rect 175129 529066 175141 529100
rect 175175 529066 175185 529100
rect 175129 529033 175185 529066
rect 175215 529100 175281 529117
rect 175215 529066 175227 529100
rect 175261 529066 175281 529100
rect 175215 529033 175281 529066
rect 175311 529033 175353 529117
rect 175383 529100 175567 529117
rect 175383 529066 175424 529100
rect 175458 529066 175499 529100
rect 175533 529066 175567 529100
rect 175383 529033 175567 529066
rect 175597 529033 175670 529117
rect 175700 529108 175779 529117
rect 175700 529074 175735 529108
rect 175769 529074 175779 529108
rect 175700 529040 175779 529074
rect 175700 529033 175735 529040
rect 174613 528994 174665 529006
rect 175727 529006 175735 529033
rect 175769 529006 175779 529040
rect 175727 528994 175779 529006
rect 175809 529176 175861 529194
rect 175809 529142 175819 529176
rect 175853 529142 175861 529176
rect 175809 529108 175861 529142
rect 175809 529074 175819 529108
rect 175853 529074 175861 529108
rect 175809 529040 175861 529074
rect 175809 529006 175819 529040
rect 175853 529006 175861 529040
rect 175809 528994 175861 529006
rect 175932 529064 175985 529194
rect 175932 529030 175940 529064
rect 175974 529030 175985 529064
rect 175932 528994 175985 529030
rect 176015 529170 176071 529194
rect 176015 529136 176026 529170
rect 176060 529136 176071 529170
rect 176015 529084 176071 529136
rect 176015 529050 176026 529084
rect 176060 529050 176071 529084
rect 176015 528994 176071 529050
rect 176101 529064 176157 529194
rect 176101 529030 176112 529064
rect 176146 529030 176157 529064
rect 176101 528994 176157 529030
rect 176187 529170 176243 529194
rect 176187 529136 176198 529170
rect 176232 529136 176243 529170
rect 176187 529084 176243 529136
rect 176187 529050 176198 529084
rect 176232 529050 176243 529084
rect 176187 528994 176243 529050
rect 176273 529064 176329 529194
rect 176273 529030 176284 529064
rect 176318 529030 176329 529064
rect 176273 528994 176329 529030
rect 176359 529170 176415 529194
rect 176359 529136 176370 529170
rect 176404 529136 176415 529170
rect 176359 529084 176415 529136
rect 176359 529050 176370 529084
rect 176404 529050 176415 529084
rect 176359 528994 176415 529050
rect 176445 529064 176501 529194
rect 176445 529030 176456 529064
rect 176490 529030 176501 529064
rect 176445 528994 176501 529030
rect 176531 529170 176587 529194
rect 176531 529136 176542 529170
rect 176576 529136 176587 529170
rect 176531 529084 176587 529136
rect 176531 529050 176542 529084
rect 176576 529050 176587 529084
rect 176531 528994 176587 529050
rect 176617 529064 176672 529194
rect 176617 529030 176627 529064
rect 176661 529030 176672 529064
rect 176617 528994 176672 529030
rect 176702 529170 176758 529194
rect 176702 529136 176713 529170
rect 176747 529136 176758 529170
rect 176702 529084 176758 529136
rect 176702 529050 176713 529084
rect 176747 529050 176758 529084
rect 176702 528994 176758 529050
rect 176788 529064 176844 529194
rect 176788 529030 176799 529064
rect 176833 529030 176844 529064
rect 176788 528994 176844 529030
rect 176874 529170 176930 529194
rect 176874 529136 176885 529170
rect 176919 529136 176930 529170
rect 176874 529084 176930 529136
rect 176874 529050 176885 529084
rect 176919 529050 176930 529084
rect 176874 528994 176930 529050
rect 176960 529064 177016 529194
rect 176960 529030 176971 529064
rect 177005 529030 177016 529064
rect 176960 528994 177016 529030
rect 177046 529170 177102 529194
rect 177046 529136 177057 529170
rect 177091 529136 177102 529170
rect 177046 529084 177102 529136
rect 177046 529050 177057 529084
rect 177091 529050 177102 529084
rect 177046 528994 177102 529050
rect 177132 529064 177188 529194
rect 177132 529030 177143 529064
rect 177177 529030 177188 529064
rect 177132 528994 177188 529030
rect 177218 529170 177274 529194
rect 177218 529136 177229 529170
rect 177263 529136 177274 529170
rect 177218 529084 177274 529136
rect 177218 529050 177229 529084
rect 177263 529050 177274 529084
rect 177218 528994 177274 529050
rect 177304 529108 177360 529194
rect 177304 529074 177315 529108
rect 177349 529074 177360 529108
rect 177304 529040 177360 529074
rect 177304 529006 177315 529040
rect 177349 529006 177360 529040
rect 177304 528994 177360 529006
rect 177390 529124 177446 529194
rect 177390 529090 177401 529124
rect 177435 529090 177446 529124
rect 177390 529056 177446 529090
rect 177390 529022 177401 529056
rect 177435 529022 177446 529056
rect 177390 528994 177446 529022
rect 177476 529108 177532 529194
rect 177476 529074 177487 529108
rect 177521 529074 177532 529108
rect 177476 529040 177532 529074
rect 177476 529006 177487 529040
rect 177521 529006 177532 529040
rect 177476 528994 177532 529006
rect 177562 529116 177618 529194
rect 177562 529082 177573 529116
rect 177607 529082 177618 529116
rect 177562 529048 177618 529082
rect 177562 529014 177573 529048
rect 177607 529014 177618 529048
rect 177562 528994 177618 529014
rect 177648 529108 177701 529194
rect 177648 529074 177659 529108
rect 177693 529074 177701 529108
rect 177648 529040 177701 529074
rect 177648 529006 177659 529040
rect 177693 529006 177701 529040
rect 177648 528994 177701 529006
rect 177755 529116 177807 529128
rect 177755 529082 177763 529116
rect 177797 529082 177807 529116
rect 177755 529048 177807 529082
rect 177755 529014 177763 529048
rect 177797 529014 177807 529048
rect 177755 529000 177807 529014
rect 177837 529064 177891 529128
rect 177837 529030 177847 529064
rect 177881 529030 177891 529064
rect 177837 529000 177891 529030
rect 177921 529116 177973 529128
rect 177921 529082 177931 529116
rect 177965 529082 177973 529116
rect 177921 529048 177973 529082
rect 177921 529014 177931 529048
rect 177965 529014 177973 529048
rect 177921 529000 177973 529014
rect 178106 529040 178158 529078
rect 178106 529006 178114 529040
rect 178148 529006 178158 529040
rect 178106 528994 178158 529006
rect 178188 529048 178250 529078
rect 178188 529014 178198 529048
rect 178232 529014 178250 529048
rect 178188 528994 178250 529014
rect 178280 529042 178349 529078
rect 178280 529008 178291 529042
rect 178325 529008 178349 529042
rect 178280 528994 178349 529008
rect 178379 529066 178489 529078
rect 178379 529032 178445 529066
rect 178479 529032 178489 529066
rect 178379 528994 178489 529032
rect 178519 529050 178586 529078
rect 178519 529016 178542 529050
rect 178576 529016 178586 529050
rect 178519 528994 178586 529016
rect 178616 529066 178668 529078
rect 178616 529032 178626 529066
rect 178660 529032 178668 529066
rect 178616 528994 178668 529032
rect 178731 529040 178783 529162
rect 178731 529006 178739 529040
rect 178773 529006 178783 529040
rect 178731 528994 178783 529006
rect 178813 529078 178867 529162
rect 179409 529122 179459 529194
rect 179393 529108 179459 529122
rect 178813 529048 178882 529078
rect 178813 529014 178827 529048
rect 178861 529014 178882 529048
rect 178813 528994 178882 529014
rect 178912 529041 178968 529078
rect 178912 529007 178924 529041
rect 178958 529007 178968 529041
rect 178912 528994 178968 529007
rect 178998 528994 179052 529078
rect 179082 529040 179160 529078
rect 179082 529006 179116 529040
rect 179150 529006 179160 529040
rect 179082 528994 179160 529006
rect 179190 529066 179244 529078
rect 179190 529032 179200 529066
rect 179234 529032 179244 529066
rect 179190 528994 179244 529032
rect 179274 529040 179328 529078
rect 179274 529006 179286 529040
rect 179320 529006 179328 529040
rect 179274 528994 179328 529006
rect 179393 529074 179415 529108
rect 179449 529074 179459 529108
rect 179393 529040 179459 529074
rect 179393 529006 179415 529040
rect 179449 529006 179459 529040
rect 179393 528994 179459 529006
rect 179489 529144 179541 529194
rect 179489 529110 179499 529144
rect 179533 529110 179541 529144
rect 179489 529076 179541 529110
rect 179489 529042 179499 529076
rect 179533 529042 179541 529076
rect 179489 528994 179541 529042
rect 179687 529116 179739 529152
rect 179687 529082 179695 529116
rect 179729 529082 179739 529116
rect 179687 529048 179739 529082
rect 179687 529014 179695 529048
rect 179729 529014 179739 529048
rect 179687 528994 179739 529014
rect 179769 529116 179827 529152
rect 179769 529082 179781 529116
rect 179815 529082 179827 529116
rect 179769 529048 179827 529082
rect 179769 529014 179781 529048
rect 179815 529014 179827 529048
rect 179769 528994 179827 529014
rect 179857 529129 179909 529152
rect 179857 529095 179867 529129
rect 179901 529095 179909 529129
rect 179857 529048 179909 529095
rect 179857 529014 179867 529048
rect 179901 529014 179909 529048
rect 179857 528994 179909 529014
rect 180055 529142 180107 529168
rect 180055 529108 180063 529142
rect 180097 529108 180107 529142
rect 180055 529040 180107 529108
rect 180055 529006 180063 529040
rect 180097 529006 180107 529040
rect 180055 528994 180107 529006
rect 180501 529142 180553 529168
rect 180501 529108 180511 529142
rect 180545 529108 180553 529142
rect 180501 529040 180553 529108
rect 180501 529006 180511 529040
rect 180545 529006 180553 529040
rect 180501 528994 180553 529006
rect 180699 529108 180752 529194
rect 180699 529074 180707 529108
rect 180741 529074 180752 529108
rect 180699 529040 180752 529074
rect 180699 529006 180707 529040
rect 180741 529006 180752 529040
rect 180699 528994 180752 529006
rect 180782 529116 180838 529194
rect 180782 529082 180793 529116
rect 180827 529082 180838 529116
rect 180782 529048 180838 529082
rect 180782 529014 180793 529048
rect 180827 529014 180838 529048
rect 180782 528994 180838 529014
rect 180868 529108 180924 529194
rect 180868 529074 180879 529108
rect 180913 529074 180924 529108
rect 180868 529040 180924 529074
rect 180868 529006 180879 529040
rect 180913 529006 180924 529040
rect 180868 528994 180924 529006
rect 180954 529124 181010 529194
rect 180954 529090 180965 529124
rect 180999 529090 181010 529124
rect 180954 529056 181010 529090
rect 180954 529022 180965 529056
rect 180999 529022 181010 529056
rect 180954 528994 181010 529022
rect 181040 529108 181096 529194
rect 181040 529074 181051 529108
rect 181085 529074 181096 529108
rect 181040 529040 181096 529074
rect 181040 529006 181051 529040
rect 181085 529006 181096 529040
rect 181040 528994 181096 529006
rect 181126 529170 181182 529194
rect 181126 529136 181137 529170
rect 181171 529136 181182 529170
rect 181126 529084 181182 529136
rect 181126 529050 181137 529084
rect 181171 529050 181182 529084
rect 181126 528994 181182 529050
rect 181212 529064 181268 529194
rect 181212 529030 181223 529064
rect 181257 529030 181268 529064
rect 181212 528994 181268 529030
rect 181298 529170 181354 529194
rect 181298 529136 181309 529170
rect 181343 529136 181354 529170
rect 181298 529084 181354 529136
rect 181298 529050 181309 529084
rect 181343 529050 181354 529084
rect 181298 528994 181354 529050
rect 181384 529064 181440 529194
rect 181384 529030 181395 529064
rect 181429 529030 181440 529064
rect 181384 528994 181440 529030
rect 181470 529170 181526 529194
rect 181470 529136 181481 529170
rect 181515 529136 181526 529170
rect 181470 529084 181526 529136
rect 181470 529050 181481 529084
rect 181515 529050 181526 529084
rect 181470 528994 181526 529050
rect 181556 529064 181612 529194
rect 181556 529030 181567 529064
rect 181601 529030 181612 529064
rect 181556 528994 181612 529030
rect 181642 529170 181698 529194
rect 181642 529136 181653 529170
rect 181687 529136 181698 529170
rect 181642 529084 181698 529136
rect 181642 529050 181653 529084
rect 181687 529050 181698 529084
rect 181642 528994 181698 529050
rect 181728 529064 181783 529194
rect 181728 529030 181739 529064
rect 181773 529030 181783 529064
rect 181728 528994 181783 529030
rect 181813 529170 181869 529194
rect 181813 529136 181824 529170
rect 181858 529136 181869 529170
rect 181813 529084 181869 529136
rect 181813 529050 181824 529084
rect 181858 529050 181869 529084
rect 181813 528994 181869 529050
rect 181899 529064 181955 529194
rect 181899 529030 181910 529064
rect 181944 529030 181955 529064
rect 181899 528994 181955 529030
rect 181985 529170 182041 529194
rect 181985 529136 181996 529170
rect 182030 529136 182041 529170
rect 181985 529084 182041 529136
rect 181985 529050 181996 529084
rect 182030 529050 182041 529084
rect 181985 528994 182041 529050
rect 182071 529064 182127 529194
rect 182071 529030 182082 529064
rect 182116 529030 182127 529064
rect 182071 528994 182127 529030
rect 182157 529170 182213 529194
rect 182157 529136 182168 529170
rect 182202 529136 182213 529170
rect 182157 529084 182213 529136
rect 182157 529050 182168 529084
rect 182202 529050 182213 529084
rect 182157 528994 182213 529050
rect 182243 529064 182299 529194
rect 182243 529030 182254 529064
rect 182288 529030 182299 529064
rect 182243 528994 182299 529030
rect 182329 529170 182385 529194
rect 182329 529136 182340 529170
rect 182374 529136 182385 529170
rect 182329 529084 182385 529136
rect 182329 529050 182340 529084
rect 182374 529050 182385 529084
rect 182329 528994 182385 529050
rect 182415 529064 182468 529194
rect 182415 529030 182426 529064
rect 182460 529030 182468 529064
rect 182415 528994 182468 529030
rect 182539 529129 182591 529152
rect 182539 529095 182547 529129
rect 182581 529095 182591 529129
rect 182539 529048 182591 529095
rect 182539 529014 182547 529048
rect 182581 529014 182591 529048
rect 182539 528994 182591 529014
rect 182621 529116 182679 529152
rect 182621 529082 182633 529116
rect 182667 529082 182679 529116
rect 182621 529048 182679 529082
rect 182621 529014 182633 529048
rect 182667 529014 182679 529048
rect 182621 528994 182679 529014
rect 182709 529116 182761 529152
rect 182709 529082 182719 529116
rect 182753 529082 182761 529116
rect 182709 529048 182761 529082
rect 182709 529014 182719 529048
rect 182753 529014 182761 529048
rect 182709 528994 182761 529014
rect 182815 529040 182867 529168
rect 182815 529006 182823 529040
rect 182857 529006 182867 529040
rect 182815 528994 182867 529006
rect 183813 529040 183865 529168
rect 183813 529006 183823 529040
rect 183857 529006 183865 529040
rect 183813 528994 183865 529006
rect 183919 529040 183971 529168
rect 183919 529006 183927 529040
rect 183961 529006 183971 529040
rect 183919 528994 183971 529006
rect 184917 529040 184969 529168
rect 184917 529006 184927 529040
rect 184961 529006 184969 529040
rect 185207 529040 185259 529168
rect 184917 528994 184969 529006
rect 185207 529006 185215 529040
rect 185249 529006 185259 529040
rect 185207 528994 185259 529006
rect 186205 529040 186257 529168
rect 186205 529006 186215 529040
rect 186249 529006 186257 529040
rect 186205 528994 186257 529006
rect 186311 529142 186363 529168
rect 186311 529108 186319 529142
rect 186353 529108 186363 529142
rect 186311 529040 186363 529108
rect 186311 529006 186319 529040
rect 186353 529006 186363 529040
rect 186311 528994 186363 529006
rect 186941 529142 186993 529168
rect 186941 529108 186951 529142
rect 186985 529108 186993 529142
rect 186941 529040 186993 529108
rect 186941 529006 186951 529040
rect 186985 529006 186993 529040
rect 186941 528994 186993 529006
rect 187231 529135 187283 529168
rect 187231 529101 187239 529135
rect 187273 529101 187283 529135
rect 187231 529040 187283 529101
rect 187231 529006 187239 529040
rect 187273 529006 187283 529040
rect 187231 528994 187283 529006
rect 187401 529135 187453 529168
rect 187401 529101 187411 529135
rect 187445 529101 187453 529135
rect 187401 529040 187453 529101
rect 187401 529006 187411 529040
rect 187445 529006 187453 529040
rect 187401 528994 187453 529006
rect 172235 528888 172287 528900
rect 172235 528854 172243 528888
rect 172277 528854 172287 528888
rect 172235 528793 172287 528854
rect 172235 528759 172243 528793
rect 172277 528759 172287 528793
rect 172235 528726 172287 528759
rect 172405 528888 172457 528900
rect 172405 528854 172415 528888
rect 172449 528854 172457 528888
rect 172405 528793 172457 528854
rect 172405 528759 172415 528793
rect 172449 528759 172457 528793
rect 172405 528726 172457 528759
rect 172511 528888 172563 528900
rect 172511 528854 172519 528888
rect 172553 528854 172563 528888
rect 172511 528726 172563 528854
rect 173509 528888 173561 528900
rect 173509 528854 173519 528888
rect 173553 528854 173561 528888
rect 173509 528726 173561 528854
rect 173615 528888 173667 528900
rect 173615 528854 173623 528888
rect 173657 528854 173667 528888
rect 173615 528726 173667 528854
rect 174613 528888 174665 528900
rect 174613 528854 174623 528888
rect 174657 528854 174665 528888
rect 174613 528726 174665 528854
rect 174719 528888 174771 528900
rect 174719 528854 174727 528888
rect 174761 528854 174771 528888
rect 174719 528726 174771 528854
rect 175717 528888 175769 528900
rect 175717 528854 175727 528888
rect 175761 528854 175769 528888
rect 175717 528726 175769 528854
rect 175915 528880 175967 528900
rect 175915 528846 175923 528880
rect 175957 528846 175967 528880
rect 175915 528812 175967 528846
rect 175915 528778 175923 528812
rect 175957 528778 175967 528812
rect 175915 528742 175967 528778
rect 175997 528880 176055 528900
rect 175997 528846 176009 528880
rect 176043 528846 176055 528880
rect 175997 528812 176055 528846
rect 175997 528778 176009 528812
rect 176043 528778 176055 528812
rect 175997 528742 176055 528778
rect 176085 528880 176137 528900
rect 176085 528846 176095 528880
rect 176129 528846 176137 528880
rect 176085 528799 176137 528846
rect 176085 528765 176095 528799
rect 176129 528765 176137 528799
rect 176085 528742 176137 528765
rect 176191 528880 176243 528900
rect 176191 528846 176199 528880
rect 176233 528846 176243 528880
rect 176191 528812 176243 528846
rect 176191 528778 176199 528812
rect 176233 528778 176243 528812
rect 176191 528742 176243 528778
rect 176273 528880 176331 528900
rect 176273 528846 176285 528880
rect 176319 528846 176331 528880
rect 176273 528812 176331 528846
rect 176273 528778 176285 528812
rect 176319 528778 176331 528812
rect 176273 528742 176331 528778
rect 176361 528880 176413 528900
rect 177107 528888 177159 528900
rect 176361 528846 176371 528880
rect 176405 528846 176413 528880
rect 177107 528861 177115 528888
rect 176361 528799 176413 528846
rect 176361 528765 176371 528799
rect 176405 528765 176413 528799
rect 176509 528828 176565 528861
rect 176509 528794 176521 528828
rect 176555 528794 176565 528828
rect 176509 528777 176565 528794
rect 176595 528828 176661 528861
rect 176595 528794 176607 528828
rect 176641 528794 176661 528828
rect 176595 528777 176661 528794
rect 176691 528777 176733 528861
rect 176763 528828 176947 528861
rect 176763 528794 176804 528828
rect 176838 528794 176879 528828
rect 176913 528794 176947 528828
rect 176763 528777 176947 528794
rect 176977 528777 177050 528861
rect 177080 528854 177115 528861
rect 177149 528854 177159 528888
rect 177080 528820 177159 528854
rect 177080 528786 177115 528820
rect 177149 528786 177159 528820
rect 177080 528777 177159 528786
rect 176361 528742 176413 528765
rect 177107 528752 177159 528777
rect 177107 528718 177115 528752
rect 177149 528718 177159 528752
rect 177107 528700 177159 528718
rect 177189 528888 177241 528900
rect 177189 528854 177199 528888
rect 177233 528854 177241 528888
rect 177189 528820 177241 528854
rect 177189 528786 177199 528820
rect 177233 528786 177241 528820
rect 177189 528752 177241 528786
rect 177189 528718 177199 528752
rect 177233 528718 177241 528752
rect 177189 528700 177241 528718
rect 177498 528862 177550 528900
rect 177498 528828 177506 528862
rect 177540 528828 177550 528862
rect 177498 528700 177550 528828
rect 177580 528888 177645 528900
rect 177580 528854 177596 528888
rect 177630 528854 177645 528888
rect 177580 528816 177645 528854
rect 177745 528862 177797 528900
rect 177745 528828 177755 528862
rect 177789 528828 177797 528862
rect 177745 528816 177797 528828
rect 177851 528862 177903 528900
rect 177851 528828 177859 528862
rect 177893 528828 177903 528862
rect 177851 528816 177903 528828
rect 178003 528888 178057 528900
rect 178003 528854 178013 528888
rect 178047 528854 178057 528888
rect 178003 528816 178057 528854
rect 178087 528862 178139 528900
rect 178087 528828 178097 528862
rect 178131 528828 178139 528862
rect 178087 528816 178139 528828
rect 178399 528888 178452 528900
rect 178399 528854 178407 528888
rect 178441 528854 178452 528888
rect 178399 528820 178452 528854
rect 177580 528700 177630 528816
rect 178399 528786 178407 528820
rect 178441 528786 178452 528820
rect 178399 528700 178452 528786
rect 178482 528880 178538 528900
rect 178482 528846 178493 528880
rect 178527 528846 178538 528880
rect 178482 528812 178538 528846
rect 178482 528778 178493 528812
rect 178527 528778 178538 528812
rect 178482 528700 178538 528778
rect 178568 528888 178624 528900
rect 178568 528854 178579 528888
rect 178613 528854 178624 528888
rect 178568 528820 178624 528854
rect 178568 528786 178579 528820
rect 178613 528786 178624 528820
rect 178568 528700 178624 528786
rect 178654 528872 178710 528900
rect 178654 528838 178665 528872
rect 178699 528838 178710 528872
rect 178654 528804 178710 528838
rect 178654 528770 178665 528804
rect 178699 528770 178710 528804
rect 178654 528700 178710 528770
rect 178740 528888 178796 528900
rect 178740 528854 178751 528888
rect 178785 528854 178796 528888
rect 178740 528820 178796 528854
rect 178740 528786 178751 528820
rect 178785 528786 178796 528820
rect 178740 528700 178796 528786
rect 178826 528844 178882 528900
rect 178826 528810 178837 528844
rect 178871 528810 178882 528844
rect 178826 528758 178882 528810
rect 178826 528724 178837 528758
rect 178871 528724 178882 528758
rect 178826 528700 178882 528724
rect 178912 528864 178968 528900
rect 178912 528830 178923 528864
rect 178957 528830 178968 528864
rect 178912 528700 178968 528830
rect 178998 528844 179054 528900
rect 178998 528810 179009 528844
rect 179043 528810 179054 528844
rect 178998 528758 179054 528810
rect 178998 528724 179009 528758
rect 179043 528724 179054 528758
rect 178998 528700 179054 528724
rect 179084 528864 179140 528900
rect 179084 528830 179095 528864
rect 179129 528830 179140 528864
rect 179084 528700 179140 528830
rect 179170 528844 179226 528900
rect 179170 528810 179181 528844
rect 179215 528810 179226 528844
rect 179170 528758 179226 528810
rect 179170 528724 179181 528758
rect 179215 528724 179226 528758
rect 179170 528700 179226 528724
rect 179256 528864 179312 528900
rect 179256 528830 179267 528864
rect 179301 528830 179312 528864
rect 179256 528700 179312 528830
rect 179342 528844 179398 528900
rect 179342 528810 179353 528844
rect 179387 528810 179398 528844
rect 179342 528758 179398 528810
rect 179342 528724 179353 528758
rect 179387 528724 179398 528758
rect 179342 528700 179398 528724
rect 179428 528864 179483 528900
rect 179428 528830 179439 528864
rect 179473 528830 179483 528864
rect 179428 528700 179483 528830
rect 179513 528844 179569 528900
rect 179513 528810 179524 528844
rect 179558 528810 179569 528844
rect 179513 528758 179569 528810
rect 179513 528724 179524 528758
rect 179558 528724 179569 528758
rect 179513 528700 179569 528724
rect 179599 528864 179655 528900
rect 179599 528830 179610 528864
rect 179644 528830 179655 528864
rect 179599 528700 179655 528830
rect 179685 528844 179741 528900
rect 179685 528810 179696 528844
rect 179730 528810 179741 528844
rect 179685 528758 179741 528810
rect 179685 528724 179696 528758
rect 179730 528724 179741 528758
rect 179685 528700 179741 528724
rect 179771 528864 179827 528900
rect 179771 528830 179782 528864
rect 179816 528830 179827 528864
rect 179771 528700 179827 528830
rect 179857 528844 179913 528900
rect 179857 528810 179868 528844
rect 179902 528810 179913 528844
rect 179857 528758 179913 528810
rect 179857 528724 179868 528758
rect 179902 528724 179913 528758
rect 179857 528700 179913 528724
rect 179943 528864 179999 528900
rect 179943 528830 179954 528864
rect 179988 528830 179999 528864
rect 179943 528700 179999 528830
rect 180029 528844 180085 528900
rect 180029 528810 180040 528844
rect 180074 528810 180085 528844
rect 180029 528758 180085 528810
rect 180029 528724 180040 528758
rect 180074 528724 180085 528758
rect 180029 528700 180085 528724
rect 180115 528864 180168 528900
rect 180115 528830 180126 528864
rect 180160 528830 180168 528864
rect 180115 528700 180168 528830
rect 180239 528880 180291 528900
rect 180239 528846 180247 528880
rect 180281 528846 180291 528880
rect 180239 528812 180291 528846
rect 180239 528778 180247 528812
rect 180281 528778 180291 528812
rect 180239 528742 180291 528778
rect 180321 528880 180379 528900
rect 180321 528846 180333 528880
rect 180367 528846 180379 528880
rect 180321 528812 180379 528846
rect 180321 528778 180333 528812
rect 180367 528778 180379 528812
rect 180321 528742 180379 528778
rect 180409 528880 180461 528900
rect 180409 528846 180419 528880
rect 180453 528846 180461 528880
rect 180409 528799 180461 528846
rect 180409 528765 180419 528799
rect 180453 528765 180461 528799
rect 180515 528880 180567 528894
rect 180515 528846 180523 528880
rect 180557 528846 180567 528880
rect 180515 528812 180567 528846
rect 180515 528778 180523 528812
rect 180557 528778 180567 528812
rect 180515 528766 180567 528778
rect 180597 528864 180651 528894
rect 180597 528830 180607 528864
rect 180641 528830 180651 528864
rect 180597 528766 180651 528830
rect 180681 528880 180733 528894
rect 180681 528846 180691 528880
rect 180725 528846 180733 528880
rect 180681 528812 180733 528846
rect 180866 528888 180918 528900
rect 180866 528854 180874 528888
rect 180908 528854 180918 528888
rect 180866 528816 180918 528854
rect 180948 528880 181010 528900
rect 180948 528846 180958 528880
rect 180992 528846 181010 528880
rect 180948 528816 181010 528846
rect 181040 528886 181109 528900
rect 181040 528852 181051 528886
rect 181085 528852 181109 528886
rect 181040 528816 181109 528852
rect 181139 528862 181249 528900
rect 181139 528828 181205 528862
rect 181239 528828 181249 528862
rect 181139 528816 181249 528828
rect 181279 528878 181346 528900
rect 181279 528844 181302 528878
rect 181336 528844 181346 528878
rect 181279 528816 181346 528844
rect 181376 528862 181428 528900
rect 181376 528828 181386 528862
rect 181420 528828 181428 528862
rect 181376 528816 181428 528828
rect 181491 528888 181543 528900
rect 181491 528854 181499 528888
rect 181533 528854 181543 528888
rect 180681 528778 180691 528812
rect 180725 528778 180733 528812
rect 180681 528766 180733 528778
rect 180409 528742 180461 528765
rect 181491 528732 181543 528854
rect 181573 528880 181642 528900
rect 181573 528846 181587 528880
rect 181621 528846 181642 528880
rect 181573 528816 181642 528846
rect 181672 528887 181728 528900
rect 181672 528853 181684 528887
rect 181718 528853 181728 528887
rect 181672 528816 181728 528853
rect 181758 528816 181812 528900
rect 181842 528888 181920 528900
rect 181842 528854 181876 528888
rect 181910 528854 181920 528888
rect 181842 528816 181920 528854
rect 181950 528862 182004 528900
rect 181950 528828 181960 528862
rect 181994 528828 182004 528862
rect 181950 528816 182004 528828
rect 182034 528888 182088 528900
rect 182034 528854 182046 528888
rect 182080 528854 182088 528888
rect 182034 528816 182088 528854
rect 182153 528888 182219 528900
rect 182153 528854 182175 528888
rect 182209 528854 182219 528888
rect 182153 528820 182219 528854
rect 181573 528732 181627 528816
rect 182153 528786 182175 528820
rect 182209 528786 182219 528820
rect 182153 528772 182219 528786
rect 182169 528700 182219 528772
rect 182249 528852 182301 528900
rect 182631 528888 182683 528900
rect 182249 528818 182259 528852
rect 182293 528818 182301 528852
rect 182249 528784 182301 528818
rect 182249 528750 182259 528784
rect 182293 528750 182301 528784
rect 182249 528700 182301 528750
rect 182631 528854 182639 528888
rect 182673 528854 182683 528888
rect 182631 528726 182683 528854
rect 183629 528888 183681 528900
rect 183629 528854 183639 528888
rect 183673 528854 183681 528888
rect 183629 528726 183681 528854
rect 183735 528888 183787 528900
rect 183735 528854 183743 528888
rect 183777 528854 183787 528888
rect 183735 528726 183787 528854
rect 184733 528888 184785 528900
rect 184733 528854 184743 528888
rect 184777 528854 184785 528888
rect 184733 528726 184785 528854
rect 184839 528888 184891 528900
rect 184839 528854 184847 528888
rect 184881 528854 184891 528888
rect 184839 528726 184891 528854
rect 185837 528888 185889 528900
rect 185837 528854 185847 528888
rect 185881 528854 185889 528888
rect 185837 528726 185889 528854
rect 185943 528888 185995 528900
rect 185943 528854 185951 528888
rect 185985 528854 185995 528888
rect 185943 528726 185995 528854
rect 186941 528888 186993 528900
rect 186941 528854 186951 528888
rect 186985 528854 186993 528888
rect 186941 528726 186993 528854
rect 187231 528888 187283 528900
rect 187231 528854 187239 528888
rect 187273 528854 187283 528888
rect 187231 528793 187283 528854
rect 187231 528759 187239 528793
rect 187273 528759 187283 528793
rect 187231 528726 187283 528759
rect 187401 528888 187453 528900
rect 187401 528854 187411 528888
rect 187445 528854 187453 528888
rect 187401 528793 187453 528854
rect 187401 528759 187411 528793
rect 187445 528759 187453 528793
rect 187401 528726 187453 528759
rect 172235 528047 172287 528080
rect 172235 528013 172243 528047
rect 172277 528013 172287 528047
rect 172235 527952 172287 528013
rect 172235 527918 172243 527952
rect 172277 527918 172287 527952
rect 172235 527906 172287 527918
rect 172405 528047 172457 528080
rect 172405 528013 172415 528047
rect 172449 528013 172457 528047
rect 172405 527952 172457 528013
rect 172405 527918 172415 527952
rect 172449 527918 172457 527952
rect 172405 527906 172457 527918
rect 172511 527952 172563 528080
rect 172511 527918 172519 527952
rect 172553 527918 172563 527952
rect 172511 527906 172563 527918
rect 173509 527952 173561 528080
rect 173509 527918 173519 527952
rect 173553 527918 173561 527952
rect 173509 527906 173561 527918
rect 173615 527952 173667 528080
rect 173615 527918 173623 527952
rect 173657 527918 173667 527952
rect 173615 527906 173667 527918
rect 174613 527952 174665 528080
rect 174613 527918 174623 527952
rect 174657 527918 174665 527952
rect 174903 527952 174955 528080
rect 174613 527906 174665 527918
rect 174903 527918 174911 527952
rect 174945 527918 174955 527952
rect 174903 527906 174955 527918
rect 175901 527952 175953 528080
rect 175901 527918 175911 527952
rect 175945 527918 175953 527952
rect 175901 527906 175953 527918
rect 176099 528028 176151 528040
rect 176099 527994 176107 528028
rect 176141 527994 176151 528028
rect 176099 527960 176151 527994
rect 176099 527926 176107 527960
rect 176141 527926 176151 527960
rect 176099 527912 176151 527926
rect 176181 527976 176235 528040
rect 176181 527942 176191 527976
rect 176225 527942 176235 527976
rect 176181 527912 176235 527942
rect 176265 528028 176317 528040
rect 176265 527994 176275 528028
rect 176309 527994 176317 528028
rect 176265 527960 176317 527994
rect 176265 527926 176275 527960
rect 176309 527926 176317 527960
rect 176265 527912 176317 527926
rect 176450 527952 176502 527990
rect 176450 527918 176458 527952
rect 176492 527918 176502 527952
rect 176450 527906 176502 527918
rect 176532 527960 176594 527990
rect 176532 527926 176542 527960
rect 176576 527926 176594 527960
rect 176532 527906 176594 527926
rect 176624 527954 176693 527990
rect 176624 527920 176635 527954
rect 176669 527920 176693 527954
rect 176624 527906 176693 527920
rect 176723 527978 176833 527990
rect 176723 527944 176789 527978
rect 176823 527944 176833 527978
rect 176723 527906 176833 527944
rect 176863 527962 176930 527990
rect 176863 527928 176886 527962
rect 176920 527928 176930 527962
rect 176863 527906 176930 527928
rect 176960 527978 177012 527990
rect 176960 527944 176970 527978
rect 177004 527944 177012 527978
rect 176960 527906 177012 527944
rect 177075 527952 177127 528074
rect 177075 527918 177083 527952
rect 177117 527918 177127 527952
rect 177075 527906 177127 527918
rect 177157 527990 177211 528074
rect 177753 528034 177803 528106
rect 177737 528020 177803 528034
rect 177157 527960 177226 527990
rect 177157 527926 177171 527960
rect 177205 527926 177226 527960
rect 177157 527906 177226 527926
rect 177256 527953 177312 527990
rect 177256 527919 177268 527953
rect 177302 527919 177312 527953
rect 177256 527906 177312 527919
rect 177342 527906 177396 527990
rect 177426 527952 177504 527990
rect 177426 527918 177460 527952
rect 177494 527918 177504 527952
rect 177426 527906 177504 527918
rect 177534 527978 177588 527990
rect 177534 527944 177544 527978
rect 177578 527944 177588 527978
rect 177534 527906 177588 527944
rect 177618 527952 177672 527990
rect 177618 527918 177630 527952
rect 177664 527918 177672 527952
rect 177618 527906 177672 527918
rect 177737 527986 177759 528020
rect 177793 527986 177803 528020
rect 177737 527952 177803 527986
rect 177737 527918 177759 527952
rect 177793 527918 177803 527952
rect 177737 527906 177803 527918
rect 177833 528056 177885 528106
rect 178951 528088 179003 528106
rect 177833 528022 177843 528056
rect 177877 528022 177885 528056
rect 177833 527988 177885 528022
rect 177833 527954 177843 527988
rect 177877 527954 177885 527988
rect 177833 527906 177885 527954
rect 177939 528041 177991 528064
rect 177939 528007 177947 528041
rect 177981 528007 177991 528041
rect 177939 527960 177991 528007
rect 177939 527926 177947 527960
rect 177981 527926 177991 527960
rect 177939 527906 177991 527926
rect 178021 528028 178079 528064
rect 178021 527994 178033 528028
rect 178067 527994 178079 528028
rect 178021 527960 178079 527994
rect 178021 527926 178033 527960
rect 178067 527926 178079 527960
rect 178021 527906 178079 527926
rect 178109 528028 178161 528064
rect 178109 527994 178119 528028
rect 178153 527994 178161 528028
rect 178109 527960 178161 527994
rect 178109 527926 178119 527960
rect 178153 527926 178161 527960
rect 178109 527906 178161 527926
rect 178215 528054 178267 528080
rect 178215 528020 178223 528054
rect 178257 528020 178267 528054
rect 178215 527952 178267 528020
rect 178215 527918 178223 527952
rect 178257 527918 178267 527952
rect 178215 527906 178267 527918
rect 178845 528054 178897 528080
rect 178845 528020 178855 528054
rect 178889 528020 178897 528054
rect 178845 527952 178897 528020
rect 178845 527918 178855 527952
rect 178889 527918 178897 527952
rect 178845 527906 178897 527918
rect 178951 528054 178959 528088
rect 178993 528054 179003 528088
rect 178951 528020 179003 528054
rect 178951 527986 178959 528020
rect 178993 527986 179003 528020
rect 178951 527952 179003 527986
rect 178951 527918 178959 527952
rect 178993 527918 179003 527952
rect 178951 527906 179003 527918
rect 179033 528088 179085 528106
rect 179033 528054 179043 528088
rect 179077 528054 179085 528088
rect 179033 528029 179085 528054
rect 180975 528088 181027 528106
rect 179033 528020 179112 528029
rect 179033 527986 179043 528020
rect 179077 527986 179112 528020
rect 179033 527952 179112 527986
rect 179033 527918 179043 527952
rect 179077 527945 179112 527952
rect 179142 527945 179215 528029
rect 179245 528012 179429 528029
rect 179245 527978 179279 528012
rect 179313 527978 179354 528012
rect 179388 527978 179429 528012
rect 179245 527945 179429 527978
rect 179459 527945 179501 528029
rect 179531 528012 179597 528029
rect 179531 527978 179551 528012
rect 179585 527978 179597 528012
rect 179531 527945 179597 527978
rect 179627 528012 179683 528029
rect 179627 527978 179637 528012
rect 179671 527978 179683 528012
rect 179627 527945 179683 527978
rect 179077 527918 179085 527945
rect 180055 528054 180107 528080
rect 180055 528020 180063 528054
rect 180097 528020 180107 528054
rect 180055 527952 180107 528020
rect 179033 527906 179085 527918
rect 180055 527918 180063 527952
rect 180097 527918 180107 527952
rect 180055 527906 180107 527918
rect 180685 528054 180737 528080
rect 180685 528020 180695 528054
rect 180729 528020 180737 528054
rect 180685 527952 180737 528020
rect 180685 527918 180695 527952
rect 180729 527918 180737 527952
rect 180685 527906 180737 527918
rect 180975 528054 180983 528088
rect 181017 528054 181027 528088
rect 180975 528020 181027 528054
rect 180975 527986 180983 528020
rect 181017 527986 181027 528020
rect 180975 527952 181027 527986
rect 180975 527918 180983 527952
rect 181017 527918 181027 527952
rect 180975 527906 181027 527918
rect 181057 528088 181109 528106
rect 181057 528054 181067 528088
rect 181101 528054 181109 528088
rect 181057 528029 181109 528054
rect 181057 528020 181136 528029
rect 181057 527986 181067 528020
rect 181101 527986 181136 528020
rect 181057 527952 181136 527986
rect 181057 527918 181067 527952
rect 181101 527945 181136 527952
rect 181166 527945 181239 528029
rect 181269 528012 181453 528029
rect 181269 527978 181303 528012
rect 181337 527978 181378 528012
rect 181412 527978 181453 528012
rect 181269 527945 181453 527978
rect 181483 527945 181525 528029
rect 181555 528012 181621 528029
rect 181555 527978 181575 528012
rect 181609 527978 181621 528012
rect 181555 527945 181621 527978
rect 181651 528012 181707 528029
rect 181651 527978 181661 528012
rect 181695 527978 181707 528012
rect 181651 527945 181707 527978
rect 181803 527952 181855 528080
rect 181101 527918 181109 527945
rect 181057 527906 181109 527918
rect 181803 527918 181811 527952
rect 181845 527918 181855 527952
rect 181803 527906 181855 527918
rect 182801 527952 182853 528080
rect 182801 527918 182811 527952
rect 182845 527918 182853 527952
rect 182801 527906 182853 527918
rect 182907 527952 182959 528080
rect 182907 527918 182915 527952
rect 182949 527918 182959 527952
rect 182907 527906 182959 527918
rect 183905 527952 183957 528080
rect 183905 527918 183915 527952
rect 183949 527918 183957 527952
rect 183905 527906 183957 527918
rect 184011 527952 184063 528080
rect 184011 527918 184019 527952
rect 184053 527918 184063 527952
rect 184011 527906 184063 527918
rect 185009 527952 185061 528080
rect 185009 527918 185019 527952
rect 185053 527918 185061 527952
rect 185207 527952 185259 528080
rect 185009 527906 185061 527918
rect 185207 527918 185215 527952
rect 185249 527918 185259 527952
rect 185207 527906 185259 527918
rect 186205 527952 186257 528080
rect 186205 527918 186215 527952
rect 186249 527918 186257 527952
rect 186205 527906 186257 527918
rect 186311 528054 186363 528080
rect 186311 528020 186319 528054
rect 186353 528020 186363 528054
rect 186311 527952 186363 528020
rect 186311 527918 186319 527952
rect 186353 527918 186363 527952
rect 186311 527906 186363 527918
rect 186941 528054 186993 528080
rect 186941 528020 186951 528054
rect 186985 528020 186993 528054
rect 186941 527952 186993 528020
rect 186941 527918 186951 527952
rect 186985 527918 186993 527952
rect 186941 527906 186993 527918
rect 187231 528047 187283 528080
rect 187231 528013 187239 528047
rect 187273 528013 187283 528047
rect 187231 527952 187283 528013
rect 187231 527918 187239 527952
rect 187273 527918 187283 527952
rect 187231 527906 187283 527918
rect 187401 528047 187453 528080
rect 187401 528013 187411 528047
rect 187445 528013 187453 528047
rect 187401 527952 187453 528013
rect 187401 527918 187411 527952
rect 187445 527918 187453 527952
rect 187401 527906 187453 527918
rect 172235 527800 172287 527812
rect 172235 527766 172243 527800
rect 172277 527766 172287 527800
rect 172235 527705 172287 527766
rect 172235 527671 172243 527705
rect 172277 527671 172287 527705
rect 172235 527638 172287 527671
rect 172405 527800 172457 527812
rect 172405 527766 172415 527800
rect 172449 527766 172457 527800
rect 172405 527705 172457 527766
rect 172405 527671 172415 527705
rect 172449 527671 172457 527705
rect 172405 527638 172457 527671
rect 172511 527800 172563 527812
rect 172511 527766 172519 527800
rect 172553 527766 172563 527800
rect 172511 527638 172563 527766
rect 173509 527800 173561 527812
rect 173509 527766 173519 527800
rect 173553 527766 173561 527800
rect 173509 527638 173561 527766
rect 173615 527800 173667 527812
rect 173615 527766 173623 527800
rect 173657 527766 173667 527800
rect 173615 527638 173667 527766
rect 174613 527800 174665 527812
rect 174613 527766 174623 527800
rect 174657 527766 174665 527800
rect 174613 527638 174665 527766
rect 174719 527800 174771 527812
rect 174719 527766 174727 527800
rect 174761 527766 174771 527800
rect 174719 527638 174771 527766
rect 175717 527800 175769 527812
rect 175717 527766 175727 527800
rect 175761 527766 175769 527800
rect 175717 527638 175769 527766
rect 175823 527800 175875 527812
rect 175823 527766 175831 527800
rect 175865 527766 175875 527800
rect 175823 527698 175875 527766
rect 175823 527664 175831 527698
rect 175865 527664 175875 527698
rect 175823 527638 175875 527664
rect 176269 527800 176321 527812
rect 176269 527766 176279 527800
rect 176313 527766 176321 527800
rect 176269 527698 176321 527766
rect 176269 527664 176279 527698
rect 176313 527664 176321 527698
rect 176269 527638 176321 527664
rect 176394 527774 176446 527812
rect 176394 527740 176402 527774
rect 176436 527740 176446 527774
rect 176394 527612 176446 527740
rect 176476 527800 176541 527812
rect 176476 527766 176492 527800
rect 176526 527766 176541 527800
rect 176476 527728 176541 527766
rect 176641 527774 176693 527812
rect 176641 527740 176651 527774
rect 176685 527740 176693 527774
rect 176641 527728 176693 527740
rect 176747 527774 176799 527812
rect 176747 527740 176755 527774
rect 176789 527740 176799 527774
rect 176747 527728 176799 527740
rect 176899 527800 176953 527812
rect 176899 527766 176909 527800
rect 176943 527766 176953 527800
rect 176899 527728 176953 527766
rect 176983 527774 177035 527812
rect 176983 527740 176993 527774
rect 177027 527740 177035 527774
rect 176983 527728 177035 527740
rect 177111 527800 177163 527812
rect 177111 527766 177119 527800
rect 177153 527766 177163 527800
rect 176476 527612 176526 527728
rect 177111 527705 177163 527766
rect 177111 527671 177119 527705
rect 177153 527671 177163 527705
rect 177111 527638 177163 527671
rect 177281 527800 177333 527812
rect 177281 527766 177291 527800
rect 177325 527766 177333 527800
rect 177479 527800 177531 527812
rect 177281 527705 177333 527766
rect 177281 527671 177291 527705
rect 177325 527671 177333 527705
rect 177281 527638 177333 527671
rect 177479 527766 177487 527800
rect 177521 527766 177531 527800
rect 177479 527638 177531 527766
rect 178477 527800 178529 527812
rect 178477 527766 178487 527800
rect 178521 527766 178529 527800
rect 178477 527638 178529 527766
rect 178583 527800 178635 527812
rect 178583 527766 178591 527800
rect 178625 527766 178635 527800
rect 178583 527698 178635 527766
rect 178583 527664 178591 527698
rect 178625 527664 178635 527698
rect 178583 527638 178635 527664
rect 178845 527800 178897 527812
rect 178845 527766 178855 527800
rect 178889 527766 178897 527800
rect 178845 527698 178897 527766
rect 178845 527664 178855 527698
rect 178889 527664 178897 527698
rect 178845 527638 178897 527664
rect 178970 527774 179022 527812
rect 178970 527740 178978 527774
rect 179012 527740 179022 527774
rect 178970 527612 179022 527740
rect 179052 527800 179117 527812
rect 179052 527766 179068 527800
rect 179102 527766 179117 527800
rect 179052 527728 179117 527766
rect 179217 527774 179269 527812
rect 179217 527740 179227 527774
rect 179261 527740 179269 527774
rect 179217 527728 179269 527740
rect 179323 527774 179375 527812
rect 179323 527740 179331 527774
rect 179365 527740 179375 527774
rect 179323 527728 179375 527740
rect 179475 527800 179529 527812
rect 179475 527766 179485 527800
rect 179519 527766 179529 527800
rect 179475 527728 179529 527766
rect 179559 527774 179611 527812
rect 179559 527740 179569 527774
rect 179603 527740 179611 527774
rect 179559 527728 179611 527740
rect 179687 527800 179739 527812
rect 179687 527766 179695 527800
rect 179729 527766 179739 527800
rect 179052 527612 179102 527728
rect 179687 527638 179739 527766
rect 180685 527800 180737 527812
rect 180685 527766 180695 527800
rect 180729 527766 180737 527800
rect 180685 527638 180737 527766
rect 180791 527800 180843 527812
rect 180791 527766 180799 527800
rect 180833 527766 180843 527800
rect 180791 527638 180843 527766
rect 181789 527800 181841 527812
rect 181789 527766 181799 527800
rect 181833 527766 181841 527800
rect 181789 527638 181841 527766
rect 181895 527800 181947 527812
rect 181895 527766 181903 527800
rect 181937 527766 181947 527800
rect 181895 527698 181947 527766
rect 181895 527664 181903 527698
rect 181937 527664 181947 527698
rect 181895 527638 181947 527664
rect 182341 527800 182393 527812
rect 182341 527766 182351 527800
rect 182385 527766 182393 527800
rect 182631 527800 182683 527812
rect 182341 527698 182393 527766
rect 182341 527664 182351 527698
rect 182385 527664 182393 527698
rect 182341 527638 182393 527664
rect 182631 527766 182639 527800
rect 182673 527766 182683 527800
rect 182631 527638 182683 527766
rect 183629 527800 183681 527812
rect 183629 527766 183639 527800
rect 183673 527766 183681 527800
rect 183629 527638 183681 527766
rect 183735 527800 183787 527812
rect 183735 527766 183743 527800
rect 183777 527766 183787 527800
rect 183735 527638 183787 527766
rect 184733 527800 184785 527812
rect 184733 527766 184743 527800
rect 184777 527766 184785 527800
rect 184733 527638 184785 527766
rect 184839 527800 184891 527812
rect 184839 527766 184847 527800
rect 184881 527766 184891 527800
rect 184839 527638 184891 527766
rect 185837 527800 185889 527812
rect 185837 527766 185847 527800
rect 185881 527766 185889 527800
rect 185837 527638 185889 527766
rect 185943 527800 185995 527812
rect 185943 527766 185951 527800
rect 185985 527766 185995 527800
rect 185943 527638 185995 527766
rect 186941 527800 186993 527812
rect 186941 527766 186951 527800
rect 186985 527766 186993 527800
rect 186941 527638 186993 527766
rect 187231 527800 187283 527812
rect 187231 527766 187239 527800
rect 187273 527766 187283 527800
rect 187231 527705 187283 527766
rect 187231 527671 187239 527705
rect 187273 527671 187283 527705
rect 187231 527638 187283 527671
rect 187401 527800 187453 527812
rect 187401 527766 187411 527800
rect 187445 527766 187453 527800
rect 187401 527705 187453 527766
rect 187401 527671 187411 527705
rect 187445 527671 187453 527705
rect 187401 527638 187453 527671
rect 172235 526959 172287 526992
rect 172235 526925 172243 526959
rect 172277 526925 172287 526959
rect 172235 526864 172287 526925
rect 172235 526830 172243 526864
rect 172277 526830 172287 526864
rect 172235 526818 172287 526830
rect 172405 526959 172457 526992
rect 172405 526925 172415 526959
rect 172449 526925 172457 526959
rect 172405 526864 172457 526925
rect 172405 526830 172415 526864
rect 172449 526830 172457 526864
rect 172405 526818 172457 526830
rect 172511 526864 172563 526992
rect 172511 526830 172519 526864
rect 172553 526830 172563 526864
rect 172511 526818 172563 526830
rect 173509 526864 173561 526992
rect 173509 526830 173519 526864
rect 173553 526830 173561 526864
rect 173509 526818 173561 526830
rect 173615 526864 173667 526992
rect 173615 526830 173623 526864
rect 173657 526830 173667 526864
rect 173615 526818 173667 526830
rect 174613 526864 174665 526992
rect 174613 526830 174623 526864
rect 174657 526830 174665 526864
rect 174903 526864 174955 526992
rect 174613 526818 174665 526830
rect 174903 526830 174911 526864
rect 174945 526830 174955 526864
rect 174903 526818 174955 526830
rect 175901 526864 175953 526992
rect 175901 526830 175911 526864
rect 175945 526830 175953 526864
rect 175901 526818 175953 526830
rect 176007 526864 176059 526992
rect 176007 526830 176015 526864
rect 176049 526830 176059 526864
rect 176007 526818 176059 526830
rect 177005 526864 177057 526992
rect 177005 526830 177015 526864
rect 177049 526830 177057 526864
rect 177005 526818 177057 526830
rect 177111 526864 177163 526992
rect 177111 526830 177119 526864
rect 177153 526830 177163 526864
rect 177111 526818 177163 526830
rect 178109 526864 178161 526992
rect 178109 526830 178119 526864
rect 178153 526830 178161 526864
rect 178109 526818 178161 526830
rect 178215 526864 178267 526992
rect 178215 526830 178223 526864
rect 178257 526830 178267 526864
rect 178215 526818 178267 526830
rect 179213 526864 179265 526992
rect 179213 526830 179223 526864
rect 179257 526830 179265 526864
rect 179213 526818 179265 526830
rect 179319 526966 179371 526992
rect 179319 526932 179327 526966
rect 179361 526932 179371 526966
rect 179319 526864 179371 526932
rect 179319 526830 179327 526864
rect 179361 526830 179371 526864
rect 179319 526818 179371 526830
rect 179765 526966 179817 526992
rect 179765 526932 179775 526966
rect 179809 526932 179817 526966
rect 179765 526864 179817 526932
rect 179765 526830 179775 526864
rect 179809 526830 179817 526864
rect 180055 526864 180107 526992
rect 179765 526818 179817 526830
rect 180055 526830 180063 526864
rect 180097 526830 180107 526864
rect 180055 526818 180107 526830
rect 181053 526864 181105 526992
rect 181053 526830 181063 526864
rect 181097 526830 181105 526864
rect 181053 526818 181105 526830
rect 181159 526864 181211 526992
rect 181159 526830 181167 526864
rect 181201 526830 181211 526864
rect 181159 526818 181211 526830
rect 182157 526864 182209 526992
rect 182157 526830 182167 526864
rect 182201 526830 182209 526864
rect 182157 526818 182209 526830
rect 182263 526864 182315 526992
rect 182263 526830 182271 526864
rect 182305 526830 182315 526864
rect 182263 526818 182315 526830
rect 183261 526864 183313 526992
rect 183261 526830 183271 526864
rect 183305 526830 183313 526864
rect 183261 526818 183313 526830
rect 183367 526864 183419 526992
rect 183367 526830 183375 526864
rect 183409 526830 183419 526864
rect 183367 526818 183419 526830
rect 184365 526864 184417 526992
rect 184365 526830 184375 526864
rect 184409 526830 184417 526864
rect 184365 526818 184417 526830
rect 184471 526966 184523 526992
rect 184471 526932 184479 526966
rect 184513 526932 184523 526966
rect 184471 526864 184523 526932
rect 184471 526830 184479 526864
rect 184513 526830 184523 526864
rect 184471 526818 184523 526830
rect 184917 526966 184969 526992
rect 184917 526932 184927 526966
rect 184961 526932 184969 526966
rect 184917 526864 184969 526932
rect 184917 526830 184927 526864
rect 184961 526830 184969 526864
rect 185207 526864 185259 526992
rect 184917 526818 184969 526830
rect 185207 526830 185215 526864
rect 185249 526830 185259 526864
rect 185207 526818 185259 526830
rect 186205 526864 186257 526992
rect 186205 526830 186215 526864
rect 186249 526830 186257 526864
rect 186205 526818 186257 526830
rect 186311 526966 186363 526992
rect 186311 526932 186319 526966
rect 186353 526932 186363 526966
rect 186311 526864 186363 526932
rect 186311 526830 186319 526864
rect 186353 526830 186363 526864
rect 186311 526818 186363 526830
rect 186941 526966 186993 526992
rect 186941 526932 186951 526966
rect 186985 526932 186993 526966
rect 186941 526864 186993 526932
rect 186941 526830 186951 526864
rect 186985 526830 186993 526864
rect 186941 526818 186993 526830
rect 187231 526959 187283 526992
rect 187231 526925 187239 526959
rect 187273 526925 187283 526959
rect 187231 526864 187283 526925
rect 187231 526830 187239 526864
rect 187273 526830 187283 526864
rect 187231 526818 187283 526830
rect 187401 526959 187453 526992
rect 187401 526925 187411 526959
rect 187445 526925 187453 526959
rect 187401 526864 187453 526925
rect 187401 526830 187411 526864
rect 187445 526830 187453 526864
rect 187401 526818 187453 526830
rect 172235 526712 172287 526724
rect 172235 526678 172243 526712
rect 172277 526678 172287 526712
rect 172235 526617 172287 526678
rect 172235 526583 172243 526617
rect 172277 526583 172287 526617
rect 172235 526550 172287 526583
rect 172405 526712 172457 526724
rect 172405 526678 172415 526712
rect 172449 526678 172457 526712
rect 172405 526617 172457 526678
rect 172405 526583 172415 526617
rect 172449 526583 172457 526617
rect 172405 526550 172457 526583
rect 172511 526712 172563 526724
rect 172511 526678 172519 526712
rect 172553 526678 172563 526712
rect 172511 526550 172563 526678
rect 173509 526712 173561 526724
rect 173509 526678 173519 526712
rect 173553 526678 173561 526712
rect 173509 526550 173561 526678
rect 173615 526712 173667 526724
rect 173615 526678 173623 526712
rect 173657 526678 173667 526712
rect 173615 526550 173667 526678
rect 174613 526712 174665 526724
rect 174613 526678 174623 526712
rect 174657 526678 174665 526712
rect 174613 526550 174665 526678
rect 174719 526712 174771 526724
rect 174719 526678 174727 526712
rect 174761 526678 174771 526712
rect 174719 526550 174771 526678
rect 175717 526712 175769 526724
rect 175717 526678 175727 526712
rect 175761 526678 175769 526712
rect 175717 526550 175769 526678
rect 175823 526712 175875 526724
rect 175823 526678 175831 526712
rect 175865 526678 175875 526712
rect 175823 526550 175875 526678
rect 176821 526712 176873 526724
rect 176821 526678 176831 526712
rect 176865 526678 176873 526712
rect 176821 526550 176873 526678
rect 176927 526712 176979 526724
rect 176927 526678 176935 526712
rect 176969 526678 176979 526712
rect 176927 526610 176979 526678
rect 176927 526576 176935 526610
rect 176969 526576 176979 526610
rect 176927 526550 176979 526576
rect 177189 526712 177241 526724
rect 177189 526678 177199 526712
rect 177233 526678 177241 526712
rect 177479 526712 177531 526724
rect 177189 526610 177241 526678
rect 177189 526576 177199 526610
rect 177233 526576 177241 526610
rect 177189 526550 177241 526576
rect 177479 526678 177487 526712
rect 177521 526678 177531 526712
rect 177479 526550 177531 526678
rect 178477 526712 178529 526724
rect 178477 526678 178487 526712
rect 178521 526678 178529 526712
rect 178477 526550 178529 526678
rect 178583 526712 178635 526724
rect 178583 526678 178591 526712
rect 178625 526678 178635 526712
rect 178583 526550 178635 526678
rect 179581 526712 179633 526724
rect 179581 526678 179591 526712
rect 179625 526678 179633 526712
rect 179581 526550 179633 526678
rect 179687 526712 179739 526724
rect 179687 526678 179695 526712
rect 179729 526678 179739 526712
rect 179687 526550 179739 526678
rect 180685 526712 180737 526724
rect 180685 526678 180695 526712
rect 180729 526678 180737 526712
rect 180685 526550 180737 526678
rect 180791 526712 180843 526724
rect 180791 526678 180799 526712
rect 180833 526678 180843 526712
rect 180791 526550 180843 526678
rect 181789 526712 181841 526724
rect 181789 526678 181799 526712
rect 181833 526678 181841 526712
rect 181789 526550 181841 526678
rect 181895 526712 181947 526724
rect 181895 526678 181903 526712
rect 181937 526678 181947 526712
rect 181895 526610 181947 526678
rect 181895 526576 181903 526610
rect 181937 526576 181947 526610
rect 181895 526550 181947 526576
rect 182341 526712 182393 526724
rect 182341 526678 182351 526712
rect 182385 526678 182393 526712
rect 182631 526712 182683 526724
rect 182341 526610 182393 526678
rect 182341 526576 182351 526610
rect 182385 526576 182393 526610
rect 182341 526550 182393 526576
rect 182631 526678 182639 526712
rect 182673 526678 182683 526712
rect 182631 526550 182683 526678
rect 183629 526712 183681 526724
rect 183629 526678 183639 526712
rect 183673 526678 183681 526712
rect 183629 526550 183681 526678
rect 183735 526712 183787 526724
rect 183735 526678 183743 526712
rect 183777 526678 183787 526712
rect 183735 526550 183787 526678
rect 184733 526712 184785 526724
rect 184733 526678 184743 526712
rect 184777 526678 184785 526712
rect 184733 526550 184785 526678
rect 184839 526712 184891 526724
rect 184839 526678 184847 526712
rect 184881 526678 184891 526712
rect 184839 526550 184891 526678
rect 185837 526712 185889 526724
rect 185837 526678 185847 526712
rect 185881 526678 185889 526712
rect 185837 526550 185889 526678
rect 185943 526712 185995 526724
rect 185943 526678 185951 526712
rect 185985 526678 185995 526712
rect 185943 526550 185995 526678
rect 186941 526712 186993 526724
rect 186941 526678 186951 526712
rect 186985 526678 186993 526712
rect 186941 526550 186993 526678
rect 187231 526712 187283 526724
rect 187231 526678 187239 526712
rect 187273 526678 187283 526712
rect 187231 526617 187283 526678
rect 187231 526583 187239 526617
rect 187273 526583 187283 526617
rect 187231 526550 187283 526583
rect 187401 526712 187453 526724
rect 187401 526678 187411 526712
rect 187445 526678 187453 526712
rect 187401 526617 187453 526678
rect 187401 526583 187411 526617
rect 187445 526583 187453 526617
rect 187401 526550 187453 526583
rect 172235 525871 172287 525904
rect 172235 525837 172243 525871
rect 172277 525837 172287 525871
rect 172235 525776 172287 525837
rect 172235 525742 172243 525776
rect 172277 525742 172287 525776
rect 172235 525730 172287 525742
rect 172405 525871 172457 525904
rect 172405 525837 172415 525871
rect 172449 525837 172457 525871
rect 172405 525776 172457 525837
rect 172405 525742 172415 525776
rect 172449 525742 172457 525776
rect 172405 525730 172457 525742
rect 172511 525776 172563 525904
rect 172511 525742 172519 525776
rect 172553 525742 172563 525776
rect 172511 525730 172563 525742
rect 173509 525776 173561 525904
rect 173509 525742 173519 525776
rect 173553 525742 173561 525776
rect 173509 525730 173561 525742
rect 173615 525776 173667 525904
rect 173615 525742 173623 525776
rect 173657 525742 173667 525776
rect 173615 525730 173667 525742
rect 174613 525776 174665 525904
rect 174613 525742 174623 525776
rect 174657 525742 174665 525776
rect 174903 525776 174955 525904
rect 174613 525730 174665 525742
rect 174903 525742 174911 525776
rect 174945 525742 174955 525776
rect 174903 525730 174955 525742
rect 175901 525776 175953 525904
rect 175901 525742 175911 525776
rect 175945 525742 175953 525776
rect 175901 525730 175953 525742
rect 176007 525776 176059 525904
rect 176007 525742 176015 525776
rect 176049 525742 176059 525776
rect 176007 525730 176059 525742
rect 177005 525776 177057 525904
rect 177005 525742 177015 525776
rect 177049 525742 177057 525776
rect 177005 525730 177057 525742
rect 177111 525776 177163 525904
rect 177111 525742 177119 525776
rect 177153 525742 177163 525776
rect 177111 525730 177163 525742
rect 178109 525776 178161 525904
rect 178109 525742 178119 525776
rect 178153 525742 178161 525776
rect 178109 525730 178161 525742
rect 178215 525776 178267 525904
rect 178215 525742 178223 525776
rect 178257 525742 178267 525776
rect 178215 525730 178267 525742
rect 179213 525776 179265 525904
rect 179213 525742 179223 525776
rect 179257 525742 179265 525776
rect 179213 525730 179265 525742
rect 179319 525878 179371 525904
rect 179319 525844 179327 525878
rect 179361 525844 179371 525878
rect 179319 525776 179371 525844
rect 179319 525742 179327 525776
rect 179361 525742 179371 525776
rect 179319 525730 179371 525742
rect 179765 525878 179817 525904
rect 179765 525844 179775 525878
rect 179809 525844 179817 525878
rect 179765 525776 179817 525844
rect 179765 525742 179775 525776
rect 179809 525742 179817 525776
rect 180055 525776 180107 525904
rect 179765 525730 179817 525742
rect 180055 525742 180063 525776
rect 180097 525742 180107 525776
rect 180055 525730 180107 525742
rect 181053 525776 181105 525904
rect 181053 525742 181063 525776
rect 181097 525742 181105 525776
rect 181053 525730 181105 525742
rect 181159 525776 181211 525904
rect 181159 525742 181167 525776
rect 181201 525742 181211 525776
rect 181159 525730 181211 525742
rect 182157 525776 182209 525904
rect 182157 525742 182167 525776
rect 182201 525742 182209 525776
rect 182157 525730 182209 525742
rect 182263 525776 182315 525904
rect 182263 525742 182271 525776
rect 182305 525742 182315 525776
rect 182263 525730 182315 525742
rect 183261 525776 183313 525904
rect 183261 525742 183271 525776
rect 183305 525742 183313 525776
rect 183261 525730 183313 525742
rect 183367 525776 183419 525904
rect 183367 525742 183375 525776
rect 183409 525742 183419 525776
rect 183367 525730 183419 525742
rect 184365 525776 184417 525904
rect 184365 525742 184375 525776
rect 184409 525742 184417 525776
rect 184365 525730 184417 525742
rect 184471 525878 184523 525904
rect 184471 525844 184479 525878
rect 184513 525844 184523 525878
rect 184471 525776 184523 525844
rect 184471 525742 184479 525776
rect 184513 525742 184523 525776
rect 184471 525730 184523 525742
rect 184917 525878 184969 525904
rect 184917 525844 184927 525878
rect 184961 525844 184969 525878
rect 184917 525776 184969 525844
rect 184917 525742 184927 525776
rect 184961 525742 184969 525776
rect 185207 525776 185259 525904
rect 184917 525730 184969 525742
rect 185207 525742 185215 525776
rect 185249 525742 185259 525776
rect 185207 525730 185259 525742
rect 186205 525776 186257 525904
rect 186205 525742 186215 525776
rect 186249 525742 186257 525776
rect 186205 525730 186257 525742
rect 186311 525878 186363 525904
rect 186311 525844 186319 525878
rect 186353 525844 186363 525878
rect 186311 525776 186363 525844
rect 186311 525742 186319 525776
rect 186353 525742 186363 525776
rect 186311 525730 186363 525742
rect 186941 525878 186993 525904
rect 186941 525844 186951 525878
rect 186985 525844 186993 525878
rect 186941 525776 186993 525844
rect 186941 525742 186951 525776
rect 186985 525742 186993 525776
rect 186941 525730 186993 525742
rect 187231 525871 187283 525904
rect 187231 525837 187239 525871
rect 187273 525837 187283 525871
rect 187231 525776 187283 525837
rect 187231 525742 187239 525776
rect 187273 525742 187283 525776
rect 187231 525730 187283 525742
rect 187401 525871 187453 525904
rect 187401 525837 187411 525871
rect 187445 525837 187453 525871
rect 187401 525776 187453 525837
rect 187401 525742 187411 525776
rect 187445 525742 187453 525776
rect 187401 525730 187453 525742
rect 172235 525624 172287 525636
rect 172235 525590 172243 525624
rect 172277 525590 172287 525624
rect 172235 525529 172287 525590
rect 172235 525495 172243 525529
rect 172277 525495 172287 525529
rect 172235 525462 172287 525495
rect 172405 525624 172457 525636
rect 172405 525590 172415 525624
rect 172449 525590 172457 525624
rect 172405 525529 172457 525590
rect 172405 525495 172415 525529
rect 172449 525495 172457 525529
rect 172405 525462 172457 525495
rect 172511 525624 172563 525636
rect 172511 525590 172519 525624
rect 172553 525590 172563 525624
rect 172511 525462 172563 525590
rect 173509 525624 173561 525636
rect 173509 525590 173519 525624
rect 173553 525590 173561 525624
rect 173509 525462 173561 525590
rect 173615 525624 173667 525636
rect 173615 525590 173623 525624
rect 173657 525590 173667 525624
rect 173615 525462 173667 525590
rect 174613 525624 174665 525636
rect 174613 525590 174623 525624
rect 174657 525590 174665 525624
rect 174613 525462 174665 525590
rect 174719 525624 174771 525636
rect 174719 525590 174727 525624
rect 174761 525590 174771 525624
rect 174719 525462 174771 525590
rect 175717 525624 175769 525636
rect 175717 525590 175727 525624
rect 175761 525590 175769 525624
rect 175717 525462 175769 525590
rect 175823 525624 175875 525636
rect 175823 525590 175831 525624
rect 175865 525590 175875 525624
rect 175823 525462 175875 525590
rect 176821 525624 176873 525636
rect 176821 525590 176831 525624
rect 176865 525590 176873 525624
rect 176821 525462 176873 525590
rect 176927 525624 176979 525636
rect 176927 525590 176935 525624
rect 176969 525590 176979 525624
rect 176927 525522 176979 525590
rect 176927 525488 176935 525522
rect 176969 525488 176979 525522
rect 176927 525462 176979 525488
rect 177189 525624 177241 525636
rect 177189 525590 177199 525624
rect 177233 525590 177241 525624
rect 177479 525624 177531 525636
rect 177189 525522 177241 525590
rect 177189 525488 177199 525522
rect 177233 525488 177241 525522
rect 177189 525462 177241 525488
rect 177479 525590 177487 525624
rect 177521 525590 177531 525624
rect 177479 525462 177531 525590
rect 178477 525624 178529 525636
rect 178477 525590 178487 525624
rect 178521 525590 178529 525624
rect 178477 525462 178529 525590
rect 178583 525624 178635 525636
rect 178583 525590 178591 525624
rect 178625 525590 178635 525624
rect 178583 525462 178635 525590
rect 179581 525624 179633 525636
rect 179581 525590 179591 525624
rect 179625 525590 179633 525624
rect 179581 525462 179633 525590
rect 179687 525624 179739 525636
rect 179687 525590 179695 525624
rect 179729 525590 179739 525624
rect 179687 525462 179739 525590
rect 180685 525624 180737 525636
rect 180685 525590 180695 525624
rect 180729 525590 180737 525624
rect 180685 525462 180737 525590
rect 180791 525624 180843 525636
rect 180791 525590 180799 525624
rect 180833 525590 180843 525624
rect 180791 525462 180843 525590
rect 181789 525624 181841 525636
rect 181789 525590 181799 525624
rect 181833 525590 181841 525624
rect 181789 525462 181841 525590
rect 181895 525624 181947 525636
rect 181895 525590 181903 525624
rect 181937 525590 181947 525624
rect 181895 525522 181947 525590
rect 181895 525488 181903 525522
rect 181937 525488 181947 525522
rect 181895 525462 181947 525488
rect 182341 525624 182393 525636
rect 182341 525590 182351 525624
rect 182385 525590 182393 525624
rect 182631 525624 182683 525636
rect 182341 525522 182393 525590
rect 182341 525488 182351 525522
rect 182385 525488 182393 525522
rect 182341 525462 182393 525488
rect 182631 525590 182639 525624
rect 182673 525590 182683 525624
rect 182631 525462 182683 525590
rect 183629 525624 183681 525636
rect 183629 525590 183639 525624
rect 183673 525590 183681 525624
rect 183629 525462 183681 525590
rect 183735 525624 183787 525636
rect 183735 525590 183743 525624
rect 183777 525590 183787 525624
rect 183735 525462 183787 525590
rect 184733 525624 184785 525636
rect 184733 525590 184743 525624
rect 184777 525590 184785 525624
rect 184733 525462 184785 525590
rect 184839 525624 184891 525636
rect 184839 525590 184847 525624
rect 184881 525590 184891 525624
rect 184839 525462 184891 525590
rect 185837 525624 185889 525636
rect 185837 525590 185847 525624
rect 185881 525590 185889 525624
rect 185837 525462 185889 525590
rect 185943 525624 185995 525636
rect 185943 525590 185951 525624
rect 185985 525590 185995 525624
rect 185943 525462 185995 525590
rect 186941 525624 186993 525636
rect 186941 525590 186951 525624
rect 186985 525590 186993 525624
rect 186941 525462 186993 525590
rect 187231 525624 187283 525636
rect 187231 525590 187239 525624
rect 187273 525590 187283 525624
rect 187231 525529 187283 525590
rect 187231 525495 187239 525529
rect 187273 525495 187283 525529
rect 187231 525462 187283 525495
rect 187401 525624 187453 525636
rect 187401 525590 187411 525624
rect 187445 525590 187453 525624
rect 187401 525529 187453 525590
rect 187401 525495 187411 525529
rect 187445 525495 187453 525529
rect 187401 525462 187453 525495
rect 172235 524783 172287 524816
rect 172235 524749 172243 524783
rect 172277 524749 172287 524783
rect 172235 524688 172287 524749
rect 172235 524654 172243 524688
rect 172277 524654 172287 524688
rect 172235 524642 172287 524654
rect 172405 524783 172457 524816
rect 172405 524749 172415 524783
rect 172449 524749 172457 524783
rect 172405 524688 172457 524749
rect 172405 524654 172415 524688
rect 172449 524654 172457 524688
rect 172405 524642 172457 524654
rect 172511 524688 172563 524816
rect 172511 524654 172519 524688
rect 172553 524654 172563 524688
rect 172511 524642 172563 524654
rect 173509 524688 173561 524816
rect 173509 524654 173519 524688
rect 173553 524654 173561 524688
rect 173509 524642 173561 524654
rect 173615 524688 173667 524816
rect 173615 524654 173623 524688
rect 173657 524654 173667 524688
rect 173615 524642 173667 524654
rect 174613 524688 174665 524816
rect 174613 524654 174623 524688
rect 174657 524654 174665 524688
rect 174903 524688 174955 524816
rect 174613 524642 174665 524654
rect 174903 524654 174911 524688
rect 174945 524654 174955 524688
rect 174903 524642 174955 524654
rect 175901 524688 175953 524816
rect 175901 524654 175911 524688
rect 175945 524654 175953 524688
rect 175901 524642 175953 524654
rect 176007 524688 176059 524816
rect 176007 524654 176015 524688
rect 176049 524654 176059 524688
rect 176007 524642 176059 524654
rect 177005 524688 177057 524816
rect 177005 524654 177015 524688
rect 177049 524654 177057 524688
rect 177005 524642 177057 524654
rect 177111 524688 177163 524816
rect 177111 524654 177119 524688
rect 177153 524654 177163 524688
rect 177111 524642 177163 524654
rect 178109 524688 178161 524816
rect 178109 524654 178119 524688
rect 178153 524654 178161 524688
rect 178109 524642 178161 524654
rect 178215 524688 178267 524816
rect 178215 524654 178223 524688
rect 178257 524654 178267 524688
rect 178215 524642 178267 524654
rect 179213 524688 179265 524816
rect 179213 524654 179223 524688
rect 179257 524654 179265 524688
rect 179213 524642 179265 524654
rect 179319 524790 179371 524816
rect 179319 524756 179327 524790
rect 179361 524756 179371 524790
rect 179319 524688 179371 524756
rect 179319 524654 179327 524688
rect 179361 524654 179371 524688
rect 179319 524642 179371 524654
rect 179765 524790 179817 524816
rect 179765 524756 179775 524790
rect 179809 524756 179817 524790
rect 179765 524688 179817 524756
rect 179765 524654 179775 524688
rect 179809 524654 179817 524688
rect 180055 524688 180107 524816
rect 179765 524642 179817 524654
rect 180055 524654 180063 524688
rect 180097 524654 180107 524688
rect 180055 524642 180107 524654
rect 181053 524688 181105 524816
rect 181053 524654 181063 524688
rect 181097 524654 181105 524688
rect 181053 524642 181105 524654
rect 181159 524688 181211 524816
rect 181159 524654 181167 524688
rect 181201 524654 181211 524688
rect 181159 524642 181211 524654
rect 182157 524688 182209 524816
rect 182157 524654 182167 524688
rect 182201 524654 182209 524688
rect 182157 524642 182209 524654
rect 182263 524688 182315 524816
rect 182263 524654 182271 524688
rect 182305 524654 182315 524688
rect 182263 524642 182315 524654
rect 183261 524688 183313 524816
rect 183261 524654 183271 524688
rect 183305 524654 183313 524688
rect 183261 524642 183313 524654
rect 183367 524688 183419 524816
rect 183367 524654 183375 524688
rect 183409 524654 183419 524688
rect 183367 524642 183419 524654
rect 184365 524688 184417 524816
rect 184365 524654 184375 524688
rect 184409 524654 184417 524688
rect 184365 524642 184417 524654
rect 184471 524790 184523 524816
rect 184471 524756 184479 524790
rect 184513 524756 184523 524790
rect 184471 524688 184523 524756
rect 184471 524654 184479 524688
rect 184513 524654 184523 524688
rect 184471 524642 184523 524654
rect 184917 524790 184969 524816
rect 184917 524756 184927 524790
rect 184961 524756 184969 524790
rect 184917 524688 184969 524756
rect 184917 524654 184927 524688
rect 184961 524654 184969 524688
rect 185207 524688 185259 524816
rect 184917 524642 184969 524654
rect 185207 524654 185215 524688
rect 185249 524654 185259 524688
rect 185207 524642 185259 524654
rect 186205 524688 186257 524816
rect 186205 524654 186215 524688
rect 186249 524654 186257 524688
rect 186205 524642 186257 524654
rect 186311 524790 186363 524816
rect 186311 524756 186319 524790
rect 186353 524756 186363 524790
rect 186311 524688 186363 524756
rect 186311 524654 186319 524688
rect 186353 524654 186363 524688
rect 186311 524642 186363 524654
rect 186941 524790 186993 524816
rect 186941 524756 186951 524790
rect 186985 524756 186993 524790
rect 186941 524688 186993 524756
rect 186941 524654 186951 524688
rect 186985 524654 186993 524688
rect 186941 524642 186993 524654
rect 187231 524783 187283 524816
rect 187231 524749 187239 524783
rect 187273 524749 187283 524783
rect 187231 524688 187283 524749
rect 187231 524654 187239 524688
rect 187273 524654 187283 524688
rect 187231 524642 187283 524654
rect 187401 524783 187453 524816
rect 187401 524749 187411 524783
rect 187445 524749 187453 524783
rect 187401 524688 187453 524749
rect 187401 524654 187411 524688
rect 187445 524654 187453 524688
rect 187401 524642 187453 524654
rect 172235 524536 172287 524548
rect 172235 524502 172243 524536
rect 172277 524502 172287 524536
rect 172235 524441 172287 524502
rect 172235 524407 172243 524441
rect 172277 524407 172287 524441
rect 172235 524374 172287 524407
rect 172405 524536 172457 524548
rect 172405 524502 172415 524536
rect 172449 524502 172457 524536
rect 172405 524441 172457 524502
rect 172405 524407 172415 524441
rect 172449 524407 172457 524441
rect 172405 524374 172457 524407
rect 172511 524536 172563 524548
rect 172511 524502 172519 524536
rect 172553 524502 172563 524536
rect 172511 524374 172563 524502
rect 173509 524536 173561 524548
rect 173509 524502 173519 524536
rect 173553 524502 173561 524536
rect 173509 524374 173561 524502
rect 173615 524536 173667 524548
rect 173615 524502 173623 524536
rect 173657 524502 173667 524536
rect 173615 524374 173667 524502
rect 174613 524536 174665 524548
rect 174613 524502 174623 524536
rect 174657 524502 174665 524536
rect 174613 524374 174665 524502
rect 174719 524536 174771 524548
rect 174719 524502 174727 524536
rect 174761 524502 174771 524536
rect 174719 524374 174771 524502
rect 175717 524536 175769 524548
rect 175717 524502 175727 524536
rect 175761 524502 175769 524536
rect 175717 524374 175769 524502
rect 175823 524536 175875 524548
rect 175823 524502 175831 524536
rect 175865 524502 175875 524536
rect 175823 524374 175875 524502
rect 176821 524536 176873 524548
rect 176821 524502 176831 524536
rect 176865 524502 176873 524536
rect 176821 524374 176873 524502
rect 176927 524536 176979 524548
rect 176927 524502 176935 524536
rect 176969 524502 176979 524536
rect 176927 524434 176979 524502
rect 176927 524400 176935 524434
rect 176969 524400 176979 524434
rect 176927 524374 176979 524400
rect 177189 524536 177241 524548
rect 177189 524502 177199 524536
rect 177233 524502 177241 524536
rect 177479 524536 177531 524548
rect 177189 524434 177241 524502
rect 177189 524400 177199 524434
rect 177233 524400 177241 524434
rect 177189 524374 177241 524400
rect 177479 524502 177487 524536
rect 177521 524502 177531 524536
rect 177479 524374 177531 524502
rect 178477 524536 178529 524548
rect 178477 524502 178487 524536
rect 178521 524502 178529 524536
rect 178477 524374 178529 524502
rect 178583 524536 178635 524548
rect 178583 524502 178591 524536
rect 178625 524502 178635 524536
rect 178583 524374 178635 524502
rect 179581 524536 179633 524548
rect 179581 524502 179591 524536
rect 179625 524502 179633 524536
rect 179581 524374 179633 524502
rect 179687 524536 179739 524548
rect 179687 524502 179695 524536
rect 179729 524502 179739 524536
rect 179687 524374 179739 524502
rect 180685 524536 180737 524548
rect 180685 524502 180695 524536
rect 180729 524502 180737 524536
rect 180685 524374 180737 524502
rect 180791 524536 180843 524548
rect 180791 524502 180799 524536
rect 180833 524502 180843 524536
rect 180791 524374 180843 524502
rect 181789 524536 181841 524548
rect 181789 524502 181799 524536
rect 181833 524502 181841 524536
rect 181789 524374 181841 524502
rect 181895 524536 181947 524548
rect 181895 524502 181903 524536
rect 181937 524502 181947 524536
rect 181895 524434 181947 524502
rect 181895 524400 181903 524434
rect 181937 524400 181947 524434
rect 181895 524374 181947 524400
rect 182341 524536 182393 524548
rect 182341 524502 182351 524536
rect 182385 524502 182393 524536
rect 182631 524536 182683 524548
rect 182341 524434 182393 524502
rect 182341 524400 182351 524434
rect 182385 524400 182393 524434
rect 182341 524374 182393 524400
rect 182631 524502 182639 524536
rect 182673 524502 182683 524536
rect 182631 524374 182683 524502
rect 183629 524536 183681 524548
rect 183629 524502 183639 524536
rect 183673 524502 183681 524536
rect 183629 524374 183681 524502
rect 183735 524536 183787 524548
rect 183735 524502 183743 524536
rect 183777 524502 183787 524536
rect 183735 524374 183787 524502
rect 184733 524536 184785 524548
rect 184733 524502 184743 524536
rect 184777 524502 184785 524536
rect 184733 524374 184785 524502
rect 184839 524536 184891 524548
rect 184839 524502 184847 524536
rect 184881 524502 184891 524536
rect 184839 524374 184891 524502
rect 185837 524536 185889 524548
rect 185837 524502 185847 524536
rect 185881 524502 185889 524536
rect 185837 524374 185889 524502
rect 185943 524536 185995 524548
rect 185943 524502 185951 524536
rect 185985 524502 185995 524536
rect 185943 524374 185995 524502
rect 186941 524536 186993 524548
rect 186941 524502 186951 524536
rect 186985 524502 186993 524536
rect 186941 524374 186993 524502
rect 187231 524536 187283 524548
rect 187231 524502 187239 524536
rect 187273 524502 187283 524536
rect 187231 524441 187283 524502
rect 187231 524407 187239 524441
rect 187273 524407 187283 524441
rect 187231 524374 187283 524407
rect 187401 524536 187453 524548
rect 187401 524502 187411 524536
rect 187445 524502 187453 524536
rect 187401 524441 187453 524502
rect 187401 524407 187411 524441
rect 187445 524407 187453 524441
rect 187401 524374 187453 524407
rect 172235 523695 172287 523728
rect 172235 523661 172243 523695
rect 172277 523661 172287 523695
rect 172235 523600 172287 523661
rect 172235 523566 172243 523600
rect 172277 523566 172287 523600
rect 172235 523554 172287 523566
rect 172405 523695 172457 523728
rect 172405 523661 172415 523695
rect 172449 523661 172457 523695
rect 172405 523600 172457 523661
rect 172405 523566 172415 523600
rect 172449 523566 172457 523600
rect 172405 523554 172457 523566
rect 172511 523600 172563 523728
rect 172511 523566 172519 523600
rect 172553 523566 172563 523600
rect 172511 523554 172563 523566
rect 173509 523600 173561 523728
rect 173509 523566 173519 523600
rect 173553 523566 173561 523600
rect 173509 523554 173561 523566
rect 173615 523600 173667 523728
rect 173615 523566 173623 523600
rect 173657 523566 173667 523600
rect 173615 523554 173667 523566
rect 174613 523600 174665 523728
rect 174613 523566 174623 523600
rect 174657 523566 174665 523600
rect 174903 523600 174955 523728
rect 174613 523554 174665 523566
rect 174903 523566 174911 523600
rect 174945 523566 174955 523600
rect 174903 523554 174955 523566
rect 175901 523600 175953 523728
rect 175901 523566 175911 523600
rect 175945 523566 175953 523600
rect 175901 523554 175953 523566
rect 176007 523600 176059 523728
rect 176007 523566 176015 523600
rect 176049 523566 176059 523600
rect 176007 523554 176059 523566
rect 177005 523600 177057 523728
rect 177005 523566 177015 523600
rect 177049 523566 177057 523600
rect 177005 523554 177057 523566
rect 177111 523600 177163 523728
rect 177111 523566 177119 523600
rect 177153 523566 177163 523600
rect 177111 523554 177163 523566
rect 178109 523600 178161 523728
rect 178109 523566 178119 523600
rect 178153 523566 178161 523600
rect 178109 523554 178161 523566
rect 178215 523600 178267 523728
rect 178215 523566 178223 523600
rect 178257 523566 178267 523600
rect 178215 523554 178267 523566
rect 179213 523600 179265 523728
rect 179213 523566 179223 523600
rect 179257 523566 179265 523600
rect 179213 523554 179265 523566
rect 179319 523702 179371 523728
rect 179319 523668 179327 523702
rect 179361 523668 179371 523702
rect 179319 523600 179371 523668
rect 179319 523566 179327 523600
rect 179361 523566 179371 523600
rect 179319 523554 179371 523566
rect 179765 523702 179817 523728
rect 179765 523668 179775 523702
rect 179809 523668 179817 523702
rect 179765 523600 179817 523668
rect 179765 523566 179775 523600
rect 179809 523566 179817 523600
rect 180055 523600 180107 523728
rect 179765 523554 179817 523566
rect 180055 523566 180063 523600
rect 180097 523566 180107 523600
rect 180055 523554 180107 523566
rect 181053 523600 181105 523728
rect 181053 523566 181063 523600
rect 181097 523566 181105 523600
rect 181053 523554 181105 523566
rect 181159 523600 181211 523728
rect 181159 523566 181167 523600
rect 181201 523566 181211 523600
rect 181159 523554 181211 523566
rect 182157 523600 182209 523728
rect 182157 523566 182167 523600
rect 182201 523566 182209 523600
rect 182157 523554 182209 523566
rect 182263 523600 182315 523728
rect 182263 523566 182271 523600
rect 182305 523566 182315 523600
rect 182263 523554 182315 523566
rect 183261 523600 183313 523728
rect 183261 523566 183271 523600
rect 183305 523566 183313 523600
rect 183261 523554 183313 523566
rect 183367 523600 183419 523728
rect 183367 523566 183375 523600
rect 183409 523566 183419 523600
rect 183367 523554 183419 523566
rect 184365 523600 184417 523728
rect 184365 523566 184375 523600
rect 184409 523566 184417 523600
rect 184365 523554 184417 523566
rect 184471 523702 184523 523728
rect 184471 523668 184479 523702
rect 184513 523668 184523 523702
rect 184471 523600 184523 523668
rect 184471 523566 184479 523600
rect 184513 523566 184523 523600
rect 184471 523554 184523 523566
rect 184917 523702 184969 523728
rect 184917 523668 184927 523702
rect 184961 523668 184969 523702
rect 184917 523600 184969 523668
rect 184917 523566 184927 523600
rect 184961 523566 184969 523600
rect 185207 523600 185259 523728
rect 184917 523554 184969 523566
rect 185207 523566 185215 523600
rect 185249 523566 185259 523600
rect 185207 523554 185259 523566
rect 186205 523600 186257 523728
rect 186205 523566 186215 523600
rect 186249 523566 186257 523600
rect 186205 523554 186257 523566
rect 186311 523702 186363 523728
rect 186311 523668 186319 523702
rect 186353 523668 186363 523702
rect 186311 523600 186363 523668
rect 186311 523566 186319 523600
rect 186353 523566 186363 523600
rect 186311 523554 186363 523566
rect 186941 523702 186993 523728
rect 186941 523668 186951 523702
rect 186985 523668 186993 523702
rect 186941 523600 186993 523668
rect 186941 523566 186951 523600
rect 186985 523566 186993 523600
rect 186941 523554 186993 523566
rect 187231 523695 187283 523728
rect 187231 523661 187239 523695
rect 187273 523661 187283 523695
rect 187231 523600 187283 523661
rect 187231 523566 187239 523600
rect 187273 523566 187283 523600
rect 187231 523554 187283 523566
rect 187401 523695 187453 523728
rect 187401 523661 187411 523695
rect 187445 523661 187453 523695
rect 187401 523600 187453 523661
rect 187401 523566 187411 523600
rect 187445 523566 187453 523600
rect 187401 523554 187453 523566
rect 172235 523448 172287 523460
rect 172235 523414 172243 523448
rect 172277 523414 172287 523448
rect 172235 523353 172287 523414
rect 172235 523319 172243 523353
rect 172277 523319 172287 523353
rect 172235 523286 172287 523319
rect 172405 523448 172457 523460
rect 172405 523414 172415 523448
rect 172449 523414 172457 523448
rect 172405 523353 172457 523414
rect 172405 523319 172415 523353
rect 172449 523319 172457 523353
rect 172405 523286 172457 523319
rect 172511 523448 172563 523460
rect 172511 523414 172519 523448
rect 172553 523414 172563 523448
rect 172511 523286 172563 523414
rect 173509 523448 173561 523460
rect 173509 523414 173519 523448
rect 173553 523414 173561 523448
rect 173509 523286 173561 523414
rect 173615 523448 173667 523460
rect 173615 523414 173623 523448
rect 173657 523414 173667 523448
rect 173615 523286 173667 523414
rect 174613 523448 174665 523460
rect 174613 523414 174623 523448
rect 174657 523414 174665 523448
rect 174613 523286 174665 523414
rect 174719 523448 174771 523460
rect 174719 523414 174727 523448
rect 174761 523414 174771 523448
rect 174719 523286 174771 523414
rect 175717 523448 175769 523460
rect 175717 523414 175727 523448
rect 175761 523414 175769 523448
rect 175717 523286 175769 523414
rect 175823 523448 175875 523460
rect 175823 523414 175831 523448
rect 175865 523414 175875 523448
rect 175823 523286 175875 523414
rect 176821 523448 176873 523460
rect 176821 523414 176831 523448
rect 176865 523414 176873 523448
rect 176821 523286 176873 523414
rect 176927 523448 176979 523460
rect 176927 523414 176935 523448
rect 176969 523414 176979 523448
rect 176927 523346 176979 523414
rect 176927 523312 176935 523346
rect 176969 523312 176979 523346
rect 176927 523286 176979 523312
rect 177189 523448 177241 523460
rect 177189 523414 177199 523448
rect 177233 523414 177241 523448
rect 177479 523448 177531 523460
rect 177189 523346 177241 523414
rect 177189 523312 177199 523346
rect 177233 523312 177241 523346
rect 177189 523286 177241 523312
rect 177479 523414 177487 523448
rect 177521 523414 177531 523448
rect 177479 523286 177531 523414
rect 178477 523448 178529 523460
rect 178477 523414 178487 523448
rect 178521 523414 178529 523448
rect 178477 523286 178529 523414
rect 178583 523448 178635 523460
rect 178583 523414 178591 523448
rect 178625 523414 178635 523448
rect 178583 523286 178635 523414
rect 179581 523448 179633 523460
rect 179581 523414 179591 523448
rect 179625 523414 179633 523448
rect 179581 523286 179633 523414
rect 179687 523448 179739 523460
rect 179687 523414 179695 523448
rect 179729 523414 179739 523448
rect 179687 523286 179739 523414
rect 180685 523448 180737 523460
rect 180685 523414 180695 523448
rect 180729 523414 180737 523448
rect 180685 523286 180737 523414
rect 180791 523448 180843 523460
rect 180791 523414 180799 523448
rect 180833 523414 180843 523448
rect 180791 523286 180843 523414
rect 181789 523448 181841 523460
rect 181789 523414 181799 523448
rect 181833 523414 181841 523448
rect 181789 523286 181841 523414
rect 181895 523448 181947 523460
rect 181895 523414 181903 523448
rect 181937 523414 181947 523448
rect 181895 523346 181947 523414
rect 181895 523312 181903 523346
rect 181937 523312 181947 523346
rect 181895 523286 181947 523312
rect 182341 523448 182393 523460
rect 182341 523414 182351 523448
rect 182385 523414 182393 523448
rect 182631 523448 182683 523460
rect 182341 523346 182393 523414
rect 182341 523312 182351 523346
rect 182385 523312 182393 523346
rect 182341 523286 182393 523312
rect 182631 523414 182639 523448
rect 182673 523414 182683 523448
rect 182631 523286 182683 523414
rect 183629 523448 183681 523460
rect 183629 523414 183639 523448
rect 183673 523414 183681 523448
rect 183629 523286 183681 523414
rect 183735 523448 183787 523460
rect 183735 523414 183743 523448
rect 183777 523414 183787 523448
rect 183735 523286 183787 523414
rect 184733 523448 184785 523460
rect 184733 523414 184743 523448
rect 184777 523414 184785 523448
rect 184733 523286 184785 523414
rect 184839 523448 184891 523460
rect 184839 523414 184847 523448
rect 184881 523414 184891 523448
rect 184839 523286 184891 523414
rect 185837 523448 185889 523460
rect 185837 523414 185847 523448
rect 185881 523414 185889 523448
rect 185837 523286 185889 523414
rect 185943 523448 185995 523460
rect 185943 523414 185951 523448
rect 185985 523414 185995 523448
rect 185943 523286 185995 523414
rect 186941 523448 186993 523460
rect 186941 523414 186951 523448
rect 186985 523414 186993 523448
rect 186941 523286 186993 523414
rect 187231 523448 187283 523460
rect 187231 523414 187239 523448
rect 187273 523414 187283 523448
rect 187231 523353 187283 523414
rect 187231 523319 187239 523353
rect 187273 523319 187283 523353
rect 187231 523286 187283 523319
rect 187401 523448 187453 523460
rect 187401 523414 187411 523448
rect 187445 523414 187453 523448
rect 187401 523353 187453 523414
rect 187401 523319 187411 523353
rect 187445 523319 187453 523353
rect 187401 523286 187453 523319
rect 172235 522607 172287 522640
rect 172235 522573 172243 522607
rect 172277 522573 172287 522607
rect 172235 522512 172287 522573
rect 172235 522478 172243 522512
rect 172277 522478 172287 522512
rect 172235 522466 172287 522478
rect 172405 522607 172457 522640
rect 172405 522573 172415 522607
rect 172449 522573 172457 522607
rect 172405 522512 172457 522573
rect 172405 522478 172415 522512
rect 172449 522478 172457 522512
rect 172405 522466 172457 522478
rect 172511 522512 172563 522640
rect 172511 522478 172519 522512
rect 172553 522478 172563 522512
rect 172511 522466 172563 522478
rect 173509 522512 173561 522640
rect 173509 522478 173519 522512
rect 173553 522478 173561 522512
rect 173509 522466 173561 522478
rect 173615 522512 173667 522640
rect 173615 522478 173623 522512
rect 173657 522478 173667 522512
rect 173615 522466 173667 522478
rect 174613 522512 174665 522640
rect 174613 522478 174623 522512
rect 174657 522478 174665 522512
rect 174903 522512 174955 522640
rect 174613 522466 174665 522478
rect 174903 522478 174911 522512
rect 174945 522478 174955 522512
rect 174903 522466 174955 522478
rect 175901 522512 175953 522640
rect 175901 522478 175911 522512
rect 175945 522478 175953 522512
rect 175901 522466 175953 522478
rect 176007 522512 176059 522640
rect 176007 522478 176015 522512
rect 176049 522478 176059 522512
rect 176007 522466 176059 522478
rect 177005 522512 177057 522640
rect 177005 522478 177015 522512
rect 177049 522478 177057 522512
rect 177005 522466 177057 522478
rect 177111 522512 177163 522640
rect 177111 522478 177119 522512
rect 177153 522478 177163 522512
rect 177111 522466 177163 522478
rect 178109 522512 178161 522640
rect 178109 522478 178119 522512
rect 178153 522478 178161 522512
rect 178109 522466 178161 522478
rect 178215 522512 178267 522640
rect 178215 522478 178223 522512
rect 178257 522478 178267 522512
rect 178215 522466 178267 522478
rect 179213 522512 179265 522640
rect 179213 522478 179223 522512
rect 179257 522478 179265 522512
rect 179213 522466 179265 522478
rect 179319 522614 179371 522640
rect 179319 522580 179327 522614
rect 179361 522580 179371 522614
rect 179319 522512 179371 522580
rect 179319 522478 179327 522512
rect 179361 522478 179371 522512
rect 179319 522466 179371 522478
rect 179765 522614 179817 522640
rect 179765 522580 179775 522614
rect 179809 522580 179817 522614
rect 179765 522512 179817 522580
rect 179765 522478 179775 522512
rect 179809 522478 179817 522512
rect 180055 522512 180107 522640
rect 179765 522466 179817 522478
rect 180055 522478 180063 522512
rect 180097 522478 180107 522512
rect 180055 522466 180107 522478
rect 181053 522512 181105 522640
rect 181053 522478 181063 522512
rect 181097 522478 181105 522512
rect 181053 522466 181105 522478
rect 181159 522512 181211 522640
rect 181159 522478 181167 522512
rect 181201 522478 181211 522512
rect 181159 522466 181211 522478
rect 182157 522512 182209 522640
rect 182157 522478 182167 522512
rect 182201 522478 182209 522512
rect 182157 522466 182209 522478
rect 182263 522512 182315 522640
rect 182263 522478 182271 522512
rect 182305 522478 182315 522512
rect 182263 522466 182315 522478
rect 183261 522512 183313 522640
rect 183261 522478 183271 522512
rect 183305 522478 183313 522512
rect 183261 522466 183313 522478
rect 183367 522512 183419 522640
rect 183367 522478 183375 522512
rect 183409 522478 183419 522512
rect 183367 522466 183419 522478
rect 184365 522512 184417 522640
rect 184365 522478 184375 522512
rect 184409 522478 184417 522512
rect 184365 522466 184417 522478
rect 184471 522614 184523 522640
rect 184471 522580 184479 522614
rect 184513 522580 184523 522614
rect 184471 522512 184523 522580
rect 184471 522478 184479 522512
rect 184513 522478 184523 522512
rect 184471 522466 184523 522478
rect 184917 522614 184969 522640
rect 184917 522580 184927 522614
rect 184961 522580 184969 522614
rect 184917 522512 184969 522580
rect 184917 522478 184927 522512
rect 184961 522478 184969 522512
rect 185207 522512 185259 522640
rect 184917 522466 184969 522478
rect 185207 522478 185215 522512
rect 185249 522478 185259 522512
rect 185207 522466 185259 522478
rect 186205 522512 186257 522640
rect 186205 522478 186215 522512
rect 186249 522478 186257 522512
rect 186205 522466 186257 522478
rect 186311 522614 186363 522640
rect 186311 522580 186319 522614
rect 186353 522580 186363 522614
rect 186311 522512 186363 522580
rect 186311 522478 186319 522512
rect 186353 522478 186363 522512
rect 186311 522466 186363 522478
rect 186941 522614 186993 522640
rect 186941 522580 186951 522614
rect 186985 522580 186993 522614
rect 186941 522512 186993 522580
rect 186941 522478 186951 522512
rect 186985 522478 186993 522512
rect 186941 522466 186993 522478
rect 187231 522607 187283 522640
rect 187231 522573 187239 522607
rect 187273 522573 187283 522607
rect 187231 522512 187283 522573
rect 187231 522478 187239 522512
rect 187273 522478 187283 522512
rect 187231 522466 187283 522478
rect 187401 522607 187453 522640
rect 187401 522573 187411 522607
rect 187445 522573 187453 522607
rect 187401 522512 187453 522573
rect 187401 522478 187411 522512
rect 187445 522478 187453 522512
rect 187401 522466 187453 522478
rect 172235 522360 172287 522372
rect 172235 522326 172243 522360
rect 172277 522326 172287 522360
rect 172235 522265 172287 522326
rect 172235 522231 172243 522265
rect 172277 522231 172287 522265
rect 172235 522198 172287 522231
rect 172405 522360 172457 522372
rect 172405 522326 172415 522360
rect 172449 522326 172457 522360
rect 172405 522265 172457 522326
rect 172405 522231 172415 522265
rect 172449 522231 172457 522265
rect 172405 522198 172457 522231
rect 172511 522360 172563 522372
rect 172511 522326 172519 522360
rect 172553 522326 172563 522360
rect 172511 522198 172563 522326
rect 173509 522360 173561 522372
rect 173509 522326 173519 522360
rect 173553 522326 173561 522360
rect 173509 522198 173561 522326
rect 173615 522360 173667 522372
rect 173615 522326 173623 522360
rect 173657 522326 173667 522360
rect 173615 522198 173667 522326
rect 174613 522360 174665 522372
rect 174613 522326 174623 522360
rect 174657 522326 174665 522360
rect 174613 522198 174665 522326
rect 174719 522360 174771 522372
rect 174719 522326 174727 522360
rect 174761 522326 174771 522360
rect 174719 522198 174771 522326
rect 175717 522360 175769 522372
rect 175717 522326 175727 522360
rect 175761 522326 175769 522360
rect 175717 522198 175769 522326
rect 175823 522360 175875 522372
rect 175823 522326 175831 522360
rect 175865 522326 175875 522360
rect 175823 522198 175875 522326
rect 176821 522360 176873 522372
rect 176821 522326 176831 522360
rect 176865 522326 176873 522360
rect 176821 522198 176873 522326
rect 176927 522360 176979 522372
rect 176927 522326 176935 522360
rect 176969 522326 176979 522360
rect 176927 522258 176979 522326
rect 176927 522224 176935 522258
rect 176969 522224 176979 522258
rect 176927 522198 176979 522224
rect 177189 522360 177241 522372
rect 177189 522326 177199 522360
rect 177233 522326 177241 522360
rect 177479 522360 177531 522372
rect 177189 522258 177241 522326
rect 177189 522224 177199 522258
rect 177233 522224 177241 522258
rect 177189 522198 177241 522224
rect 177479 522326 177487 522360
rect 177521 522326 177531 522360
rect 177479 522198 177531 522326
rect 178477 522360 178529 522372
rect 178477 522326 178487 522360
rect 178521 522326 178529 522360
rect 178477 522198 178529 522326
rect 178583 522360 178635 522372
rect 178583 522326 178591 522360
rect 178625 522326 178635 522360
rect 178583 522198 178635 522326
rect 179581 522360 179633 522372
rect 179581 522326 179591 522360
rect 179625 522326 179633 522360
rect 179581 522198 179633 522326
rect 179687 522360 179739 522372
rect 179687 522326 179695 522360
rect 179729 522326 179739 522360
rect 179687 522198 179739 522326
rect 180685 522360 180737 522372
rect 180685 522326 180695 522360
rect 180729 522326 180737 522360
rect 180685 522198 180737 522326
rect 180791 522360 180843 522372
rect 180791 522326 180799 522360
rect 180833 522326 180843 522360
rect 180791 522198 180843 522326
rect 181789 522360 181841 522372
rect 181789 522326 181799 522360
rect 181833 522326 181841 522360
rect 181789 522198 181841 522326
rect 181895 522360 181947 522372
rect 181895 522326 181903 522360
rect 181937 522326 181947 522360
rect 181895 522258 181947 522326
rect 181895 522224 181903 522258
rect 181937 522224 181947 522258
rect 181895 522198 181947 522224
rect 182341 522360 182393 522372
rect 182341 522326 182351 522360
rect 182385 522326 182393 522360
rect 182631 522360 182683 522372
rect 182341 522258 182393 522326
rect 182341 522224 182351 522258
rect 182385 522224 182393 522258
rect 182341 522198 182393 522224
rect 182631 522326 182639 522360
rect 182673 522326 182683 522360
rect 182631 522198 182683 522326
rect 183629 522360 183681 522372
rect 183629 522326 183639 522360
rect 183673 522326 183681 522360
rect 183629 522198 183681 522326
rect 183735 522360 183787 522372
rect 183735 522326 183743 522360
rect 183777 522326 183787 522360
rect 183735 522198 183787 522326
rect 184733 522360 184785 522372
rect 184733 522326 184743 522360
rect 184777 522326 184785 522360
rect 184733 522198 184785 522326
rect 184839 522360 184891 522372
rect 184839 522326 184847 522360
rect 184881 522326 184891 522360
rect 184839 522198 184891 522326
rect 185837 522360 185889 522372
rect 185837 522326 185847 522360
rect 185881 522326 185889 522360
rect 185837 522198 185889 522326
rect 185943 522360 185995 522372
rect 185943 522326 185951 522360
rect 185985 522326 185995 522360
rect 185943 522198 185995 522326
rect 186941 522360 186993 522372
rect 186941 522326 186951 522360
rect 186985 522326 186993 522360
rect 186941 522198 186993 522326
rect 187231 522360 187283 522372
rect 187231 522326 187239 522360
rect 187273 522326 187283 522360
rect 187231 522265 187283 522326
rect 187231 522231 187239 522265
rect 187273 522231 187283 522265
rect 187231 522198 187283 522231
rect 187401 522360 187453 522372
rect 187401 522326 187411 522360
rect 187445 522326 187453 522360
rect 187401 522265 187453 522326
rect 187401 522231 187411 522265
rect 187445 522231 187453 522265
rect 187401 522198 187453 522231
rect 172235 521519 172287 521552
rect 172235 521485 172243 521519
rect 172277 521485 172287 521519
rect 172235 521424 172287 521485
rect 172235 521390 172243 521424
rect 172277 521390 172287 521424
rect 172235 521378 172287 521390
rect 172405 521519 172457 521552
rect 172405 521485 172415 521519
rect 172449 521485 172457 521519
rect 172405 521424 172457 521485
rect 172405 521390 172415 521424
rect 172449 521390 172457 521424
rect 172405 521378 172457 521390
rect 172511 521424 172563 521552
rect 172511 521390 172519 521424
rect 172553 521390 172563 521424
rect 172511 521378 172563 521390
rect 173509 521424 173561 521552
rect 173509 521390 173519 521424
rect 173553 521390 173561 521424
rect 173509 521378 173561 521390
rect 173615 521424 173667 521552
rect 173615 521390 173623 521424
rect 173657 521390 173667 521424
rect 173615 521378 173667 521390
rect 174613 521424 174665 521552
rect 174613 521390 174623 521424
rect 174657 521390 174665 521424
rect 174903 521424 174955 521552
rect 174613 521378 174665 521390
rect 174903 521390 174911 521424
rect 174945 521390 174955 521424
rect 174903 521378 174955 521390
rect 175901 521424 175953 521552
rect 175901 521390 175911 521424
rect 175945 521390 175953 521424
rect 175901 521378 175953 521390
rect 176007 521424 176059 521552
rect 176007 521390 176015 521424
rect 176049 521390 176059 521424
rect 176007 521378 176059 521390
rect 177005 521424 177057 521552
rect 177005 521390 177015 521424
rect 177049 521390 177057 521424
rect 177005 521378 177057 521390
rect 177111 521424 177163 521552
rect 177111 521390 177119 521424
rect 177153 521390 177163 521424
rect 177111 521378 177163 521390
rect 178109 521424 178161 521552
rect 178109 521390 178119 521424
rect 178153 521390 178161 521424
rect 178109 521378 178161 521390
rect 178215 521424 178267 521552
rect 178215 521390 178223 521424
rect 178257 521390 178267 521424
rect 178215 521378 178267 521390
rect 179213 521424 179265 521552
rect 179213 521390 179223 521424
rect 179257 521390 179265 521424
rect 179213 521378 179265 521390
rect 179319 521526 179371 521552
rect 179319 521492 179327 521526
rect 179361 521492 179371 521526
rect 179319 521424 179371 521492
rect 179319 521390 179327 521424
rect 179361 521390 179371 521424
rect 179319 521378 179371 521390
rect 179765 521526 179817 521552
rect 179765 521492 179775 521526
rect 179809 521492 179817 521526
rect 179765 521424 179817 521492
rect 179765 521390 179775 521424
rect 179809 521390 179817 521424
rect 180055 521424 180107 521552
rect 179765 521378 179817 521390
rect 180055 521390 180063 521424
rect 180097 521390 180107 521424
rect 180055 521378 180107 521390
rect 181053 521424 181105 521552
rect 181053 521390 181063 521424
rect 181097 521390 181105 521424
rect 181053 521378 181105 521390
rect 181159 521424 181211 521552
rect 181159 521390 181167 521424
rect 181201 521390 181211 521424
rect 181159 521378 181211 521390
rect 182157 521424 182209 521552
rect 182157 521390 182167 521424
rect 182201 521390 182209 521424
rect 182157 521378 182209 521390
rect 182263 521424 182315 521552
rect 182263 521390 182271 521424
rect 182305 521390 182315 521424
rect 182263 521378 182315 521390
rect 183261 521424 183313 521552
rect 183261 521390 183271 521424
rect 183305 521390 183313 521424
rect 183261 521378 183313 521390
rect 183367 521424 183419 521552
rect 183367 521390 183375 521424
rect 183409 521390 183419 521424
rect 183367 521378 183419 521390
rect 184365 521424 184417 521552
rect 184365 521390 184375 521424
rect 184409 521390 184417 521424
rect 184365 521378 184417 521390
rect 184471 521526 184523 521552
rect 184471 521492 184479 521526
rect 184513 521492 184523 521526
rect 184471 521424 184523 521492
rect 184471 521390 184479 521424
rect 184513 521390 184523 521424
rect 184471 521378 184523 521390
rect 184917 521526 184969 521552
rect 184917 521492 184927 521526
rect 184961 521492 184969 521526
rect 184917 521424 184969 521492
rect 184917 521390 184927 521424
rect 184961 521390 184969 521424
rect 185207 521424 185259 521552
rect 184917 521378 184969 521390
rect 185207 521390 185215 521424
rect 185249 521390 185259 521424
rect 185207 521378 185259 521390
rect 186205 521424 186257 521552
rect 186205 521390 186215 521424
rect 186249 521390 186257 521424
rect 186205 521378 186257 521390
rect 186311 521526 186363 521552
rect 186311 521492 186319 521526
rect 186353 521492 186363 521526
rect 186311 521424 186363 521492
rect 186311 521390 186319 521424
rect 186353 521390 186363 521424
rect 186311 521378 186363 521390
rect 186941 521526 186993 521552
rect 186941 521492 186951 521526
rect 186985 521492 186993 521526
rect 186941 521424 186993 521492
rect 186941 521390 186951 521424
rect 186985 521390 186993 521424
rect 186941 521378 186993 521390
rect 187231 521519 187283 521552
rect 187231 521485 187239 521519
rect 187273 521485 187283 521519
rect 187231 521424 187283 521485
rect 187231 521390 187239 521424
rect 187273 521390 187283 521424
rect 187231 521378 187283 521390
rect 187401 521519 187453 521552
rect 187401 521485 187411 521519
rect 187445 521485 187453 521519
rect 187401 521424 187453 521485
rect 187401 521390 187411 521424
rect 187445 521390 187453 521424
rect 187401 521378 187453 521390
rect 172235 521272 172287 521284
rect 172235 521238 172243 521272
rect 172277 521238 172287 521272
rect 172235 521177 172287 521238
rect 172235 521143 172243 521177
rect 172277 521143 172287 521177
rect 172235 521110 172287 521143
rect 172405 521272 172457 521284
rect 172405 521238 172415 521272
rect 172449 521238 172457 521272
rect 172405 521177 172457 521238
rect 172405 521143 172415 521177
rect 172449 521143 172457 521177
rect 172405 521110 172457 521143
rect 172511 521272 172563 521284
rect 172511 521238 172519 521272
rect 172553 521238 172563 521272
rect 172511 521110 172563 521238
rect 173509 521272 173561 521284
rect 173509 521238 173519 521272
rect 173553 521238 173561 521272
rect 173509 521110 173561 521238
rect 173615 521272 173667 521284
rect 173615 521238 173623 521272
rect 173657 521238 173667 521272
rect 173615 521110 173667 521238
rect 174613 521272 174665 521284
rect 174613 521238 174623 521272
rect 174657 521238 174665 521272
rect 174613 521110 174665 521238
rect 174719 521272 174771 521284
rect 174719 521238 174727 521272
rect 174761 521238 174771 521272
rect 174719 521110 174771 521238
rect 175717 521272 175769 521284
rect 175717 521238 175727 521272
rect 175761 521238 175769 521272
rect 175717 521110 175769 521238
rect 175823 521272 175875 521284
rect 175823 521238 175831 521272
rect 175865 521238 175875 521272
rect 175823 521110 175875 521238
rect 176821 521272 176873 521284
rect 176821 521238 176831 521272
rect 176865 521238 176873 521272
rect 176821 521110 176873 521238
rect 176927 521272 176979 521284
rect 176927 521238 176935 521272
rect 176969 521238 176979 521272
rect 176927 521170 176979 521238
rect 176927 521136 176935 521170
rect 176969 521136 176979 521170
rect 176927 521110 176979 521136
rect 177189 521272 177241 521284
rect 177189 521238 177199 521272
rect 177233 521238 177241 521272
rect 177479 521272 177531 521284
rect 177189 521170 177241 521238
rect 177189 521136 177199 521170
rect 177233 521136 177241 521170
rect 177189 521110 177241 521136
rect 177479 521238 177487 521272
rect 177521 521238 177531 521272
rect 177479 521110 177531 521238
rect 178477 521272 178529 521284
rect 178477 521238 178487 521272
rect 178521 521238 178529 521272
rect 178477 521110 178529 521238
rect 178583 521272 178635 521284
rect 178583 521238 178591 521272
rect 178625 521238 178635 521272
rect 178583 521110 178635 521238
rect 179581 521272 179633 521284
rect 179581 521238 179591 521272
rect 179625 521238 179633 521272
rect 179581 521110 179633 521238
rect 179687 521272 179739 521284
rect 179687 521238 179695 521272
rect 179729 521238 179739 521272
rect 179687 521110 179739 521238
rect 180685 521272 180737 521284
rect 180685 521238 180695 521272
rect 180729 521238 180737 521272
rect 180685 521110 180737 521238
rect 180791 521272 180843 521284
rect 180791 521238 180799 521272
rect 180833 521238 180843 521272
rect 180791 521110 180843 521238
rect 181789 521272 181841 521284
rect 181789 521238 181799 521272
rect 181833 521238 181841 521272
rect 181789 521110 181841 521238
rect 181895 521272 181947 521284
rect 181895 521238 181903 521272
rect 181937 521238 181947 521272
rect 181895 521170 181947 521238
rect 181895 521136 181903 521170
rect 181937 521136 181947 521170
rect 181895 521110 181947 521136
rect 182341 521272 182393 521284
rect 182341 521238 182351 521272
rect 182385 521238 182393 521272
rect 182631 521272 182683 521284
rect 182341 521170 182393 521238
rect 182341 521136 182351 521170
rect 182385 521136 182393 521170
rect 182341 521110 182393 521136
rect 182631 521238 182639 521272
rect 182673 521238 182683 521272
rect 182631 521110 182683 521238
rect 183629 521272 183681 521284
rect 183629 521238 183639 521272
rect 183673 521238 183681 521272
rect 183629 521110 183681 521238
rect 183735 521272 183787 521284
rect 183735 521238 183743 521272
rect 183777 521238 183787 521272
rect 183735 521110 183787 521238
rect 184733 521272 184785 521284
rect 184733 521238 184743 521272
rect 184777 521238 184785 521272
rect 184733 521110 184785 521238
rect 184839 521272 184891 521284
rect 184839 521238 184847 521272
rect 184881 521238 184891 521272
rect 184839 521110 184891 521238
rect 185837 521272 185889 521284
rect 185837 521238 185847 521272
rect 185881 521238 185889 521272
rect 185837 521110 185889 521238
rect 185943 521272 185995 521284
rect 185943 521238 185951 521272
rect 185985 521238 185995 521272
rect 185943 521110 185995 521238
rect 186941 521272 186993 521284
rect 186941 521238 186951 521272
rect 186985 521238 186993 521272
rect 186941 521110 186993 521238
rect 187231 521272 187283 521284
rect 187231 521238 187239 521272
rect 187273 521238 187283 521272
rect 187231 521177 187283 521238
rect 187231 521143 187239 521177
rect 187273 521143 187283 521177
rect 187231 521110 187283 521143
rect 187401 521272 187453 521284
rect 187401 521238 187411 521272
rect 187445 521238 187453 521272
rect 187401 521177 187453 521238
rect 187401 521143 187411 521177
rect 187445 521143 187453 521177
rect 187401 521110 187453 521143
rect 172235 520431 172287 520464
rect 172235 520397 172243 520431
rect 172277 520397 172287 520431
rect 172235 520336 172287 520397
rect 172235 520302 172243 520336
rect 172277 520302 172287 520336
rect 172235 520290 172287 520302
rect 172405 520431 172457 520464
rect 172405 520397 172415 520431
rect 172449 520397 172457 520431
rect 172405 520336 172457 520397
rect 172405 520302 172415 520336
rect 172449 520302 172457 520336
rect 172405 520290 172457 520302
rect 172511 520336 172563 520464
rect 172511 520302 172519 520336
rect 172553 520302 172563 520336
rect 172511 520290 172563 520302
rect 173509 520336 173561 520464
rect 173509 520302 173519 520336
rect 173553 520302 173561 520336
rect 173509 520290 173561 520302
rect 173615 520336 173667 520464
rect 173615 520302 173623 520336
rect 173657 520302 173667 520336
rect 173615 520290 173667 520302
rect 174613 520336 174665 520464
rect 174613 520302 174623 520336
rect 174657 520302 174665 520336
rect 174903 520336 174955 520464
rect 174613 520290 174665 520302
rect 174903 520302 174911 520336
rect 174945 520302 174955 520336
rect 174903 520290 174955 520302
rect 175901 520336 175953 520464
rect 175901 520302 175911 520336
rect 175945 520302 175953 520336
rect 175901 520290 175953 520302
rect 176007 520336 176059 520464
rect 176007 520302 176015 520336
rect 176049 520302 176059 520336
rect 176007 520290 176059 520302
rect 177005 520336 177057 520464
rect 177005 520302 177015 520336
rect 177049 520302 177057 520336
rect 177005 520290 177057 520302
rect 177111 520336 177163 520464
rect 177111 520302 177119 520336
rect 177153 520302 177163 520336
rect 177111 520290 177163 520302
rect 178109 520336 178161 520464
rect 178109 520302 178119 520336
rect 178153 520302 178161 520336
rect 178109 520290 178161 520302
rect 178215 520336 178267 520464
rect 178215 520302 178223 520336
rect 178257 520302 178267 520336
rect 178215 520290 178267 520302
rect 179213 520336 179265 520464
rect 179213 520302 179223 520336
rect 179257 520302 179265 520336
rect 179213 520290 179265 520302
rect 179319 520438 179371 520464
rect 179319 520404 179327 520438
rect 179361 520404 179371 520438
rect 179319 520336 179371 520404
rect 179319 520302 179327 520336
rect 179361 520302 179371 520336
rect 179319 520290 179371 520302
rect 179765 520438 179817 520464
rect 179765 520404 179775 520438
rect 179809 520404 179817 520438
rect 179765 520336 179817 520404
rect 179765 520302 179775 520336
rect 179809 520302 179817 520336
rect 180055 520336 180107 520464
rect 179765 520290 179817 520302
rect 180055 520302 180063 520336
rect 180097 520302 180107 520336
rect 180055 520290 180107 520302
rect 181053 520336 181105 520464
rect 181053 520302 181063 520336
rect 181097 520302 181105 520336
rect 181053 520290 181105 520302
rect 181159 520336 181211 520464
rect 181159 520302 181167 520336
rect 181201 520302 181211 520336
rect 181159 520290 181211 520302
rect 182157 520336 182209 520464
rect 182157 520302 182167 520336
rect 182201 520302 182209 520336
rect 182157 520290 182209 520302
rect 182263 520336 182315 520464
rect 182263 520302 182271 520336
rect 182305 520302 182315 520336
rect 182263 520290 182315 520302
rect 183261 520336 183313 520464
rect 183261 520302 183271 520336
rect 183305 520302 183313 520336
rect 183261 520290 183313 520302
rect 183367 520336 183419 520464
rect 183367 520302 183375 520336
rect 183409 520302 183419 520336
rect 183367 520290 183419 520302
rect 184365 520336 184417 520464
rect 184365 520302 184375 520336
rect 184409 520302 184417 520336
rect 184365 520290 184417 520302
rect 184471 520438 184523 520464
rect 184471 520404 184479 520438
rect 184513 520404 184523 520438
rect 184471 520336 184523 520404
rect 184471 520302 184479 520336
rect 184513 520302 184523 520336
rect 184471 520290 184523 520302
rect 184917 520438 184969 520464
rect 184917 520404 184927 520438
rect 184961 520404 184969 520438
rect 184917 520336 184969 520404
rect 184917 520302 184927 520336
rect 184961 520302 184969 520336
rect 185207 520336 185259 520464
rect 184917 520290 184969 520302
rect 185207 520302 185215 520336
rect 185249 520302 185259 520336
rect 185207 520290 185259 520302
rect 186205 520336 186257 520464
rect 186205 520302 186215 520336
rect 186249 520302 186257 520336
rect 186205 520290 186257 520302
rect 186311 520438 186363 520464
rect 186311 520404 186319 520438
rect 186353 520404 186363 520438
rect 186311 520336 186363 520404
rect 186311 520302 186319 520336
rect 186353 520302 186363 520336
rect 186311 520290 186363 520302
rect 186941 520438 186993 520464
rect 186941 520404 186951 520438
rect 186985 520404 186993 520438
rect 186941 520336 186993 520404
rect 186941 520302 186951 520336
rect 186985 520302 186993 520336
rect 186941 520290 186993 520302
rect 187231 520431 187283 520464
rect 187231 520397 187239 520431
rect 187273 520397 187283 520431
rect 187231 520336 187283 520397
rect 187231 520302 187239 520336
rect 187273 520302 187283 520336
rect 187231 520290 187283 520302
rect 187401 520431 187453 520464
rect 187401 520397 187411 520431
rect 187445 520397 187453 520431
rect 187401 520336 187453 520397
rect 187401 520302 187411 520336
rect 187445 520302 187453 520336
rect 187401 520290 187453 520302
rect 172235 520184 172287 520196
rect 172235 520150 172243 520184
rect 172277 520150 172287 520184
rect 172235 520089 172287 520150
rect 172235 520055 172243 520089
rect 172277 520055 172287 520089
rect 172235 520022 172287 520055
rect 172405 520184 172457 520196
rect 172405 520150 172415 520184
rect 172449 520150 172457 520184
rect 172405 520089 172457 520150
rect 172405 520055 172415 520089
rect 172449 520055 172457 520089
rect 172405 520022 172457 520055
rect 172511 520184 172563 520196
rect 172511 520150 172519 520184
rect 172553 520150 172563 520184
rect 172511 520022 172563 520150
rect 173509 520184 173561 520196
rect 173509 520150 173519 520184
rect 173553 520150 173561 520184
rect 173509 520022 173561 520150
rect 173615 520184 173667 520196
rect 173615 520150 173623 520184
rect 173657 520150 173667 520184
rect 173615 520022 173667 520150
rect 174613 520184 174665 520196
rect 174613 520150 174623 520184
rect 174657 520150 174665 520184
rect 174613 520022 174665 520150
rect 174719 520184 174771 520196
rect 174719 520150 174727 520184
rect 174761 520150 174771 520184
rect 174719 520022 174771 520150
rect 175717 520184 175769 520196
rect 175717 520150 175727 520184
rect 175761 520150 175769 520184
rect 175717 520022 175769 520150
rect 175823 520184 175875 520196
rect 175823 520150 175831 520184
rect 175865 520150 175875 520184
rect 175823 520022 175875 520150
rect 176821 520184 176873 520196
rect 176821 520150 176831 520184
rect 176865 520150 176873 520184
rect 176821 520022 176873 520150
rect 176927 520184 176979 520196
rect 176927 520150 176935 520184
rect 176969 520150 176979 520184
rect 176927 520082 176979 520150
rect 176927 520048 176935 520082
rect 176969 520048 176979 520082
rect 176927 520022 176979 520048
rect 177189 520184 177241 520196
rect 177189 520150 177199 520184
rect 177233 520150 177241 520184
rect 177479 520184 177531 520196
rect 177189 520082 177241 520150
rect 177189 520048 177199 520082
rect 177233 520048 177241 520082
rect 177189 520022 177241 520048
rect 177479 520150 177487 520184
rect 177521 520150 177531 520184
rect 177479 520022 177531 520150
rect 178477 520184 178529 520196
rect 178477 520150 178487 520184
rect 178521 520150 178529 520184
rect 178477 520022 178529 520150
rect 178583 520184 178635 520196
rect 178583 520150 178591 520184
rect 178625 520150 178635 520184
rect 178583 520022 178635 520150
rect 179581 520184 179633 520196
rect 179581 520150 179591 520184
rect 179625 520150 179633 520184
rect 179581 520022 179633 520150
rect 179687 520184 179739 520196
rect 179687 520150 179695 520184
rect 179729 520150 179739 520184
rect 179687 520022 179739 520150
rect 180685 520184 180737 520196
rect 180685 520150 180695 520184
rect 180729 520150 180737 520184
rect 180685 520022 180737 520150
rect 180791 520184 180843 520196
rect 180791 520150 180799 520184
rect 180833 520150 180843 520184
rect 180791 520022 180843 520150
rect 181789 520184 181841 520196
rect 181789 520150 181799 520184
rect 181833 520150 181841 520184
rect 181789 520022 181841 520150
rect 181895 520184 181947 520196
rect 181895 520150 181903 520184
rect 181937 520150 181947 520184
rect 181895 520082 181947 520150
rect 181895 520048 181903 520082
rect 181937 520048 181947 520082
rect 181895 520022 181947 520048
rect 182341 520184 182393 520196
rect 182341 520150 182351 520184
rect 182385 520150 182393 520184
rect 182631 520184 182683 520196
rect 182341 520082 182393 520150
rect 182341 520048 182351 520082
rect 182385 520048 182393 520082
rect 182341 520022 182393 520048
rect 182631 520150 182639 520184
rect 182673 520150 182683 520184
rect 182631 520022 182683 520150
rect 183629 520184 183681 520196
rect 183629 520150 183639 520184
rect 183673 520150 183681 520184
rect 183629 520022 183681 520150
rect 183735 520184 183787 520196
rect 183735 520150 183743 520184
rect 183777 520150 183787 520184
rect 183735 520022 183787 520150
rect 184733 520184 184785 520196
rect 184733 520150 184743 520184
rect 184777 520150 184785 520184
rect 184733 520022 184785 520150
rect 184839 520184 184891 520196
rect 184839 520150 184847 520184
rect 184881 520150 184891 520184
rect 184839 520022 184891 520150
rect 185837 520184 185889 520196
rect 185837 520150 185847 520184
rect 185881 520150 185889 520184
rect 185837 520022 185889 520150
rect 185943 520184 185995 520196
rect 185943 520150 185951 520184
rect 185985 520150 185995 520184
rect 185943 520022 185995 520150
rect 186941 520184 186993 520196
rect 186941 520150 186951 520184
rect 186985 520150 186993 520184
rect 186941 520022 186993 520150
rect 187231 520184 187283 520196
rect 187231 520150 187239 520184
rect 187273 520150 187283 520184
rect 187231 520089 187283 520150
rect 187231 520055 187239 520089
rect 187273 520055 187283 520089
rect 187231 520022 187283 520055
rect 187401 520184 187453 520196
rect 187401 520150 187411 520184
rect 187445 520150 187453 520184
rect 187401 520089 187453 520150
rect 187401 520055 187411 520089
rect 187445 520055 187453 520089
rect 187401 520022 187453 520055
rect 172235 519343 172287 519376
rect 172235 519309 172243 519343
rect 172277 519309 172287 519343
rect 172235 519248 172287 519309
rect 172235 519214 172243 519248
rect 172277 519214 172287 519248
rect 172235 519202 172287 519214
rect 172405 519343 172457 519376
rect 172405 519309 172415 519343
rect 172449 519309 172457 519343
rect 172405 519248 172457 519309
rect 172405 519214 172415 519248
rect 172449 519214 172457 519248
rect 172405 519202 172457 519214
rect 172511 519248 172563 519376
rect 172511 519214 172519 519248
rect 172553 519214 172563 519248
rect 172511 519202 172563 519214
rect 173509 519248 173561 519376
rect 173509 519214 173519 519248
rect 173553 519214 173561 519248
rect 173509 519202 173561 519214
rect 173615 519248 173667 519376
rect 173615 519214 173623 519248
rect 173657 519214 173667 519248
rect 173615 519202 173667 519214
rect 174613 519248 174665 519376
rect 174613 519214 174623 519248
rect 174657 519214 174665 519248
rect 174903 519248 174955 519376
rect 174613 519202 174665 519214
rect 174903 519214 174911 519248
rect 174945 519214 174955 519248
rect 174903 519202 174955 519214
rect 175901 519248 175953 519376
rect 175901 519214 175911 519248
rect 175945 519214 175953 519248
rect 175901 519202 175953 519214
rect 176007 519248 176059 519376
rect 176007 519214 176015 519248
rect 176049 519214 176059 519248
rect 176007 519202 176059 519214
rect 177005 519248 177057 519376
rect 177005 519214 177015 519248
rect 177049 519214 177057 519248
rect 177005 519202 177057 519214
rect 177111 519248 177163 519376
rect 177111 519214 177119 519248
rect 177153 519214 177163 519248
rect 177111 519202 177163 519214
rect 178109 519248 178161 519376
rect 178109 519214 178119 519248
rect 178153 519214 178161 519248
rect 178109 519202 178161 519214
rect 178215 519248 178267 519376
rect 178215 519214 178223 519248
rect 178257 519214 178267 519248
rect 178215 519202 178267 519214
rect 179213 519248 179265 519376
rect 179213 519214 179223 519248
rect 179257 519214 179265 519248
rect 179213 519202 179265 519214
rect 179319 519350 179371 519376
rect 179319 519316 179327 519350
rect 179361 519316 179371 519350
rect 179319 519248 179371 519316
rect 179319 519214 179327 519248
rect 179361 519214 179371 519248
rect 179319 519202 179371 519214
rect 179765 519350 179817 519376
rect 179765 519316 179775 519350
rect 179809 519316 179817 519350
rect 179765 519248 179817 519316
rect 179765 519214 179775 519248
rect 179809 519214 179817 519248
rect 180055 519248 180107 519376
rect 179765 519202 179817 519214
rect 180055 519214 180063 519248
rect 180097 519214 180107 519248
rect 180055 519202 180107 519214
rect 181053 519248 181105 519376
rect 181053 519214 181063 519248
rect 181097 519214 181105 519248
rect 181053 519202 181105 519214
rect 181159 519248 181211 519376
rect 181159 519214 181167 519248
rect 181201 519214 181211 519248
rect 181159 519202 181211 519214
rect 182157 519248 182209 519376
rect 182157 519214 182167 519248
rect 182201 519214 182209 519248
rect 182157 519202 182209 519214
rect 182263 519248 182315 519376
rect 182263 519214 182271 519248
rect 182305 519214 182315 519248
rect 182263 519202 182315 519214
rect 183261 519248 183313 519376
rect 183261 519214 183271 519248
rect 183305 519214 183313 519248
rect 183261 519202 183313 519214
rect 183367 519248 183419 519376
rect 183367 519214 183375 519248
rect 183409 519214 183419 519248
rect 183367 519202 183419 519214
rect 184365 519248 184417 519376
rect 184365 519214 184375 519248
rect 184409 519214 184417 519248
rect 184365 519202 184417 519214
rect 184471 519350 184523 519376
rect 184471 519316 184479 519350
rect 184513 519316 184523 519350
rect 184471 519248 184523 519316
rect 184471 519214 184479 519248
rect 184513 519214 184523 519248
rect 184471 519202 184523 519214
rect 184917 519350 184969 519376
rect 184917 519316 184927 519350
rect 184961 519316 184969 519350
rect 184917 519248 184969 519316
rect 184917 519214 184927 519248
rect 184961 519214 184969 519248
rect 185207 519248 185259 519376
rect 184917 519202 184969 519214
rect 185207 519214 185215 519248
rect 185249 519214 185259 519248
rect 185207 519202 185259 519214
rect 186205 519248 186257 519376
rect 186205 519214 186215 519248
rect 186249 519214 186257 519248
rect 186205 519202 186257 519214
rect 186311 519350 186363 519376
rect 186311 519316 186319 519350
rect 186353 519316 186363 519350
rect 186311 519248 186363 519316
rect 186311 519214 186319 519248
rect 186353 519214 186363 519248
rect 186311 519202 186363 519214
rect 186941 519350 186993 519376
rect 186941 519316 186951 519350
rect 186985 519316 186993 519350
rect 186941 519248 186993 519316
rect 186941 519214 186951 519248
rect 186985 519214 186993 519248
rect 186941 519202 186993 519214
rect 187231 519343 187283 519376
rect 187231 519309 187239 519343
rect 187273 519309 187283 519343
rect 187231 519248 187283 519309
rect 187231 519214 187239 519248
rect 187273 519214 187283 519248
rect 187231 519202 187283 519214
rect 187401 519343 187453 519376
rect 187401 519309 187411 519343
rect 187445 519309 187453 519343
rect 187401 519248 187453 519309
rect 187401 519214 187411 519248
rect 187445 519214 187453 519248
rect 187401 519202 187453 519214
rect 172235 519096 172287 519108
rect 172235 519062 172243 519096
rect 172277 519062 172287 519096
rect 172235 519001 172287 519062
rect 172235 518967 172243 519001
rect 172277 518967 172287 519001
rect 172235 518934 172287 518967
rect 172405 519096 172457 519108
rect 172405 519062 172415 519096
rect 172449 519062 172457 519096
rect 172405 519001 172457 519062
rect 172405 518967 172415 519001
rect 172449 518967 172457 519001
rect 172405 518934 172457 518967
rect 172511 519096 172563 519108
rect 172511 519062 172519 519096
rect 172553 519062 172563 519096
rect 172511 518934 172563 519062
rect 173509 519096 173561 519108
rect 173509 519062 173519 519096
rect 173553 519062 173561 519096
rect 173509 518934 173561 519062
rect 173615 519096 173667 519108
rect 173615 519062 173623 519096
rect 173657 519062 173667 519096
rect 173615 518934 173667 519062
rect 174613 519096 174665 519108
rect 174613 519062 174623 519096
rect 174657 519062 174665 519096
rect 174613 518934 174665 519062
rect 174719 519096 174771 519108
rect 174719 519062 174727 519096
rect 174761 519062 174771 519096
rect 174719 518934 174771 519062
rect 175717 519096 175769 519108
rect 175717 519062 175727 519096
rect 175761 519062 175769 519096
rect 175717 518934 175769 519062
rect 175823 519096 175875 519108
rect 175823 519062 175831 519096
rect 175865 519062 175875 519096
rect 175823 518934 175875 519062
rect 176821 519096 176873 519108
rect 176821 519062 176831 519096
rect 176865 519062 176873 519096
rect 176821 518934 176873 519062
rect 176927 519096 176979 519108
rect 176927 519062 176935 519096
rect 176969 519062 176979 519096
rect 176927 518994 176979 519062
rect 176927 518960 176935 518994
rect 176969 518960 176979 518994
rect 176927 518934 176979 518960
rect 177189 519096 177241 519108
rect 177189 519062 177199 519096
rect 177233 519062 177241 519096
rect 177479 519096 177531 519108
rect 177189 518994 177241 519062
rect 177189 518960 177199 518994
rect 177233 518960 177241 518994
rect 177189 518934 177241 518960
rect 177479 519062 177487 519096
rect 177521 519062 177531 519096
rect 177479 518934 177531 519062
rect 178477 519096 178529 519108
rect 178477 519062 178487 519096
rect 178521 519062 178529 519096
rect 178477 518934 178529 519062
rect 178583 519096 178635 519108
rect 178583 519062 178591 519096
rect 178625 519062 178635 519096
rect 178583 518934 178635 519062
rect 179581 519096 179633 519108
rect 179581 519062 179591 519096
rect 179625 519062 179633 519096
rect 179581 518934 179633 519062
rect 179687 519096 179739 519108
rect 179687 519062 179695 519096
rect 179729 519062 179739 519096
rect 179687 518934 179739 519062
rect 180685 519096 180737 519108
rect 180685 519062 180695 519096
rect 180729 519062 180737 519096
rect 180685 518934 180737 519062
rect 180791 519096 180843 519108
rect 180791 519062 180799 519096
rect 180833 519062 180843 519096
rect 180791 518934 180843 519062
rect 181789 519096 181841 519108
rect 181789 519062 181799 519096
rect 181833 519062 181841 519096
rect 181789 518934 181841 519062
rect 181895 519096 181947 519108
rect 181895 519062 181903 519096
rect 181937 519062 181947 519096
rect 181895 518994 181947 519062
rect 181895 518960 181903 518994
rect 181937 518960 181947 518994
rect 181895 518934 181947 518960
rect 182341 519096 182393 519108
rect 182341 519062 182351 519096
rect 182385 519062 182393 519096
rect 182631 519096 182683 519108
rect 182341 518994 182393 519062
rect 182341 518960 182351 518994
rect 182385 518960 182393 518994
rect 182341 518934 182393 518960
rect 182631 519062 182639 519096
rect 182673 519062 182683 519096
rect 182631 518934 182683 519062
rect 183629 519096 183681 519108
rect 183629 519062 183639 519096
rect 183673 519062 183681 519096
rect 183629 518934 183681 519062
rect 183735 519096 183787 519108
rect 183735 519062 183743 519096
rect 183777 519062 183787 519096
rect 183735 518934 183787 519062
rect 184733 519096 184785 519108
rect 184733 519062 184743 519096
rect 184777 519062 184785 519096
rect 184733 518934 184785 519062
rect 184839 519096 184891 519108
rect 184839 519062 184847 519096
rect 184881 519062 184891 519096
rect 184839 518934 184891 519062
rect 185837 519096 185889 519108
rect 185837 519062 185847 519096
rect 185881 519062 185889 519096
rect 185837 518934 185889 519062
rect 185943 519096 185995 519108
rect 185943 519062 185951 519096
rect 185985 519062 185995 519096
rect 185943 518934 185995 519062
rect 186941 519096 186993 519108
rect 186941 519062 186951 519096
rect 186985 519062 186993 519096
rect 186941 518934 186993 519062
rect 187231 519096 187283 519108
rect 187231 519062 187239 519096
rect 187273 519062 187283 519096
rect 187231 519001 187283 519062
rect 187231 518967 187239 519001
rect 187273 518967 187283 519001
rect 187231 518934 187283 518967
rect 187401 519096 187453 519108
rect 187401 519062 187411 519096
rect 187445 519062 187453 519096
rect 187401 519001 187453 519062
rect 187401 518967 187411 519001
rect 187445 518967 187453 519001
rect 187401 518934 187453 518967
rect 172235 518255 172287 518288
rect 172235 518221 172243 518255
rect 172277 518221 172287 518255
rect 172235 518160 172287 518221
rect 172235 518126 172243 518160
rect 172277 518126 172287 518160
rect 172235 518114 172287 518126
rect 172405 518255 172457 518288
rect 172405 518221 172415 518255
rect 172449 518221 172457 518255
rect 172405 518160 172457 518221
rect 172405 518126 172415 518160
rect 172449 518126 172457 518160
rect 172405 518114 172457 518126
rect 172511 518160 172563 518288
rect 172511 518126 172519 518160
rect 172553 518126 172563 518160
rect 172511 518114 172563 518126
rect 173509 518160 173561 518288
rect 173509 518126 173519 518160
rect 173553 518126 173561 518160
rect 173509 518114 173561 518126
rect 173615 518160 173667 518288
rect 173615 518126 173623 518160
rect 173657 518126 173667 518160
rect 173615 518114 173667 518126
rect 174613 518160 174665 518288
rect 174613 518126 174623 518160
rect 174657 518126 174665 518160
rect 174903 518160 174955 518288
rect 174613 518114 174665 518126
rect 174903 518126 174911 518160
rect 174945 518126 174955 518160
rect 174903 518114 174955 518126
rect 175901 518160 175953 518288
rect 175901 518126 175911 518160
rect 175945 518126 175953 518160
rect 175901 518114 175953 518126
rect 176007 518160 176059 518288
rect 176007 518126 176015 518160
rect 176049 518126 176059 518160
rect 176007 518114 176059 518126
rect 177005 518160 177057 518288
rect 177005 518126 177015 518160
rect 177049 518126 177057 518160
rect 177005 518114 177057 518126
rect 177111 518160 177163 518288
rect 177111 518126 177119 518160
rect 177153 518126 177163 518160
rect 177111 518114 177163 518126
rect 178109 518160 178161 518288
rect 178109 518126 178119 518160
rect 178153 518126 178161 518160
rect 178109 518114 178161 518126
rect 178215 518160 178267 518288
rect 178215 518126 178223 518160
rect 178257 518126 178267 518160
rect 178215 518114 178267 518126
rect 179213 518160 179265 518288
rect 179213 518126 179223 518160
rect 179257 518126 179265 518160
rect 179213 518114 179265 518126
rect 179319 518262 179371 518288
rect 179319 518228 179327 518262
rect 179361 518228 179371 518262
rect 179319 518160 179371 518228
rect 179319 518126 179327 518160
rect 179361 518126 179371 518160
rect 179319 518114 179371 518126
rect 179765 518262 179817 518288
rect 179765 518228 179775 518262
rect 179809 518228 179817 518262
rect 179765 518160 179817 518228
rect 179765 518126 179775 518160
rect 179809 518126 179817 518160
rect 180055 518160 180107 518288
rect 179765 518114 179817 518126
rect 180055 518126 180063 518160
rect 180097 518126 180107 518160
rect 180055 518114 180107 518126
rect 181053 518160 181105 518288
rect 181053 518126 181063 518160
rect 181097 518126 181105 518160
rect 181053 518114 181105 518126
rect 181159 518160 181211 518288
rect 181159 518126 181167 518160
rect 181201 518126 181211 518160
rect 181159 518114 181211 518126
rect 182157 518160 182209 518288
rect 182157 518126 182167 518160
rect 182201 518126 182209 518160
rect 182157 518114 182209 518126
rect 182263 518160 182315 518288
rect 182263 518126 182271 518160
rect 182305 518126 182315 518160
rect 182263 518114 182315 518126
rect 183261 518160 183313 518288
rect 183261 518126 183271 518160
rect 183305 518126 183313 518160
rect 183261 518114 183313 518126
rect 183367 518160 183419 518288
rect 183367 518126 183375 518160
rect 183409 518126 183419 518160
rect 183367 518114 183419 518126
rect 184365 518160 184417 518288
rect 184365 518126 184375 518160
rect 184409 518126 184417 518160
rect 184365 518114 184417 518126
rect 184471 518262 184523 518288
rect 184471 518228 184479 518262
rect 184513 518228 184523 518262
rect 184471 518160 184523 518228
rect 184471 518126 184479 518160
rect 184513 518126 184523 518160
rect 184471 518114 184523 518126
rect 184917 518262 184969 518288
rect 184917 518228 184927 518262
rect 184961 518228 184969 518262
rect 184917 518160 184969 518228
rect 184917 518126 184927 518160
rect 184961 518126 184969 518160
rect 185207 518160 185259 518288
rect 184917 518114 184969 518126
rect 185207 518126 185215 518160
rect 185249 518126 185259 518160
rect 185207 518114 185259 518126
rect 186205 518160 186257 518288
rect 186205 518126 186215 518160
rect 186249 518126 186257 518160
rect 186205 518114 186257 518126
rect 186311 518262 186363 518288
rect 186311 518228 186319 518262
rect 186353 518228 186363 518262
rect 186311 518160 186363 518228
rect 186311 518126 186319 518160
rect 186353 518126 186363 518160
rect 186311 518114 186363 518126
rect 186941 518262 186993 518288
rect 186941 518228 186951 518262
rect 186985 518228 186993 518262
rect 186941 518160 186993 518228
rect 186941 518126 186951 518160
rect 186985 518126 186993 518160
rect 186941 518114 186993 518126
rect 187231 518255 187283 518288
rect 187231 518221 187239 518255
rect 187273 518221 187283 518255
rect 187231 518160 187283 518221
rect 187231 518126 187239 518160
rect 187273 518126 187283 518160
rect 187231 518114 187283 518126
rect 187401 518255 187453 518288
rect 187401 518221 187411 518255
rect 187445 518221 187453 518255
rect 187401 518160 187453 518221
rect 187401 518126 187411 518160
rect 187445 518126 187453 518160
rect 187401 518114 187453 518126
rect 172235 518008 172287 518020
rect 172235 517974 172243 518008
rect 172277 517974 172287 518008
rect 172235 517913 172287 517974
rect 172235 517879 172243 517913
rect 172277 517879 172287 517913
rect 172235 517846 172287 517879
rect 172405 518008 172457 518020
rect 172405 517974 172415 518008
rect 172449 517974 172457 518008
rect 172405 517913 172457 517974
rect 172405 517879 172415 517913
rect 172449 517879 172457 517913
rect 172405 517846 172457 517879
rect 172511 518008 172563 518020
rect 172511 517974 172519 518008
rect 172553 517974 172563 518008
rect 172511 517846 172563 517974
rect 173509 518008 173561 518020
rect 173509 517974 173519 518008
rect 173553 517974 173561 518008
rect 173509 517846 173561 517974
rect 173615 518008 173667 518020
rect 173615 517974 173623 518008
rect 173657 517974 173667 518008
rect 173615 517846 173667 517974
rect 174613 518008 174665 518020
rect 174613 517974 174623 518008
rect 174657 517974 174665 518008
rect 174613 517846 174665 517974
rect 174719 518008 174771 518020
rect 174719 517974 174727 518008
rect 174761 517974 174771 518008
rect 174719 517846 174771 517974
rect 175717 518008 175769 518020
rect 175717 517974 175727 518008
rect 175761 517974 175769 518008
rect 175717 517846 175769 517974
rect 175823 518008 175875 518020
rect 175823 517974 175831 518008
rect 175865 517974 175875 518008
rect 175823 517846 175875 517974
rect 176821 518008 176873 518020
rect 176821 517974 176831 518008
rect 176865 517974 176873 518008
rect 176821 517846 176873 517974
rect 176927 518008 176979 518020
rect 176927 517974 176935 518008
rect 176969 517974 176979 518008
rect 176927 517906 176979 517974
rect 176927 517872 176935 517906
rect 176969 517872 176979 517906
rect 176927 517846 176979 517872
rect 177189 518008 177241 518020
rect 177189 517974 177199 518008
rect 177233 517974 177241 518008
rect 177479 518008 177531 518020
rect 177189 517906 177241 517974
rect 177189 517872 177199 517906
rect 177233 517872 177241 517906
rect 177189 517846 177241 517872
rect 177479 517974 177487 518008
rect 177521 517974 177531 518008
rect 177479 517846 177531 517974
rect 178477 518008 178529 518020
rect 178477 517974 178487 518008
rect 178521 517974 178529 518008
rect 178477 517846 178529 517974
rect 178583 518008 178635 518020
rect 178583 517974 178591 518008
rect 178625 517974 178635 518008
rect 178583 517846 178635 517974
rect 179581 518008 179633 518020
rect 179581 517974 179591 518008
rect 179625 517974 179633 518008
rect 179581 517846 179633 517974
rect 179687 518008 179739 518020
rect 179687 517974 179695 518008
rect 179729 517974 179739 518008
rect 179687 517846 179739 517974
rect 180685 518008 180737 518020
rect 180685 517974 180695 518008
rect 180729 517974 180737 518008
rect 180685 517846 180737 517974
rect 180791 518008 180843 518020
rect 180791 517974 180799 518008
rect 180833 517974 180843 518008
rect 180791 517846 180843 517974
rect 181789 518008 181841 518020
rect 181789 517974 181799 518008
rect 181833 517974 181841 518008
rect 181789 517846 181841 517974
rect 181895 518008 181947 518020
rect 181895 517974 181903 518008
rect 181937 517974 181947 518008
rect 181895 517906 181947 517974
rect 181895 517872 181903 517906
rect 181937 517872 181947 517906
rect 181895 517846 181947 517872
rect 182341 518008 182393 518020
rect 182341 517974 182351 518008
rect 182385 517974 182393 518008
rect 182631 518008 182683 518020
rect 182341 517906 182393 517974
rect 182341 517872 182351 517906
rect 182385 517872 182393 517906
rect 182341 517846 182393 517872
rect 182631 517974 182639 518008
rect 182673 517974 182683 518008
rect 182631 517846 182683 517974
rect 183629 518008 183681 518020
rect 183629 517974 183639 518008
rect 183673 517974 183681 518008
rect 183629 517846 183681 517974
rect 183735 518008 183787 518020
rect 183735 517974 183743 518008
rect 183777 517974 183787 518008
rect 183735 517846 183787 517974
rect 184733 518008 184785 518020
rect 184733 517974 184743 518008
rect 184777 517974 184785 518008
rect 184733 517846 184785 517974
rect 184839 518008 184891 518020
rect 184839 517974 184847 518008
rect 184881 517974 184891 518008
rect 184839 517846 184891 517974
rect 185837 518008 185889 518020
rect 185837 517974 185847 518008
rect 185881 517974 185889 518008
rect 185837 517846 185889 517974
rect 185943 518008 185995 518020
rect 185943 517974 185951 518008
rect 185985 517974 185995 518008
rect 185943 517846 185995 517974
rect 186941 518008 186993 518020
rect 186941 517974 186951 518008
rect 186985 517974 186993 518008
rect 186941 517846 186993 517974
rect 187231 518008 187283 518020
rect 187231 517974 187239 518008
rect 187273 517974 187283 518008
rect 187231 517913 187283 517974
rect 187231 517879 187239 517913
rect 187273 517879 187283 517913
rect 187231 517846 187283 517879
rect 187401 518008 187453 518020
rect 187401 517974 187411 518008
rect 187445 517974 187453 518008
rect 187401 517913 187453 517974
rect 187401 517879 187411 517913
rect 187445 517879 187453 517913
rect 187401 517846 187453 517879
rect 172235 517167 172287 517200
rect 172235 517133 172243 517167
rect 172277 517133 172287 517167
rect 172235 517072 172287 517133
rect 172235 517038 172243 517072
rect 172277 517038 172287 517072
rect 172235 517026 172287 517038
rect 172405 517167 172457 517200
rect 172405 517133 172415 517167
rect 172449 517133 172457 517167
rect 172405 517072 172457 517133
rect 172405 517038 172415 517072
rect 172449 517038 172457 517072
rect 172405 517026 172457 517038
rect 172511 517072 172563 517200
rect 172511 517038 172519 517072
rect 172553 517038 172563 517072
rect 172511 517026 172563 517038
rect 173509 517072 173561 517200
rect 173509 517038 173519 517072
rect 173553 517038 173561 517072
rect 173509 517026 173561 517038
rect 173615 517072 173667 517200
rect 173615 517038 173623 517072
rect 173657 517038 173667 517072
rect 173615 517026 173667 517038
rect 174613 517072 174665 517200
rect 174613 517038 174623 517072
rect 174657 517038 174665 517072
rect 174903 517072 174955 517200
rect 174613 517026 174665 517038
rect 174903 517038 174911 517072
rect 174945 517038 174955 517072
rect 174903 517026 174955 517038
rect 175901 517072 175953 517200
rect 175901 517038 175911 517072
rect 175945 517038 175953 517072
rect 175901 517026 175953 517038
rect 176007 517072 176059 517200
rect 176007 517038 176015 517072
rect 176049 517038 176059 517072
rect 176007 517026 176059 517038
rect 177005 517072 177057 517200
rect 177005 517038 177015 517072
rect 177049 517038 177057 517072
rect 177005 517026 177057 517038
rect 177111 517072 177163 517200
rect 177111 517038 177119 517072
rect 177153 517038 177163 517072
rect 177111 517026 177163 517038
rect 178109 517072 178161 517200
rect 178109 517038 178119 517072
rect 178153 517038 178161 517072
rect 178109 517026 178161 517038
rect 178215 517072 178267 517200
rect 178215 517038 178223 517072
rect 178257 517038 178267 517072
rect 178215 517026 178267 517038
rect 179213 517072 179265 517200
rect 179213 517038 179223 517072
rect 179257 517038 179265 517072
rect 179213 517026 179265 517038
rect 179319 517174 179371 517200
rect 179319 517140 179327 517174
rect 179361 517140 179371 517174
rect 179319 517072 179371 517140
rect 179319 517038 179327 517072
rect 179361 517038 179371 517072
rect 179319 517026 179371 517038
rect 179765 517174 179817 517200
rect 179765 517140 179775 517174
rect 179809 517140 179817 517174
rect 179765 517072 179817 517140
rect 179765 517038 179775 517072
rect 179809 517038 179817 517072
rect 180055 517072 180107 517200
rect 179765 517026 179817 517038
rect 180055 517038 180063 517072
rect 180097 517038 180107 517072
rect 180055 517026 180107 517038
rect 181053 517072 181105 517200
rect 181053 517038 181063 517072
rect 181097 517038 181105 517072
rect 181053 517026 181105 517038
rect 181159 517072 181211 517200
rect 181159 517038 181167 517072
rect 181201 517038 181211 517072
rect 181159 517026 181211 517038
rect 182157 517072 182209 517200
rect 182157 517038 182167 517072
rect 182201 517038 182209 517072
rect 182157 517026 182209 517038
rect 182263 517072 182315 517200
rect 182263 517038 182271 517072
rect 182305 517038 182315 517072
rect 182263 517026 182315 517038
rect 183261 517072 183313 517200
rect 183261 517038 183271 517072
rect 183305 517038 183313 517072
rect 183261 517026 183313 517038
rect 183367 517072 183419 517200
rect 183367 517038 183375 517072
rect 183409 517038 183419 517072
rect 183367 517026 183419 517038
rect 184365 517072 184417 517200
rect 184365 517038 184375 517072
rect 184409 517038 184417 517072
rect 184365 517026 184417 517038
rect 184471 517174 184523 517200
rect 184471 517140 184479 517174
rect 184513 517140 184523 517174
rect 184471 517072 184523 517140
rect 184471 517038 184479 517072
rect 184513 517038 184523 517072
rect 184471 517026 184523 517038
rect 184917 517174 184969 517200
rect 184917 517140 184927 517174
rect 184961 517140 184969 517174
rect 184917 517072 184969 517140
rect 184917 517038 184927 517072
rect 184961 517038 184969 517072
rect 185207 517072 185259 517200
rect 184917 517026 184969 517038
rect 185207 517038 185215 517072
rect 185249 517038 185259 517072
rect 185207 517026 185259 517038
rect 186205 517072 186257 517200
rect 186205 517038 186215 517072
rect 186249 517038 186257 517072
rect 186205 517026 186257 517038
rect 186311 517174 186363 517200
rect 186311 517140 186319 517174
rect 186353 517140 186363 517174
rect 186311 517072 186363 517140
rect 186311 517038 186319 517072
rect 186353 517038 186363 517072
rect 186311 517026 186363 517038
rect 186941 517174 186993 517200
rect 186941 517140 186951 517174
rect 186985 517140 186993 517174
rect 186941 517072 186993 517140
rect 186941 517038 186951 517072
rect 186985 517038 186993 517072
rect 186941 517026 186993 517038
rect 187231 517167 187283 517200
rect 187231 517133 187239 517167
rect 187273 517133 187283 517167
rect 187231 517072 187283 517133
rect 187231 517038 187239 517072
rect 187273 517038 187283 517072
rect 187231 517026 187283 517038
rect 187401 517167 187453 517200
rect 187401 517133 187411 517167
rect 187445 517133 187453 517167
rect 187401 517072 187453 517133
rect 187401 517038 187411 517072
rect 187445 517038 187453 517072
rect 187401 517026 187453 517038
rect 172235 516920 172287 516932
rect 172235 516886 172243 516920
rect 172277 516886 172287 516920
rect 172235 516825 172287 516886
rect 172235 516791 172243 516825
rect 172277 516791 172287 516825
rect 172235 516758 172287 516791
rect 172405 516920 172457 516932
rect 172405 516886 172415 516920
rect 172449 516886 172457 516920
rect 172405 516825 172457 516886
rect 172405 516791 172415 516825
rect 172449 516791 172457 516825
rect 172405 516758 172457 516791
rect 172511 516920 172563 516932
rect 172511 516886 172519 516920
rect 172553 516886 172563 516920
rect 172511 516758 172563 516886
rect 173509 516920 173561 516932
rect 173509 516886 173519 516920
rect 173553 516886 173561 516920
rect 173509 516758 173561 516886
rect 173615 516920 173667 516932
rect 173615 516886 173623 516920
rect 173657 516886 173667 516920
rect 173615 516758 173667 516886
rect 174613 516920 174665 516932
rect 174613 516886 174623 516920
rect 174657 516886 174665 516920
rect 174613 516758 174665 516886
rect 174719 516920 174771 516932
rect 174719 516886 174727 516920
rect 174761 516886 174771 516920
rect 174719 516758 174771 516886
rect 175717 516920 175769 516932
rect 175717 516886 175727 516920
rect 175761 516886 175769 516920
rect 175717 516758 175769 516886
rect 175823 516920 175875 516932
rect 175823 516886 175831 516920
rect 175865 516886 175875 516920
rect 175823 516758 175875 516886
rect 176821 516920 176873 516932
rect 176821 516886 176831 516920
rect 176865 516886 176873 516920
rect 176821 516758 176873 516886
rect 176927 516920 176979 516932
rect 176927 516886 176935 516920
rect 176969 516886 176979 516920
rect 176927 516818 176979 516886
rect 176927 516784 176935 516818
rect 176969 516784 176979 516818
rect 176927 516758 176979 516784
rect 177189 516920 177241 516932
rect 177189 516886 177199 516920
rect 177233 516886 177241 516920
rect 177479 516920 177531 516932
rect 177189 516818 177241 516886
rect 177189 516784 177199 516818
rect 177233 516784 177241 516818
rect 177189 516758 177241 516784
rect 177479 516886 177487 516920
rect 177521 516886 177531 516920
rect 177479 516758 177531 516886
rect 178477 516920 178529 516932
rect 178477 516886 178487 516920
rect 178521 516886 178529 516920
rect 178477 516758 178529 516886
rect 178583 516920 178635 516932
rect 178583 516886 178591 516920
rect 178625 516886 178635 516920
rect 178583 516758 178635 516886
rect 179581 516920 179633 516932
rect 179581 516886 179591 516920
rect 179625 516886 179633 516920
rect 179581 516758 179633 516886
rect 179687 516920 179739 516932
rect 179687 516886 179695 516920
rect 179729 516886 179739 516920
rect 179687 516758 179739 516886
rect 180685 516920 180737 516932
rect 180685 516886 180695 516920
rect 180729 516886 180737 516920
rect 180685 516758 180737 516886
rect 180791 516920 180843 516932
rect 180791 516886 180799 516920
rect 180833 516886 180843 516920
rect 180791 516758 180843 516886
rect 181789 516920 181841 516932
rect 181789 516886 181799 516920
rect 181833 516886 181841 516920
rect 181789 516758 181841 516886
rect 181895 516920 181947 516932
rect 181895 516886 181903 516920
rect 181937 516886 181947 516920
rect 181895 516818 181947 516886
rect 181895 516784 181903 516818
rect 181937 516784 181947 516818
rect 181895 516758 181947 516784
rect 182341 516920 182393 516932
rect 182341 516886 182351 516920
rect 182385 516886 182393 516920
rect 182631 516920 182683 516932
rect 182341 516818 182393 516886
rect 182341 516784 182351 516818
rect 182385 516784 182393 516818
rect 182341 516758 182393 516784
rect 182631 516886 182639 516920
rect 182673 516886 182683 516920
rect 182631 516758 182683 516886
rect 183629 516920 183681 516932
rect 183629 516886 183639 516920
rect 183673 516886 183681 516920
rect 183629 516758 183681 516886
rect 183735 516920 183787 516932
rect 183735 516886 183743 516920
rect 183777 516886 183787 516920
rect 183735 516758 183787 516886
rect 184733 516920 184785 516932
rect 184733 516886 184743 516920
rect 184777 516886 184785 516920
rect 184733 516758 184785 516886
rect 184839 516920 184891 516932
rect 184839 516886 184847 516920
rect 184881 516886 184891 516920
rect 184839 516758 184891 516886
rect 185837 516920 185889 516932
rect 185837 516886 185847 516920
rect 185881 516886 185889 516920
rect 185837 516758 185889 516886
rect 185943 516920 185995 516932
rect 185943 516886 185951 516920
rect 185985 516886 185995 516920
rect 185943 516758 185995 516886
rect 186941 516920 186993 516932
rect 186941 516886 186951 516920
rect 186985 516886 186993 516920
rect 186941 516758 186993 516886
rect 187231 516920 187283 516932
rect 187231 516886 187239 516920
rect 187273 516886 187283 516920
rect 187231 516825 187283 516886
rect 187231 516791 187239 516825
rect 187273 516791 187283 516825
rect 187231 516758 187283 516791
rect 187401 516920 187453 516932
rect 187401 516886 187411 516920
rect 187445 516886 187453 516920
rect 187401 516825 187453 516886
rect 187401 516791 187411 516825
rect 187445 516791 187453 516825
rect 187401 516758 187453 516791
rect 172235 516079 172287 516112
rect 172235 516045 172243 516079
rect 172277 516045 172287 516079
rect 172235 515984 172287 516045
rect 172235 515950 172243 515984
rect 172277 515950 172287 515984
rect 172235 515938 172287 515950
rect 172405 516079 172457 516112
rect 172405 516045 172415 516079
rect 172449 516045 172457 516079
rect 172405 515984 172457 516045
rect 172405 515950 172415 515984
rect 172449 515950 172457 515984
rect 172405 515938 172457 515950
rect 172511 515984 172563 516112
rect 172511 515950 172519 515984
rect 172553 515950 172563 515984
rect 172511 515938 172563 515950
rect 173509 515984 173561 516112
rect 173509 515950 173519 515984
rect 173553 515950 173561 515984
rect 173509 515938 173561 515950
rect 173615 515984 173667 516112
rect 173615 515950 173623 515984
rect 173657 515950 173667 515984
rect 173615 515938 173667 515950
rect 174613 515984 174665 516112
rect 174613 515950 174623 515984
rect 174657 515950 174665 515984
rect 174903 515984 174955 516112
rect 174613 515938 174665 515950
rect 174903 515950 174911 515984
rect 174945 515950 174955 515984
rect 174903 515938 174955 515950
rect 175901 515984 175953 516112
rect 175901 515950 175911 515984
rect 175945 515950 175953 515984
rect 175901 515938 175953 515950
rect 176007 515984 176059 516112
rect 176007 515950 176015 515984
rect 176049 515950 176059 515984
rect 176007 515938 176059 515950
rect 177005 515984 177057 516112
rect 177005 515950 177015 515984
rect 177049 515950 177057 515984
rect 177005 515938 177057 515950
rect 177111 515984 177163 516112
rect 177111 515950 177119 515984
rect 177153 515950 177163 515984
rect 177111 515938 177163 515950
rect 178109 515984 178161 516112
rect 178109 515950 178119 515984
rect 178153 515950 178161 515984
rect 178109 515938 178161 515950
rect 178215 515984 178267 516112
rect 178215 515950 178223 515984
rect 178257 515950 178267 515984
rect 178215 515938 178267 515950
rect 179213 515984 179265 516112
rect 179213 515950 179223 515984
rect 179257 515950 179265 515984
rect 179213 515938 179265 515950
rect 179319 516086 179371 516112
rect 179319 516052 179327 516086
rect 179361 516052 179371 516086
rect 179319 515984 179371 516052
rect 179319 515950 179327 515984
rect 179361 515950 179371 515984
rect 179319 515938 179371 515950
rect 179765 516086 179817 516112
rect 179765 516052 179775 516086
rect 179809 516052 179817 516086
rect 179765 515984 179817 516052
rect 179765 515950 179775 515984
rect 179809 515950 179817 515984
rect 180055 515984 180107 516112
rect 179765 515938 179817 515950
rect 180055 515950 180063 515984
rect 180097 515950 180107 515984
rect 180055 515938 180107 515950
rect 181053 515984 181105 516112
rect 181053 515950 181063 515984
rect 181097 515950 181105 515984
rect 181053 515938 181105 515950
rect 181159 515984 181211 516112
rect 181159 515950 181167 515984
rect 181201 515950 181211 515984
rect 181159 515938 181211 515950
rect 182157 515984 182209 516112
rect 182157 515950 182167 515984
rect 182201 515950 182209 515984
rect 182157 515938 182209 515950
rect 182263 515984 182315 516112
rect 182263 515950 182271 515984
rect 182305 515950 182315 515984
rect 182263 515938 182315 515950
rect 183261 515984 183313 516112
rect 183261 515950 183271 515984
rect 183305 515950 183313 515984
rect 183261 515938 183313 515950
rect 183367 515984 183419 516112
rect 183367 515950 183375 515984
rect 183409 515950 183419 515984
rect 183367 515938 183419 515950
rect 184365 515984 184417 516112
rect 184365 515950 184375 515984
rect 184409 515950 184417 515984
rect 184365 515938 184417 515950
rect 184471 516086 184523 516112
rect 184471 516052 184479 516086
rect 184513 516052 184523 516086
rect 184471 515984 184523 516052
rect 184471 515950 184479 515984
rect 184513 515950 184523 515984
rect 184471 515938 184523 515950
rect 184917 516086 184969 516112
rect 184917 516052 184927 516086
rect 184961 516052 184969 516086
rect 184917 515984 184969 516052
rect 184917 515950 184927 515984
rect 184961 515950 184969 515984
rect 185207 515984 185259 516112
rect 184917 515938 184969 515950
rect 185207 515950 185215 515984
rect 185249 515950 185259 515984
rect 185207 515938 185259 515950
rect 186205 515984 186257 516112
rect 186205 515950 186215 515984
rect 186249 515950 186257 515984
rect 186205 515938 186257 515950
rect 186311 516086 186363 516112
rect 186311 516052 186319 516086
rect 186353 516052 186363 516086
rect 186311 515984 186363 516052
rect 186311 515950 186319 515984
rect 186353 515950 186363 515984
rect 186311 515938 186363 515950
rect 186941 516086 186993 516112
rect 186941 516052 186951 516086
rect 186985 516052 186993 516086
rect 186941 515984 186993 516052
rect 186941 515950 186951 515984
rect 186985 515950 186993 515984
rect 186941 515938 186993 515950
rect 187231 516079 187283 516112
rect 187231 516045 187239 516079
rect 187273 516045 187283 516079
rect 187231 515984 187283 516045
rect 187231 515950 187239 515984
rect 187273 515950 187283 515984
rect 187231 515938 187283 515950
rect 187401 516079 187453 516112
rect 187401 516045 187411 516079
rect 187445 516045 187453 516079
rect 187401 515984 187453 516045
rect 187401 515950 187411 515984
rect 187445 515950 187453 515984
rect 187401 515938 187453 515950
rect 172235 515832 172287 515844
rect 172235 515798 172243 515832
rect 172277 515798 172287 515832
rect 172235 515737 172287 515798
rect 172235 515703 172243 515737
rect 172277 515703 172287 515737
rect 172235 515670 172287 515703
rect 172405 515832 172457 515844
rect 172405 515798 172415 515832
rect 172449 515798 172457 515832
rect 172405 515737 172457 515798
rect 172405 515703 172415 515737
rect 172449 515703 172457 515737
rect 172405 515670 172457 515703
rect 172511 515832 172563 515844
rect 172511 515798 172519 515832
rect 172553 515798 172563 515832
rect 172511 515730 172563 515798
rect 172511 515696 172519 515730
rect 172553 515696 172563 515730
rect 172511 515670 172563 515696
rect 173141 515832 173193 515844
rect 173141 515798 173151 515832
rect 173185 515798 173193 515832
rect 173141 515730 173193 515798
rect 173141 515696 173151 515730
rect 173185 515696 173193 515730
rect 173141 515670 173193 515696
rect 173431 515824 173484 515844
rect 173431 515790 173439 515824
rect 173473 515790 173484 515824
rect 173431 515702 173484 515790
rect 173431 515668 173439 515702
rect 173473 515668 173484 515702
rect 173431 515644 173484 515668
rect 173514 515832 173580 515844
rect 173514 515798 173525 515832
rect 173559 515798 173580 515832
rect 173514 515764 173580 515798
rect 173514 515730 173525 515764
rect 173559 515730 173580 515764
rect 173514 515644 173580 515730
rect 173610 515797 173666 515844
rect 173610 515763 173621 515797
rect 173655 515763 173666 515797
rect 173610 515644 173666 515763
rect 173696 515832 173752 515844
rect 173696 515798 173707 515832
rect 173741 515798 173752 515832
rect 173696 515644 173752 515798
rect 173782 515824 173838 515844
rect 173782 515790 173793 515824
rect 173827 515790 173838 515824
rect 173782 515756 173838 515790
rect 173782 515722 173793 515756
rect 173827 515722 173838 515756
rect 173782 515688 173838 515722
rect 173782 515654 173793 515688
rect 173827 515654 173838 515688
rect 173782 515644 173838 515654
rect 173868 515818 173928 515844
rect 173868 515784 173879 515818
rect 173913 515784 173928 515818
rect 173868 515750 173928 515784
rect 173868 515716 173879 515750
rect 173913 515716 173928 515750
rect 173868 515644 173928 515716
rect 173983 515832 174035 515844
rect 173983 515798 173991 515832
rect 174025 515798 174035 515832
rect 173983 515730 174035 515798
rect 173983 515696 173991 515730
rect 174025 515696 174035 515730
rect 173983 515670 174035 515696
rect 174613 515832 174665 515844
rect 174613 515798 174623 515832
rect 174657 515798 174665 515832
rect 174903 515832 174955 515844
rect 174613 515730 174665 515798
rect 174613 515696 174623 515730
rect 174657 515696 174665 515730
rect 174613 515670 174665 515696
rect 174903 515798 174911 515832
rect 174945 515798 174955 515832
rect 174903 515670 174955 515798
rect 175901 515832 175953 515844
rect 175901 515798 175911 515832
rect 175945 515798 175953 515832
rect 175901 515670 175953 515798
rect 176007 515832 176059 515844
rect 176007 515798 176015 515832
rect 176049 515798 176059 515832
rect 176007 515670 176059 515798
rect 177005 515832 177057 515844
rect 177005 515798 177015 515832
rect 177049 515798 177057 515832
rect 177005 515670 177057 515798
rect 177111 515832 177163 515844
rect 177111 515798 177119 515832
rect 177153 515798 177163 515832
rect 177111 515737 177163 515798
rect 177111 515703 177119 515737
rect 177153 515703 177163 515737
rect 177111 515670 177163 515703
rect 177281 515832 177333 515844
rect 177281 515798 177291 515832
rect 177325 515798 177333 515832
rect 177479 515832 177531 515844
rect 177281 515737 177333 515798
rect 177281 515703 177291 515737
rect 177325 515703 177333 515737
rect 177281 515670 177333 515703
rect 177479 515798 177487 515832
rect 177521 515798 177531 515832
rect 177479 515670 177531 515798
rect 178477 515832 178529 515844
rect 178477 515798 178487 515832
rect 178521 515798 178529 515832
rect 178477 515670 178529 515798
rect 178583 515832 178635 515844
rect 178583 515798 178591 515832
rect 178625 515798 178635 515832
rect 178583 515670 178635 515798
rect 179581 515832 179633 515844
rect 179581 515798 179591 515832
rect 179625 515798 179633 515832
rect 179581 515670 179633 515798
rect 179687 515832 179739 515844
rect 179687 515798 179695 515832
rect 179729 515798 179739 515832
rect 179687 515737 179739 515798
rect 179687 515703 179695 515737
rect 179729 515703 179739 515737
rect 179687 515670 179739 515703
rect 179857 515832 179909 515844
rect 179857 515798 179867 515832
rect 179901 515798 179909 515832
rect 180055 515832 180107 515844
rect 179857 515737 179909 515798
rect 179857 515703 179867 515737
rect 179901 515703 179909 515737
rect 179857 515670 179909 515703
rect 180055 515798 180063 515832
rect 180097 515798 180107 515832
rect 180055 515670 180107 515798
rect 181053 515832 181105 515844
rect 181053 515798 181063 515832
rect 181097 515798 181105 515832
rect 181053 515670 181105 515798
rect 181159 515832 181211 515844
rect 181159 515798 181167 515832
rect 181201 515798 181211 515832
rect 181159 515730 181211 515798
rect 181159 515696 181167 515730
rect 181201 515696 181211 515730
rect 181159 515670 181211 515696
rect 181789 515832 181841 515844
rect 181789 515798 181799 515832
rect 181833 515798 181841 515832
rect 181789 515730 181841 515798
rect 181789 515696 181799 515730
rect 181833 515696 181841 515730
rect 181789 515670 181841 515696
rect 182079 515824 182131 515844
rect 182079 515790 182087 515824
rect 182121 515790 182131 515824
rect 182079 515743 182131 515790
rect 182079 515709 182087 515743
rect 182121 515709 182131 515743
rect 182079 515686 182131 515709
rect 182161 515824 182219 515844
rect 182161 515790 182173 515824
rect 182207 515790 182219 515824
rect 182161 515756 182219 515790
rect 182161 515722 182173 515756
rect 182207 515722 182219 515756
rect 182161 515686 182219 515722
rect 182249 515824 182301 515844
rect 182631 515832 182683 515844
rect 182249 515790 182259 515824
rect 182293 515790 182301 515824
rect 182249 515756 182301 515790
rect 182249 515722 182259 515756
rect 182293 515722 182301 515756
rect 182249 515686 182301 515722
rect 182631 515798 182639 515832
rect 182673 515798 182683 515832
rect 182631 515670 182683 515798
rect 183629 515832 183681 515844
rect 183629 515798 183639 515832
rect 183673 515798 183681 515832
rect 183629 515670 183681 515798
rect 183735 515832 183787 515844
rect 183735 515798 183743 515832
rect 183777 515798 183787 515832
rect 183735 515670 183787 515798
rect 184733 515832 184785 515844
rect 184733 515798 184743 515832
rect 184777 515798 184785 515832
rect 184733 515670 184785 515798
rect 184839 515832 184891 515844
rect 184839 515798 184847 515832
rect 184881 515798 184891 515832
rect 184839 515737 184891 515798
rect 184839 515703 184847 515737
rect 184881 515703 184891 515737
rect 184839 515670 184891 515703
rect 185009 515832 185061 515844
rect 185009 515798 185019 515832
rect 185053 515798 185061 515832
rect 185207 515832 185259 515844
rect 185009 515737 185061 515798
rect 185009 515703 185019 515737
rect 185053 515703 185061 515737
rect 185009 515670 185061 515703
rect 185207 515798 185215 515832
rect 185249 515798 185259 515832
rect 185207 515670 185259 515798
rect 186205 515832 186257 515844
rect 186205 515798 186215 515832
rect 186249 515798 186257 515832
rect 186205 515670 186257 515798
rect 186403 515824 186456 515844
rect 186403 515790 186411 515824
rect 186445 515790 186456 515824
rect 186403 515702 186456 515790
rect 186403 515668 186411 515702
rect 186445 515668 186456 515702
rect 186403 515644 186456 515668
rect 186486 515832 186552 515844
rect 186486 515798 186497 515832
rect 186531 515798 186552 515832
rect 186486 515764 186552 515798
rect 186486 515730 186497 515764
rect 186531 515730 186552 515764
rect 186486 515644 186552 515730
rect 186582 515797 186638 515844
rect 186582 515763 186593 515797
rect 186627 515763 186638 515797
rect 186582 515644 186638 515763
rect 186668 515832 186724 515844
rect 186668 515798 186679 515832
rect 186713 515798 186724 515832
rect 186668 515644 186724 515798
rect 186754 515824 186810 515844
rect 186754 515790 186765 515824
rect 186799 515790 186810 515824
rect 186754 515756 186810 515790
rect 186754 515722 186765 515756
rect 186799 515722 186810 515756
rect 186754 515688 186810 515722
rect 186754 515654 186765 515688
rect 186799 515654 186810 515688
rect 186754 515644 186810 515654
rect 186840 515818 186900 515844
rect 186840 515784 186851 515818
rect 186885 515784 186900 515818
rect 186840 515750 186900 515784
rect 186840 515716 186851 515750
rect 186885 515716 186900 515750
rect 186840 515644 186900 515716
rect 186955 515832 187007 515844
rect 186955 515798 186963 515832
rect 186997 515798 187007 515832
rect 186955 515737 187007 515798
rect 186955 515703 186963 515737
rect 186997 515703 187007 515737
rect 186955 515670 187007 515703
rect 187125 515832 187177 515844
rect 187125 515798 187135 515832
rect 187169 515798 187177 515832
rect 187125 515737 187177 515798
rect 187125 515703 187135 515737
rect 187169 515703 187177 515737
rect 187125 515670 187177 515703
rect 187231 515832 187283 515844
rect 187231 515798 187239 515832
rect 187273 515798 187283 515832
rect 187231 515737 187283 515798
rect 187231 515703 187239 515737
rect 187273 515703 187283 515737
rect 187231 515670 187283 515703
rect 187401 515832 187453 515844
rect 187401 515798 187411 515832
rect 187445 515798 187453 515832
rect 187401 515737 187453 515798
rect 187401 515703 187411 515737
rect 187445 515703 187453 515737
rect 187401 515670 187453 515703
<< ndiffc >>
rect 164684 540059 164718 541035
rect 164772 540059 164806 541035
rect 164887 540066 164921 541042
rect 164983 540066 165017 541042
rect 165079 540066 165113 541042
rect 165175 540066 165209 541042
rect 165271 540066 165305 541042
rect 165367 540066 165401 541042
rect 165463 540066 165497 541042
rect 165559 540066 165593 541042
rect 165655 540066 165689 541042
rect 165751 540066 165785 541042
rect 165847 540066 165881 541042
rect 165943 540066 165977 541042
rect 166039 540066 166073 541042
rect 166164 540059 166198 540235
rect 166252 540059 166286 540235
rect 166364 540059 166398 541035
rect 166452 540059 166486 541035
rect 168484 540059 168518 541035
rect 168572 540059 168606 541035
rect 168687 540066 168721 541042
rect 168783 540066 168817 541042
rect 168879 540066 168913 541042
rect 168975 540066 169009 541042
rect 169071 540066 169105 541042
rect 169167 540066 169201 541042
rect 169263 540066 169297 541042
rect 169359 540066 169393 541042
rect 169455 540066 169489 541042
rect 169551 540066 169585 541042
rect 169647 540066 169681 541042
rect 169743 540066 169777 541042
rect 169839 540066 169873 541042
rect 169964 540059 169998 540235
rect 170052 540059 170086 540235
rect 170164 540059 170198 541035
rect 170252 540059 170286 541035
rect 172184 540059 172218 541035
rect 172272 540059 172306 541035
rect 172387 540066 172421 541042
rect 172483 540066 172517 541042
rect 172579 540066 172613 541042
rect 172675 540066 172709 541042
rect 172771 540066 172805 541042
rect 172867 540066 172901 541042
rect 172963 540066 172997 541042
rect 173059 540066 173093 541042
rect 173155 540066 173189 541042
rect 173251 540066 173285 541042
rect 173347 540066 173381 541042
rect 173443 540066 173477 541042
rect 173539 540066 173573 541042
rect 173664 540059 173698 540235
rect 173752 540059 173786 540235
rect 173864 540059 173898 541035
rect 173952 540059 173986 541035
rect 175684 540059 175718 541035
rect 175772 540059 175806 541035
rect 175887 540066 175921 541042
rect 175983 540066 176017 541042
rect 176079 540066 176113 541042
rect 176175 540066 176209 541042
rect 176271 540066 176305 541042
rect 176367 540066 176401 541042
rect 176463 540066 176497 541042
rect 176559 540066 176593 541042
rect 176655 540066 176689 541042
rect 176751 540066 176785 541042
rect 176847 540066 176881 541042
rect 176943 540066 176977 541042
rect 177039 540066 177073 541042
rect 177164 540059 177198 540235
rect 177252 540059 177286 540235
rect 177364 540059 177398 541035
rect 177452 540059 177486 541035
rect 179284 540059 179318 541035
rect 179372 540059 179406 541035
rect 179487 540066 179521 541042
rect 179583 540066 179617 541042
rect 179679 540066 179713 541042
rect 179775 540066 179809 541042
rect 179871 540066 179905 541042
rect 179967 540066 180001 541042
rect 180063 540066 180097 541042
rect 180159 540066 180193 541042
rect 180255 540066 180289 541042
rect 180351 540066 180385 541042
rect 180447 540066 180481 541042
rect 180543 540066 180577 541042
rect 180639 540066 180673 541042
rect 180764 540059 180798 540235
rect 180852 540059 180886 540235
rect 180964 540059 180998 541035
rect 181052 540059 181086 541035
rect 182584 540059 182618 541035
rect 182672 540059 182706 541035
rect 182787 540066 182821 541042
rect 182883 540066 182917 541042
rect 182979 540066 183013 541042
rect 183075 540066 183109 541042
rect 183171 540066 183205 541042
rect 183267 540066 183301 541042
rect 183363 540066 183397 541042
rect 183459 540066 183493 541042
rect 183555 540066 183589 541042
rect 183651 540066 183685 541042
rect 183747 540066 183781 541042
rect 183843 540066 183877 541042
rect 183939 540066 183973 541042
rect 184064 540059 184098 540235
rect 184152 540059 184186 540235
rect 184264 540059 184298 541035
rect 184352 540059 184386 541035
rect 185884 540059 185918 541035
rect 185972 540059 186006 541035
rect 186087 540066 186121 541042
rect 186183 540066 186217 541042
rect 186279 540066 186313 541042
rect 186375 540066 186409 541042
rect 186471 540066 186505 541042
rect 186567 540066 186601 541042
rect 186663 540066 186697 541042
rect 186759 540066 186793 541042
rect 186855 540066 186889 541042
rect 186951 540066 186985 541042
rect 187047 540066 187081 541042
rect 187143 540066 187177 541042
rect 187239 540066 187273 541042
rect 187364 540059 187398 540235
rect 187452 540059 187486 540235
rect 187564 540059 187598 541035
rect 187652 540059 187686 541035
rect 189184 540059 189218 541035
rect 189272 540059 189306 541035
rect 189387 540066 189421 541042
rect 189483 540066 189517 541042
rect 189579 540066 189613 541042
rect 189675 540066 189709 541042
rect 189771 540066 189805 541042
rect 189867 540066 189901 541042
rect 189963 540066 189997 541042
rect 190059 540066 190093 541042
rect 190155 540066 190189 541042
rect 190251 540066 190285 541042
rect 190347 540066 190381 541042
rect 190443 540066 190477 541042
rect 190539 540066 190573 541042
rect 190664 540059 190698 540235
rect 190752 540059 190786 540235
rect 190864 540059 190898 541035
rect 190952 540059 190986 541035
rect 158664 538209 158698 538385
rect 158922 538209 158956 538385
rect 159040 538209 159074 538385
rect 159298 538209 159332 538385
rect 159556 538209 159590 538385
rect 159814 538209 159848 538385
rect 160072 538209 160106 538385
rect 160330 538209 160364 538385
rect 160588 538209 160622 538385
rect 160846 538209 160880 538385
rect 161104 538209 161138 538385
rect 161362 538209 161396 538385
rect 161484 538209 161518 538385
rect 161742 538209 161776 538385
rect 161884 538209 161918 538385
rect 162142 538209 162176 538385
rect 162264 538209 162298 538385
rect 162522 538209 162556 538385
rect 172243 530465 172277 530499
rect 172415 530465 172449 530499
rect 172526 530482 172560 530516
rect 172612 530460 172646 530494
rect 172698 530482 172732 530516
rect 172784 530460 172818 530494
rect 172881 530482 172915 530516
rect 172967 530478 173001 530512
rect 173071 530467 173105 530501
rect 174071 530467 174105 530501
rect 174175 530467 174209 530501
rect 174623 530467 174657 530501
rect 174918 530482 174952 530516
rect 175004 530460 175038 530494
rect 175090 530482 175124 530516
rect 175176 530460 175210 530494
rect 175273 530482 175307 530516
rect 175359 530478 175393 530512
rect 175555 530436 175589 530470
rect 175639 530486 175673 530520
rect 175763 530470 175797 530504
rect 175981 530490 176015 530524
rect 176193 530486 176227 530520
rect 176303 530490 176337 530524
rect 176415 530486 176449 530520
rect 176761 530484 176795 530518
rect 176868 530484 176902 530518
rect 177001 530490 177035 530524
rect 177123 530460 177157 530494
rect 177207 530486 177241 530520
rect 177291 530460 177325 530494
rect 177690 530460 177724 530494
rect 177780 530486 177814 530520
rect 177939 530460 177973 530494
rect 178043 530460 178077 530494
rect 178197 530486 178231 530520
rect 178281 530460 178315 530494
rect 178407 530456 178441 530490
rect 178493 530486 178527 530520
rect 178579 530473 178613 530507
rect 178690 530482 178724 530516
rect 178776 530460 178810 530494
rect 178862 530482 178896 530516
rect 178948 530460 178982 530494
rect 179045 530482 179079 530516
rect 179131 530478 179165 530512
rect 179235 530478 179269 530512
rect 179321 530482 179355 530516
rect 179418 530460 179452 530494
rect 179504 530482 179538 530516
rect 179590 530460 179624 530494
rect 179676 530482 179710 530516
rect 180247 530467 180281 530501
rect 180331 530486 180365 530520
rect 180538 530471 180572 530505
rect 180773 530471 180807 530505
rect 180841 530471 180875 530505
rect 180925 530471 180959 530505
rect 181213 530471 181247 530505
rect 181297 530471 181331 530505
rect 181365 530471 181399 530505
rect 181600 530471 181634 530505
rect 181807 530486 181841 530520
rect 181891 530467 181925 530501
rect 181995 530478 182029 530512
rect 182081 530482 182115 530516
rect 182178 530460 182212 530494
rect 182264 530482 182298 530516
rect 182350 530460 182384 530494
rect 182436 530482 182470 530516
rect 182639 530460 182673 530494
rect 182903 530460 182937 530494
rect 183099 530478 183133 530512
rect 183185 530482 183219 530516
rect 183282 530460 183316 530494
rect 183368 530482 183402 530516
rect 183454 530460 183488 530494
rect 183540 530482 183574 530516
rect 183651 530467 183685 530501
rect 184651 530467 184685 530501
rect 184755 530460 184789 530494
rect 185019 530460 185053 530494
rect 185215 530478 185249 530512
rect 185301 530482 185335 530516
rect 185398 530460 185432 530494
rect 185484 530482 185518 530516
rect 185570 530460 185604 530494
rect 185656 530482 185690 530516
rect 185767 530467 185801 530501
rect 186767 530467 186801 530501
rect 187239 530465 187273 530499
rect 187411 530465 187445 530499
rect 172243 529571 172277 529605
rect 172415 529571 172449 529605
rect 172519 529569 172553 529603
rect 173519 529569 173553 529603
rect 173623 529569 173657 529603
rect 174623 529569 174657 529603
rect 174841 529576 174875 529610
rect 174925 529550 174959 529584
rect 175079 529576 175113 529610
rect 175183 529576 175217 529610
rect 175342 529550 175376 529584
rect 175432 529576 175466 529610
rect 175555 529576 175589 529610
rect 175639 529550 175673 529584
rect 175723 529576 175757 529610
rect 175845 529546 175879 529580
rect 175978 529552 176012 529586
rect 176085 529552 176119 529586
rect 176431 529550 176465 529584
rect 176543 529546 176577 529580
rect 176653 529550 176687 529584
rect 176865 529546 176899 529580
rect 177083 529566 177117 529600
rect 177207 529550 177241 529584
rect 177291 529600 177325 529634
rect 177625 529565 177659 529599
rect 177709 529565 177743 529599
rect 177777 529565 177811 529599
rect 178012 529565 178046 529599
rect 178219 529550 178253 529584
rect 178303 529569 178337 529603
rect 178407 529600 178441 529634
rect 178491 529550 178525 529584
rect 178615 529566 178649 529600
rect 178833 529546 178867 529580
rect 179045 529550 179079 529584
rect 179155 529546 179189 529580
rect 179267 529550 179301 529584
rect 179613 529552 179647 529586
rect 179720 529552 179754 529586
rect 179853 529546 179887 529580
rect 179975 529576 180009 529610
rect 180059 529550 180093 529584
rect 180143 529576 180177 529610
rect 180247 529576 180281 529610
rect 180331 529550 180365 529584
rect 180415 529576 180449 529610
rect 180537 529546 180571 529580
rect 180670 529552 180704 529586
rect 180777 529552 180811 529586
rect 181123 529550 181157 529584
rect 181235 529546 181269 529580
rect 181345 529550 181379 529584
rect 181557 529546 181591 529580
rect 181775 529566 181809 529600
rect 181899 529550 181933 529584
rect 181983 529600 182017 529634
rect 182087 529576 182121 529610
rect 182351 529576 182385 529610
rect 182658 529576 182692 529610
rect 182748 529550 182782 529584
rect 182907 529576 182941 529610
rect 183011 529576 183045 529610
rect 183165 529550 183199 529584
rect 183249 529576 183283 529610
rect 183375 529569 183409 529603
rect 184375 529569 184409 529603
rect 184479 529569 184513 529603
rect 185479 529569 185513 529603
rect 185583 529569 185617 529603
rect 186583 529569 186617 529603
rect 186687 529569 186721 529603
rect 187135 529569 187169 529603
rect 187239 529571 187273 529605
rect 187411 529571 187445 529605
rect 172243 529377 172277 529411
rect 172415 529377 172449 529411
rect 172519 529379 172553 529413
rect 173519 529379 173553 529413
rect 173623 529379 173657 529413
rect 174623 529379 174657 529413
rect 175141 529383 175175 529417
rect 175225 529383 175259 529417
rect 175293 529383 175327 529417
rect 175528 529383 175562 529417
rect 175735 529398 175769 529432
rect 175819 529379 175853 529413
rect 175940 529394 175974 529428
rect 176026 529385 176060 529419
rect 176112 529394 176146 529428
rect 176198 529385 176232 529419
rect 176284 529394 176318 529428
rect 176370 529385 176404 529419
rect 176456 529394 176490 529428
rect 176542 529385 176576 529419
rect 176627 529394 176661 529428
rect 176713 529385 176747 529419
rect 176799 529394 176833 529428
rect 176885 529385 176919 529419
rect 176971 529394 177005 529428
rect 177057 529385 177091 529419
rect 177143 529394 177177 529428
rect 177229 529385 177263 529419
rect 177315 529385 177349 529419
rect 177401 529385 177435 529419
rect 177487 529385 177521 529419
rect 177573 529385 177607 529419
rect 177659 529398 177693 529432
rect 177763 529372 177797 529406
rect 177847 529398 177881 529432
rect 177931 529372 177965 529406
rect 178053 529402 178087 529436
rect 178186 529396 178220 529430
rect 178293 529396 178327 529430
rect 178639 529398 178673 529432
rect 178751 529402 178785 529436
rect 178861 529398 178895 529432
rect 179073 529402 179107 529436
rect 179291 529382 179325 529416
rect 179415 529398 179449 529432
rect 179499 529348 179533 529382
rect 179695 529385 179729 529419
rect 179781 529398 179815 529432
rect 179867 529368 179901 529402
rect 180063 529379 180097 529413
rect 180511 529379 180545 529413
rect 180707 529398 180741 529432
rect 180793 529385 180827 529419
rect 180879 529385 180913 529419
rect 180965 529385 180999 529419
rect 181051 529385 181085 529419
rect 181137 529385 181171 529419
rect 181223 529394 181257 529428
rect 181309 529385 181343 529419
rect 181395 529394 181429 529428
rect 181481 529385 181515 529419
rect 181567 529394 181601 529428
rect 181653 529385 181687 529419
rect 181739 529394 181773 529428
rect 181824 529385 181858 529419
rect 181910 529394 181944 529428
rect 181996 529385 182030 529419
rect 182082 529394 182116 529428
rect 182168 529385 182202 529419
rect 182254 529394 182288 529428
rect 182340 529385 182374 529419
rect 182426 529394 182460 529428
rect 182547 529368 182581 529402
rect 182633 529398 182667 529432
rect 182719 529385 182753 529419
rect 182823 529379 182857 529413
rect 183823 529379 183857 529413
rect 183927 529379 183961 529413
rect 184927 529379 184961 529413
rect 185215 529379 185249 529413
rect 186215 529379 186249 529413
rect 186319 529379 186353 529413
rect 186951 529379 186985 529413
rect 187239 529377 187273 529411
rect 187411 529377 187445 529411
rect 172243 528483 172277 528517
rect 172415 528483 172449 528517
rect 172519 528481 172553 528515
rect 173519 528481 173553 528515
rect 173623 528481 173657 528515
rect 174623 528481 174657 528515
rect 174727 528481 174761 528515
rect 175727 528481 175761 528515
rect 175923 528475 175957 528509
rect 176009 528462 176043 528496
rect 176095 528492 176129 528526
rect 176199 528475 176233 528509
rect 176285 528462 176319 528496
rect 176371 528492 176405 528526
rect 176521 528477 176555 528511
rect 176605 528477 176639 528511
rect 176673 528477 176707 528511
rect 176908 528477 176942 528511
rect 177115 528462 177149 528496
rect 177199 528481 177233 528515
rect 177506 528488 177540 528522
rect 177596 528462 177630 528496
rect 177755 528488 177789 528522
rect 177859 528488 177893 528522
rect 178013 528462 178047 528496
rect 178097 528488 178131 528522
rect 178407 528462 178441 528496
rect 178493 528475 178527 528509
rect 178579 528475 178613 528509
rect 178665 528475 178699 528509
rect 178751 528475 178785 528509
rect 178837 528475 178871 528509
rect 178923 528466 178957 528500
rect 179009 528475 179043 528509
rect 179095 528466 179129 528500
rect 179181 528475 179215 528509
rect 179267 528466 179301 528500
rect 179353 528475 179387 528509
rect 179439 528466 179473 528500
rect 179524 528475 179558 528509
rect 179610 528466 179644 528500
rect 179696 528475 179730 528509
rect 179782 528466 179816 528500
rect 179868 528475 179902 528509
rect 179954 528466 179988 528500
rect 180040 528475 180074 528509
rect 180126 528466 180160 528500
rect 180247 528475 180281 528509
rect 180333 528462 180367 528496
rect 180419 528492 180453 528526
rect 180523 528488 180557 528522
rect 180607 528462 180641 528496
rect 180691 528488 180725 528522
rect 180813 528458 180847 528492
rect 180946 528464 180980 528498
rect 181053 528464 181087 528498
rect 181399 528462 181433 528496
rect 181511 528458 181545 528492
rect 181621 528462 181655 528496
rect 181833 528458 181867 528492
rect 182051 528478 182085 528512
rect 182175 528462 182209 528496
rect 182259 528512 182293 528546
rect 182639 528481 182673 528515
rect 183639 528481 183673 528515
rect 183743 528481 183777 528515
rect 184743 528481 184777 528515
rect 184847 528481 184881 528515
rect 185847 528481 185881 528515
rect 185951 528481 185985 528515
rect 186951 528481 186985 528515
rect 187239 528483 187273 528517
rect 187411 528483 187445 528517
rect 172243 528289 172277 528323
rect 172415 528289 172449 528323
rect 172519 528291 172553 528325
rect 173519 528291 173553 528325
rect 173623 528291 173657 528325
rect 174623 528291 174657 528325
rect 174911 528291 174945 528325
rect 175911 528291 175945 528325
rect 176107 528284 176141 528318
rect 176191 528310 176225 528344
rect 176275 528284 176309 528318
rect 176397 528314 176431 528348
rect 176530 528308 176564 528342
rect 176637 528308 176671 528342
rect 176983 528310 177017 528344
rect 177095 528314 177129 528348
rect 177205 528310 177239 528344
rect 177417 528314 177451 528348
rect 177635 528294 177669 528328
rect 177759 528310 177793 528344
rect 177843 528260 177877 528294
rect 177947 528280 177981 528314
rect 178033 528310 178067 528344
rect 178119 528297 178153 528331
rect 178223 528291 178257 528325
rect 178855 528291 178889 528325
rect 178959 528291 178993 528325
rect 179043 528310 179077 528344
rect 179250 528295 179284 528329
rect 179485 528295 179519 528329
rect 179553 528295 179587 528329
rect 179637 528295 179671 528329
rect 180063 528291 180097 528325
rect 180695 528291 180729 528325
rect 180983 528291 181017 528325
rect 181067 528310 181101 528344
rect 181274 528295 181308 528329
rect 181509 528295 181543 528329
rect 181577 528295 181611 528329
rect 181661 528295 181695 528329
rect 181811 528291 181845 528325
rect 182811 528291 182845 528325
rect 182915 528291 182949 528325
rect 183915 528291 183949 528325
rect 184019 528291 184053 528325
rect 185019 528291 185053 528325
rect 185215 528291 185249 528325
rect 186215 528291 186249 528325
rect 186319 528291 186353 528325
rect 186951 528291 186985 528325
rect 187239 528289 187273 528323
rect 187411 528289 187445 528323
rect 172243 527395 172277 527429
rect 172415 527395 172449 527429
rect 172519 527393 172553 527427
rect 173519 527393 173553 527427
rect 173623 527393 173657 527427
rect 174623 527393 174657 527427
rect 174727 527393 174761 527427
rect 175727 527393 175761 527427
rect 175831 527393 175865 527427
rect 176279 527393 176313 527427
rect 176402 527400 176436 527434
rect 176492 527374 176526 527408
rect 176651 527400 176685 527434
rect 176755 527400 176789 527434
rect 176909 527374 176943 527408
rect 176993 527400 177027 527434
rect 177119 527395 177153 527429
rect 177291 527395 177325 527429
rect 177487 527393 177521 527427
rect 178487 527393 178521 527427
rect 178591 527400 178625 527434
rect 178855 527400 178889 527434
rect 178978 527400 179012 527434
rect 179068 527374 179102 527408
rect 179227 527400 179261 527434
rect 179331 527400 179365 527434
rect 179485 527374 179519 527408
rect 179569 527400 179603 527434
rect 179695 527393 179729 527427
rect 180695 527393 180729 527427
rect 180799 527393 180833 527427
rect 181799 527393 181833 527427
rect 181903 527393 181937 527427
rect 182351 527393 182385 527427
rect 182639 527393 182673 527427
rect 183639 527393 183673 527427
rect 183743 527393 183777 527427
rect 184743 527393 184777 527427
rect 184847 527393 184881 527427
rect 185847 527393 185881 527427
rect 185951 527393 185985 527427
rect 186951 527393 186985 527427
rect 187239 527395 187273 527429
rect 187411 527395 187445 527429
rect 172243 527201 172277 527235
rect 172415 527201 172449 527235
rect 172519 527203 172553 527237
rect 173519 527203 173553 527237
rect 173623 527203 173657 527237
rect 174623 527203 174657 527237
rect 174911 527203 174945 527237
rect 175911 527203 175945 527237
rect 176015 527203 176049 527237
rect 177015 527203 177049 527237
rect 177119 527203 177153 527237
rect 178119 527203 178153 527237
rect 178223 527203 178257 527237
rect 179223 527203 179257 527237
rect 179327 527203 179361 527237
rect 179775 527203 179809 527237
rect 180063 527203 180097 527237
rect 181063 527203 181097 527237
rect 181167 527203 181201 527237
rect 182167 527203 182201 527237
rect 182271 527203 182305 527237
rect 183271 527203 183305 527237
rect 183375 527203 183409 527237
rect 184375 527203 184409 527237
rect 184479 527203 184513 527237
rect 184927 527203 184961 527237
rect 185215 527203 185249 527237
rect 186215 527203 186249 527237
rect 186319 527203 186353 527237
rect 186951 527203 186985 527237
rect 187239 527201 187273 527235
rect 187411 527201 187445 527235
rect 172243 526307 172277 526341
rect 172415 526307 172449 526341
rect 172519 526305 172553 526339
rect 173519 526305 173553 526339
rect 173623 526305 173657 526339
rect 174623 526305 174657 526339
rect 174727 526305 174761 526339
rect 175727 526305 175761 526339
rect 175831 526305 175865 526339
rect 176831 526305 176865 526339
rect 176935 526312 176969 526346
rect 177199 526312 177233 526346
rect 177487 526305 177521 526339
rect 178487 526305 178521 526339
rect 178591 526305 178625 526339
rect 179591 526305 179625 526339
rect 179695 526305 179729 526339
rect 180695 526305 180729 526339
rect 180799 526305 180833 526339
rect 181799 526305 181833 526339
rect 181903 526305 181937 526339
rect 182351 526305 182385 526339
rect 182639 526305 182673 526339
rect 183639 526305 183673 526339
rect 183743 526305 183777 526339
rect 184743 526305 184777 526339
rect 184847 526305 184881 526339
rect 185847 526305 185881 526339
rect 185951 526305 185985 526339
rect 186951 526305 186985 526339
rect 187239 526307 187273 526341
rect 187411 526307 187445 526341
rect 172243 526113 172277 526147
rect 172415 526113 172449 526147
rect 172519 526115 172553 526149
rect 173519 526115 173553 526149
rect 173623 526115 173657 526149
rect 174623 526115 174657 526149
rect 174911 526115 174945 526149
rect 175911 526115 175945 526149
rect 176015 526115 176049 526149
rect 177015 526115 177049 526149
rect 177119 526115 177153 526149
rect 178119 526115 178153 526149
rect 178223 526115 178257 526149
rect 179223 526115 179257 526149
rect 179327 526115 179361 526149
rect 179775 526115 179809 526149
rect 180063 526115 180097 526149
rect 181063 526115 181097 526149
rect 181167 526115 181201 526149
rect 182167 526115 182201 526149
rect 182271 526115 182305 526149
rect 183271 526115 183305 526149
rect 183375 526115 183409 526149
rect 184375 526115 184409 526149
rect 184479 526115 184513 526149
rect 184927 526115 184961 526149
rect 185215 526115 185249 526149
rect 186215 526115 186249 526149
rect 186319 526115 186353 526149
rect 186951 526115 186985 526149
rect 187239 526113 187273 526147
rect 187411 526113 187445 526147
rect 172243 525219 172277 525253
rect 172415 525219 172449 525253
rect 172519 525217 172553 525251
rect 173519 525217 173553 525251
rect 173623 525217 173657 525251
rect 174623 525217 174657 525251
rect 174727 525217 174761 525251
rect 175727 525217 175761 525251
rect 175831 525217 175865 525251
rect 176831 525217 176865 525251
rect 176935 525224 176969 525258
rect 177199 525224 177233 525258
rect 177487 525217 177521 525251
rect 178487 525217 178521 525251
rect 178591 525217 178625 525251
rect 179591 525217 179625 525251
rect 179695 525217 179729 525251
rect 180695 525217 180729 525251
rect 180799 525217 180833 525251
rect 181799 525217 181833 525251
rect 181903 525217 181937 525251
rect 182351 525217 182385 525251
rect 182639 525217 182673 525251
rect 183639 525217 183673 525251
rect 183743 525217 183777 525251
rect 184743 525217 184777 525251
rect 184847 525217 184881 525251
rect 185847 525217 185881 525251
rect 185951 525217 185985 525251
rect 186951 525217 186985 525251
rect 187239 525219 187273 525253
rect 187411 525219 187445 525253
rect 172243 525025 172277 525059
rect 172415 525025 172449 525059
rect 172519 525027 172553 525061
rect 173519 525027 173553 525061
rect 173623 525027 173657 525061
rect 174623 525027 174657 525061
rect 174911 525027 174945 525061
rect 175911 525027 175945 525061
rect 176015 525027 176049 525061
rect 177015 525027 177049 525061
rect 177119 525027 177153 525061
rect 178119 525027 178153 525061
rect 178223 525027 178257 525061
rect 179223 525027 179257 525061
rect 179327 525027 179361 525061
rect 179775 525027 179809 525061
rect 180063 525027 180097 525061
rect 181063 525027 181097 525061
rect 181167 525027 181201 525061
rect 182167 525027 182201 525061
rect 182271 525027 182305 525061
rect 183271 525027 183305 525061
rect 183375 525027 183409 525061
rect 184375 525027 184409 525061
rect 184479 525027 184513 525061
rect 184927 525027 184961 525061
rect 185215 525027 185249 525061
rect 186215 525027 186249 525061
rect 186319 525027 186353 525061
rect 186951 525027 186985 525061
rect 187239 525025 187273 525059
rect 187411 525025 187445 525059
rect 172243 524131 172277 524165
rect 172415 524131 172449 524165
rect 172519 524129 172553 524163
rect 173519 524129 173553 524163
rect 173623 524129 173657 524163
rect 174623 524129 174657 524163
rect 174727 524129 174761 524163
rect 175727 524129 175761 524163
rect 175831 524129 175865 524163
rect 176831 524129 176865 524163
rect 176935 524136 176969 524170
rect 177199 524136 177233 524170
rect 177487 524129 177521 524163
rect 178487 524129 178521 524163
rect 178591 524129 178625 524163
rect 179591 524129 179625 524163
rect 179695 524129 179729 524163
rect 180695 524129 180729 524163
rect 180799 524129 180833 524163
rect 181799 524129 181833 524163
rect 181903 524129 181937 524163
rect 182351 524129 182385 524163
rect 182639 524129 182673 524163
rect 183639 524129 183673 524163
rect 183743 524129 183777 524163
rect 184743 524129 184777 524163
rect 184847 524129 184881 524163
rect 185847 524129 185881 524163
rect 185951 524129 185985 524163
rect 186951 524129 186985 524163
rect 187239 524131 187273 524165
rect 187411 524131 187445 524165
rect 172243 523937 172277 523971
rect 172415 523937 172449 523971
rect 172519 523939 172553 523973
rect 173519 523939 173553 523973
rect 173623 523939 173657 523973
rect 174623 523939 174657 523973
rect 174911 523939 174945 523973
rect 175911 523939 175945 523973
rect 176015 523939 176049 523973
rect 177015 523939 177049 523973
rect 177119 523939 177153 523973
rect 178119 523939 178153 523973
rect 178223 523939 178257 523973
rect 179223 523939 179257 523973
rect 179327 523939 179361 523973
rect 179775 523939 179809 523973
rect 180063 523939 180097 523973
rect 181063 523939 181097 523973
rect 181167 523939 181201 523973
rect 182167 523939 182201 523973
rect 182271 523939 182305 523973
rect 183271 523939 183305 523973
rect 183375 523939 183409 523973
rect 184375 523939 184409 523973
rect 184479 523939 184513 523973
rect 184927 523939 184961 523973
rect 185215 523939 185249 523973
rect 186215 523939 186249 523973
rect 186319 523939 186353 523973
rect 186951 523939 186985 523973
rect 187239 523937 187273 523971
rect 187411 523937 187445 523971
rect 172243 523043 172277 523077
rect 172415 523043 172449 523077
rect 172519 523041 172553 523075
rect 173519 523041 173553 523075
rect 173623 523041 173657 523075
rect 174623 523041 174657 523075
rect 174727 523041 174761 523075
rect 175727 523041 175761 523075
rect 175831 523041 175865 523075
rect 176831 523041 176865 523075
rect 176935 523048 176969 523082
rect 177199 523048 177233 523082
rect 177487 523041 177521 523075
rect 178487 523041 178521 523075
rect 178591 523041 178625 523075
rect 179591 523041 179625 523075
rect 179695 523041 179729 523075
rect 180695 523041 180729 523075
rect 180799 523041 180833 523075
rect 181799 523041 181833 523075
rect 181903 523041 181937 523075
rect 182351 523041 182385 523075
rect 182639 523041 182673 523075
rect 183639 523041 183673 523075
rect 183743 523041 183777 523075
rect 184743 523041 184777 523075
rect 184847 523041 184881 523075
rect 185847 523041 185881 523075
rect 185951 523041 185985 523075
rect 186951 523041 186985 523075
rect 187239 523043 187273 523077
rect 187411 523043 187445 523077
rect 172243 522849 172277 522883
rect 172415 522849 172449 522883
rect 172519 522851 172553 522885
rect 173519 522851 173553 522885
rect 173623 522851 173657 522885
rect 174623 522851 174657 522885
rect 174911 522851 174945 522885
rect 175911 522851 175945 522885
rect 176015 522851 176049 522885
rect 177015 522851 177049 522885
rect 177119 522851 177153 522885
rect 178119 522851 178153 522885
rect 178223 522851 178257 522885
rect 179223 522851 179257 522885
rect 179327 522851 179361 522885
rect 179775 522851 179809 522885
rect 180063 522851 180097 522885
rect 181063 522851 181097 522885
rect 181167 522851 181201 522885
rect 182167 522851 182201 522885
rect 182271 522851 182305 522885
rect 183271 522851 183305 522885
rect 183375 522851 183409 522885
rect 184375 522851 184409 522885
rect 184479 522851 184513 522885
rect 184927 522851 184961 522885
rect 185215 522851 185249 522885
rect 186215 522851 186249 522885
rect 186319 522851 186353 522885
rect 186951 522851 186985 522885
rect 187239 522849 187273 522883
rect 187411 522849 187445 522883
rect 172243 521955 172277 521989
rect 172415 521955 172449 521989
rect 172519 521953 172553 521987
rect 173519 521953 173553 521987
rect 173623 521953 173657 521987
rect 174623 521953 174657 521987
rect 174727 521953 174761 521987
rect 175727 521953 175761 521987
rect 175831 521953 175865 521987
rect 176831 521953 176865 521987
rect 176935 521960 176969 521994
rect 177199 521960 177233 521994
rect 177487 521953 177521 521987
rect 178487 521953 178521 521987
rect 178591 521953 178625 521987
rect 179591 521953 179625 521987
rect 179695 521953 179729 521987
rect 180695 521953 180729 521987
rect 180799 521953 180833 521987
rect 181799 521953 181833 521987
rect 181903 521953 181937 521987
rect 182351 521953 182385 521987
rect 182639 521953 182673 521987
rect 183639 521953 183673 521987
rect 183743 521953 183777 521987
rect 184743 521953 184777 521987
rect 184847 521953 184881 521987
rect 185847 521953 185881 521987
rect 185951 521953 185985 521987
rect 186951 521953 186985 521987
rect 187239 521955 187273 521989
rect 187411 521955 187445 521989
rect 172243 521761 172277 521795
rect 172415 521761 172449 521795
rect 172519 521763 172553 521797
rect 173519 521763 173553 521797
rect 173623 521763 173657 521797
rect 174623 521763 174657 521797
rect 174911 521763 174945 521797
rect 175911 521763 175945 521797
rect 176015 521763 176049 521797
rect 177015 521763 177049 521797
rect 177119 521763 177153 521797
rect 178119 521763 178153 521797
rect 178223 521763 178257 521797
rect 179223 521763 179257 521797
rect 179327 521763 179361 521797
rect 179775 521763 179809 521797
rect 180063 521763 180097 521797
rect 181063 521763 181097 521797
rect 181167 521763 181201 521797
rect 182167 521763 182201 521797
rect 182271 521763 182305 521797
rect 183271 521763 183305 521797
rect 183375 521763 183409 521797
rect 184375 521763 184409 521797
rect 184479 521763 184513 521797
rect 184927 521763 184961 521797
rect 185215 521763 185249 521797
rect 186215 521763 186249 521797
rect 186319 521763 186353 521797
rect 186951 521763 186985 521797
rect 187239 521761 187273 521795
rect 187411 521761 187445 521795
rect 172243 520867 172277 520901
rect 172415 520867 172449 520901
rect 172519 520865 172553 520899
rect 173519 520865 173553 520899
rect 173623 520865 173657 520899
rect 174623 520865 174657 520899
rect 174727 520865 174761 520899
rect 175727 520865 175761 520899
rect 175831 520865 175865 520899
rect 176831 520865 176865 520899
rect 176935 520872 176969 520906
rect 177199 520872 177233 520906
rect 177487 520865 177521 520899
rect 178487 520865 178521 520899
rect 178591 520865 178625 520899
rect 179591 520865 179625 520899
rect 179695 520865 179729 520899
rect 180695 520865 180729 520899
rect 180799 520865 180833 520899
rect 181799 520865 181833 520899
rect 181903 520865 181937 520899
rect 182351 520865 182385 520899
rect 182639 520865 182673 520899
rect 183639 520865 183673 520899
rect 183743 520865 183777 520899
rect 184743 520865 184777 520899
rect 184847 520865 184881 520899
rect 185847 520865 185881 520899
rect 185951 520865 185985 520899
rect 186951 520865 186985 520899
rect 187239 520867 187273 520901
rect 187411 520867 187445 520901
rect 172243 520673 172277 520707
rect 172415 520673 172449 520707
rect 172519 520675 172553 520709
rect 173519 520675 173553 520709
rect 173623 520675 173657 520709
rect 174623 520675 174657 520709
rect 174911 520675 174945 520709
rect 175911 520675 175945 520709
rect 176015 520675 176049 520709
rect 177015 520675 177049 520709
rect 177119 520675 177153 520709
rect 178119 520675 178153 520709
rect 178223 520675 178257 520709
rect 179223 520675 179257 520709
rect 179327 520675 179361 520709
rect 179775 520675 179809 520709
rect 180063 520675 180097 520709
rect 181063 520675 181097 520709
rect 181167 520675 181201 520709
rect 182167 520675 182201 520709
rect 182271 520675 182305 520709
rect 183271 520675 183305 520709
rect 183375 520675 183409 520709
rect 184375 520675 184409 520709
rect 184479 520675 184513 520709
rect 184927 520675 184961 520709
rect 185215 520675 185249 520709
rect 186215 520675 186249 520709
rect 186319 520675 186353 520709
rect 186951 520675 186985 520709
rect 187239 520673 187273 520707
rect 187411 520673 187445 520707
rect 172243 519779 172277 519813
rect 172415 519779 172449 519813
rect 172519 519777 172553 519811
rect 173519 519777 173553 519811
rect 173623 519777 173657 519811
rect 174623 519777 174657 519811
rect 174727 519777 174761 519811
rect 175727 519777 175761 519811
rect 175831 519777 175865 519811
rect 176831 519777 176865 519811
rect 176935 519784 176969 519818
rect 177199 519784 177233 519818
rect 177487 519777 177521 519811
rect 178487 519777 178521 519811
rect 178591 519777 178625 519811
rect 179591 519777 179625 519811
rect 179695 519777 179729 519811
rect 180695 519777 180729 519811
rect 180799 519777 180833 519811
rect 181799 519777 181833 519811
rect 181903 519777 181937 519811
rect 182351 519777 182385 519811
rect 182639 519777 182673 519811
rect 183639 519777 183673 519811
rect 183743 519777 183777 519811
rect 184743 519777 184777 519811
rect 184847 519777 184881 519811
rect 185847 519777 185881 519811
rect 185951 519777 185985 519811
rect 186951 519777 186985 519811
rect 187239 519779 187273 519813
rect 187411 519779 187445 519813
rect 172243 519585 172277 519619
rect 172415 519585 172449 519619
rect 172519 519587 172553 519621
rect 173519 519587 173553 519621
rect 173623 519587 173657 519621
rect 174623 519587 174657 519621
rect 174911 519587 174945 519621
rect 175911 519587 175945 519621
rect 176015 519587 176049 519621
rect 177015 519587 177049 519621
rect 177119 519587 177153 519621
rect 178119 519587 178153 519621
rect 178223 519587 178257 519621
rect 179223 519587 179257 519621
rect 179327 519587 179361 519621
rect 179775 519587 179809 519621
rect 180063 519587 180097 519621
rect 181063 519587 181097 519621
rect 181167 519587 181201 519621
rect 182167 519587 182201 519621
rect 182271 519587 182305 519621
rect 183271 519587 183305 519621
rect 183375 519587 183409 519621
rect 184375 519587 184409 519621
rect 184479 519587 184513 519621
rect 184927 519587 184961 519621
rect 185215 519587 185249 519621
rect 186215 519587 186249 519621
rect 186319 519587 186353 519621
rect 186951 519587 186985 519621
rect 187239 519585 187273 519619
rect 187411 519585 187445 519619
rect 172243 518691 172277 518725
rect 172415 518691 172449 518725
rect 172519 518689 172553 518723
rect 173519 518689 173553 518723
rect 173623 518689 173657 518723
rect 174623 518689 174657 518723
rect 174727 518689 174761 518723
rect 175727 518689 175761 518723
rect 175831 518689 175865 518723
rect 176831 518689 176865 518723
rect 176935 518696 176969 518730
rect 177199 518696 177233 518730
rect 177487 518689 177521 518723
rect 178487 518689 178521 518723
rect 178591 518689 178625 518723
rect 179591 518689 179625 518723
rect 179695 518689 179729 518723
rect 180695 518689 180729 518723
rect 180799 518689 180833 518723
rect 181799 518689 181833 518723
rect 181903 518689 181937 518723
rect 182351 518689 182385 518723
rect 182639 518689 182673 518723
rect 183639 518689 183673 518723
rect 183743 518689 183777 518723
rect 184743 518689 184777 518723
rect 184847 518689 184881 518723
rect 185847 518689 185881 518723
rect 185951 518689 185985 518723
rect 186951 518689 186985 518723
rect 187239 518691 187273 518725
rect 187411 518691 187445 518725
rect 172243 518497 172277 518531
rect 172415 518497 172449 518531
rect 172519 518499 172553 518533
rect 173519 518499 173553 518533
rect 173623 518499 173657 518533
rect 174623 518499 174657 518533
rect 174911 518499 174945 518533
rect 175911 518499 175945 518533
rect 176015 518499 176049 518533
rect 177015 518499 177049 518533
rect 177119 518499 177153 518533
rect 178119 518499 178153 518533
rect 178223 518499 178257 518533
rect 179223 518499 179257 518533
rect 179327 518499 179361 518533
rect 179775 518499 179809 518533
rect 180063 518499 180097 518533
rect 181063 518499 181097 518533
rect 181167 518499 181201 518533
rect 182167 518499 182201 518533
rect 182271 518499 182305 518533
rect 183271 518499 183305 518533
rect 183375 518499 183409 518533
rect 184375 518499 184409 518533
rect 184479 518499 184513 518533
rect 184927 518499 184961 518533
rect 185215 518499 185249 518533
rect 186215 518499 186249 518533
rect 186319 518499 186353 518533
rect 186951 518499 186985 518533
rect 187239 518497 187273 518531
rect 187411 518497 187445 518531
rect 172243 517603 172277 517637
rect 172415 517603 172449 517637
rect 172519 517601 172553 517635
rect 173519 517601 173553 517635
rect 173623 517601 173657 517635
rect 174623 517601 174657 517635
rect 174727 517601 174761 517635
rect 175727 517601 175761 517635
rect 175831 517601 175865 517635
rect 176831 517601 176865 517635
rect 176935 517608 176969 517642
rect 177199 517608 177233 517642
rect 177487 517601 177521 517635
rect 178487 517601 178521 517635
rect 178591 517601 178625 517635
rect 179591 517601 179625 517635
rect 179695 517601 179729 517635
rect 180695 517601 180729 517635
rect 180799 517601 180833 517635
rect 181799 517601 181833 517635
rect 181903 517601 181937 517635
rect 182351 517601 182385 517635
rect 182639 517601 182673 517635
rect 183639 517601 183673 517635
rect 183743 517601 183777 517635
rect 184743 517601 184777 517635
rect 184847 517601 184881 517635
rect 185847 517601 185881 517635
rect 185951 517601 185985 517635
rect 186951 517601 186985 517635
rect 187239 517603 187273 517637
rect 187411 517603 187445 517637
rect 172243 517409 172277 517443
rect 172415 517409 172449 517443
rect 172519 517411 172553 517445
rect 173519 517411 173553 517445
rect 173623 517411 173657 517445
rect 174623 517411 174657 517445
rect 174911 517411 174945 517445
rect 175911 517411 175945 517445
rect 176015 517411 176049 517445
rect 177015 517411 177049 517445
rect 177119 517411 177153 517445
rect 178119 517411 178153 517445
rect 178223 517411 178257 517445
rect 179223 517411 179257 517445
rect 179327 517411 179361 517445
rect 179775 517411 179809 517445
rect 180063 517411 180097 517445
rect 181063 517411 181097 517445
rect 181167 517411 181201 517445
rect 182167 517411 182201 517445
rect 182271 517411 182305 517445
rect 183271 517411 183305 517445
rect 183375 517411 183409 517445
rect 184375 517411 184409 517445
rect 184479 517411 184513 517445
rect 184927 517411 184961 517445
rect 185215 517411 185249 517445
rect 186215 517411 186249 517445
rect 186319 517411 186353 517445
rect 186951 517411 186985 517445
rect 187239 517409 187273 517443
rect 187411 517409 187445 517443
rect 172243 516515 172277 516549
rect 172415 516515 172449 516549
rect 172519 516513 172553 516547
rect 173519 516513 173553 516547
rect 173623 516513 173657 516547
rect 174623 516513 174657 516547
rect 174727 516513 174761 516547
rect 175727 516513 175761 516547
rect 175831 516513 175865 516547
rect 176831 516513 176865 516547
rect 176935 516520 176969 516554
rect 177199 516520 177233 516554
rect 177487 516513 177521 516547
rect 178487 516513 178521 516547
rect 178591 516513 178625 516547
rect 179591 516513 179625 516547
rect 179695 516513 179729 516547
rect 180695 516513 180729 516547
rect 180799 516513 180833 516547
rect 181799 516513 181833 516547
rect 181903 516513 181937 516547
rect 182351 516513 182385 516547
rect 182639 516513 182673 516547
rect 183639 516513 183673 516547
rect 183743 516513 183777 516547
rect 184743 516513 184777 516547
rect 184847 516513 184881 516547
rect 185847 516513 185881 516547
rect 185951 516513 185985 516547
rect 186951 516513 186985 516547
rect 187239 516515 187273 516549
rect 187411 516515 187445 516549
rect 172243 516321 172277 516355
rect 172415 516321 172449 516355
rect 172519 516323 172553 516357
rect 173519 516323 173553 516357
rect 173623 516323 173657 516357
rect 174623 516323 174657 516357
rect 174911 516323 174945 516357
rect 175911 516323 175945 516357
rect 176015 516323 176049 516357
rect 177015 516323 177049 516357
rect 177119 516323 177153 516357
rect 178119 516323 178153 516357
rect 178223 516323 178257 516357
rect 179223 516323 179257 516357
rect 179327 516323 179361 516357
rect 179775 516323 179809 516357
rect 180063 516323 180097 516357
rect 181063 516323 181097 516357
rect 181167 516323 181201 516357
rect 182167 516323 182201 516357
rect 182271 516323 182305 516357
rect 183271 516323 183305 516357
rect 183375 516323 183409 516357
rect 184375 516323 184409 516357
rect 184479 516323 184513 516357
rect 184927 516323 184961 516357
rect 185215 516323 185249 516357
rect 186215 516323 186249 516357
rect 186319 516323 186353 516357
rect 186951 516323 186985 516357
rect 187239 516321 187273 516355
rect 187411 516321 187445 516355
rect 172243 515427 172277 515461
rect 172415 515427 172449 515461
rect 172519 515425 172553 515459
rect 173151 515425 173185 515459
rect 173439 515414 173473 515448
rect 173525 515410 173559 515444
rect 173622 515432 173656 515466
rect 173708 515410 173742 515444
rect 173794 515432 173828 515466
rect 173880 515410 173914 515444
rect 173991 515425 174025 515459
rect 174623 515425 174657 515459
rect 174911 515425 174945 515459
rect 175911 515425 175945 515459
rect 176015 515425 176049 515459
rect 177015 515425 177049 515459
rect 177119 515427 177153 515461
rect 177291 515427 177325 515461
rect 177487 515425 177521 515459
rect 178487 515425 178521 515459
rect 178591 515425 178625 515459
rect 179591 515425 179625 515459
rect 179695 515427 179729 515461
rect 179867 515427 179901 515461
rect 180063 515425 180097 515459
rect 181063 515425 181097 515459
rect 181167 515425 181201 515459
rect 181799 515425 181833 515459
rect 182087 515436 182121 515470
rect 182173 515406 182207 515440
rect 182259 515419 182293 515453
rect 182639 515425 182673 515459
rect 183639 515425 183673 515459
rect 183743 515425 183777 515459
rect 184743 515425 184777 515459
rect 184847 515427 184881 515461
rect 185019 515427 185053 515461
rect 185215 515425 185249 515459
rect 186215 515425 186249 515459
rect 186411 515414 186445 515448
rect 186497 515410 186531 515444
rect 186594 515432 186628 515466
rect 186680 515410 186714 515444
rect 186766 515432 186800 515466
rect 186852 515410 186886 515444
rect 186963 515427 186997 515461
rect 187135 515427 187169 515461
rect 187239 515427 187273 515461
rect 187411 515427 187445 515461
<< pdiffc >>
rect 164668 538537 164702 539513
rect 164756 538537 164790 539513
rect 164891 538544 164925 539520
rect 164987 538544 165021 539520
rect 165083 538544 165117 539520
rect 165179 538544 165213 539520
rect 165275 538544 165309 539520
rect 165371 538544 165405 539520
rect 165467 538544 165501 539520
rect 165563 538544 165597 539520
rect 165659 538544 165693 539520
rect 165755 538544 165789 539520
rect 165851 538544 165885 539520
rect 165947 538544 165981 539520
rect 166043 538544 166077 539520
rect 166168 538937 166202 539513
rect 166256 538937 166290 539513
rect 166368 538537 166402 539513
rect 166456 538537 166490 539513
rect 168468 538537 168502 539513
rect 168556 538537 168590 539513
rect 168691 538544 168725 539520
rect 168787 538544 168821 539520
rect 168883 538544 168917 539520
rect 168979 538544 169013 539520
rect 169075 538544 169109 539520
rect 169171 538544 169205 539520
rect 169267 538544 169301 539520
rect 169363 538544 169397 539520
rect 169459 538544 169493 539520
rect 169555 538544 169589 539520
rect 169651 538544 169685 539520
rect 169747 538544 169781 539520
rect 169843 538544 169877 539520
rect 169968 538937 170002 539513
rect 170056 538937 170090 539513
rect 170168 538537 170202 539513
rect 170256 538537 170290 539513
rect 172168 538537 172202 539513
rect 172256 538537 172290 539513
rect 172391 538544 172425 539520
rect 172487 538544 172521 539520
rect 172583 538544 172617 539520
rect 172679 538544 172713 539520
rect 172775 538544 172809 539520
rect 172871 538544 172905 539520
rect 172967 538544 173001 539520
rect 173063 538544 173097 539520
rect 173159 538544 173193 539520
rect 173255 538544 173289 539520
rect 173351 538544 173385 539520
rect 173447 538544 173481 539520
rect 173543 538544 173577 539520
rect 173668 538937 173702 539513
rect 173756 538937 173790 539513
rect 173868 538537 173902 539513
rect 173956 538537 173990 539513
rect 175668 538537 175702 539513
rect 175756 538537 175790 539513
rect 175891 538544 175925 539520
rect 175987 538544 176021 539520
rect 176083 538544 176117 539520
rect 176179 538544 176213 539520
rect 176275 538544 176309 539520
rect 176371 538544 176405 539520
rect 176467 538544 176501 539520
rect 176563 538544 176597 539520
rect 176659 538544 176693 539520
rect 176755 538544 176789 539520
rect 176851 538544 176885 539520
rect 176947 538544 176981 539520
rect 177043 538544 177077 539520
rect 177168 538937 177202 539513
rect 177256 538937 177290 539513
rect 177368 538537 177402 539513
rect 177456 538537 177490 539513
rect 179268 538537 179302 539513
rect 179356 538537 179390 539513
rect 179491 538544 179525 539520
rect 179587 538544 179621 539520
rect 179683 538544 179717 539520
rect 179779 538544 179813 539520
rect 179875 538544 179909 539520
rect 179971 538544 180005 539520
rect 180067 538544 180101 539520
rect 180163 538544 180197 539520
rect 180259 538544 180293 539520
rect 180355 538544 180389 539520
rect 180451 538544 180485 539520
rect 180547 538544 180581 539520
rect 180643 538544 180677 539520
rect 180768 538937 180802 539513
rect 180856 538937 180890 539513
rect 180968 538537 181002 539513
rect 181056 538537 181090 539513
rect 182568 538537 182602 539513
rect 182656 538537 182690 539513
rect 182791 538544 182825 539520
rect 182887 538544 182921 539520
rect 182983 538544 183017 539520
rect 183079 538544 183113 539520
rect 183175 538544 183209 539520
rect 183271 538544 183305 539520
rect 183367 538544 183401 539520
rect 183463 538544 183497 539520
rect 183559 538544 183593 539520
rect 183655 538544 183689 539520
rect 183751 538544 183785 539520
rect 183847 538544 183881 539520
rect 183943 538544 183977 539520
rect 184068 538937 184102 539513
rect 184156 538937 184190 539513
rect 184268 538537 184302 539513
rect 184356 538537 184390 539513
rect 185868 538537 185902 539513
rect 185956 538537 185990 539513
rect 186091 538544 186125 539520
rect 186187 538544 186221 539520
rect 186283 538544 186317 539520
rect 186379 538544 186413 539520
rect 186475 538544 186509 539520
rect 186571 538544 186605 539520
rect 186667 538544 186701 539520
rect 186763 538544 186797 539520
rect 186859 538544 186893 539520
rect 186955 538544 186989 539520
rect 187051 538544 187085 539520
rect 187147 538544 187181 539520
rect 187243 538544 187277 539520
rect 187368 538937 187402 539513
rect 187456 538937 187490 539513
rect 187568 538537 187602 539513
rect 187656 538537 187690 539513
rect 189168 538537 189202 539513
rect 189256 538537 189290 539513
rect 189391 538544 189425 539520
rect 189487 538544 189521 539520
rect 189583 538544 189617 539520
rect 189679 538544 189713 539520
rect 189775 538544 189809 539520
rect 189871 538544 189905 539520
rect 189967 538544 190001 539520
rect 190063 538544 190097 539520
rect 190159 538544 190193 539520
rect 190255 538544 190289 539520
rect 190351 538544 190385 539520
rect 190447 538544 190481 539520
rect 190543 538544 190577 539520
rect 190668 538937 190702 539513
rect 190756 538937 190790 539513
rect 190868 538537 190902 539513
rect 190956 538537 190990 539513
rect 161258 537037 161292 537613
rect 161346 537037 161380 537613
rect 161458 537037 161492 537613
rect 161554 537037 161588 537613
rect 161650 537037 161684 537613
rect 161746 537037 161780 537613
rect 161858 537037 161892 537613
rect 161954 537037 161988 537613
rect 162050 537037 162084 537613
rect 162146 537037 162180 537613
rect 162278 537037 162312 537613
rect 162366 537037 162400 537613
rect 157748 536017 157782 536593
rect 158006 536017 158040 536593
rect 158126 536017 158160 536593
rect 158384 536017 158418 536593
rect 158642 536017 158676 536593
rect 158900 536017 158934 536593
rect 159158 536017 159192 536593
rect 159416 536017 159450 536593
rect 159674 536017 159708 536593
rect 159932 536017 159966 536593
rect 160190 536017 160224 536593
rect 160448 536017 160482 536593
rect 160706 536017 160740 536593
rect 160832 536017 160866 536593
rect 161090 536017 161124 536593
rect 161348 536017 161382 536593
rect 161606 536017 161640 536593
rect 161730 536017 161764 536593
rect 161988 536017 162022 536593
rect 162246 536017 162280 536593
rect 162368 536017 162402 536593
rect 162626 536017 162660 536593
rect 172243 530189 172277 530223
rect 172243 530094 172277 530128
rect 172415 530189 172449 530223
rect 172415 530094 172449 530128
rect 172527 530176 172561 530210
rect 172527 530108 172561 530142
rect 172613 530238 172647 530272
rect 172613 530170 172647 530204
rect 172613 530102 172647 530136
rect 172699 530094 172733 530128
rect 172785 530129 172819 530163
rect 172881 530162 172915 530196
rect 172881 530094 172915 530128
rect 172967 530224 173001 530258
rect 172967 530102 173001 530136
rect 173071 530094 173105 530128
rect 174071 530094 174105 530128
rect 174175 530196 174209 530230
rect 174175 530094 174209 530128
rect 174623 530196 174657 530230
rect 174623 530094 174657 530128
rect 174919 530176 174953 530210
rect 174919 530108 174953 530142
rect 175005 530238 175039 530272
rect 175005 530170 175039 530204
rect 175005 530102 175039 530136
rect 175091 530094 175125 530128
rect 175177 530129 175211 530163
rect 175273 530162 175307 530196
rect 175273 530094 175307 530128
rect 175359 530224 175393 530258
rect 175359 530102 175393 530136
rect 175555 530198 175589 530232
rect 175555 530130 175589 530164
rect 175639 530162 175673 530196
rect 175639 530094 175673 530128
rect 175768 530094 175802 530128
rect 175854 530120 175888 530154
rect 175938 530094 175972 530128
rect 176130 530095 176164 530129
rect 176227 530102 176261 530136
rect 177123 530170 177157 530204
rect 176315 530094 176349 530128
rect 176428 530120 176462 530154
rect 176512 530104 176546 530138
rect 176609 530120 176643 530154
rect 176763 530096 176797 530130
rect 176856 530102 176890 530136
rect 176940 530094 176974 530128
rect 177123 530102 177157 530136
rect 177207 530118 177241 530152
rect 177291 530170 177325 530204
rect 177291 530102 177325 530136
rect 177690 530120 177724 530154
rect 178407 530183 178441 530217
rect 177780 530094 177814 530128
rect 177939 530120 177973 530154
rect 178043 530120 178077 530154
rect 178197 530094 178231 530128
rect 178281 530120 178315 530154
rect 178407 530102 178441 530136
rect 178493 530170 178527 530204
rect 178493 530102 178527 530136
rect 178579 530170 178613 530204
rect 178579 530102 178613 530136
rect 178691 530176 178725 530210
rect 178691 530108 178725 530142
rect 178777 530238 178811 530272
rect 178777 530170 178811 530204
rect 178777 530102 178811 530136
rect 178863 530094 178897 530128
rect 178949 530129 178983 530163
rect 179045 530162 179079 530196
rect 179045 530094 179079 530128
rect 179131 530224 179165 530258
rect 179131 530102 179165 530136
rect 179235 530224 179269 530258
rect 179235 530102 179269 530136
rect 179321 530162 179355 530196
rect 179321 530094 179355 530128
rect 179417 530129 179451 530163
rect 179503 530094 179537 530128
rect 179589 530238 179623 530272
rect 179589 530170 179623 530204
rect 179589 530102 179623 530136
rect 179675 530176 179709 530210
rect 179675 530108 179709 530142
rect 180247 530230 180281 530264
rect 180247 530162 180281 530196
rect 180247 530094 180281 530128
rect 180331 530230 180365 530264
rect 181807 530230 181841 530264
rect 180331 530162 180365 530196
rect 180331 530094 180365 530128
rect 180567 530154 180601 530188
rect 180642 530154 180676 530188
rect 180839 530154 180873 530188
rect 180925 530154 180959 530188
rect 181213 530154 181247 530188
rect 181299 530154 181333 530188
rect 181496 530154 181530 530188
rect 181571 530154 181605 530188
rect 181807 530162 181841 530196
rect 181807 530094 181841 530128
rect 181891 530230 181925 530264
rect 181891 530162 181925 530196
rect 181891 530094 181925 530128
rect 181995 530224 182029 530258
rect 181995 530102 182029 530136
rect 182081 530162 182115 530196
rect 182081 530094 182115 530128
rect 182177 530129 182211 530163
rect 182263 530094 182297 530128
rect 182349 530238 182383 530272
rect 182349 530170 182383 530204
rect 182349 530102 182383 530136
rect 182435 530176 182469 530210
rect 182435 530108 182469 530142
rect 182639 530196 182673 530230
rect 182639 530094 182673 530128
rect 182903 530196 182937 530230
rect 182903 530094 182937 530128
rect 183099 530224 183133 530258
rect 183099 530102 183133 530136
rect 183185 530162 183219 530196
rect 183185 530094 183219 530128
rect 183281 530129 183315 530163
rect 183367 530094 183401 530128
rect 183453 530238 183487 530272
rect 183453 530170 183487 530204
rect 183453 530102 183487 530136
rect 183539 530176 183573 530210
rect 183539 530108 183573 530142
rect 183651 530094 183685 530128
rect 184651 530094 184685 530128
rect 184755 530196 184789 530230
rect 184755 530094 184789 530128
rect 185019 530196 185053 530230
rect 185019 530094 185053 530128
rect 185215 530224 185249 530258
rect 185215 530102 185249 530136
rect 185301 530162 185335 530196
rect 185301 530094 185335 530128
rect 185397 530129 185431 530163
rect 185483 530094 185517 530128
rect 185569 530238 185603 530272
rect 185569 530170 185603 530204
rect 185569 530102 185603 530136
rect 185655 530176 185689 530210
rect 185655 530108 185689 530142
rect 185767 530094 185801 530128
rect 186767 530094 186801 530128
rect 187239 530189 187273 530223
rect 187239 530094 187273 530128
rect 187411 530189 187445 530223
rect 187411 530094 187445 530128
rect 172243 529942 172277 529976
rect 172243 529847 172277 529881
rect 172415 529942 172449 529976
rect 172415 529847 172449 529881
rect 172519 529942 172553 529976
rect 173519 529942 173553 529976
rect 173623 529942 173657 529976
rect 174623 529942 174657 529976
rect 174841 529916 174875 529950
rect 174925 529942 174959 529976
rect 175079 529916 175113 529950
rect 175183 529916 175217 529950
rect 175342 529942 175376 529976
rect 175432 529916 175466 529950
rect 175555 529934 175589 529968
rect 175555 529866 175589 529900
rect 175639 529918 175673 529952
rect 175723 529934 175757 529968
rect 175906 529942 175940 529976
rect 175990 529934 176024 529968
rect 176083 529940 176117 529974
rect 176237 529916 176271 529950
rect 176334 529932 176368 529966
rect 176418 529916 176452 529950
rect 176531 529942 176565 529976
rect 175723 529866 175757 529900
rect 176619 529934 176653 529968
rect 176716 529941 176750 529975
rect 176908 529942 176942 529976
rect 176992 529916 177026 529950
rect 177078 529942 177112 529976
rect 177207 529942 177241 529976
rect 177207 529874 177241 529908
rect 177291 529906 177325 529940
rect 177291 529838 177325 529872
rect 177625 529882 177659 529916
rect 177711 529882 177745 529916
rect 177908 529882 177942 529916
rect 177983 529882 178017 529916
rect 178219 529942 178253 529976
rect 178219 529874 178253 529908
rect 178219 529806 178253 529840
rect 178303 529942 178337 529976
rect 178303 529874 178337 529908
rect 178303 529806 178337 529840
rect 178407 529906 178441 529940
rect 178407 529838 178441 529872
rect 178491 529942 178525 529976
rect 178491 529874 178525 529908
rect 178620 529942 178654 529976
rect 178706 529916 178740 529950
rect 178790 529942 178824 529976
rect 178982 529941 179016 529975
rect 179079 529934 179113 529968
rect 179167 529942 179201 529976
rect 179280 529916 179314 529950
rect 179364 529932 179398 529966
rect 179461 529916 179495 529950
rect 179615 529940 179649 529974
rect 179708 529934 179742 529968
rect 179792 529942 179826 529976
rect 179975 529934 180009 529968
rect 179975 529866 180009 529900
rect 180059 529918 180093 529952
rect 180143 529934 180177 529968
rect 180143 529866 180177 529900
rect 180247 529934 180281 529968
rect 180247 529866 180281 529900
rect 180331 529918 180365 529952
rect 180415 529934 180449 529968
rect 180598 529942 180632 529976
rect 180682 529934 180716 529968
rect 180775 529940 180809 529974
rect 180929 529916 180963 529950
rect 181026 529932 181060 529966
rect 181110 529916 181144 529950
rect 181223 529942 181257 529976
rect 180415 529866 180449 529900
rect 181311 529934 181345 529968
rect 181408 529941 181442 529975
rect 181600 529942 181634 529976
rect 181684 529916 181718 529950
rect 181770 529942 181804 529976
rect 181899 529942 181933 529976
rect 181899 529874 181933 529908
rect 181983 529906 182017 529940
rect 181983 529838 182017 529872
rect 182087 529942 182121 529976
rect 182087 529840 182121 529874
rect 182351 529942 182385 529976
rect 182351 529840 182385 529874
rect 182658 529916 182692 529950
rect 182748 529942 182782 529976
rect 182907 529916 182941 529950
rect 183011 529916 183045 529950
rect 183165 529942 183199 529976
rect 183249 529916 183283 529950
rect 183375 529942 183409 529976
rect 184375 529942 184409 529976
rect 184479 529942 184513 529976
rect 185479 529942 185513 529976
rect 185583 529942 185617 529976
rect 186583 529942 186617 529976
rect 186687 529942 186721 529976
rect 186687 529840 186721 529874
rect 187135 529942 187169 529976
rect 187135 529840 187169 529874
rect 187239 529942 187273 529976
rect 187239 529847 187273 529881
rect 187411 529942 187445 529976
rect 187411 529847 187445 529881
rect 172243 529101 172277 529135
rect 172243 529006 172277 529040
rect 172415 529101 172449 529135
rect 172415 529006 172449 529040
rect 172519 529006 172553 529040
rect 173519 529006 173553 529040
rect 173623 529006 173657 529040
rect 174623 529006 174657 529040
rect 175735 529142 175769 529176
rect 175141 529066 175175 529100
rect 175227 529066 175261 529100
rect 175424 529066 175458 529100
rect 175499 529066 175533 529100
rect 175735 529074 175769 529108
rect 175735 529006 175769 529040
rect 175819 529142 175853 529176
rect 175819 529074 175853 529108
rect 175819 529006 175853 529040
rect 175940 529030 175974 529064
rect 176026 529136 176060 529170
rect 176026 529050 176060 529084
rect 176112 529030 176146 529064
rect 176198 529136 176232 529170
rect 176198 529050 176232 529084
rect 176284 529030 176318 529064
rect 176370 529136 176404 529170
rect 176370 529050 176404 529084
rect 176456 529030 176490 529064
rect 176542 529136 176576 529170
rect 176542 529050 176576 529084
rect 176627 529030 176661 529064
rect 176713 529136 176747 529170
rect 176713 529050 176747 529084
rect 176799 529030 176833 529064
rect 176885 529136 176919 529170
rect 176885 529050 176919 529084
rect 176971 529030 177005 529064
rect 177057 529136 177091 529170
rect 177057 529050 177091 529084
rect 177143 529030 177177 529064
rect 177229 529136 177263 529170
rect 177229 529050 177263 529084
rect 177315 529074 177349 529108
rect 177315 529006 177349 529040
rect 177401 529090 177435 529124
rect 177401 529022 177435 529056
rect 177487 529074 177521 529108
rect 177487 529006 177521 529040
rect 177573 529082 177607 529116
rect 177573 529014 177607 529048
rect 177659 529074 177693 529108
rect 177659 529006 177693 529040
rect 177763 529082 177797 529116
rect 177763 529014 177797 529048
rect 177847 529030 177881 529064
rect 177931 529082 177965 529116
rect 177931 529014 177965 529048
rect 178114 529006 178148 529040
rect 178198 529014 178232 529048
rect 178291 529008 178325 529042
rect 178445 529032 178479 529066
rect 178542 529016 178576 529050
rect 178626 529032 178660 529066
rect 178739 529006 178773 529040
rect 178827 529014 178861 529048
rect 178924 529007 178958 529041
rect 179116 529006 179150 529040
rect 179200 529032 179234 529066
rect 179286 529006 179320 529040
rect 179415 529074 179449 529108
rect 179415 529006 179449 529040
rect 179499 529110 179533 529144
rect 179499 529042 179533 529076
rect 179695 529082 179729 529116
rect 179695 529014 179729 529048
rect 179781 529082 179815 529116
rect 179781 529014 179815 529048
rect 179867 529095 179901 529129
rect 179867 529014 179901 529048
rect 180063 529108 180097 529142
rect 180063 529006 180097 529040
rect 180511 529108 180545 529142
rect 180511 529006 180545 529040
rect 180707 529074 180741 529108
rect 180707 529006 180741 529040
rect 180793 529082 180827 529116
rect 180793 529014 180827 529048
rect 180879 529074 180913 529108
rect 180879 529006 180913 529040
rect 180965 529090 180999 529124
rect 180965 529022 180999 529056
rect 181051 529074 181085 529108
rect 181051 529006 181085 529040
rect 181137 529136 181171 529170
rect 181137 529050 181171 529084
rect 181223 529030 181257 529064
rect 181309 529136 181343 529170
rect 181309 529050 181343 529084
rect 181395 529030 181429 529064
rect 181481 529136 181515 529170
rect 181481 529050 181515 529084
rect 181567 529030 181601 529064
rect 181653 529136 181687 529170
rect 181653 529050 181687 529084
rect 181739 529030 181773 529064
rect 181824 529136 181858 529170
rect 181824 529050 181858 529084
rect 181910 529030 181944 529064
rect 181996 529136 182030 529170
rect 181996 529050 182030 529084
rect 182082 529030 182116 529064
rect 182168 529136 182202 529170
rect 182168 529050 182202 529084
rect 182254 529030 182288 529064
rect 182340 529136 182374 529170
rect 182340 529050 182374 529084
rect 182426 529030 182460 529064
rect 182547 529095 182581 529129
rect 182547 529014 182581 529048
rect 182633 529082 182667 529116
rect 182633 529014 182667 529048
rect 182719 529082 182753 529116
rect 182719 529014 182753 529048
rect 182823 529006 182857 529040
rect 183823 529006 183857 529040
rect 183927 529006 183961 529040
rect 184927 529006 184961 529040
rect 185215 529006 185249 529040
rect 186215 529006 186249 529040
rect 186319 529108 186353 529142
rect 186319 529006 186353 529040
rect 186951 529108 186985 529142
rect 186951 529006 186985 529040
rect 187239 529101 187273 529135
rect 187239 529006 187273 529040
rect 187411 529101 187445 529135
rect 187411 529006 187445 529040
rect 172243 528854 172277 528888
rect 172243 528759 172277 528793
rect 172415 528854 172449 528888
rect 172415 528759 172449 528793
rect 172519 528854 172553 528888
rect 173519 528854 173553 528888
rect 173623 528854 173657 528888
rect 174623 528854 174657 528888
rect 174727 528854 174761 528888
rect 175727 528854 175761 528888
rect 175923 528846 175957 528880
rect 175923 528778 175957 528812
rect 176009 528846 176043 528880
rect 176009 528778 176043 528812
rect 176095 528846 176129 528880
rect 176095 528765 176129 528799
rect 176199 528846 176233 528880
rect 176199 528778 176233 528812
rect 176285 528846 176319 528880
rect 176285 528778 176319 528812
rect 176371 528846 176405 528880
rect 176371 528765 176405 528799
rect 176521 528794 176555 528828
rect 176607 528794 176641 528828
rect 176804 528794 176838 528828
rect 176879 528794 176913 528828
rect 177115 528854 177149 528888
rect 177115 528786 177149 528820
rect 177115 528718 177149 528752
rect 177199 528854 177233 528888
rect 177199 528786 177233 528820
rect 177199 528718 177233 528752
rect 177506 528828 177540 528862
rect 177596 528854 177630 528888
rect 177755 528828 177789 528862
rect 177859 528828 177893 528862
rect 178013 528854 178047 528888
rect 178097 528828 178131 528862
rect 178407 528854 178441 528888
rect 178407 528786 178441 528820
rect 178493 528846 178527 528880
rect 178493 528778 178527 528812
rect 178579 528854 178613 528888
rect 178579 528786 178613 528820
rect 178665 528838 178699 528872
rect 178665 528770 178699 528804
rect 178751 528854 178785 528888
rect 178751 528786 178785 528820
rect 178837 528810 178871 528844
rect 178837 528724 178871 528758
rect 178923 528830 178957 528864
rect 179009 528810 179043 528844
rect 179009 528724 179043 528758
rect 179095 528830 179129 528864
rect 179181 528810 179215 528844
rect 179181 528724 179215 528758
rect 179267 528830 179301 528864
rect 179353 528810 179387 528844
rect 179353 528724 179387 528758
rect 179439 528830 179473 528864
rect 179524 528810 179558 528844
rect 179524 528724 179558 528758
rect 179610 528830 179644 528864
rect 179696 528810 179730 528844
rect 179696 528724 179730 528758
rect 179782 528830 179816 528864
rect 179868 528810 179902 528844
rect 179868 528724 179902 528758
rect 179954 528830 179988 528864
rect 180040 528810 180074 528844
rect 180040 528724 180074 528758
rect 180126 528830 180160 528864
rect 180247 528846 180281 528880
rect 180247 528778 180281 528812
rect 180333 528846 180367 528880
rect 180333 528778 180367 528812
rect 180419 528846 180453 528880
rect 180419 528765 180453 528799
rect 180523 528846 180557 528880
rect 180523 528778 180557 528812
rect 180607 528830 180641 528864
rect 180691 528846 180725 528880
rect 180874 528854 180908 528888
rect 180958 528846 180992 528880
rect 181051 528852 181085 528886
rect 181205 528828 181239 528862
rect 181302 528844 181336 528878
rect 181386 528828 181420 528862
rect 181499 528854 181533 528888
rect 180691 528778 180725 528812
rect 181587 528846 181621 528880
rect 181684 528853 181718 528887
rect 181876 528854 181910 528888
rect 181960 528828 181994 528862
rect 182046 528854 182080 528888
rect 182175 528854 182209 528888
rect 182175 528786 182209 528820
rect 182259 528818 182293 528852
rect 182259 528750 182293 528784
rect 182639 528854 182673 528888
rect 183639 528854 183673 528888
rect 183743 528854 183777 528888
rect 184743 528854 184777 528888
rect 184847 528854 184881 528888
rect 185847 528854 185881 528888
rect 185951 528854 185985 528888
rect 186951 528854 186985 528888
rect 187239 528854 187273 528888
rect 187239 528759 187273 528793
rect 187411 528854 187445 528888
rect 187411 528759 187445 528793
rect 172243 528013 172277 528047
rect 172243 527918 172277 527952
rect 172415 528013 172449 528047
rect 172415 527918 172449 527952
rect 172519 527918 172553 527952
rect 173519 527918 173553 527952
rect 173623 527918 173657 527952
rect 174623 527918 174657 527952
rect 174911 527918 174945 527952
rect 175911 527918 175945 527952
rect 176107 527994 176141 528028
rect 176107 527926 176141 527960
rect 176191 527942 176225 527976
rect 176275 527994 176309 528028
rect 176275 527926 176309 527960
rect 176458 527918 176492 527952
rect 176542 527926 176576 527960
rect 176635 527920 176669 527954
rect 176789 527944 176823 527978
rect 176886 527928 176920 527962
rect 176970 527944 177004 527978
rect 177083 527918 177117 527952
rect 177171 527926 177205 527960
rect 177268 527919 177302 527953
rect 177460 527918 177494 527952
rect 177544 527944 177578 527978
rect 177630 527918 177664 527952
rect 177759 527986 177793 528020
rect 177759 527918 177793 527952
rect 177843 528022 177877 528056
rect 177843 527954 177877 527988
rect 177947 528007 177981 528041
rect 177947 527926 177981 527960
rect 178033 527994 178067 528028
rect 178033 527926 178067 527960
rect 178119 527994 178153 528028
rect 178119 527926 178153 527960
rect 178223 528020 178257 528054
rect 178223 527918 178257 527952
rect 178855 528020 178889 528054
rect 178855 527918 178889 527952
rect 178959 528054 178993 528088
rect 178959 527986 178993 528020
rect 178959 527918 178993 527952
rect 179043 528054 179077 528088
rect 179043 527986 179077 528020
rect 179043 527918 179077 527952
rect 179279 527978 179313 528012
rect 179354 527978 179388 528012
rect 179551 527978 179585 528012
rect 179637 527978 179671 528012
rect 180063 528020 180097 528054
rect 180063 527918 180097 527952
rect 180695 528020 180729 528054
rect 180695 527918 180729 527952
rect 180983 528054 181017 528088
rect 180983 527986 181017 528020
rect 180983 527918 181017 527952
rect 181067 528054 181101 528088
rect 181067 527986 181101 528020
rect 181067 527918 181101 527952
rect 181303 527978 181337 528012
rect 181378 527978 181412 528012
rect 181575 527978 181609 528012
rect 181661 527978 181695 528012
rect 181811 527918 181845 527952
rect 182811 527918 182845 527952
rect 182915 527918 182949 527952
rect 183915 527918 183949 527952
rect 184019 527918 184053 527952
rect 185019 527918 185053 527952
rect 185215 527918 185249 527952
rect 186215 527918 186249 527952
rect 186319 528020 186353 528054
rect 186319 527918 186353 527952
rect 186951 528020 186985 528054
rect 186951 527918 186985 527952
rect 187239 528013 187273 528047
rect 187239 527918 187273 527952
rect 187411 528013 187445 528047
rect 187411 527918 187445 527952
rect 172243 527766 172277 527800
rect 172243 527671 172277 527705
rect 172415 527766 172449 527800
rect 172415 527671 172449 527705
rect 172519 527766 172553 527800
rect 173519 527766 173553 527800
rect 173623 527766 173657 527800
rect 174623 527766 174657 527800
rect 174727 527766 174761 527800
rect 175727 527766 175761 527800
rect 175831 527766 175865 527800
rect 175831 527664 175865 527698
rect 176279 527766 176313 527800
rect 176279 527664 176313 527698
rect 176402 527740 176436 527774
rect 176492 527766 176526 527800
rect 176651 527740 176685 527774
rect 176755 527740 176789 527774
rect 176909 527766 176943 527800
rect 176993 527740 177027 527774
rect 177119 527766 177153 527800
rect 177119 527671 177153 527705
rect 177291 527766 177325 527800
rect 177291 527671 177325 527705
rect 177487 527766 177521 527800
rect 178487 527766 178521 527800
rect 178591 527766 178625 527800
rect 178591 527664 178625 527698
rect 178855 527766 178889 527800
rect 178855 527664 178889 527698
rect 178978 527740 179012 527774
rect 179068 527766 179102 527800
rect 179227 527740 179261 527774
rect 179331 527740 179365 527774
rect 179485 527766 179519 527800
rect 179569 527740 179603 527774
rect 179695 527766 179729 527800
rect 180695 527766 180729 527800
rect 180799 527766 180833 527800
rect 181799 527766 181833 527800
rect 181903 527766 181937 527800
rect 181903 527664 181937 527698
rect 182351 527766 182385 527800
rect 182351 527664 182385 527698
rect 182639 527766 182673 527800
rect 183639 527766 183673 527800
rect 183743 527766 183777 527800
rect 184743 527766 184777 527800
rect 184847 527766 184881 527800
rect 185847 527766 185881 527800
rect 185951 527766 185985 527800
rect 186951 527766 186985 527800
rect 187239 527766 187273 527800
rect 187239 527671 187273 527705
rect 187411 527766 187445 527800
rect 187411 527671 187445 527705
rect 172243 526925 172277 526959
rect 172243 526830 172277 526864
rect 172415 526925 172449 526959
rect 172415 526830 172449 526864
rect 172519 526830 172553 526864
rect 173519 526830 173553 526864
rect 173623 526830 173657 526864
rect 174623 526830 174657 526864
rect 174911 526830 174945 526864
rect 175911 526830 175945 526864
rect 176015 526830 176049 526864
rect 177015 526830 177049 526864
rect 177119 526830 177153 526864
rect 178119 526830 178153 526864
rect 178223 526830 178257 526864
rect 179223 526830 179257 526864
rect 179327 526932 179361 526966
rect 179327 526830 179361 526864
rect 179775 526932 179809 526966
rect 179775 526830 179809 526864
rect 180063 526830 180097 526864
rect 181063 526830 181097 526864
rect 181167 526830 181201 526864
rect 182167 526830 182201 526864
rect 182271 526830 182305 526864
rect 183271 526830 183305 526864
rect 183375 526830 183409 526864
rect 184375 526830 184409 526864
rect 184479 526932 184513 526966
rect 184479 526830 184513 526864
rect 184927 526932 184961 526966
rect 184927 526830 184961 526864
rect 185215 526830 185249 526864
rect 186215 526830 186249 526864
rect 186319 526932 186353 526966
rect 186319 526830 186353 526864
rect 186951 526932 186985 526966
rect 186951 526830 186985 526864
rect 187239 526925 187273 526959
rect 187239 526830 187273 526864
rect 187411 526925 187445 526959
rect 187411 526830 187445 526864
rect 172243 526678 172277 526712
rect 172243 526583 172277 526617
rect 172415 526678 172449 526712
rect 172415 526583 172449 526617
rect 172519 526678 172553 526712
rect 173519 526678 173553 526712
rect 173623 526678 173657 526712
rect 174623 526678 174657 526712
rect 174727 526678 174761 526712
rect 175727 526678 175761 526712
rect 175831 526678 175865 526712
rect 176831 526678 176865 526712
rect 176935 526678 176969 526712
rect 176935 526576 176969 526610
rect 177199 526678 177233 526712
rect 177199 526576 177233 526610
rect 177487 526678 177521 526712
rect 178487 526678 178521 526712
rect 178591 526678 178625 526712
rect 179591 526678 179625 526712
rect 179695 526678 179729 526712
rect 180695 526678 180729 526712
rect 180799 526678 180833 526712
rect 181799 526678 181833 526712
rect 181903 526678 181937 526712
rect 181903 526576 181937 526610
rect 182351 526678 182385 526712
rect 182351 526576 182385 526610
rect 182639 526678 182673 526712
rect 183639 526678 183673 526712
rect 183743 526678 183777 526712
rect 184743 526678 184777 526712
rect 184847 526678 184881 526712
rect 185847 526678 185881 526712
rect 185951 526678 185985 526712
rect 186951 526678 186985 526712
rect 187239 526678 187273 526712
rect 187239 526583 187273 526617
rect 187411 526678 187445 526712
rect 187411 526583 187445 526617
rect 172243 525837 172277 525871
rect 172243 525742 172277 525776
rect 172415 525837 172449 525871
rect 172415 525742 172449 525776
rect 172519 525742 172553 525776
rect 173519 525742 173553 525776
rect 173623 525742 173657 525776
rect 174623 525742 174657 525776
rect 174911 525742 174945 525776
rect 175911 525742 175945 525776
rect 176015 525742 176049 525776
rect 177015 525742 177049 525776
rect 177119 525742 177153 525776
rect 178119 525742 178153 525776
rect 178223 525742 178257 525776
rect 179223 525742 179257 525776
rect 179327 525844 179361 525878
rect 179327 525742 179361 525776
rect 179775 525844 179809 525878
rect 179775 525742 179809 525776
rect 180063 525742 180097 525776
rect 181063 525742 181097 525776
rect 181167 525742 181201 525776
rect 182167 525742 182201 525776
rect 182271 525742 182305 525776
rect 183271 525742 183305 525776
rect 183375 525742 183409 525776
rect 184375 525742 184409 525776
rect 184479 525844 184513 525878
rect 184479 525742 184513 525776
rect 184927 525844 184961 525878
rect 184927 525742 184961 525776
rect 185215 525742 185249 525776
rect 186215 525742 186249 525776
rect 186319 525844 186353 525878
rect 186319 525742 186353 525776
rect 186951 525844 186985 525878
rect 186951 525742 186985 525776
rect 187239 525837 187273 525871
rect 187239 525742 187273 525776
rect 187411 525837 187445 525871
rect 187411 525742 187445 525776
rect 172243 525590 172277 525624
rect 172243 525495 172277 525529
rect 172415 525590 172449 525624
rect 172415 525495 172449 525529
rect 172519 525590 172553 525624
rect 173519 525590 173553 525624
rect 173623 525590 173657 525624
rect 174623 525590 174657 525624
rect 174727 525590 174761 525624
rect 175727 525590 175761 525624
rect 175831 525590 175865 525624
rect 176831 525590 176865 525624
rect 176935 525590 176969 525624
rect 176935 525488 176969 525522
rect 177199 525590 177233 525624
rect 177199 525488 177233 525522
rect 177487 525590 177521 525624
rect 178487 525590 178521 525624
rect 178591 525590 178625 525624
rect 179591 525590 179625 525624
rect 179695 525590 179729 525624
rect 180695 525590 180729 525624
rect 180799 525590 180833 525624
rect 181799 525590 181833 525624
rect 181903 525590 181937 525624
rect 181903 525488 181937 525522
rect 182351 525590 182385 525624
rect 182351 525488 182385 525522
rect 182639 525590 182673 525624
rect 183639 525590 183673 525624
rect 183743 525590 183777 525624
rect 184743 525590 184777 525624
rect 184847 525590 184881 525624
rect 185847 525590 185881 525624
rect 185951 525590 185985 525624
rect 186951 525590 186985 525624
rect 187239 525590 187273 525624
rect 187239 525495 187273 525529
rect 187411 525590 187445 525624
rect 187411 525495 187445 525529
rect 172243 524749 172277 524783
rect 172243 524654 172277 524688
rect 172415 524749 172449 524783
rect 172415 524654 172449 524688
rect 172519 524654 172553 524688
rect 173519 524654 173553 524688
rect 173623 524654 173657 524688
rect 174623 524654 174657 524688
rect 174911 524654 174945 524688
rect 175911 524654 175945 524688
rect 176015 524654 176049 524688
rect 177015 524654 177049 524688
rect 177119 524654 177153 524688
rect 178119 524654 178153 524688
rect 178223 524654 178257 524688
rect 179223 524654 179257 524688
rect 179327 524756 179361 524790
rect 179327 524654 179361 524688
rect 179775 524756 179809 524790
rect 179775 524654 179809 524688
rect 180063 524654 180097 524688
rect 181063 524654 181097 524688
rect 181167 524654 181201 524688
rect 182167 524654 182201 524688
rect 182271 524654 182305 524688
rect 183271 524654 183305 524688
rect 183375 524654 183409 524688
rect 184375 524654 184409 524688
rect 184479 524756 184513 524790
rect 184479 524654 184513 524688
rect 184927 524756 184961 524790
rect 184927 524654 184961 524688
rect 185215 524654 185249 524688
rect 186215 524654 186249 524688
rect 186319 524756 186353 524790
rect 186319 524654 186353 524688
rect 186951 524756 186985 524790
rect 186951 524654 186985 524688
rect 187239 524749 187273 524783
rect 187239 524654 187273 524688
rect 187411 524749 187445 524783
rect 187411 524654 187445 524688
rect 172243 524502 172277 524536
rect 172243 524407 172277 524441
rect 172415 524502 172449 524536
rect 172415 524407 172449 524441
rect 172519 524502 172553 524536
rect 173519 524502 173553 524536
rect 173623 524502 173657 524536
rect 174623 524502 174657 524536
rect 174727 524502 174761 524536
rect 175727 524502 175761 524536
rect 175831 524502 175865 524536
rect 176831 524502 176865 524536
rect 176935 524502 176969 524536
rect 176935 524400 176969 524434
rect 177199 524502 177233 524536
rect 177199 524400 177233 524434
rect 177487 524502 177521 524536
rect 178487 524502 178521 524536
rect 178591 524502 178625 524536
rect 179591 524502 179625 524536
rect 179695 524502 179729 524536
rect 180695 524502 180729 524536
rect 180799 524502 180833 524536
rect 181799 524502 181833 524536
rect 181903 524502 181937 524536
rect 181903 524400 181937 524434
rect 182351 524502 182385 524536
rect 182351 524400 182385 524434
rect 182639 524502 182673 524536
rect 183639 524502 183673 524536
rect 183743 524502 183777 524536
rect 184743 524502 184777 524536
rect 184847 524502 184881 524536
rect 185847 524502 185881 524536
rect 185951 524502 185985 524536
rect 186951 524502 186985 524536
rect 187239 524502 187273 524536
rect 187239 524407 187273 524441
rect 187411 524502 187445 524536
rect 187411 524407 187445 524441
rect 172243 523661 172277 523695
rect 172243 523566 172277 523600
rect 172415 523661 172449 523695
rect 172415 523566 172449 523600
rect 172519 523566 172553 523600
rect 173519 523566 173553 523600
rect 173623 523566 173657 523600
rect 174623 523566 174657 523600
rect 174911 523566 174945 523600
rect 175911 523566 175945 523600
rect 176015 523566 176049 523600
rect 177015 523566 177049 523600
rect 177119 523566 177153 523600
rect 178119 523566 178153 523600
rect 178223 523566 178257 523600
rect 179223 523566 179257 523600
rect 179327 523668 179361 523702
rect 179327 523566 179361 523600
rect 179775 523668 179809 523702
rect 179775 523566 179809 523600
rect 180063 523566 180097 523600
rect 181063 523566 181097 523600
rect 181167 523566 181201 523600
rect 182167 523566 182201 523600
rect 182271 523566 182305 523600
rect 183271 523566 183305 523600
rect 183375 523566 183409 523600
rect 184375 523566 184409 523600
rect 184479 523668 184513 523702
rect 184479 523566 184513 523600
rect 184927 523668 184961 523702
rect 184927 523566 184961 523600
rect 185215 523566 185249 523600
rect 186215 523566 186249 523600
rect 186319 523668 186353 523702
rect 186319 523566 186353 523600
rect 186951 523668 186985 523702
rect 186951 523566 186985 523600
rect 187239 523661 187273 523695
rect 187239 523566 187273 523600
rect 187411 523661 187445 523695
rect 187411 523566 187445 523600
rect 172243 523414 172277 523448
rect 172243 523319 172277 523353
rect 172415 523414 172449 523448
rect 172415 523319 172449 523353
rect 172519 523414 172553 523448
rect 173519 523414 173553 523448
rect 173623 523414 173657 523448
rect 174623 523414 174657 523448
rect 174727 523414 174761 523448
rect 175727 523414 175761 523448
rect 175831 523414 175865 523448
rect 176831 523414 176865 523448
rect 176935 523414 176969 523448
rect 176935 523312 176969 523346
rect 177199 523414 177233 523448
rect 177199 523312 177233 523346
rect 177487 523414 177521 523448
rect 178487 523414 178521 523448
rect 178591 523414 178625 523448
rect 179591 523414 179625 523448
rect 179695 523414 179729 523448
rect 180695 523414 180729 523448
rect 180799 523414 180833 523448
rect 181799 523414 181833 523448
rect 181903 523414 181937 523448
rect 181903 523312 181937 523346
rect 182351 523414 182385 523448
rect 182351 523312 182385 523346
rect 182639 523414 182673 523448
rect 183639 523414 183673 523448
rect 183743 523414 183777 523448
rect 184743 523414 184777 523448
rect 184847 523414 184881 523448
rect 185847 523414 185881 523448
rect 185951 523414 185985 523448
rect 186951 523414 186985 523448
rect 187239 523414 187273 523448
rect 187239 523319 187273 523353
rect 187411 523414 187445 523448
rect 187411 523319 187445 523353
rect 172243 522573 172277 522607
rect 172243 522478 172277 522512
rect 172415 522573 172449 522607
rect 172415 522478 172449 522512
rect 172519 522478 172553 522512
rect 173519 522478 173553 522512
rect 173623 522478 173657 522512
rect 174623 522478 174657 522512
rect 174911 522478 174945 522512
rect 175911 522478 175945 522512
rect 176015 522478 176049 522512
rect 177015 522478 177049 522512
rect 177119 522478 177153 522512
rect 178119 522478 178153 522512
rect 178223 522478 178257 522512
rect 179223 522478 179257 522512
rect 179327 522580 179361 522614
rect 179327 522478 179361 522512
rect 179775 522580 179809 522614
rect 179775 522478 179809 522512
rect 180063 522478 180097 522512
rect 181063 522478 181097 522512
rect 181167 522478 181201 522512
rect 182167 522478 182201 522512
rect 182271 522478 182305 522512
rect 183271 522478 183305 522512
rect 183375 522478 183409 522512
rect 184375 522478 184409 522512
rect 184479 522580 184513 522614
rect 184479 522478 184513 522512
rect 184927 522580 184961 522614
rect 184927 522478 184961 522512
rect 185215 522478 185249 522512
rect 186215 522478 186249 522512
rect 186319 522580 186353 522614
rect 186319 522478 186353 522512
rect 186951 522580 186985 522614
rect 186951 522478 186985 522512
rect 187239 522573 187273 522607
rect 187239 522478 187273 522512
rect 187411 522573 187445 522607
rect 187411 522478 187445 522512
rect 172243 522326 172277 522360
rect 172243 522231 172277 522265
rect 172415 522326 172449 522360
rect 172415 522231 172449 522265
rect 172519 522326 172553 522360
rect 173519 522326 173553 522360
rect 173623 522326 173657 522360
rect 174623 522326 174657 522360
rect 174727 522326 174761 522360
rect 175727 522326 175761 522360
rect 175831 522326 175865 522360
rect 176831 522326 176865 522360
rect 176935 522326 176969 522360
rect 176935 522224 176969 522258
rect 177199 522326 177233 522360
rect 177199 522224 177233 522258
rect 177487 522326 177521 522360
rect 178487 522326 178521 522360
rect 178591 522326 178625 522360
rect 179591 522326 179625 522360
rect 179695 522326 179729 522360
rect 180695 522326 180729 522360
rect 180799 522326 180833 522360
rect 181799 522326 181833 522360
rect 181903 522326 181937 522360
rect 181903 522224 181937 522258
rect 182351 522326 182385 522360
rect 182351 522224 182385 522258
rect 182639 522326 182673 522360
rect 183639 522326 183673 522360
rect 183743 522326 183777 522360
rect 184743 522326 184777 522360
rect 184847 522326 184881 522360
rect 185847 522326 185881 522360
rect 185951 522326 185985 522360
rect 186951 522326 186985 522360
rect 187239 522326 187273 522360
rect 187239 522231 187273 522265
rect 187411 522326 187445 522360
rect 187411 522231 187445 522265
rect 172243 521485 172277 521519
rect 172243 521390 172277 521424
rect 172415 521485 172449 521519
rect 172415 521390 172449 521424
rect 172519 521390 172553 521424
rect 173519 521390 173553 521424
rect 173623 521390 173657 521424
rect 174623 521390 174657 521424
rect 174911 521390 174945 521424
rect 175911 521390 175945 521424
rect 176015 521390 176049 521424
rect 177015 521390 177049 521424
rect 177119 521390 177153 521424
rect 178119 521390 178153 521424
rect 178223 521390 178257 521424
rect 179223 521390 179257 521424
rect 179327 521492 179361 521526
rect 179327 521390 179361 521424
rect 179775 521492 179809 521526
rect 179775 521390 179809 521424
rect 180063 521390 180097 521424
rect 181063 521390 181097 521424
rect 181167 521390 181201 521424
rect 182167 521390 182201 521424
rect 182271 521390 182305 521424
rect 183271 521390 183305 521424
rect 183375 521390 183409 521424
rect 184375 521390 184409 521424
rect 184479 521492 184513 521526
rect 184479 521390 184513 521424
rect 184927 521492 184961 521526
rect 184927 521390 184961 521424
rect 185215 521390 185249 521424
rect 186215 521390 186249 521424
rect 186319 521492 186353 521526
rect 186319 521390 186353 521424
rect 186951 521492 186985 521526
rect 186951 521390 186985 521424
rect 187239 521485 187273 521519
rect 187239 521390 187273 521424
rect 187411 521485 187445 521519
rect 187411 521390 187445 521424
rect 172243 521238 172277 521272
rect 172243 521143 172277 521177
rect 172415 521238 172449 521272
rect 172415 521143 172449 521177
rect 172519 521238 172553 521272
rect 173519 521238 173553 521272
rect 173623 521238 173657 521272
rect 174623 521238 174657 521272
rect 174727 521238 174761 521272
rect 175727 521238 175761 521272
rect 175831 521238 175865 521272
rect 176831 521238 176865 521272
rect 176935 521238 176969 521272
rect 176935 521136 176969 521170
rect 177199 521238 177233 521272
rect 177199 521136 177233 521170
rect 177487 521238 177521 521272
rect 178487 521238 178521 521272
rect 178591 521238 178625 521272
rect 179591 521238 179625 521272
rect 179695 521238 179729 521272
rect 180695 521238 180729 521272
rect 180799 521238 180833 521272
rect 181799 521238 181833 521272
rect 181903 521238 181937 521272
rect 181903 521136 181937 521170
rect 182351 521238 182385 521272
rect 182351 521136 182385 521170
rect 182639 521238 182673 521272
rect 183639 521238 183673 521272
rect 183743 521238 183777 521272
rect 184743 521238 184777 521272
rect 184847 521238 184881 521272
rect 185847 521238 185881 521272
rect 185951 521238 185985 521272
rect 186951 521238 186985 521272
rect 187239 521238 187273 521272
rect 187239 521143 187273 521177
rect 187411 521238 187445 521272
rect 187411 521143 187445 521177
rect 172243 520397 172277 520431
rect 172243 520302 172277 520336
rect 172415 520397 172449 520431
rect 172415 520302 172449 520336
rect 172519 520302 172553 520336
rect 173519 520302 173553 520336
rect 173623 520302 173657 520336
rect 174623 520302 174657 520336
rect 174911 520302 174945 520336
rect 175911 520302 175945 520336
rect 176015 520302 176049 520336
rect 177015 520302 177049 520336
rect 177119 520302 177153 520336
rect 178119 520302 178153 520336
rect 178223 520302 178257 520336
rect 179223 520302 179257 520336
rect 179327 520404 179361 520438
rect 179327 520302 179361 520336
rect 179775 520404 179809 520438
rect 179775 520302 179809 520336
rect 180063 520302 180097 520336
rect 181063 520302 181097 520336
rect 181167 520302 181201 520336
rect 182167 520302 182201 520336
rect 182271 520302 182305 520336
rect 183271 520302 183305 520336
rect 183375 520302 183409 520336
rect 184375 520302 184409 520336
rect 184479 520404 184513 520438
rect 184479 520302 184513 520336
rect 184927 520404 184961 520438
rect 184927 520302 184961 520336
rect 185215 520302 185249 520336
rect 186215 520302 186249 520336
rect 186319 520404 186353 520438
rect 186319 520302 186353 520336
rect 186951 520404 186985 520438
rect 186951 520302 186985 520336
rect 187239 520397 187273 520431
rect 187239 520302 187273 520336
rect 187411 520397 187445 520431
rect 187411 520302 187445 520336
rect 172243 520150 172277 520184
rect 172243 520055 172277 520089
rect 172415 520150 172449 520184
rect 172415 520055 172449 520089
rect 172519 520150 172553 520184
rect 173519 520150 173553 520184
rect 173623 520150 173657 520184
rect 174623 520150 174657 520184
rect 174727 520150 174761 520184
rect 175727 520150 175761 520184
rect 175831 520150 175865 520184
rect 176831 520150 176865 520184
rect 176935 520150 176969 520184
rect 176935 520048 176969 520082
rect 177199 520150 177233 520184
rect 177199 520048 177233 520082
rect 177487 520150 177521 520184
rect 178487 520150 178521 520184
rect 178591 520150 178625 520184
rect 179591 520150 179625 520184
rect 179695 520150 179729 520184
rect 180695 520150 180729 520184
rect 180799 520150 180833 520184
rect 181799 520150 181833 520184
rect 181903 520150 181937 520184
rect 181903 520048 181937 520082
rect 182351 520150 182385 520184
rect 182351 520048 182385 520082
rect 182639 520150 182673 520184
rect 183639 520150 183673 520184
rect 183743 520150 183777 520184
rect 184743 520150 184777 520184
rect 184847 520150 184881 520184
rect 185847 520150 185881 520184
rect 185951 520150 185985 520184
rect 186951 520150 186985 520184
rect 187239 520150 187273 520184
rect 187239 520055 187273 520089
rect 187411 520150 187445 520184
rect 187411 520055 187445 520089
rect 172243 519309 172277 519343
rect 172243 519214 172277 519248
rect 172415 519309 172449 519343
rect 172415 519214 172449 519248
rect 172519 519214 172553 519248
rect 173519 519214 173553 519248
rect 173623 519214 173657 519248
rect 174623 519214 174657 519248
rect 174911 519214 174945 519248
rect 175911 519214 175945 519248
rect 176015 519214 176049 519248
rect 177015 519214 177049 519248
rect 177119 519214 177153 519248
rect 178119 519214 178153 519248
rect 178223 519214 178257 519248
rect 179223 519214 179257 519248
rect 179327 519316 179361 519350
rect 179327 519214 179361 519248
rect 179775 519316 179809 519350
rect 179775 519214 179809 519248
rect 180063 519214 180097 519248
rect 181063 519214 181097 519248
rect 181167 519214 181201 519248
rect 182167 519214 182201 519248
rect 182271 519214 182305 519248
rect 183271 519214 183305 519248
rect 183375 519214 183409 519248
rect 184375 519214 184409 519248
rect 184479 519316 184513 519350
rect 184479 519214 184513 519248
rect 184927 519316 184961 519350
rect 184927 519214 184961 519248
rect 185215 519214 185249 519248
rect 186215 519214 186249 519248
rect 186319 519316 186353 519350
rect 186319 519214 186353 519248
rect 186951 519316 186985 519350
rect 186951 519214 186985 519248
rect 187239 519309 187273 519343
rect 187239 519214 187273 519248
rect 187411 519309 187445 519343
rect 187411 519214 187445 519248
rect 172243 519062 172277 519096
rect 172243 518967 172277 519001
rect 172415 519062 172449 519096
rect 172415 518967 172449 519001
rect 172519 519062 172553 519096
rect 173519 519062 173553 519096
rect 173623 519062 173657 519096
rect 174623 519062 174657 519096
rect 174727 519062 174761 519096
rect 175727 519062 175761 519096
rect 175831 519062 175865 519096
rect 176831 519062 176865 519096
rect 176935 519062 176969 519096
rect 176935 518960 176969 518994
rect 177199 519062 177233 519096
rect 177199 518960 177233 518994
rect 177487 519062 177521 519096
rect 178487 519062 178521 519096
rect 178591 519062 178625 519096
rect 179591 519062 179625 519096
rect 179695 519062 179729 519096
rect 180695 519062 180729 519096
rect 180799 519062 180833 519096
rect 181799 519062 181833 519096
rect 181903 519062 181937 519096
rect 181903 518960 181937 518994
rect 182351 519062 182385 519096
rect 182351 518960 182385 518994
rect 182639 519062 182673 519096
rect 183639 519062 183673 519096
rect 183743 519062 183777 519096
rect 184743 519062 184777 519096
rect 184847 519062 184881 519096
rect 185847 519062 185881 519096
rect 185951 519062 185985 519096
rect 186951 519062 186985 519096
rect 187239 519062 187273 519096
rect 187239 518967 187273 519001
rect 187411 519062 187445 519096
rect 187411 518967 187445 519001
rect 172243 518221 172277 518255
rect 172243 518126 172277 518160
rect 172415 518221 172449 518255
rect 172415 518126 172449 518160
rect 172519 518126 172553 518160
rect 173519 518126 173553 518160
rect 173623 518126 173657 518160
rect 174623 518126 174657 518160
rect 174911 518126 174945 518160
rect 175911 518126 175945 518160
rect 176015 518126 176049 518160
rect 177015 518126 177049 518160
rect 177119 518126 177153 518160
rect 178119 518126 178153 518160
rect 178223 518126 178257 518160
rect 179223 518126 179257 518160
rect 179327 518228 179361 518262
rect 179327 518126 179361 518160
rect 179775 518228 179809 518262
rect 179775 518126 179809 518160
rect 180063 518126 180097 518160
rect 181063 518126 181097 518160
rect 181167 518126 181201 518160
rect 182167 518126 182201 518160
rect 182271 518126 182305 518160
rect 183271 518126 183305 518160
rect 183375 518126 183409 518160
rect 184375 518126 184409 518160
rect 184479 518228 184513 518262
rect 184479 518126 184513 518160
rect 184927 518228 184961 518262
rect 184927 518126 184961 518160
rect 185215 518126 185249 518160
rect 186215 518126 186249 518160
rect 186319 518228 186353 518262
rect 186319 518126 186353 518160
rect 186951 518228 186985 518262
rect 186951 518126 186985 518160
rect 187239 518221 187273 518255
rect 187239 518126 187273 518160
rect 187411 518221 187445 518255
rect 187411 518126 187445 518160
rect 172243 517974 172277 518008
rect 172243 517879 172277 517913
rect 172415 517974 172449 518008
rect 172415 517879 172449 517913
rect 172519 517974 172553 518008
rect 173519 517974 173553 518008
rect 173623 517974 173657 518008
rect 174623 517974 174657 518008
rect 174727 517974 174761 518008
rect 175727 517974 175761 518008
rect 175831 517974 175865 518008
rect 176831 517974 176865 518008
rect 176935 517974 176969 518008
rect 176935 517872 176969 517906
rect 177199 517974 177233 518008
rect 177199 517872 177233 517906
rect 177487 517974 177521 518008
rect 178487 517974 178521 518008
rect 178591 517974 178625 518008
rect 179591 517974 179625 518008
rect 179695 517974 179729 518008
rect 180695 517974 180729 518008
rect 180799 517974 180833 518008
rect 181799 517974 181833 518008
rect 181903 517974 181937 518008
rect 181903 517872 181937 517906
rect 182351 517974 182385 518008
rect 182351 517872 182385 517906
rect 182639 517974 182673 518008
rect 183639 517974 183673 518008
rect 183743 517974 183777 518008
rect 184743 517974 184777 518008
rect 184847 517974 184881 518008
rect 185847 517974 185881 518008
rect 185951 517974 185985 518008
rect 186951 517974 186985 518008
rect 187239 517974 187273 518008
rect 187239 517879 187273 517913
rect 187411 517974 187445 518008
rect 187411 517879 187445 517913
rect 172243 517133 172277 517167
rect 172243 517038 172277 517072
rect 172415 517133 172449 517167
rect 172415 517038 172449 517072
rect 172519 517038 172553 517072
rect 173519 517038 173553 517072
rect 173623 517038 173657 517072
rect 174623 517038 174657 517072
rect 174911 517038 174945 517072
rect 175911 517038 175945 517072
rect 176015 517038 176049 517072
rect 177015 517038 177049 517072
rect 177119 517038 177153 517072
rect 178119 517038 178153 517072
rect 178223 517038 178257 517072
rect 179223 517038 179257 517072
rect 179327 517140 179361 517174
rect 179327 517038 179361 517072
rect 179775 517140 179809 517174
rect 179775 517038 179809 517072
rect 180063 517038 180097 517072
rect 181063 517038 181097 517072
rect 181167 517038 181201 517072
rect 182167 517038 182201 517072
rect 182271 517038 182305 517072
rect 183271 517038 183305 517072
rect 183375 517038 183409 517072
rect 184375 517038 184409 517072
rect 184479 517140 184513 517174
rect 184479 517038 184513 517072
rect 184927 517140 184961 517174
rect 184927 517038 184961 517072
rect 185215 517038 185249 517072
rect 186215 517038 186249 517072
rect 186319 517140 186353 517174
rect 186319 517038 186353 517072
rect 186951 517140 186985 517174
rect 186951 517038 186985 517072
rect 187239 517133 187273 517167
rect 187239 517038 187273 517072
rect 187411 517133 187445 517167
rect 187411 517038 187445 517072
rect 172243 516886 172277 516920
rect 172243 516791 172277 516825
rect 172415 516886 172449 516920
rect 172415 516791 172449 516825
rect 172519 516886 172553 516920
rect 173519 516886 173553 516920
rect 173623 516886 173657 516920
rect 174623 516886 174657 516920
rect 174727 516886 174761 516920
rect 175727 516886 175761 516920
rect 175831 516886 175865 516920
rect 176831 516886 176865 516920
rect 176935 516886 176969 516920
rect 176935 516784 176969 516818
rect 177199 516886 177233 516920
rect 177199 516784 177233 516818
rect 177487 516886 177521 516920
rect 178487 516886 178521 516920
rect 178591 516886 178625 516920
rect 179591 516886 179625 516920
rect 179695 516886 179729 516920
rect 180695 516886 180729 516920
rect 180799 516886 180833 516920
rect 181799 516886 181833 516920
rect 181903 516886 181937 516920
rect 181903 516784 181937 516818
rect 182351 516886 182385 516920
rect 182351 516784 182385 516818
rect 182639 516886 182673 516920
rect 183639 516886 183673 516920
rect 183743 516886 183777 516920
rect 184743 516886 184777 516920
rect 184847 516886 184881 516920
rect 185847 516886 185881 516920
rect 185951 516886 185985 516920
rect 186951 516886 186985 516920
rect 187239 516886 187273 516920
rect 187239 516791 187273 516825
rect 187411 516886 187445 516920
rect 187411 516791 187445 516825
rect 172243 516045 172277 516079
rect 172243 515950 172277 515984
rect 172415 516045 172449 516079
rect 172415 515950 172449 515984
rect 172519 515950 172553 515984
rect 173519 515950 173553 515984
rect 173623 515950 173657 515984
rect 174623 515950 174657 515984
rect 174911 515950 174945 515984
rect 175911 515950 175945 515984
rect 176015 515950 176049 515984
rect 177015 515950 177049 515984
rect 177119 515950 177153 515984
rect 178119 515950 178153 515984
rect 178223 515950 178257 515984
rect 179223 515950 179257 515984
rect 179327 516052 179361 516086
rect 179327 515950 179361 515984
rect 179775 516052 179809 516086
rect 179775 515950 179809 515984
rect 180063 515950 180097 515984
rect 181063 515950 181097 515984
rect 181167 515950 181201 515984
rect 182167 515950 182201 515984
rect 182271 515950 182305 515984
rect 183271 515950 183305 515984
rect 183375 515950 183409 515984
rect 184375 515950 184409 515984
rect 184479 516052 184513 516086
rect 184479 515950 184513 515984
rect 184927 516052 184961 516086
rect 184927 515950 184961 515984
rect 185215 515950 185249 515984
rect 186215 515950 186249 515984
rect 186319 516052 186353 516086
rect 186319 515950 186353 515984
rect 186951 516052 186985 516086
rect 186951 515950 186985 515984
rect 187239 516045 187273 516079
rect 187239 515950 187273 515984
rect 187411 516045 187445 516079
rect 187411 515950 187445 515984
rect 172243 515798 172277 515832
rect 172243 515703 172277 515737
rect 172415 515798 172449 515832
rect 172415 515703 172449 515737
rect 172519 515798 172553 515832
rect 172519 515696 172553 515730
rect 173151 515798 173185 515832
rect 173151 515696 173185 515730
rect 173439 515790 173473 515824
rect 173439 515668 173473 515702
rect 173525 515798 173559 515832
rect 173525 515730 173559 515764
rect 173621 515763 173655 515797
rect 173707 515798 173741 515832
rect 173793 515790 173827 515824
rect 173793 515722 173827 515756
rect 173793 515654 173827 515688
rect 173879 515784 173913 515818
rect 173879 515716 173913 515750
rect 173991 515798 174025 515832
rect 173991 515696 174025 515730
rect 174623 515798 174657 515832
rect 174623 515696 174657 515730
rect 174911 515798 174945 515832
rect 175911 515798 175945 515832
rect 176015 515798 176049 515832
rect 177015 515798 177049 515832
rect 177119 515798 177153 515832
rect 177119 515703 177153 515737
rect 177291 515798 177325 515832
rect 177291 515703 177325 515737
rect 177487 515798 177521 515832
rect 178487 515798 178521 515832
rect 178591 515798 178625 515832
rect 179591 515798 179625 515832
rect 179695 515798 179729 515832
rect 179695 515703 179729 515737
rect 179867 515798 179901 515832
rect 179867 515703 179901 515737
rect 180063 515798 180097 515832
rect 181063 515798 181097 515832
rect 181167 515798 181201 515832
rect 181167 515696 181201 515730
rect 181799 515798 181833 515832
rect 181799 515696 181833 515730
rect 182087 515790 182121 515824
rect 182087 515709 182121 515743
rect 182173 515790 182207 515824
rect 182173 515722 182207 515756
rect 182259 515790 182293 515824
rect 182259 515722 182293 515756
rect 182639 515798 182673 515832
rect 183639 515798 183673 515832
rect 183743 515798 183777 515832
rect 184743 515798 184777 515832
rect 184847 515798 184881 515832
rect 184847 515703 184881 515737
rect 185019 515798 185053 515832
rect 185019 515703 185053 515737
rect 185215 515798 185249 515832
rect 186215 515798 186249 515832
rect 186411 515790 186445 515824
rect 186411 515668 186445 515702
rect 186497 515798 186531 515832
rect 186497 515730 186531 515764
rect 186593 515763 186627 515797
rect 186679 515798 186713 515832
rect 186765 515790 186799 515824
rect 186765 515722 186799 515756
rect 186765 515654 186799 515688
rect 186851 515784 186885 515818
rect 186851 515716 186885 515750
rect 186963 515798 186997 515832
rect 186963 515703 186997 515737
rect 187135 515798 187169 515832
rect 187135 515703 187169 515737
rect 187239 515798 187273 515832
rect 187239 515703 187273 515737
rect 187411 515798 187445 515832
rect 187411 515703 187445 515737
<< psubdiff >>
rect 164518 541255 166648 541275
rect 164518 541245 164618 541255
rect 164518 539865 164538 541245
rect 164578 541215 164618 541245
rect 166538 541235 166648 541255
rect 166538 541215 166578 541235
rect 164578 541185 166578 541215
rect 164578 539915 164598 541185
rect 166558 539915 166578 541185
rect 164578 539895 166578 539915
rect 164578 539865 164618 539895
rect 164518 539855 164618 539865
rect 166538 539855 166578 539895
rect 166618 539855 166648 541235
rect 164518 539825 166648 539855
rect 168318 541255 170448 541275
rect 168318 541245 168418 541255
rect 168318 539865 168338 541245
rect 168378 541215 168418 541245
rect 170338 541235 170448 541255
rect 170338 541215 170378 541235
rect 168378 541185 170378 541215
rect 168378 539915 168398 541185
rect 170358 539915 170378 541185
rect 168378 539895 170378 539915
rect 168378 539865 168418 539895
rect 168318 539855 168418 539865
rect 170338 539855 170378 539895
rect 170418 539855 170448 541235
rect 168318 539825 170448 539855
rect 172018 541255 174148 541275
rect 172018 541245 172118 541255
rect 172018 539865 172038 541245
rect 172078 541215 172118 541245
rect 174038 541235 174148 541255
rect 174038 541215 174078 541235
rect 172078 541185 174078 541215
rect 172078 539915 172098 541185
rect 174058 539915 174078 541185
rect 172078 539895 174078 539915
rect 172078 539865 172118 539895
rect 172018 539855 172118 539865
rect 174038 539855 174078 539895
rect 174118 539855 174148 541235
rect 172018 539825 174148 539855
rect 175518 541255 177648 541275
rect 175518 541245 175618 541255
rect 175518 539865 175538 541245
rect 175578 541215 175618 541245
rect 177538 541235 177648 541255
rect 177538 541215 177578 541235
rect 175578 541185 177578 541215
rect 175578 539915 175598 541185
rect 177558 539915 177578 541185
rect 175578 539895 177578 539915
rect 175578 539865 175618 539895
rect 175518 539855 175618 539865
rect 177538 539855 177578 539895
rect 177618 539855 177648 541235
rect 175518 539825 177648 539855
rect 179118 541255 181248 541275
rect 179118 541245 179218 541255
rect 179118 539865 179138 541245
rect 179178 541215 179218 541245
rect 181138 541235 181248 541255
rect 181138 541215 181178 541235
rect 179178 541185 181178 541215
rect 179178 539915 179198 541185
rect 181158 539915 181178 541185
rect 179178 539895 181178 539915
rect 179178 539865 179218 539895
rect 179118 539855 179218 539865
rect 181138 539855 181178 539895
rect 181218 539855 181248 541235
rect 179118 539825 181248 539855
rect 182418 541255 184548 541275
rect 182418 541245 182518 541255
rect 182418 539865 182438 541245
rect 182478 541215 182518 541245
rect 184438 541235 184548 541255
rect 184438 541215 184478 541235
rect 182478 541185 184478 541215
rect 182478 539915 182498 541185
rect 184458 539915 184478 541185
rect 182478 539895 184478 539915
rect 182478 539865 182518 539895
rect 182418 539855 182518 539865
rect 184438 539855 184478 539895
rect 184518 539855 184548 541235
rect 182418 539825 184548 539855
rect 185718 541255 187848 541275
rect 185718 541245 185818 541255
rect 185718 539865 185738 541245
rect 185778 541215 185818 541245
rect 187738 541235 187848 541255
rect 187738 541215 187778 541235
rect 185778 541185 187778 541215
rect 185778 539915 185798 541185
rect 187758 539915 187778 541185
rect 185778 539895 187778 539915
rect 185778 539865 185818 539895
rect 185718 539855 185818 539865
rect 187738 539855 187778 539895
rect 187818 539855 187848 541235
rect 185718 539825 187848 539855
rect 189018 541255 191148 541275
rect 189018 541245 189118 541255
rect 189018 539865 189038 541245
rect 189078 541215 189118 541245
rect 191038 541235 191148 541255
rect 191038 541215 191078 541235
rect 189078 541185 191078 541215
rect 189078 539915 189098 541185
rect 191058 539915 191078 541185
rect 189078 539895 191078 539915
rect 189078 539865 189118 539895
rect 189018 539855 189118 539865
rect 191038 539855 191078 539895
rect 191118 539855 191148 541235
rect 191808 540245 191988 540269
rect 191808 540041 191988 540065
rect 189018 539825 191148 539855
rect 157628 538705 162868 538725
rect 157628 538665 157708 538705
rect 162768 538665 162868 538705
rect 157628 538645 162868 538665
rect 157628 538625 157708 538645
rect 157628 537965 157648 538625
rect 157688 538005 157708 538625
rect 162788 538005 162808 538645
rect 162848 538005 162868 538645
rect 157688 537985 162868 538005
rect 157688 537965 157728 537985
rect 157628 537945 157728 537965
rect 162768 537945 162868 537985
rect 157628 537925 162868 537945
rect 164186 538045 164282 538079
rect 166646 538045 166742 538079
rect 164186 537983 164220 538045
rect 166708 537983 166742 538045
rect 164186 535905 164220 535967
rect 166708 535905 166742 535967
rect 164186 535871 164282 535905
rect 166646 535871 166742 535905
rect 167958 538045 168054 538079
rect 169146 538045 169242 538079
rect 167958 537983 167992 538045
rect 169208 537983 169242 538045
rect 167958 535905 167992 535967
rect 169208 535905 169242 535967
rect 167958 535871 168054 535905
rect 169146 535871 169242 535905
rect 171694 538045 171790 538079
rect 172246 538045 172342 538079
rect 171694 537983 171728 538045
rect 172308 537983 172342 538045
rect 171694 535905 171728 535967
rect 172308 535905 172342 535967
rect 171694 535871 171790 535905
rect 172246 535871 172342 535905
rect 175212 538045 175308 538079
rect 175446 538045 175542 538079
rect 175212 537983 175246 538045
rect 175508 537983 175542 538045
rect 175212 535905 175246 535967
rect 178812 538045 178908 538079
rect 179046 538045 179142 538079
rect 178812 537983 178846 538045
rect 179108 537983 179142 538045
rect 178812 536465 178846 536527
rect 182112 538045 182208 538079
rect 182346 538045 182442 538079
rect 182112 537983 182146 538045
rect 182408 537983 182442 538045
rect 182112 536745 182146 536807
rect 185412 538045 185508 538079
rect 185646 538045 185742 538079
rect 185412 537983 185446 538045
rect 185708 537983 185742 538045
rect 185412 536885 185446 536947
rect 185708 536885 185742 536947
rect 185412 536851 185508 536885
rect 185646 536851 185742 536885
rect 188712 538045 188808 538079
rect 188946 538045 189042 538079
rect 188712 537983 188746 538045
rect 189008 537983 189042 538045
rect 182408 536745 182442 536807
rect 188712 536789 188746 536851
rect 189008 536789 189042 536851
rect 188712 536755 188808 536789
rect 188946 536755 189042 536789
rect 182112 536711 182208 536745
rect 182346 536711 182442 536745
rect 179108 536465 179142 536527
rect 178812 536431 178908 536465
rect 179046 536431 179142 536465
rect 175508 535905 175542 535967
rect 175212 535871 175308 535905
rect 175446 535871 175542 535905
rect 164156 535705 164252 535739
rect 166616 535705 166712 535739
rect 164156 535643 164190 535705
rect 166678 535643 166712 535705
rect 164156 533565 164190 533627
rect 166678 533565 166712 533627
rect 164156 533531 164252 533565
rect 166616 533531 166712 533565
rect 174813 530468 174847 530515
rect 174813 530410 174847 530434
rect 177389 530468 177423 530515
rect 177389 530410 177423 530434
rect 179965 530468 179999 530515
rect 179965 530410 179999 530434
rect 182541 530468 182575 530515
rect 182541 530410 182575 530434
rect 185117 530468 185151 530515
rect 185117 530410 185151 530434
rect 177389 529636 177423 529660
rect 177389 529555 177423 529602
rect 182541 529636 182575 529660
rect 182541 529555 182575 529602
rect 174813 529380 174847 529427
rect 174813 529322 174847 529346
rect 179965 529380 179999 529427
rect 179965 529322 179999 529346
rect 185117 529380 185151 529427
rect 185117 529322 185151 529346
rect 177389 528548 177423 528572
rect 177389 528467 177423 528514
rect 182541 528548 182575 528572
rect 182541 528467 182575 528514
rect 174813 528292 174847 528339
rect 174813 528234 174847 528258
rect 179965 528292 179999 528339
rect 179965 528234 179999 528258
rect 185117 528292 185151 528339
rect 185117 528234 185151 528258
rect 177389 527460 177423 527484
rect 177389 527379 177423 527426
rect 182541 527460 182575 527484
rect 182541 527379 182575 527426
rect 174813 527204 174847 527251
rect 174813 527146 174847 527170
rect 179965 527204 179999 527251
rect 179965 527146 179999 527170
rect 185117 527204 185151 527251
rect 185117 527146 185151 527170
rect 177389 526372 177423 526396
rect 177389 526291 177423 526338
rect 182541 526372 182575 526396
rect 182541 526291 182575 526338
rect 174813 526116 174847 526163
rect 174813 526058 174847 526082
rect 179965 526116 179999 526163
rect 179965 526058 179999 526082
rect 185117 526116 185151 526163
rect 185117 526058 185151 526082
rect 177389 525284 177423 525308
rect 177389 525203 177423 525250
rect 182541 525284 182575 525308
rect 182541 525203 182575 525250
rect 174813 525028 174847 525075
rect 174813 524970 174847 524994
rect 179965 525028 179999 525075
rect 179965 524970 179999 524994
rect 185117 525028 185151 525075
rect 185117 524970 185151 524994
rect 177389 524196 177423 524220
rect 177389 524115 177423 524162
rect 182541 524196 182575 524220
rect 182541 524115 182575 524162
rect 174813 523940 174847 523987
rect 174813 523882 174847 523906
rect 179965 523940 179999 523987
rect 179965 523882 179999 523906
rect 185117 523940 185151 523987
rect 185117 523882 185151 523906
rect 177389 523108 177423 523132
rect 177389 523027 177423 523074
rect 182541 523108 182575 523132
rect 182541 523027 182575 523074
rect 174813 522852 174847 522899
rect 174813 522794 174847 522818
rect 179965 522852 179999 522899
rect 179965 522794 179999 522818
rect 185117 522852 185151 522899
rect 185117 522794 185151 522818
rect 177389 522020 177423 522044
rect 177389 521939 177423 521986
rect 182541 522020 182575 522044
rect 182541 521939 182575 521986
rect 174813 521764 174847 521811
rect 174813 521706 174847 521730
rect 179965 521764 179999 521811
rect 179965 521706 179999 521730
rect 185117 521764 185151 521811
rect 185117 521706 185151 521730
rect 177389 520932 177423 520956
rect 177389 520851 177423 520898
rect 182541 520932 182575 520956
rect 182541 520851 182575 520898
rect 174813 520676 174847 520723
rect 174813 520618 174847 520642
rect 179965 520676 179999 520723
rect 179965 520618 179999 520642
rect 185117 520676 185151 520723
rect 185117 520618 185151 520642
rect 177389 519844 177423 519868
rect 177389 519763 177423 519810
rect 182541 519844 182575 519868
rect 182541 519763 182575 519810
rect 174813 519588 174847 519635
rect 174813 519530 174847 519554
rect 179965 519588 179999 519635
rect 179965 519530 179999 519554
rect 185117 519588 185151 519635
rect 185117 519530 185151 519554
rect 177389 518756 177423 518780
rect 177389 518675 177423 518722
rect 182541 518756 182575 518780
rect 182541 518675 182575 518722
rect 174813 518500 174847 518547
rect 174813 518442 174847 518466
rect 179965 518500 179999 518547
rect 179965 518442 179999 518466
rect 185117 518500 185151 518547
rect 185117 518442 185151 518466
rect 177389 517668 177423 517692
rect 177389 517587 177423 517634
rect 182541 517668 182575 517692
rect 182541 517587 182575 517634
rect 174813 517412 174847 517459
rect 174813 517354 174847 517378
rect 179965 517412 179999 517459
rect 179965 517354 179999 517378
rect 185117 517412 185151 517459
rect 185117 517354 185151 517378
rect 177389 516580 177423 516604
rect 177389 516499 177423 516546
rect 182541 516580 182575 516604
rect 182541 516499 182575 516546
rect 174813 516324 174847 516371
rect 174813 516266 174847 516290
rect 179965 516324 179999 516371
rect 179965 516266 179999 516290
rect 185117 516324 185151 516371
rect 185117 516266 185151 516290
rect 174813 515492 174847 515516
rect 174813 515411 174847 515458
rect 177389 515492 177423 515516
rect 177389 515411 177423 515458
rect 179965 515492 179999 515516
rect 179965 515411 179999 515458
rect 182541 515492 182575 515516
rect 182541 515411 182575 515458
rect 185117 515492 185151 515516
rect 185117 515411 185151 515458
<< nsubdiff >>
rect 164518 539735 166638 539755
rect 164518 539715 164618 539735
rect 164518 538315 164538 539715
rect 164578 539695 164618 539715
rect 166538 539715 166638 539735
rect 166538 539695 166578 539715
rect 164578 539675 166578 539695
rect 164578 538355 164598 539675
rect 166538 539655 166578 539675
rect 166558 538355 166578 539655
rect 164578 538335 166578 538355
rect 164578 538315 164618 538335
rect 164518 538295 164618 538315
rect 166538 538315 166578 538335
rect 166618 538315 166638 539715
rect 166538 538295 166638 538315
rect 164518 538275 166638 538295
rect 168318 539735 170438 539755
rect 168318 539715 168418 539735
rect 168318 538315 168338 539715
rect 168378 539695 168418 539715
rect 170338 539715 170438 539735
rect 170338 539695 170378 539715
rect 168378 539675 170378 539695
rect 168378 538355 168398 539675
rect 170338 539655 170378 539675
rect 170358 538355 170378 539655
rect 168378 538335 170378 538355
rect 168378 538315 168418 538335
rect 168318 538295 168418 538315
rect 170338 538315 170378 538335
rect 170418 538315 170438 539715
rect 170338 538295 170438 538315
rect 168318 538275 170438 538295
rect 172018 539735 174138 539755
rect 172018 539715 172118 539735
rect 172018 538315 172038 539715
rect 172078 539695 172118 539715
rect 174038 539715 174138 539735
rect 174038 539695 174078 539715
rect 172078 539675 174078 539695
rect 172078 538355 172098 539675
rect 174038 539655 174078 539675
rect 174058 538355 174078 539655
rect 172078 538335 174078 538355
rect 172078 538315 172118 538335
rect 172018 538295 172118 538315
rect 174038 538315 174078 538335
rect 174118 538315 174138 539715
rect 174038 538295 174138 538315
rect 172018 538275 174138 538295
rect 175518 539735 177638 539755
rect 175518 539715 175618 539735
rect 175518 538315 175538 539715
rect 175578 539695 175618 539715
rect 177538 539715 177638 539735
rect 177538 539695 177578 539715
rect 175578 539675 177578 539695
rect 175578 538355 175598 539675
rect 177538 539655 177578 539675
rect 177558 538355 177578 539655
rect 175578 538335 177578 538355
rect 175578 538315 175618 538335
rect 175518 538295 175618 538315
rect 177538 538315 177578 538335
rect 177618 538315 177638 539715
rect 177538 538295 177638 538315
rect 175518 538275 177638 538295
rect 179118 539735 181238 539755
rect 179118 539715 179218 539735
rect 179118 538315 179138 539715
rect 179178 539695 179218 539715
rect 181138 539715 181238 539735
rect 181138 539695 181178 539715
rect 179178 539675 181178 539695
rect 179178 538355 179198 539675
rect 181138 539655 181178 539675
rect 181158 538355 181178 539655
rect 179178 538335 181178 538355
rect 179178 538315 179218 538335
rect 179118 538295 179218 538315
rect 181138 538315 181178 538335
rect 181218 538315 181238 539715
rect 181138 538295 181238 538315
rect 179118 538275 181238 538295
rect 182418 539735 184538 539755
rect 182418 539715 182518 539735
rect 182418 538315 182438 539715
rect 182478 539695 182518 539715
rect 184438 539715 184538 539735
rect 184438 539695 184478 539715
rect 182478 539675 184478 539695
rect 182478 538355 182498 539675
rect 184438 539655 184478 539675
rect 184458 538355 184478 539655
rect 182478 538335 184478 538355
rect 182478 538315 182518 538335
rect 182418 538295 182518 538315
rect 184438 538315 184478 538335
rect 184518 538315 184538 539715
rect 184438 538295 184538 538315
rect 182418 538275 184538 538295
rect 185718 539735 187838 539755
rect 185718 539715 185818 539735
rect 185718 538315 185738 539715
rect 185778 539695 185818 539715
rect 187738 539715 187838 539735
rect 187738 539695 187778 539715
rect 185778 539675 187778 539695
rect 185778 538355 185798 539675
rect 187738 539655 187778 539675
rect 187758 538355 187778 539655
rect 185778 538335 187778 538355
rect 185778 538315 185818 538335
rect 185718 538295 185818 538315
rect 187738 538315 187778 538335
rect 187818 538315 187838 539715
rect 187738 538295 187838 538315
rect 185718 538275 187838 538295
rect 189018 539735 191138 539755
rect 189018 539715 189118 539735
rect 189018 538315 189038 539715
rect 189078 539695 189118 539715
rect 191038 539715 191138 539735
rect 191038 539695 191078 539715
rect 189078 539675 191078 539695
rect 189078 538355 189098 539675
rect 191038 539655 191078 539675
rect 191058 538355 191078 539655
rect 189078 538335 191078 538355
rect 189078 538315 189118 538335
rect 189018 538295 189118 538315
rect 191038 538315 191078 538335
rect 191118 538315 191138 539715
rect 191038 538295 191138 538315
rect 189018 538275 191138 538295
rect 157588 537825 162848 537845
rect 157588 537785 157648 537825
rect 162748 537785 162848 537825
rect 157588 537765 162788 537785
rect 157588 537725 157668 537765
rect 157588 535785 157608 537725
rect 157648 535785 157668 537725
rect 157588 535765 157668 535785
rect 162768 535765 162788 537765
rect 162828 535765 162848 537785
rect 157588 535745 162848 535765
rect 157588 535705 157668 535745
rect 162748 535705 162848 535745
rect 157588 535685 162848 535705
rect 174813 530250 174847 530274
rect 174813 530157 174847 530216
rect 174813 530099 174847 530123
rect 177389 530250 177423 530274
rect 177389 530157 177423 530216
rect 177389 530099 177423 530123
rect 179965 530250 179999 530274
rect 179965 530157 179999 530216
rect 179965 530099 179999 530123
rect 182541 530250 182575 530274
rect 182541 530157 182575 530216
rect 182541 530099 182575 530123
rect 185117 530250 185151 530274
rect 185117 530157 185151 530216
rect 185117 530099 185151 530123
rect 177389 529947 177423 529971
rect 177389 529854 177423 529913
rect 177389 529796 177423 529820
rect 182541 529947 182575 529971
rect 182541 529854 182575 529913
rect 182541 529796 182575 529820
rect 174813 529162 174847 529186
rect 174813 529069 174847 529128
rect 174813 529011 174847 529035
rect 179965 529162 179999 529186
rect 179965 529069 179999 529128
rect 179965 529011 179999 529035
rect 185117 529162 185151 529186
rect 185117 529069 185151 529128
rect 185117 529011 185151 529035
rect 177389 528859 177423 528883
rect 177389 528766 177423 528825
rect 177389 528708 177423 528732
rect 182541 528859 182575 528883
rect 182541 528766 182575 528825
rect 182541 528708 182575 528732
rect 174813 528074 174847 528098
rect 174813 527981 174847 528040
rect 174813 527923 174847 527947
rect 179965 528074 179999 528098
rect 179965 527981 179999 528040
rect 179965 527923 179999 527947
rect 185117 528074 185151 528098
rect 185117 527981 185151 528040
rect 185117 527923 185151 527947
rect 177389 527771 177423 527795
rect 177389 527678 177423 527737
rect 177389 527620 177423 527644
rect 182541 527771 182575 527795
rect 182541 527678 182575 527737
rect 182541 527620 182575 527644
rect 174813 526986 174847 527010
rect 174813 526893 174847 526952
rect 174813 526835 174847 526859
rect 179965 526986 179999 527010
rect 179965 526893 179999 526952
rect 179965 526835 179999 526859
rect 185117 526986 185151 527010
rect 185117 526893 185151 526952
rect 185117 526835 185151 526859
rect 177389 526683 177423 526707
rect 177389 526590 177423 526649
rect 177389 526532 177423 526556
rect 182541 526683 182575 526707
rect 182541 526590 182575 526649
rect 182541 526532 182575 526556
rect 174813 525898 174847 525922
rect 174813 525805 174847 525864
rect 174813 525747 174847 525771
rect 179965 525898 179999 525922
rect 179965 525805 179999 525864
rect 179965 525747 179999 525771
rect 185117 525898 185151 525922
rect 185117 525805 185151 525864
rect 185117 525747 185151 525771
rect 177389 525595 177423 525619
rect 177389 525502 177423 525561
rect 177389 525444 177423 525468
rect 182541 525595 182575 525619
rect 182541 525502 182575 525561
rect 182541 525444 182575 525468
rect 174813 524810 174847 524834
rect 174813 524717 174847 524776
rect 174813 524659 174847 524683
rect 179965 524810 179999 524834
rect 179965 524717 179999 524776
rect 179965 524659 179999 524683
rect 185117 524810 185151 524834
rect 185117 524717 185151 524776
rect 185117 524659 185151 524683
rect 177389 524507 177423 524531
rect 177389 524414 177423 524473
rect 177389 524356 177423 524380
rect 182541 524507 182575 524531
rect 182541 524414 182575 524473
rect 182541 524356 182575 524380
rect 174813 523722 174847 523746
rect 174813 523629 174847 523688
rect 174813 523571 174847 523595
rect 179965 523722 179999 523746
rect 179965 523629 179999 523688
rect 179965 523571 179999 523595
rect 185117 523722 185151 523746
rect 185117 523629 185151 523688
rect 185117 523571 185151 523595
rect 177389 523419 177423 523443
rect 177389 523326 177423 523385
rect 177389 523268 177423 523292
rect 182541 523419 182575 523443
rect 182541 523326 182575 523385
rect 182541 523268 182575 523292
rect 174813 522634 174847 522658
rect 174813 522541 174847 522600
rect 174813 522483 174847 522507
rect 179965 522634 179999 522658
rect 179965 522541 179999 522600
rect 179965 522483 179999 522507
rect 185117 522634 185151 522658
rect 185117 522541 185151 522600
rect 185117 522483 185151 522507
rect 177389 522331 177423 522355
rect 177389 522238 177423 522297
rect 177389 522180 177423 522204
rect 182541 522331 182575 522355
rect 182541 522238 182575 522297
rect 182541 522180 182575 522204
rect 174813 521546 174847 521570
rect 174813 521453 174847 521512
rect 174813 521395 174847 521419
rect 179965 521546 179999 521570
rect 179965 521453 179999 521512
rect 179965 521395 179999 521419
rect 185117 521546 185151 521570
rect 185117 521453 185151 521512
rect 185117 521395 185151 521419
rect 177389 521243 177423 521267
rect 177389 521150 177423 521209
rect 177389 521092 177423 521116
rect 182541 521243 182575 521267
rect 182541 521150 182575 521209
rect 182541 521092 182575 521116
rect 174813 520458 174847 520482
rect 174813 520365 174847 520424
rect 174813 520307 174847 520331
rect 179965 520458 179999 520482
rect 179965 520365 179999 520424
rect 179965 520307 179999 520331
rect 185117 520458 185151 520482
rect 185117 520365 185151 520424
rect 185117 520307 185151 520331
rect 177389 520155 177423 520179
rect 177389 520062 177423 520121
rect 177389 520004 177423 520028
rect 182541 520155 182575 520179
rect 182541 520062 182575 520121
rect 182541 520004 182575 520028
rect 174813 519370 174847 519394
rect 174813 519277 174847 519336
rect 174813 519219 174847 519243
rect 179965 519370 179999 519394
rect 179965 519277 179999 519336
rect 179965 519219 179999 519243
rect 185117 519370 185151 519394
rect 185117 519277 185151 519336
rect 185117 519219 185151 519243
rect 177389 519067 177423 519091
rect 177389 518974 177423 519033
rect 177389 518916 177423 518940
rect 182541 519067 182575 519091
rect 182541 518974 182575 519033
rect 182541 518916 182575 518940
rect 174813 518282 174847 518306
rect 174813 518189 174847 518248
rect 174813 518131 174847 518155
rect 179965 518282 179999 518306
rect 179965 518189 179999 518248
rect 179965 518131 179999 518155
rect 185117 518282 185151 518306
rect 185117 518189 185151 518248
rect 185117 518131 185151 518155
rect 177389 517979 177423 518003
rect 177389 517886 177423 517945
rect 177389 517828 177423 517852
rect 182541 517979 182575 518003
rect 182541 517886 182575 517945
rect 182541 517828 182575 517852
rect 174813 517194 174847 517218
rect 174813 517101 174847 517160
rect 174813 517043 174847 517067
rect 179965 517194 179999 517218
rect 179965 517101 179999 517160
rect 179965 517043 179999 517067
rect 185117 517194 185151 517218
rect 185117 517101 185151 517160
rect 185117 517043 185151 517067
rect 177389 516891 177423 516915
rect 177389 516798 177423 516857
rect 177389 516740 177423 516764
rect 182541 516891 182575 516915
rect 182541 516798 182575 516857
rect 182541 516740 182575 516764
rect 174813 516106 174847 516130
rect 174813 516013 174847 516072
rect 174813 515955 174847 515979
rect 179965 516106 179999 516130
rect 179965 516013 179999 516072
rect 179965 515955 179999 515979
rect 185117 516106 185151 516130
rect 185117 516013 185151 516072
rect 185117 515955 185151 515979
rect 174813 515803 174847 515827
rect 174813 515710 174847 515769
rect 174813 515652 174847 515676
rect 177389 515803 177423 515827
rect 177389 515710 177423 515769
rect 177389 515652 177423 515676
rect 179965 515803 179999 515827
rect 179965 515710 179999 515769
rect 179965 515652 179999 515676
rect 182541 515803 182575 515827
rect 182541 515710 182575 515769
rect 182541 515652 182575 515676
rect 185117 515803 185151 515827
rect 185117 515710 185151 515769
rect 185117 515652 185151 515676
<< psubdiffcont >>
rect 164538 539865 164578 541245
rect 164618 541215 166538 541255
rect 164618 539855 166538 539895
rect 166578 539855 166618 541235
rect 168338 539865 168378 541245
rect 168418 541215 170338 541255
rect 168418 539855 170338 539895
rect 170378 539855 170418 541235
rect 172038 539865 172078 541245
rect 172118 541215 174038 541255
rect 172118 539855 174038 539895
rect 174078 539855 174118 541235
rect 175538 539865 175578 541245
rect 175618 541215 177538 541255
rect 175618 539855 177538 539895
rect 177578 539855 177618 541235
rect 179138 539865 179178 541245
rect 179218 541215 181138 541255
rect 179218 539855 181138 539895
rect 181178 539855 181218 541235
rect 182438 539865 182478 541245
rect 182518 541215 184438 541255
rect 182518 539855 184438 539895
rect 184478 539855 184518 541235
rect 185738 539865 185778 541245
rect 185818 541215 187738 541255
rect 185818 539855 187738 539895
rect 187778 539855 187818 541235
rect 189038 539865 189078 541245
rect 189118 541215 191038 541255
rect 189118 539855 191038 539895
rect 191078 539855 191118 541235
rect 191808 540065 191988 540245
rect 157708 538665 162768 538705
rect 157648 537965 157688 538625
rect 162808 538005 162848 538645
rect 157728 537945 162768 537985
rect 164282 538045 166646 538079
rect 164186 535967 164220 537983
rect 166708 535967 166742 537983
rect 164282 535871 166646 535905
rect 168054 538045 169146 538079
rect 167958 535967 167992 537983
rect 169208 535967 169242 537983
rect 168054 535871 169146 535905
rect 171790 538045 172246 538079
rect 171694 535967 171728 537983
rect 172308 535967 172342 537983
rect 171790 535871 172246 535905
rect 175308 538045 175446 538079
rect 175212 535967 175246 537983
rect 175508 535967 175542 537983
rect 178908 538045 179046 538079
rect 178812 536527 178846 537983
rect 179108 536527 179142 537983
rect 182208 538045 182346 538079
rect 182112 536807 182146 537983
rect 182408 536807 182442 537983
rect 185508 538045 185646 538079
rect 185412 536947 185446 537983
rect 185708 536947 185742 537983
rect 185508 536851 185646 536885
rect 188808 538045 188946 538079
rect 188712 536851 188746 537983
rect 189008 536851 189042 537983
rect 188808 536755 188946 536789
rect 182208 536711 182346 536745
rect 178908 536431 179046 536465
rect 175308 535871 175446 535905
rect 164252 535705 166616 535739
rect 164156 533627 164190 535643
rect 166678 533627 166712 535643
rect 164252 533531 166616 533565
rect 174813 530434 174847 530468
rect 177389 530434 177423 530468
rect 179965 530434 179999 530468
rect 182541 530434 182575 530468
rect 185117 530434 185151 530468
rect 177389 529602 177423 529636
rect 182541 529602 182575 529636
rect 174813 529346 174847 529380
rect 179965 529346 179999 529380
rect 185117 529346 185151 529380
rect 177389 528514 177423 528548
rect 182541 528514 182575 528548
rect 174813 528258 174847 528292
rect 179965 528258 179999 528292
rect 185117 528258 185151 528292
rect 177389 527426 177423 527460
rect 182541 527426 182575 527460
rect 174813 527170 174847 527204
rect 179965 527170 179999 527204
rect 185117 527170 185151 527204
rect 177389 526338 177423 526372
rect 182541 526338 182575 526372
rect 174813 526082 174847 526116
rect 179965 526082 179999 526116
rect 185117 526082 185151 526116
rect 177389 525250 177423 525284
rect 182541 525250 182575 525284
rect 174813 524994 174847 525028
rect 179965 524994 179999 525028
rect 185117 524994 185151 525028
rect 177389 524162 177423 524196
rect 182541 524162 182575 524196
rect 174813 523906 174847 523940
rect 179965 523906 179999 523940
rect 185117 523906 185151 523940
rect 177389 523074 177423 523108
rect 182541 523074 182575 523108
rect 174813 522818 174847 522852
rect 179965 522818 179999 522852
rect 185117 522818 185151 522852
rect 177389 521986 177423 522020
rect 182541 521986 182575 522020
rect 174813 521730 174847 521764
rect 179965 521730 179999 521764
rect 185117 521730 185151 521764
rect 177389 520898 177423 520932
rect 182541 520898 182575 520932
rect 174813 520642 174847 520676
rect 179965 520642 179999 520676
rect 185117 520642 185151 520676
rect 177389 519810 177423 519844
rect 182541 519810 182575 519844
rect 174813 519554 174847 519588
rect 179965 519554 179999 519588
rect 185117 519554 185151 519588
rect 177389 518722 177423 518756
rect 182541 518722 182575 518756
rect 174813 518466 174847 518500
rect 179965 518466 179999 518500
rect 185117 518466 185151 518500
rect 177389 517634 177423 517668
rect 182541 517634 182575 517668
rect 174813 517378 174847 517412
rect 179965 517378 179999 517412
rect 185117 517378 185151 517412
rect 177389 516546 177423 516580
rect 182541 516546 182575 516580
rect 174813 516290 174847 516324
rect 179965 516290 179999 516324
rect 185117 516290 185151 516324
rect 174813 515458 174847 515492
rect 177389 515458 177423 515492
rect 179965 515458 179999 515492
rect 182541 515458 182575 515492
rect 185117 515458 185151 515492
<< nsubdiffcont >>
rect 164538 538315 164578 539715
rect 164618 539695 166538 539735
rect 164618 538295 166538 538335
rect 166578 538315 166618 539715
rect 168338 538315 168378 539715
rect 168418 539695 170338 539735
rect 168418 538295 170338 538335
rect 170378 538315 170418 539715
rect 172038 538315 172078 539715
rect 172118 539695 174038 539735
rect 172118 538295 174038 538335
rect 174078 538315 174118 539715
rect 175538 538315 175578 539715
rect 175618 539695 177538 539735
rect 175618 538295 177538 538335
rect 177578 538315 177618 539715
rect 179138 538315 179178 539715
rect 179218 539695 181138 539735
rect 179218 538295 181138 538335
rect 181178 538315 181218 539715
rect 182438 538315 182478 539715
rect 182518 539695 184438 539735
rect 182518 538295 184438 538335
rect 184478 538315 184518 539715
rect 185738 538315 185778 539715
rect 185818 539695 187738 539735
rect 185818 538295 187738 538335
rect 187778 538315 187818 539715
rect 189038 538315 189078 539715
rect 189118 539695 191038 539735
rect 189118 538295 191038 538335
rect 191078 538315 191118 539715
rect 157648 537785 162748 537825
rect 157608 535785 157648 537725
rect 162788 535765 162828 537785
rect 157668 535705 162748 535745
rect 174813 530216 174847 530250
rect 174813 530123 174847 530157
rect 177389 530216 177423 530250
rect 177389 530123 177423 530157
rect 179965 530216 179999 530250
rect 179965 530123 179999 530157
rect 182541 530216 182575 530250
rect 182541 530123 182575 530157
rect 185117 530216 185151 530250
rect 185117 530123 185151 530157
rect 177389 529913 177423 529947
rect 177389 529820 177423 529854
rect 182541 529913 182575 529947
rect 182541 529820 182575 529854
rect 174813 529128 174847 529162
rect 174813 529035 174847 529069
rect 179965 529128 179999 529162
rect 179965 529035 179999 529069
rect 185117 529128 185151 529162
rect 185117 529035 185151 529069
rect 177389 528825 177423 528859
rect 177389 528732 177423 528766
rect 182541 528825 182575 528859
rect 182541 528732 182575 528766
rect 174813 528040 174847 528074
rect 174813 527947 174847 527981
rect 179965 528040 179999 528074
rect 179965 527947 179999 527981
rect 185117 528040 185151 528074
rect 185117 527947 185151 527981
rect 177389 527737 177423 527771
rect 177389 527644 177423 527678
rect 182541 527737 182575 527771
rect 182541 527644 182575 527678
rect 174813 526952 174847 526986
rect 174813 526859 174847 526893
rect 179965 526952 179999 526986
rect 179965 526859 179999 526893
rect 185117 526952 185151 526986
rect 185117 526859 185151 526893
rect 177389 526649 177423 526683
rect 177389 526556 177423 526590
rect 182541 526649 182575 526683
rect 182541 526556 182575 526590
rect 174813 525864 174847 525898
rect 174813 525771 174847 525805
rect 179965 525864 179999 525898
rect 179965 525771 179999 525805
rect 185117 525864 185151 525898
rect 185117 525771 185151 525805
rect 177389 525561 177423 525595
rect 177389 525468 177423 525502
rect 182541 525561 182575 525595
rect 182541 525468 182575 525502
rect 174813 524776 174847 524810
rect 174813 524683 174847 524717
rect 179965 524776 179999 524810
rect 179965 524683 179999 524717
rect 185117 524776 185151 524810
rect 185117 524683 185151 524717
rect 177389 524473 177423 524507
rect 177389 524380 177423 524414
rect 182541 524473 182575 524507
rect 182541 524380 182575 524414
rect 174813 523688 174847 523722
rect 174813 523595 174847 523629
rect 179965 523688 179999 523722
rect 179965 523595 179999 523629
rect 185117 523688 185151 523722
rect 185117 523595 185151 523629
rect 177389 523385 177423 523419
rect 177389 523292 177423 523326
rect 182541 523385 182575 523419
rect 182541 523292 182575 523326
rect 174813 522600 174847 522634
rect 174813 522507 174847 522541
rect 179965 522600 179999 522634
rect 179965 522507 179999 522541
rect 185117 522600 185151 522634
rect 185117 522507 185151 522541
rect 177389 522297 177423 522331
rect 177389 522204 177423 522238
rect 182541 522297 182575 522331
rect 182541 522204 182575 522238
rect 174813 521512 174847 521546
rect 174813 521419 174847 521453
rect 179965 521512 179999 521546
rect 179965 521419 179999 521453
rect 185117 521512 185151 521546
rect 185117 521419 185151 521453
rect 177389 521209 177423 521243
rect 177389 521116 177423 521150
rect 182541 521209 182575 521243
rect 182541 521116 182575 521150
rect 174813 520424 174847 520458
rect 174813 520331 174847 520365
rect 179965 520424 179999 520458
rect 179965 520331 179999 520365
rect 185117 520424 185151 520458
rect 185117 520331 185151 520365
rect 177389 520121 177423 520155
rect 177389 520028 177423 520062
rect 182541 520121 182575 520155
rect 182541 520028 182575 520062
rect 174813 519336 174847 519370
rect 174813 519243 174847 519277
rect 179965 519336 179999 519370
rect 179965 519243 179999 519277
rect 185117 519336 185151 519370
rect 185117 519243 185151 519277
rect 177389 519033 177423 519067
rect 177389 518940 177423 518974
rect 182541 519033 182575 519067
rect 182541 518940 182575 518974
rect 174813 518248 174847 518282
rect 174813 518155 174847 518189
rect 179965 518248 179999 518282
rect 179965 518155 179999 518189
rect 185117 518248 185151 518282
rect 185117 518155 185151 518189
rect 177389 517945 177423 517979
rect 177389 517852 177423 517886
rect 182541 517945 182575 517979
rect 182541 517852 182575 517886
rect 174813 517160 174847 517194
rect 174813 517067 174847 517101
rect 179965 517160 179999 517194
rect 179965 517067 179999 517101
rect 185117 517160 185151 517194
rect 185117 517067 185151 517101
rect 177389 516857 177423 516891
rect 177389 516764 177423 516798
rect 182541 516857 182575 516891
rect 182541 516764 182575 516798
rect 174813 516072 174847 516106
rect 174813 515979 174847 516013
rect 179965 516072 179999 516106
rect 179965 515979 179999 516013
rect 185117 516072 185151 516106
rect 185117 515979 185151 516013
rect 174813 515769 174847 515803
rect 174813 515676 174847 515710
rect 177389 515769 177423 515803
rect 177389 515676 177423 515710
rect 179965 515769 179999 515803
rect 179965 515676 179999 515710
rect 182541 515769 182575 515803
rect 182541 515676 182575 515710
rect 185117 515769 185151 515803
rect 185117 515676 185151 515710
<< poly >>
rect 164938 541142 166028 541145
rect 164938 541135 166041 541142
rect 164712 541119 164778 541135
rect 164712 541085 164728 541119
rect 164762 541085 164778 541119
rect 164712 541069 164778 541085
rect 164937 541126 166041 541135
rect 164937 541092 165031 541126
rect 165065 541092 165223 541126
rect 165257 541092 165415 541126
rect 165449 541092 165607 541126
rect 165641 541092 165799 541126
rect 165833 541092 165991 541126
rect 166025 541092 166041 541126
rect 164937 541085 166041 541092
rect 164730 541047 164760 541069
rect 164937 541054 164967 541085
rect 165015 541076 166041 541085
rect 166392 541119 166458 541135
rect 166392 541085 166408 541119
rect 166442 541085 166458 541119
rect 165032 541075 166028 541076
rect 165033 541054 165063 541075
rect 165129 541054 165159 541075
rect 165225 541054 165255 541075
rect 165321 541054 165351 541075
rect 165417 541054 165447 541075
rect 165513 541054 165543 541075
rect 165609 541054 165639 541075
rect 165705 541054 165735 541075
rect 165801 541054 165831 541075
rect 165897 541054 165927 541075
rect 165993 541054 166023 541075
rect 166392 541069 166458 541085
rect 166410 541047 166440 541069
rect 166192 540319 166258 540335
rect 166192 540285 166208 540319
rect 166242 540285 166258 540319
rect 166192 540269 166258 540285
rect 166210 540247 166240 540269
rect 164730 540025 164760 540047
rect 164937 540032 164967 540054
rect 164712 540009 164778 540025
rect 164712 539975 164728 540009
rect 164762 539975 164778 540009
rect 164712 539959 164778 539975
rect 164919 540016 164985 540032
rect 165033 540028 165063 540054
rect 165129 540032 165159 540054
rect 164919 539982 164935 540016
rect 164969 539982 164985 540016
rect 164919 539966 164985 539982
rect 165111 540016 165177 540032
rect 165225 540028 165255 540054
rect 165321 540032 165351 540054
rect 165111 539982 165127 540016
rect 165161 539982 165177 540016
rect 165111 539966 165177 539982
rect 165303 540016 165369 540032
rect 165417 540028 165447 540054
rect 165513 540032 165543 540054
rect 165303 539982 165319 540016
rect 165353 539982 165369 540016
rect 165303 539966 165369 539982
rect 165495 540016 165561 540032
rect 165609 540028 165639 540054
rect 165705 540032 165735 540054
rect 165495 539982 165511 540016
rect 165545 539982 165561 540016
rect 165495 539966 165561 539982
rect 165687 540016 165753 540032
rect 165801 540028 165831 540054
rect 165897 540032 165927 540054
rect 165687 539982 165703 540016
rect 165737 539982 165753 540016
rect 165687 539966 165753 539982
rect 165879 540016 165945 540032
rect 165993 540028 166023 540054
rect 166210 540025 166240 540047
rect 166410 540025 166440 540047
rect 165879 539982 165895 540016
rect 165929 539982 165945 540016
rect 165879 539966 165945 539982
rect 166192 540009 166258 540025
rect 166192 539975 166208 540009
rect 166242 539975 166258 540009
rect 166192 539959 166258 539975
rect 166392 540009 166458 540025
rect 166392 539975 166408 540009
rect 166442 539975 166458 540009
rect 166392 539959 166458 539975
rect 168738 541142 169828 541145
rect 168738 541135 169841 541142
rect 168512 541119 168578 541135
rect 168512 541085 168528 541119
rect 168562 541085 168578 541119
rect 168512 541069 168578 541085
rect 168737 541126 169841 541135
rect 168737 541092 168831 541126
rect 168865 541092 169023 541126
rect 169057 541092 169215 541126
rect 169249 541092 169407 541126
rect 169441 541092 169599 541126
rect 169633 541092 169791 541126
rect 169825 541092 169841 541126
rect 168737 541085 169841 541092
rect 168530 541047 168560 541069
rect 168737 541054 168767 541085
rect 168815 541076 169841 541085
rect 170192 541119 170258 541135
rect 170192 541085 170208 541119
rect 170242 541085 170258 541119
rect 168832 541075 169828 541076
rect 168833 541054 168863 541075
rect 168929 541054 168959 541075
rect 169025 541054 169055 541075
rect 169121 541054 169151 541075
rect 169217 541054 169247 541075
rect 169313 541054 169343 541075
rect 169409 541054 169439 541075
rect 169505 541054 169535 541075
rect 169601 541054 169631 541075
rect 169697 541054 169727 541075
rect 169793 541054 169823 541075
rect 170192 541069 170258 541085
rect 170210 541047 170240 541069
rect 169992 540319 170058 540335
rect 169992 540285 170008 540319
rect 170042 540285 170058 540319
rect 169992 540269 170058 540285
rect 170010 540247 170040 540269
rect 168530 540025 168560 540047
rect 168737 540032 168767 540054
rect 168512 540009 168578 540025
rect 168512 539975 168528 540009
rect 168562 539975 168578 540009
rect 168512 539959 168578 539975
rect 168719 540016 168785 540032
rect 168833 540028 168863 540054
rect 168929 540032 168959 540054
rect 168719 539982 168735 540016
rect 168769 539982 168785 540016
rect 168719 539966 168785 539982
rect 168911 540016 168977 540032
rect 169025 540028 169055 540054
rect 169121 540032 169151 540054
rect 168911 539982 168927 540016
rect 168961 539982 168977 540016
rect 168911 539966 168977 539982
rect 169103 540016 169169 540032
rect 169217 540028 169247 540054
rect 169313 540032 169343 540054
rect 169103 539982 169119 540016
rect 169153 539982 169169 540016
rect 169103 539966 169169 539982
rect 169295 540016 169361 540032
rect 169409 540028 169439 540054
rect 169505 540032 169535 540054
rect 169295 539982 169311 540016
rect 169345 539982 169361 540016
rect 169295 539966 169361 539982
rect 169487 540016 169553 540032
rect 169601 540028 169631 540054
rect 169697 540032 169727 540054
rect 169487 539982 169503 540016
rect 169537 539982 169553 540016
rect 169487 539966 169553 539982
rect 169679 540016 169745 540032
rect 169793 540028 169823 540054
rect 170010 540025 170040 540047
rect 170210 540025 170240 540047
rect 169679 539982 169695 540016
rect 169729 539982 169745 540016
rect 169679 539966 169745 539982
rect 169992 540009 170058 540025
rect 169992 539975 170008 540009
rect 170042 539975 170058 540009
rect 169992 539959 170058 539975
rect 170192 540009 170258 540025
rect 170192 539975 170208 540009
rect 170242 539975 170258 540009
rect 170192 539959 170258 539975
rect 172438 541142 173528 541145
rect 172438 541135 173541 541142
rect 172212 541119 172278 541135
rect 172212 541085 172228 541119
rect 172262 541085 172278 541119
rect 172212 541069 172278 541085
rect 172437 541126 173541 541135
rect 172437 541092 172531 541126
rect 172565 541092 172723 541126
rect 172757 541092 172915 541126
rect 172949 541092 173107 541126
rect 173141 541092 173299 541126
rect 173333 541092 173491 541126
rect 173525 541092 173541 541126
rect 172437 541085 173541 541092
rect 172230 541047 172260 541069
rect 172437 541054 172467 541085
rect 172515 541076 173541 541085
rect 173892 541119 173958 541135
rect 173892 541085 173908 541119
rect 173942 541085 173958 541119
rect 172532 541075 173528 541076
rect 172533 541054 172563 541075
rect 172629 541054 172659 541075
rect 172725 541054 172755 541075
rect 172821 541054 172851 541075
rect 172917 541054 172947 541075
rect 173013 541054 173043 541075
rect 173109 541054 173139 541075
rect 173205 541054 173235 541075
rect 173301 541054 173331 541075
rect 173397 541054 173427 541075
rect 173493 541054 173523 541075
rect 173892 541069 173958 541085
rect 173910 541047 173940 541069
rect 173692 540319 173758 540335
rect 173692 540285 173708 540319
rect 173742 540285 173758 540319
rect 173692 540269 173758 540285
rect 173710 540247 173740 540269
rect 172230 540025 172260 540047
rect 172437 540032 172467 540054
rect 172212 540009 172278 540025
rect 172212 539975 172228 540009
rect 172262 539975 172278 540009
rect 172212 539959 172278 539975
rect 172419 540016 172485 540032
rect 172533 540028 172563 540054
rect 172629 540032 172659 540054
rect 172419 539982 172435 540016
rect 172469 539982 172485 540016
rect 172419 539966 172485 539982
rect 172611 540016 172677 540032
rect 172725 540028 172755 540054
rect 172821 540032 172851 540054
rect 172611 539982 172627 540016
rect 172661 539982 172677 540016
rect 172611 539966 172677 539982
rect 172803 540016 172869 540032
rect 172917 540028 172947 540054
rect 173013 540032 173043 540054
rect 172803 539982 172819 540016
rect 172853 539982 172869 540016
rect 172803 539966 172869 539982
rect 172995 540016 173061 540032
rect 173109 540028 173139 540054
rect 173205 540032 173235 540054
rect 172995 539982 173011 540016
rect 173045 539982 173061 540016
rect 172995 539966 173061 539982
rect 173187 540016 173253 540032
rect 173301 540028 173331 540054
rect 173397 540032 173427 540054
rect 173187 539982 173203 540016
rect 173237 539982 173253 540016
rect 173187 539966 173253 539982
rect 173379 540016 173445 540032
rect 173493 540028 173523 540054
rect 173710 540025 173740 540047
rect 173910 540025 173940 540047
rect 173379 539982 173395 540016
rect 173429 539982 173445 540016
rect 173379 539966 173445 539982
rect 173692 540009 173758 540025
rect 173692 539975 173708 540009
rect 173742 539975 173758 540009
rect 173692 539959 173758 539975
rect 173892 540009 173958 540025
rect 173892 539975 173908 540009
rect 173942 539975 173958 540009
rect 173892 539959 173958 539975
rect 175938 541142 177028 541145
rect 175938 541135 177041 541142
rect 175712 541119 175778 541135
rect 175712 541085 175728 541119
rect 175762 541085 175778 541119
rect 175712 541069 175778 541085
rect 175937 541126 177041 541135
rect 175937 541092 176031 541126
rect 176065 541092 176223 541126
rect 176257 541092 176415 541126
rect 176449 541092 176607 541126
rect 176641 541092 176799 541126
rect 176833 541092 176991 541126
rect 177025 541092 177041 541126
rect 175937 541085 177041 541092
rect 175730 541047 175760 541069
rect 175937 541054 175967 541085
rect 176015 541076 177041 541085
rect 177392 541119 177458 541135
rect 177392 541085 177408 541119
rect 177442 541085 177458 541119
rect 176032 541075 177028 541076
rect 176033 541054 176063 541075
rect 176129 541054 176159 541075
rect 176225 541054 176255 541075
rect 176321 541054 176351 541075
rect 176417 541054 176447 541075
rect 176513 541054 176543 541075
rect 176609 541054 176639 541075
rect 176705 541054 176735 541075
rect 176801 541054 176831 541075
rect 176897 541054 176927 541075
rect 176993 541054 177023 541075
rect 177392 541069 177458 541085
rect 177410 541047 177440 541069
rect 177192 540319 177258 540335
rect 177192 540285 177208 540319
rect 177242 540285 177258 540319
rect 177192 540269 177258 540285
rect 177210 540247 177240 540269
rect 175730 540025 175760 540047
rect 175937 540032 175967 540054
rect 175712 540009 175778 540025
rect 175712 539975 175728 540009
rect 175762 539975 175778 540009
rect 175712 539959 175778 539975
rect 175919 540016 175985 540032
rect 176033 540028 176063 540054
rect 176129 540032 176159 540054
rect 175919 539982 175935 540016
rect 175969 539982 175985 540016
rect 175919 539966 175985 539982
rect 176111 540016 176177 540032
rect 176225 540028 176255 540054
rect 176321 540032 176351 540054
rect 176111 539982 176127 540016
rect 176161 539982 176177 540016
rect 176111 539966 176177 539982
rect 176303 540016 176369 540032
rect 176417 540028 176447 540054
rect 176513 540032 176543 540054
rect 176303 539982 176319 540016
rect 176353 539982 176369 540016
rect 176303 539966 176369 539982
rect 176495 540016 176561 540032
rect 176609 540028 176639 540054
rect 176705 540032 176735 540054
rect 176495 539982 176511 540016
rect 176545 539982 176561 540016
rect 176495 539966 176561 539982
rect 176687 540016 176753 540032
rect 176801 540028 176831 540054
rect 176897 540032 176927 540054
rect 176687 539982 176703 540016
rect 176737 539982 176753 540016
rect 176687 539966 176753 539982
rect 176879 540016 176945 540032
rect 176993 540028 177023 540054
rect 177210 540025 177240 540047
rect 177410 540025 177440 540047
rect 176879 539982 176895 540016
rect 176929 539982 176945 540016
rect 176879 539966 176945 539982
rect 177192 540009 177258 540025
rect 177192 539975 177208 540009
rect 177242 539975 177258 540009
rect 177192 539959 177258 539975
rect 177392 540009 177458 540025
rect 177392 539975 177408 540009
rect 177442 539975 177458 540009
rect 177392 539959 177458 539975
rect 179538 541142 180628 541145
rect 179538 541135 180641 541142
rect 179312 541119 179378 541135
rect 179312 541085 179328 541119
rect 179362 541085 179378 541119
rect 179312 541069 179378 541085
rect 179537 541126 180641 541135
rect 179537 541092 179631 541126
rect 179665 541092 179823 541126
rect 179857 541092 180015 541126
rect 180049 541092 180207 541126
rect 180241 541092 180399 541126
rect 180433 541092 180591 541126
rect 180625 541092 180641 541126
rect 179537 541085 180641 541092
rect 179330 541047 179360 541069
rect 179537 541054 179567 541085
rect 179615 541076 180641 541085
rect 180992 541119 181058 541135
rect 180992 541085 181008 541119
rect 181042 541085 181058 541119
rect 179632 541075 180628 541076
rect 179633 541054 179663 541075
rect 179729 541054 179759 541075
rect 179825 541054 179855 541075
rect 179921 541054 179951 541075
rect 180017 541054 180047 541075
rect 180113 541054 180143 541075
rect 180209 541054 180239 541075
rect 180305 541054 180335 541075
rect 180401 541054 180431 541075
rect 180497 541054 180527 541075
rect 180593 541054 180623 541075
rect 180992 541069 181058 541085
rect 181010 541047 181040 541069
rect 180792 540319 180858 540335
rect 180792 540285 180808 540319
rect 180842 540285 180858 540319
rect 180792 540269 180858 540285
rect 180810 540247 180840 540269
rect 179330 540025 179360 540047
rect 179537 540032 179567 540054
rect 179312 540009 179378 540025
rect 179312 539975 179328 540009
rect 179362 539975 179378 540009
rect 179312 539959 179378 539975
rect 179519 540016 179585 540032
rect 179633 540028 179663 540054
rect 179729 540032 179759 540054
rect 179519 539982 179535 540016
rect 179569 539982 179585 540016
rect 179519 539966 179585 539982
rect 179711 540016 179777 540032
rect 179825 540028 179855 540054
rect 179921 540032 179951 540054
rect 179711 539982 179727 540016
rect 179761 539982 179777 540016
rect 179711 539966 179777 539982
rect 179903 540016 179969 540032
rect 180017 540028 180047 540054
rect 180113 540032 180143 540054
rect 179903 539982 179919 540016
rect 179953 539982 179969 540016
rect 179903 539966 179969 539982
rect 180095 540016 180161 540032
rect 180209 540028 180239 540054
rect 180305 540032 180335 540054
rect 180095 539982 180111 540016
rect 180145 539982 180161 540016
rect 180095 539966 180161 539982
rect 180287 540016 180353 540032
rect 180401 540028 180431 540054
rect 180497 540032 180527 540054
rect 180287 539982 180303 540016
rect 180337 539982 180353 540016
rect 180287 539966 180353 539982
rect 180479 540016 180545 540032
rect 180593 540028 180623 540054
rect 180810 540025 180840 540047
rect 181010 540025 181040 540047
rect 180479 539982 180495 540016
rect 180529 539982 180545 540016
rect 180479 539966 180545 539982
rect 180792 540009 180858 540025
rect 180792 539975 180808 540009
rect 180842 539975 180858 540009
rect 180792 539959 180858 539975
rect 180992 540009 181058 540025
rect 180992 539975 181008 540009
rect 181042 539975 181058 540009
rect 180992 539959 181058 539975
rect 182838 541142 183928 541145
rect 182838 541135 183941 541142
rect 182612 541119 182678 541135
rect 182612 541085 182628 541119
rect 182662 541085 182678 541119
rect 182612 541069 182678 541085
rect 182837 541126 183941 541135
rect 182837 541092 182931 541126
rect 182965 541092 183123 541126
rect 183157 541092 183315 541126
rect 183349 541092 183507 541126
rect 183541 541092 183699 541126
rect 183733 541092 183891 541126
rect 183925 541092 183941 541126
rect 182837 541085 183941 541092
rect 182630 541047 182660 541069
rect 182837 541054 182867 541085
rect 182915 541076 183941 541085
rect 184292 541119 184358 541135
rect 184292 541085 184308 541119
rect 184342 541085 184358 541119
rect 182932 541075 183928 541076
rect 182933 541054 182963 541075
rect 183029 541054 183059 541075
rect 183125 541054 183155 541075
rect 183221 541054 183251 541075
rect 183317 541054 183347 541075
rect 183413 541054 183443 541075
rect 183509 541054 183539 541075
rect 183605 541054 183635 541075
rect 183701 541054 183731 541075
rect 183797 541054 183827 541075
rect 183893 541054 183923 541075
rect 184292 541069 184358 541085
rect 184310 541047 184340 541069
rect 184092 540319 184158 540335
rect 184092 540285 184108 540319
rect 184142 540285 184158 540319
rect 184092 540269 184158 540285
rect 184110 540247 184140 540269
rect 182630 540025 182660 540047
rect 182837 540032 182867 540054
rect 182612 540009 182678 540025
rect 182612 539975 182628 540009
rect 182662 539975 182678 540009
rect 182612 539959 182678 539975
rect 182819 540016 182885 540032
rect 182933 540028 182963 540054
rect 183029 540032 183059 540054
rect 182819 539982 182835 540016
rect 182869 539982 182885 540016
rect 182819 539966 182885 539982
rect 183011 540016 183077 540032
rect 183125 540028 183155 540054
rect 183221 540032 183251 540054
rect 183011 539982 183027 540016
rect 183061 539982 183077 540016
rect 183011 539966 183077 539982
rect 183203 540016 183269 540032
rect 183317 540028 183347 540054
rect 183413 540032 183443 540054
rect 183203 539982 183219 540016
rect 183253 539982 183269 540016
rect 183203 539966 183269 539982
rect 183395 540016 183461 540032
rect 183509 540028 183539 540054
rect 183605 540032 183635 540054
rect 183395 539982 183411 540016
rect 183445 539982 183461 540016
rect 183395 539966 183461 539982
rect 183587 540016 183653 540032
rect 183701 540028 183731 540054
rect 183797 540032 183827 540054
rect 183587 539982 183603 540016
rect 183637 539982 183653 540016
rect 183587 539966 183653 539982
rect 183779 540016 183845 540032
rect 183893 540028 183923 540054
rect 184110 540025 184140 540047
rect 184310 540025 184340 540047
rect 183779 539982 183795 540016
rect 183829 539982 183845 540016
rect 183779 539966 183845 539982
rect 184092 540009 184158 540025
rect 184092 539975 184108 540009
rect 184142 539975 184158 540009
rect 184092 539959 184158 539975
rect 184292 540009 184358 540025
rect 184292 539975 184308 540009
rect 184342 539975 184358 540009
rect 184292 539959 184358 539975
rect 186138 541142 187228 541145
rect 186138 541135 187241 541142
rect 185912 541119 185978 541135
rect 185912 541085 185928 541119
rect 185962 541085 185978 541119
rect 185912 541069 185978 541085
rect 186137 541126 187241 541135
rect 186137 541092 186231 541126
rect 186265 541092 186423 541126
rect 186457 541092 186615 541126
rect 186649 541092 186807 541126
rect 186841 541092 186999 541126
rect 187033 541092 187191 541126
rect 187225 541092 187241 541126
rect 186137 541085 187241 541092
rect 185930 541047 185960 541069
rect 186137 541054 186167 541085
rect 186215 541076 187241 541085
rect 187592 541119 187658 541135
rect 187592 541085 187608 541119
rect 187642 541085 187658 541119
rect 186232 541075 187228 541076
rect 186233 541054 186263 541075
rect 186329 541054 186359 541075
rect 186425 541054 186455 541075
rect 186521 541054 186551 541075
rect 186617 541054 186647 541075
rect 186713 541054 186743 541075
rect 186809 541054 186839 541075
rect 186905 541054 186935 541075
rect 187001 541054 187031 541075
rect 187097 541054 187127 541075
rect 187193 541054 187223 541075
rect 187592 541069 187658 541085
rect 187610 541047 187640 541069
rect 187392 540319 187458 540335
rect 187392 540285 187408 540319
rect 187442 540285 187458 540319
rect 187392 540269 187458 540285
rect 187410 540247 187440 540269
rect 185930 540025 185960 540047
rect 186137 540032 186167 540054
rect 185912 540009 185978 540025
rect 185912 539975 185928 540009
rect 185962 539975 185978 540009
rect 185912 539959 185978 539975
rect 186119 540016 186185 540032
rect 186233 540028 186263 540054
rect 186329 540032 186359 540054
rect 186119 539982 186135 540016
rect 186169 539982 186185 540016
rect 186119 539966 186185 539982
rect 186311 540016 186377 540032
rect 186425 540028 186455 540054
rect 186521 540032 186551 540054
rect 186311 539982 186327 540016
rect 186361 539982 186377 540016
rect 186311 539966 186377 539982
rect 186503 540016 186569 540032
rect 186617 540028 186647 540054
rect 186713 540032 186743 540054
rect 186503 539982 186519 540016
rect 186553 539982 186569 540016
rect 186503 539966 186569 539982
rect 186695 540016 186761 540032
rect 186809 540028 186839 540054
rect 186905 540032 186935 540054
rect 186695 539982 186711 540016
rect 186745 539982 186761 540016
rect 186695 539966 186761 539982
rect 186887 540016 186953 540032
rect 187001 540028 187031 540054
rect 187097 540032 187127 540054
rect 186887 539982 186903 540016
rect 186937 539982 186953 540016
rect 186887 539966 186953 539982
rect 187079 540016 187145 540032
rect 187193 540028 187223 540054
rect 187410 540025 187440 540047
rect 187610 540025 187640 540047
rect 187079 539982 187095 540016
rect 187129 539982 187145 540016
rect 187079 539966 187145 539982
rect 187392 540009 187458 540025
rect 187392 539975 187408 540009
rect 187442 539975 187458 540009
rect 187392 539959 187458 539975
rect 187592 540009 187658 540025
rect 187592 539975 187608 540009
rect 187642 539975 187658 540009
rect 187592 539959 187658 539975
rect 189438 541142 190528 541145
rect 189438 541135 190541 541142
rect 189212 541119 189278 541135
rect 189212 541085 189228 541119
rect 189262 541085 189278 541119
rect 189212 541069 189278 541085
rect 189437 541126 190541 541135
rect 189437 541092 189531 541126
rect 189565 541092 189723 541126
rect 189757 541092 189915 541126
rect 189949 541092 190107 541126
rect 190141 541092 190299 541126
rect 190333 541092 190491 541126
rect 190525 541092 190541 541126
rect 189437 541085 190541 541092
rect 189230 541047 189260 541069
rect 189437 541054 189467 541085
rect 189515 541076 190541 541085
rect 190892 541119 190958 541135
rect 190892 541085 190908 541119
rect 190942 541085 190958 541119
rect 189532 541075 190528 541076
rect 189533 541054 189563 541075
rect 189629 541054 189659 541075
rect 189725 541054 189755 541075
rect 189821 541054 189851 541075
rect 189917 541054 189947 541075
rect 190013 541054 190043 541075
rect 190109 541054 190139 541075
rect 190205 541054 190235 541075
rect 190301 541054 190331 541075
rect 190397 541054 190427 541075
rect 190493 541054 190523 541075
rect 190892 541069 190958 541085
rect 190910 541047 190940 541069
rect 190692 540319 190758 540335
rect 190692 540285 190708 540319
rect 190742 540285 190758 540319
rect 190692 540269 190758 540285
rect 190710 540247 190740 540269
rect 189230 540025 189260 540047
rect 189437 540032 189467 540054
rect 189212 540009 189278 540025
rect 189212 539975 189228 540009
rect 189262 539975 189278 540009
rect 189212 539959 189278 539975
rect 189419 540016 189485 540032
rect 189533 540028 189563 540054
rect 189629 540032 189659 540054
rect 189419 539982 189435 540016
rect 189469 539982 189485 540016
rect 189419 539966 189485 539982
rect 189611 540016 189677 540032
rect 189725 540028 189755 540054
rect 189821 540032 189851 540054
rect 189611 539982 189627 540016
rect 189661 539982 189677 540016
rect 189611 539966 189677 539982
rect 189803 540016 189869 540032
rect 189917 540028 189947 540054
rect 190013 540032 190043 540054
rect 189803 539982 189819 540016
rect 189853 539982 189869 540016
rect 189803 539966 189869 539982
rect 189995 540016 190061 540032
rect 190109 540028 190139 540054
rect 190205 540032 190235 540054
rect 189995 539982 190011 540016
rect 190045 539982 190061 540016
rect 189995 539966 190061 539982
rect 190187 540016 190253 540032
rect 190301 540028 190331 540054
rect 190397 540032 190427 540054
rect 190187 539982 190203 540016
rect 190237 539982 190253 540016
rect 190187 539966 190253 539982
rect 190379 540016 190445 540032
rect 190493 540028 190523 540054
rect 190710 540025 190740 540047
rect 190910 540025 190940 540047
rect 190379 539982 190395 540016
rect 190429 539982 190445 540016
rect 190379 539966 190445 539982
rect 190692 540009 190758 540025
rect 190692 539975 190708 540009
rect 190742 539975 190758 540009
rect 190692 539959 190758 539975
rect 190892 540009 190958 540025
rect 190892 539975 190908 540009
rect 190942 539975 190958 540009
rect 190892 539959 190958 539975
rect 158710 538469 158910 538485
rect 158710 538435 158726 538469
rect 158894 538435 158910 538469
rect 158710 538397 158910 538435
rect 159086 538469 159286 538485
rect 159086 538435 159102 538469
rect 159270 538435 159286 538469
rect 159086 538397 159286 538435
rect 159344 538469 159544 538485
rect 159344 538435 159360 538469
rect 159528 538435 159544 538469
rect 159344 538397 159544 538435
rect 159602 538469 159802 538485
rect 159602 538435 159618 538469
rect 159786 538435 159802 538469
rect 159602 538397 159802 538435
rect 159860 538469 160060 538485
rect 159860 538435 159876 538469
rect 160044 538435 160060 538469
rect 159860 538397 160060 538435
rect 160118 538469 160318 538485
rect 160118 538435 160134 538469
rect 160302 538435 160318 538469
rect 160118 538397 160318 538435
rect 160376 538469 160576 538485
rect 160376 538435 160392 538469
rect 160560 538435 160576 538469
rect 160376 538397 160576 538435
rect 160634 538469 160834 538485
rect 160634 538435 160650 538469
rect 160818 538435 160834 538469
rect 160634 538397 160834 538435
rect 160892 538469 161092 538485
rect 160892 538435 160908 538469
rect 161076 538435 161092 538469
rect 160892 538397 161092 538435
rect 161150 538469 161350 538485
rect 161150 538435 161166 538469
rect 161334 538435 161350 538469
rect 161150 538397 161350 538435
rect 161530 538469 161730 538485
rect 161530 538435 161546 538469
rect 161714 538435 161730 538469
rect 161530 538397 161730 538435
rect 161930 538469 162130 538485
rect 161930 538435 161946 538469
rect 162114 538435 162130 538469
rect 161930 538397 162130 538435
rect 162310 538469 162510 538485
rect 162310 538435 162326 538469
rect 162494 538435 162510 538469
rect 162310 538397 162510 538435
rect 158710 538159 158910 538197
rect 158710 538125 158726 538159
rect 158894 538125 158910 538159
rect 158710 538109 158910 538125
rect 159086 538159 159286 538197
rect 159086 538125 159102 538159
rect 159270 538125 159286 538159
rect 159086 538109 159286 538125
rect 159344 538159 159544 538197
rect 159344 538125 159360 538159
rect 159528 538125 159544 538159
rect 159344 538109 159544 538125
rect 159602 538159 159802 538197
rect 159602 538125 159618 538159
rect 159786 538125 159802 538159
rect 159602 538109 159802 538125
rect 159860 538159 160060 538197
rect 159860 538125 159876 538159
rect 160044 538125 160060 538159
rect 159860 538109 160060 538125
rect 160118 538159 160318 538197
rect 160118 538125 160134 538159
rect 160302 538125 160318 538159
rect 160118 538109 160318 538125
rect 160376 538159 160576 538197
rect 160376 538125 160392 538159
rect 160560 538125 160576 538159
rect 160376 538109 160576 538125
rect 160634 538159 160834 538197
rect 160634 538125 160650 538159
rect 160818 538125 160834 538159
rect 160634 538109 160834 538125
rect 160892 538159 161092 538197
rect 160892 538125 160908 538159
rect 161076 538125 161092 538159
rect 160892 538109 161092 538125
rect 161150 538159 161350 538197
rect 161150 538125 161166 538159
rect 161334 538125 161350 538159
rect 161150 538109 161350 538125
rect 161530 538159 161730 538197
rect 161530 538125 161546 538159
rect 161714 538125 161730 538159
rect 161530 538109 161730 538125
rect 161930 538159 162130 538197
rect 161930 538125 161946 538159
rect 162114 538125 162130 538159
rect 161930 538109 162130 538125
rect 162310 538159 162510 538197
rect 162310 538125 162326 538159
rect 162494 538125 162510 538159
rect 162310 538109 162510 538125
rect 164696 539606 164762 539622
rect 164696 539572 164712 539606
rect 164746 539572 164762 539606
rect 164696 539556 164762 539572
rect 165019 539613 165085 539629
rect 165019 539579 165035 539613
rect 165069 539579 165085 539613
rect 165019 539563 165085 539579
rect 165211 539613 165277 539629
rect 165211 539579 165227 539613
rect 165261 539579 165277 539613
rect 165211 539563 165277 539579
rect 165403 539613 165469 539629
rect 165403 539579 165419 539613
rect 165453 539579 165469 539613
rect 165403 539563 165469 539579
rect 165595 539613 165661 539629
rect 165595 539579 165611 539613
rect 165645 539579 165661 539613
rect 165595 539563 165661 539579
rect 165787 539613 165853 539629
rect 165787 539579 165803 539613
rect 165837 539579 165853 539613
rect 165787 539563 165853 539579
rect 165979 539613 166045 539629
rect 165979 539579 165995 539613
rect 166029 539579 166045 539613
rect 165979 539563 166045 539579
rect 166196 539606 166262 539622
rect 166196 539572 166212 539606
rect 166246 539572 166262 539606
rect 164714 539525 164744 539556
rect 164941 539532 164971 539558
rect 165037 539532 165067 539563
rect 165133 539532 165163 539558
rect 165229 539532 165259 539563
rect 165325 539532 165355 539558
rect 165421 539532 165451 539563
rect 165517 539532 165547 539558
rect 165613 539532 165643 539563
rect 165709 539532 165739 539558
rect 165805 539532 165835 539563
rect 165901 539532 165931 539558
rect 165997 539532 166027 539563
rect 166196 539556 166262 539572
rect 166396 539606 166462 539622
rect 166396 539572 166412 539606
rect 166446 539572 166462 539606
rect 166396 539556 166462 539572
rect 166214 539525 166244 539556
rect 166414 539525 166444 539556
rect 166214 538894 166244 538925
rect 166196 538878 166262 538894
rect 166196 538844 166212 538878
rect 166246 538844 166262 538878
rect 166196 538828 166262 538844
rect 164714 538494 164744 538525
rect 164941 538501 164971 538532
rect 164923 538495 164989 538501
rect 165037 538495 165067 538532
rect 165133 538501 165163 538532
rect 165115 538495 165181 538501
rect 165229 538495 165259 538532
rect 165325 538501 165355 538532
rect 165307 538495 165373 538501
rect 165421 538495 165451 538532
rect 165517 538501 165547 538532
rect 165499 538495 165565 538501
rect 165613 538495 165643 538532
rect 165709 538501 165739 538532
rect 165691 538495 165757 538501
rect 165805 538495 165835 538532
rect 165901 538501 165931 538532
rect 165997 538515 166027 538532
rect 165883 538495 165949 538501
rect 165994 538495 166028 538515
rect 164696 538478 164762 538494
rect 164696 538444 164712 538478
rect 164746 538444 164762 538478
rect 164696 538428 164762 538444
rect 164923 538485 166028 538495
rect 166414 538494 166444 538525
rect 164923 538451 164939 538485
rect 164973 538451 165131 538485
rect 165165 538451 165323 538485
rect 165357 538451 165515 538485
rect 165549 538451 165707 538485
rect 165741 538451 165899 538485
rect 165933 538451 166028 538485
rect 164923 538445 166028 538451
rect 166396 538478 166462 538494
rect 164923 538435 164989 538445
rect 165115 538435 165181 538445
rect 165307 538435 165373 538445
rect 165499 538435 165565 538445
rect 165691 538435 165757 538445
rect 165883 538435 165949 538445
rect 166396 538444 166412 538478
rect 166446 538444 166462 538478
rect 166396 538428 166462 538444
rect 168496 539606 168562 539622
rect 168496 539572 168512 539606
rect 168546 539572 168562 539606
rect 168496 539556 168562 539572
rect 168819 539613 168885 539629
rect 168819 539579 168835 539613
rect 168869 539579 168885 539613
rect 168819 539563 168885 539579
rect 169011 539613 169077 539629
rect 169011 539579 169027 539613
rect 169061 539579 169077 539613
rect 169011 539563 169077 539579
rect 169203 539613 169269 539629
rect 169203 539579 169219 539613
rect 169253 539579 169269 539613
rect 169203 539563 169269 539579
rect 169395 539613 169461 539629
rect 169395 539579 169411 539613
rect 169445 539579 169461 539613
rect 169395 539563 169461 539579
rect 169587 539613 169653 539629
rect 169587 539579 169603 539613
rect 169637 539579 169653 539613
rect 169587 539563 169653 539579
rect 169779 539613 169845 539629
rect 169779 539579 169795 539613
rect 169829 539579 169845 539613
rect 169779 539563 169845 539579
rect 169996 539606 170062 539622
rect 169996 539572 170012 539606
rect 170046 539572 170062 539606
rect 168514 539525 168544 539556
rect 168741 539532 168771 539558
rect 168837 539532 168867 539563
rect 168933 539532 168963 539558
rect 169029 539532 169059 539563
rect 169125 539532 169155 539558
rect 169221 539532 169251 539563
rect 169317 539532 169347 539558
rect 169413 539532 169443 539563
rect 169509 539532 169539 539558
rect 169605 539532 169635 539563
rect 169701 539532 169731 539558
rect 169797 539532 169827 539563
rect 169996 539556 170062 539572
rect 170196 539606 170262 539622
rect 170196 539572 170212 539606
rect 170246 539572 170262 539606
rect 170196 539556 170262 539572
rect 170014 539525 170044 539556
rect 170214 539525 170244 539556
rect 170014 538894 170044 538925
rect 169996 538878 170062 538894
rect 169996 538844 170012 538878
rect 170046 538844 170062 538878
rect 169996 538828 170062 538844
rect 168514 538494 168544 538525
rect 168741 538501 168771 538532
rect 168723 538495 168789 538501
rect 168837 538495 168867 538532
rect 168933 538501 168963 538532
rect 168915 538495 168981 538501
rect 169029 538495 169059 538532
rect 169125 538501 169155 538532
rect 169107 538495 169173 538501
rect 169221 538495 169251 538532
rect 169317 538501 169347 538532
rect 169299 538495 169365 538501
rect 169413 538495 169443 538532
rect 169509 538501 169539 538532
rect 169491 538495 169557 538501
rect 169605 538495 169635 538532
rect 169701 538501 169731 538532
rect 169797 538515 169827 538532
rect 169683 538495 169749 538501
rect 169794 538495 169828 538515
rect 168496 538478 168562 538494
rect 168496 538444 168512 538478
rect 168546 538444 168562 538478
rect 168496 538428 168562 538444
rect 168723 538485 169828 538495
rect 170214 538494 170244 538525
rect 168723 538451 168739 538485
rect 168773 538451 168931 538485
rect 168965 538451 169123 538485
rect 169157 538451 169315 538485
rect 169349 538451 169507 538485
rect 169541 538451 169699 538485
rect 169733 538451 169828 538485
rect 168723 538445 169828 538451
rect 170196 538478 170262 538494
rect 168723 538435 168789 538445
rect 168915 538435 168981 538445
rect 169107 538435 169173 538445
rect 169299 538435 169365 538445
rect 169491 538435 169557 538445
rect 169683 538435 169749 538445
rect 170196 538444 170212 538478
rect 170246 538444 170262 538478
rect 170196 538428 170262 538444
rect 172196 539606 172262 539622
rect 172196 539572 172212 539606
rect 172246 539572 172262 539606
rect 172196 539556 172262 539572
rect 172519 539613 172585 539629
rect 172519 539579 172535 539613
rect 172569 539579 172585 539613
rect 172519 539563 172585 539579
rect 172711 539613 172777 539629
rect 172711 539579 172727 539613
rect 172761 539579 172777 539613
rect 172711 539563 172777 539579
rect 172903 539613 172969 539629
rect 172903 539579 172919 539613
rect 172953 539579 172969 539613
rect 172903 539563 172969 539579
rect 173095 539613 173161 539629
rect 173095 539579 173111 539613
rect 173145 539579 173161 539613
rect 173095 539563 173161 539579
rect 173287 539613 173353 539629
rect 173287 539579 173303 539613
rect 173337 539579 173353 539613
rect 173287 539563 173353 539579
rect 173479 539613 173545 539629
rect 173479 539579 173495 539613
rect 173529 539579 173545 539613
rect 173479 539563 173545 539579
rect 173696 539606 173762 539622
rect 173696 539572 173712 539606
rect 173746 539572 173762 539606
rect 172214 539525 172244 539556
rect 172441 539532 172471 539558
rect 172537 539532 172567 539563
rect 172633 539532 172663 539558
rect 172729 539532 172759 539563
rect 172825 539532 172855 539558
rect 172921 539532 172951 539563
rect 173017 539532 173047 539558
rect 173113 539532 173143 539563
rect 173209 539532 173239 539558
rect 173305 539532 173335 539563
rect 173401 539532 173431 539558
rect 173497 539532 173527 539563
rect 173696 539556 173762 539572
rect 173896 539606 173962 539622
rect 173896 539572 173912 539606
rect 173946 539572 173962 539606
rect 173896 539556 173962 539572
rect 173714 539525 173744 539556
rect 173914 539525 173944 539556
rect 173714 538894 173744 538925
rect 173696 538878 173762 538894
rect 173696 538844 173712 538878
rect 173746 538844 173762 538878
rect 173696 538828 173762 538844
rect 172214 538494 172244 538525
rect 172441 538501 172471 538532
rect 172423 538495 172489 538501
rect 172537 538495 172567 538532
rect 172633 538501 172663 538532
rect 172615 538495 172681 538501
rect 172729 538495 172759 538532
rect 172825 538501 172855 538532
rect 172807 538495 172873 538501
rect 172921 538495 172951 538532
rect 173017 538501 173047 538532
rect 172999 538495 173065 538501
rect 173113 538495 173143 538532
rect 173209 538501 173239 538532
rect 173191 538495 173257 538501
rect 173305 538495 173335 538532
rect 173401 538501 173431 538532
rect 173497 538515 173527 538532
rect 173383 538495 173449 538501
rect 173494 538495 173528 538515
rect 172196 538478 172262 538494
rect 172196 538444 172212 538478
rect 172246 538444 172262 538478
rect 172196 538428 172262 538444
rect 172423 538485 173528 538495
rect 173914 538494 173944 538525
rect 172423 538451 172439 538485
rect 172473 538451 172631 538485
rect 172665 538451 172823 538485
rect 172857 538451 173015 538485
rect 173049 538451 173207 538485
rect 173241 538451 173399 538485
rect 173433 538451 173528 538485
rect 172423 538445 173528 538451
rect 173896 538478 173962 538494
rect 172423 538435 172489 538445
rect 172615 538435 172681 538445
rect 172807 538435 172873 538445
rect 172999 538435 173065 538445
rect 173191 538435 173257 538445
rect 173383 538435 173449 538445
rect 173896 538444 173912 538478
rect 173946 538444 173962 538478
rect 173896 538428 173962 538444
rect 175696 539606 175762 539622
rect 175696 539572 175712 539606
rect 175746 539572 175762 539606
rect 175696 539556 175762 539572
rect 176019 539613 176085 539629
rect 176019 539579 176035 539613
rect 176069 539579 176085 539613
rect 176019 539563 176085 539579
rect 176211 539613 176277 539629
rect 176211 539579 176227 539613
rect 176261 539579 176277 539613
rect 176211 539563 176277 539579
rect 176403 539613 176469 539629
rect 176403 539579 176419 539613
rect 176453 539579 176469 539613
rect 176403 539563 176469 539579
rect 176595 539613 176661 539629
rect 176595 539579 176611 539613
rect 176645 539579 176661 539613
rect 176595 539563 176661 539579
rect 176787 539613 176853 539629
rect 176787 539579 176803 539613
rect 176837 539579 176853 539613
rect 176787 539563 176853 539579
rect 176979 539613 177045 539629
rect 176979 539579 176995 539613
rect 177029 539579 177045 539613
rect 176979 539563 177045 539579
rect 177196 539606 177262 539622
rect 177196 539572 177212 539606
rect 177246 539572 177262 539606
rect 175714 539525 175744 539556
rect 175941 539532 175971 539558
rect 176037 539532 176067 539563
rect 176133 539532 176163 539558
rect 176229 539532 176259 539563
rect 176325 539532 176355 539558
rect 176421 539532 176451 539563
rect 176517 539532 176547 539558
rect 176613 539532 176643 539563
rect 176709 539532 176739 539558
rect 176805 539532 176835 539563
rect 176901 539532 176931 539558
rect 176997 539532 177027 539563
rect 177196 539556 177262 539572
rect 177396 539606 177462 539622
rect 177396 539572 177412 539606
rect 177446 539572 177462 539606
rect 177396 539556 177462 539572
rect 177214 539525 177244 539556
rect 177414 539525 177444 539556
rect 177214 538894 177244 538925
rect 177196 538878 177262 538894
rect 177196 538844 177212 538878
rect 177246 538844 177262 538878
rect 177196 538828 177262 538844
rect 175714 538494 175744 538525
rect 175941 538501 175971 538532
rect 175923 538495 175989 538501
rect 176037 538495 176067 538532
rect 176133 538501 176163 538532
rect 176115 538495 176181 538501
rect 176229 538495 176259 538532
rect 176325 538501 176355 538532
rect 176307 538495 176373 538501
rect 176421 538495 176451 538532
rect 176517 538501 176547 538532
rect 176499 538495 176565 538501
rect 176613 538495 176643 538532
rect 176709 538501 176739 538532
rect 176691 538495 176757 538501
rect 176805 538495 176835 538532
rect 176901 538501 176931 538532
rect 176997 538515 177027 538532
rect 176883 538495 176949 538501
rect 176994 538495 177028 538515
rect 175696 538478 175762 538494
rect 175696 538444 175712 538478
rect 175746 538444 175762 538478
rect 175696 538428 175762 538444
rect 175923 538485 177028 538495
rect 177414 538494 177444 538525
rect 175923 538451 175939 538485
rect 175973 538451 176131 538485
rect 176165 538451 176323 538485
rect 176357 538451 176515 538485
rect 176549 538451 176707 538485
rect 176741 538451 176899 538485
rect 176933 538451 177028 538485
rect 175923 538445 177028 538451
rect 177396 538478 177462 538494
rect 175923 538435 175989 538445
rect 176115 538435 176181 538445
rect 176307 538435 176373 538445
rect 176499 538435 176565 538445
rect 176691 538435 176757 538445
rect 176883 538435 176949 538445
rect 177396 538444 177412 538478
rect 177446 538444 177462 538478
rect 177396 538428 177462 538444
rect 179296 539606 179362 539622
rect 179296 539572 179312 539606
rect 179346 539572 179362 539606
rect 179296 539556 179362 539572
rect 179619 539613 179685 539629
rect 179619 539579 179635 539613
rect 179669 539579 179685 539613
rect 179619 539563 179685 539579
rect 179811 539613 179877 539629
rect 179811 539579 179827 539613
rect 179861 539579 179877 539613
rect 179811 539563 179877 539579
rect 180003 539613 180069 539629
rect 180003 539579 180019 539613
rect 180053 539579 180069 539613
rect 180003 539563 180069 539579
rect 180195 539613 180261 539629
rect 180195 539579 180211 539613
rect 180245 539579 180261 539613
rect 180195 539563 180261 539579
rect 180387 539613 180453 539629
rect 180387 539579 180403 539613
rect 180437 539579 180453 539613
rect 180387 539563 180453 539579
rect 180579 539613 180645 539629
rect 180579 539579 180595 539613
rect 180629 539579 180645 539613
rect 180579 539563 180645 539579
rect 180796 539606 180862 539622
rect 180796 539572 180812 539606
rect 180846 539572 180862 539606
rect 179314 539525 179344 539556
rect 179541 539532 179571 539558
rect 179637 539532 179667 539563
rect 179733 539532 179763 539558
rect 179829 539532 179859 539563
rect 179925 539532 179955 539558
rect 180021 539532 180051 539563
rect 180117 539532 180147 539558
rect 180213 539532 180243 539563
rect 180309 539532 180339 539558
rect 180405 539532 180435 539563
rect 180501 539532 180531 539558
rect 180597 539532 180627 539563
rect 180796 539556 180862 539572
rect 180996 539606 181062 539622
rect 180996 539572 181012 539606
rect 181046 539572 181062 539606
rect 180996 539556 181062 539572
rect 180814 539525 180844 539556
rect 181014 539525 181044 539556
rect 180814 538894 180844 538925
rect 180796 538878 180862 538894
rect 180796 538844 180812 538878
rect 180846 538844 180862 538878
rect 180796 538828 180862 538844
rect 179314 538494 179344 538525
rect 179541 538501 179571 538532
rect 179523 538495 179589 538501
rect 179637 538495 179667 538532
rect 179733 538501 179763 538532
rect 179715 538495 179781 538501
rect 179829 538495 179859 538532
rect 179925 538501 179955 538532
rect 179907 538495 179973 538501
rect 180021 538495 180051 538532
rect 180117 538501 180147 538532
rect 180099 538495 180165 538501
rect 180213 538495 180243 538532
rect 180309 538501 180339 538532
rect 180291 538495 180357 538501
rect 180405 538495 180435 538532
rect 180501 538501 180531 538532
rect 180597 538515 180627 538532
rect 180483 538495 180549 538501
rect 180594 538495 180628 538515
rect 179296 538478 179362 538494
rect 179296 538444 179312 538478
rect 179346 538444 179362 538478
rect 179296 538428 179362 538444
rect 179523 538485 180628 538495
rect 181014 538494 181044 538525
rect 179523 538451 179539 538485
rect 179573 538451 179731 538485
rect 179765 538451 179923 538485
rect 179957 538451 180115 538485
rect 180149 538451 180307 538485
rect 180341 538451 180499 538485
rect 180533 538451 180628 538485
rect 179523 538445 180628 538451
rect 180996 538478 181062 538494
rect 179523 538435 179589 538445
rect 179715 538435 179781 538445
rect 179907 538435 179973 538445
rect 180099 538435 180165 538445
rect 180291 538435 180357 538445
rect 180483 538435 180549 538445
rect 180996 538444 181012 538478
rect 181046 538444 181062 538478
rect 180996 538428 181062 538444
rect 182596 539606 182662 539622
rect 182596 539572 182612 539606
rect 182646 539572 182662 539606
rect 182596 539556 182662 539572
rect 182919 539613 182985 539629
rect 182919 539579 182935 539613
rect 182969 539579 182985 539613
rect 182919 539563 182985 539579
rect 183111 539613 183177 539629
rect 183111 539579 183127 539613
rect 183161 539579 183177 539613
rect 183111 539563 183177 539579
rect 183303 539613 183369 539629
rect 183303 539579 183319 539613
rect 183353 539579 183369 539613
rect 183303 539563 183369 539579
rect 183495 539613 183561 539629
rect 183495 539579 183511 539613
rect 183545 539579 183561 539613
rect 183495 539563 183561 539579
rect 183687 539613 183753 539629
rect 183687 539579 183703 539613
rect 183737 539579 183753 539613
rect 183687 539563 183753 539579
rect 183879 539613 183945 539629
rect 183879 539579 183895 539613
rect 183929 539579 183945 539613
rect 183879 539563 183945 539579
rect 184096 539606 184162 539622
rect 184096 539572 184112 539606
rect 184146 539572 184162 539606
rect 182614 539525 182644 539556
rect 182841 539532 182871 539558
rect 182937 539532 182967 539563
rect 183033 539532 183063 539558
rect 183129 539532 183159 539563
rect 183225 539532 183255 539558
rect 183321 539532 183351 539563
rect 183417 539532 183447 539558
rect 183513 539532 183543 539563
rect 183609 539532 183639 539558
rect 183705 539532 183735 539563
rect 183801 539532 183831 539558
rect 183897 539532 183927 539563
rect 184096 539556 184162 539572
rect 184296 539606 184362 539622
rect 184296 539572 184312 539606
rect 184346 539572 184362 539606
rect 184296 539556 184362 539572
rect 184114 539525 184144 539556
rect 184314 539525 184344 539556
rect 184114 538894 184144 538925
rect 184096 538878 184162 538894
rect 184096 538844 184112 538878
rect 184146 538844 184162 538878
rect 184096 538828 184162 538844
rect 182614 538494 182644 538525
rect 182841 538501 182871 538532
rect 182823 538495 182889 538501
rect 182937 538495 182967 538532
rect 183033 538501 183063 538532
rect 183015 538495 183081 538501
rect 183129 538495 183159 538532
rect 183225 538501 183255 538532
rect 183207 538495 183273 538501
rect 183321 538495 183351 538532
rect 183417 538501 183447 538532
rect 183399 538495 183465 538501
rect 183513 538495 183543 538532
rect 183609 538501 183639 538532
rect 183591 538495 183657 538501
rect 183705 538495 183735 538532
rect 183801 538501 183831 538532
rect 183897 538515 183927 538532
rect 183783 538495 183849 538501
rect 183894 538495 183928 538515
rect 182596 538478 182662 538494
rect 182596 538444 182612 538478
rect 182646 538444 182662 538478
rect 182596 538428 182662 538444
rect 182823 538485 183928 538495
rect 184314 538494 184344 538525
rect 182823 538451 182839 538485
rect 182873 538451 183031 538485
rect 183065 538451 183223 538485
rect 183257 538451 183415 538485
rect 183449 538451 183607 538485
rect 183641 538451 183799 538485
rect 183833 538451 183928 538485
rect 182823 538445 183928 538451
rect 184296 538478 184362 538494
rect 182823 538435 182889 538445
rect 183015 538435 183081 538445
rect 183207 538435 183273 538445
rect 183399 538435 183465 538445
rect 183591 538435 183657 538445
rect 183783 538435 183849 538445
rect 184296 538444 184312 538478
rect 184346 538444 184362 538478
rect 184296 538428 184362 538444
rect 185896 539606 185962 539622
rect 185896 539572 185912 539606
rect 185946 539572 185962 539606
rect 185896 539556 185962 539572
rect 186219 539613 186285 539629
rect 186219 539579 186235 539613
rect 186269 539579 186285 539613
rect 186219 539563 186285 539579
rect 186411 539613 186477 539629
rect 186411 539579 186427 539613
rect 186461 539579 186477 539613
rect 186411 539563 186477 539579
rect 186603 539613 186669 539629
rect 186603 539579 186619 539613
rect 186653 539579 186669 539613
rect 186603 539563 186669 539579
rect 186795 539613 186861 539629
rect 186795 539579 186811 539613
rect 186845 539579 186861 539613
rect 186795 539563 186861 539579
rect 186987 539613 187053 539629
rect 186987 539579 187003 539613
rect 187037 539579 187053 539613
rect 186987 539563 187053 539579
rect 187179 539613 187245 539629
rect 187179 539579 187195 539613
rect 187229 539579 187245 539613
rect 187179 539563 187245 539579
rect 187396 539606 187462 539622
rect 187396 539572 187412 539606
rect 187446 539572 187462 539606
rect 185914 539525 185944 539556
rect 186141 539532 186171 539558
rect 186237 539532 186267 539563
rect 186333 539532 186363 539558
rect 186429 539532 186459 539563
rect 186525 539532 186555 539558
rect 186621 539532 186651 539563
rect 186717 539532 186747 539558
rect 186813 539532 186843 539563
rect 186909 539532 186939 539558
rect 187005 539532 187035 539563
rect 187101 539532 187131 539558
rect 187197 539532 187227 539563
rect 187396 539556 187462 539572
rect 187596 539606 187662 539622
rect 187596 539572 187612 539606
rect 187646 539572 187662 539606
rect 187596 539556 187662 539572
rect 187414 539525 187444 539556
rect 187614 539525 187644 539556
rect 187414 538894 187444 538925
rect 187396 538878 187462 538894
rect 187396 538844 187412 538878
rect 187446 538844 187462 538878
rect 187396 538828 187462 538844
rect 185914 538494 185944 538525
rect 186141 538501 186171 538532
rect 186123 538495 186189 538501
rect 186237 538495 186267 538532
rect 186333 538501 186363 538532
rect 186315 538495 186381 538501
rect 186429 538495 186459 538532
rect 186525 538501 186555 538532
rect 186507 538495 186573 538501
rect 186621 538495 186651 538532
rect 186717 538501 186747 538532
rect 186699 538495 186765 538501
rect 186813 538495 186843 538532
rect 186909 538501 186939 538532
rect 186891 538495 186957 538501
rect 187005 538495 187035 538532
rect 187101 538501 187131 538532
rect 187197 538515 187227 538532
rect 187083 538495 187149 538501
rect 187194 538495 187228 538515
rect 185896 538478 185962 538494
rect 185896 538444 185912 538478
rect 185946 538444 185962 538478
rect 185896 538428 185962 538444
rect 186123 538485 187228 538495
rect 187614 538494 187644 538525
rect 186123 538451 186139 538485
rect 186173 538451 186331 538485
rect 186365 538451 186523 538485
rect 186557 538451 186715 538485
rect 186749 538451 186907 538485
rect 186941 538451 187099 538485
rect 187133 538451 187228 538485
rect 186123 538445 187228 538451
rect 187596 538478 187662 538494
rect 186123 538435 186189 538445
rect 186315 538435 186381 538445
rect 186507 538435 186573 538445
rect 186699 538435 186765 538445
rect 186891 538435 186957 538445
rect 187083 538435 187149 538445
rect 187596 538444 187612 538478
rect 187646 538444 187662 538478
rect 187596 538428 187662 538444
rect 189196 539606 189262 539622
rect 189196 539572 189212 539606
rect 189246 539572 189262 539606
rect 189196 539556 189262 539572
rect 189519 539613 189585 539629
rect 189519 539579 189535 539613
rect 189569 539579 189585 539613
rect 189519 539563 189585 539579
rect 189711 539613 189777 539629
rect 189711 539579 189727 539613
rect 189761 539579 189777 539613
rect 189711 539563 189777 539579
rect 189903 539613 189969 539629
rect 189903 539579 189919 539613
rect 189953 539579 189969 539613
rect 189903 539563 189969 539579
rect 190095 539613 190161 539629
rect 190095 539579 190111 539613
rect 190145 539579 190161 539613
rect 190095 539563 190161 539579
rect 190287 539613 190353 539629
rect 190287 539579 190303 539613
rect 190337 539579 190353 539613
rect 190287 539563 190353 539579
rect 190479 539613 190545 539629
rect 190479 539579 190495 539613
rect 190529 539579 190545 539613
rect 190479 539563 190545 539579
rect 190696 539606 190762 539622
rect 190696 539572 190712 539606
rect 190746 539572 190762 539606
rect 189214 539525 189244 539556
rect 189441 539532 189471 539558
rect 189537 539532 189567 539563
rect 189633 539532 189663 539558
rect 189729 539532 189759 539563
rect 189825 539532 189855 539558
rect 189921 539532 189951 539563
rect 190017 539532 190047 539558
rect 190113 539532 190143 539563
rect 190209 539532 190239 539558
rect 190305 539532 190335 539563
rect 190401 539532 190431 539558
rect 190497 539532 190527 539563
rect 190696 539556 190762 539572
rect 190896 539606 190962 539622
rect 190896 539572 190912 539606
rect 190946 539572 190962 539606
rect 190896 539556 190962 539572
rect 190714 539525 190744 539556
rect 190914 539525 190944 539556
rect 190714 538894 190744 538925
rect 190696 538878 190762 538894
rect 190696 538844 190712 538878
rect 190746 538844 190762 538878
rect 190696 538828 190762 538844
rect 189214 538494 189244 538525
rect 189441 538501 189471 538532
rect 189423 538495 189489 538501
rect 189537 538495 189567 538532
rect 189633 538501 189663 538532
rect 189615 538495 189681 538501
rect 189729 538495 189759 538532
rect 189825 538501 189855 538532
rect 189807 538495 189873 538501
rect 189921 538495 189951 538532
rect 190017 538501 190047 538532
rect 189999 538495 190065 538501
rect 190113 538495 190143 538532
rect 190209 538501 190239 538532
rect 190191 538495 190257 538501
rect 190305 538495 190335 538532
rect 190401 538501 190431 538532
rect 190497 538515 190527 538532
rect 190383 538495 190449 538501
rect 190494 538495 190528 538515
rect 189196 538478 189262 538494
rect 189196 538444 189212 538478
rect 189246 538444 189262 538478
rect 189196 538428 189262 538444
rect 189423 538485 190528 538495
rect 190914 538494 190944 538525
rect 189423 538451 189439 538485
rect 189473 538451 189631 538485
rect 189665 538451 189823 538485
rect 189857 538451 190015 538485
rect 190049 538451 190207 538485
rect 190241 538451 190399 538485
rect 190433 538451 190528 538485
rect 189423 538445 190528 538451
rect 190896 538478 190962 538494
rect 189423 538435 189489 538445
rect 189615 538435 189681 538445
rect 189807 538435 189873 538445
rect 189999 538435 190065 538445
rect 190191 538435 190257 538445
rect 190383 538435 190449 538445
rect 190896 538444 190912 538478
rect 190946 538444 190962 538478
rect 190896 538428 190962 538444
rect 161286 537706 161352 537722
rect 161286 537672 161302 537706
rect 161336 537672 161352 537706
rect 161490 537706 161556 537722
rect 161490 537705 161506 537706
rect 161286 537656 161352 537672
rect 161488 537672 161506 537705
rect 161540 537705 161556 537706
rect 161682 537706 161748 537722
rect 161682 537705 161698 537706
rect 161540 537672 161698 537705
rect 161732 537672 161748 537706
rect 161304 537625 161334 537656
rect 161488 537645 161748 537672
rect 161890 537715 161956 537722
rect 162082 537715 162148 537722
rect 161890 537706 162148 537715
rect 161890 537672 161906 537706
rect 161940 537672 162098 537706
rect 162132 537672 162148 537706
rect 161890 537656 162148 537672
rect 162306 537706 162372 537722
rect 162306 537672 162322 537706
rect 162356 537672 162372 537706
rect 162306 537656 162372 537672
rect 161908 537645 162138 537656
rect 161508 537625 161538 537645
rect 161604 537625 161634 537645
rect 161700 537625 161730 537645
rect 161908 537625 161938 537645
rect 162004 537625 162034 537645
rect 162100 537625 162130 537645
rect 162324 537625 162354 537656
rect 161304 536994 161334 537025
rect 161508 536999 161538 537025
rect 161604 536994 161634 537025
rect 161700 536999 161730 537025
rect 161908 536999 161938 537025
rect 162004 536994 162034 537025
rect 162100 536999 162130 537025
rect 162324 536994 162354 537025
rect 161286 536978 161352 536994
rect 161286 536944 161302 536978
rect 161336 536944 161352 536978
rect 161286 536928 161352 536944
rect 161586 536978 161652 536994
rect 161586 536944 161602 536978
rect 161636 536944 161652 536978
rect 161586 536928 161652 536944
rect 161986 536978 162052 536994
rect 161986 536944 162002 536978
rect 162036 536944 162052 536978
rect 161986 536928 162052 536944
rect 162306 536978 162372 536994
rect 162306 536944 162322 536978
rect 162356 536944 162372 536978
rect 162306 536928 162372 536944
rect 157794 536686 157994 536702
rect 157794 536652 157810 536686
rect 157978 536652 157994 536686
rect 157794 536605 157994 536652
rect 158172 536686 158372 536702
rect 158172 536652 158188 536686
rect 158356 536652 158372 536686
rect 158172 536605 158372 536652
rect 158430 536686 158630 536702
rect 158430 536652 158446 536686
rect 158614 536652 158630 536686
rect 158430 536605 158630 536652
rect 158688 536686 158888 536702
rect 158688 536652 158704 536686
rect 158872 536652 158888 536686
rect 158688 536605 158888 536652
rect 158946 536686 159146 536702
rect 158946 536652 158962 536686
rect 159130 536652 159146 536686
rect 158946 536605 159146 536652
rect 159204 536686 159404 536702
rect 159204 536652 159220 536686
rect 159388 536652 159404 536686
rect 159204 536605 159404 536652
rect 159462 536686 159662 536702
rect 159462 536652 159478 536686
rect 159646 536652 159662 536686
rect 159462 536605 159662 536652
rect 159720 536686 159920 536702
rect 159720 536652 159736 536686
rect 159904 536652 159920 536686
rect 159720 536605 159920 536652
rect 159978 536686 160178 536702
rect 159978 536652 159994 536686
rect 160162 536652 160178 536686
rect 159978 536605 160178 536652
rect 160236 536686 160436 536702
rect 160236 536652 160252 536686
rect 160420 536652 160436 536686
rect 160236 536605 160436 536652
rect 160494 536686 160694 536702
rect 160494 536652 160510 536686
rect 160678 536652 160694 536686
rect 160494 536605 160694 536652
rect 160878 536686 161078 536702
rect 160878 536652 160894 536686
rect 161062 536652 161078 536686
rect 160878 536605 161078 536652
rect 161136 536686 161336 536702
rect 161136 536652 161152 536686
rect 161320 536652 161336 536686
rect 161136 536605 161336 536652
rect 161394 536686 161594 536702
rect 161394 536652 161410 536686
rect 161578 536652 161594 536686
rect 161394 536605 161594 536652
rect 161776 536686 161976 536702
rect 161776 536652 161792 536686
rect 161960 536652 161976 536686
rect 161776 536605 161976 536652
rect 162034 536686 162234 536702
rect 162034 536652 162050 536686
rect 162218 536652 162234 536686
rect 162034 536605 162234 536652
rect 162414 536686 162614 536702
rect 162414 536652 162430 536686
rect 162598 536652 162614 536686
rect 162414 536605 162614 536652
rect 157794 535958 157994 536005
rect 157794 535924 157810 535958
rect 157978 535924 157994 535958
rect 157794 535908 157994 535924
rect 158172 535958 158372 536005
rect 158172 535924 158188 535958
rect 158356 535924 158372 535958
rect 158172 535908 158372 535924
rect 158430 535958 158630 536005
rect 158430 535924 158446 535958
rect 158614 535924 158630 535958
rect 158430 535908 158630 535924
rect 158688 535958 158888 536005
rect 158688 535924 158704 535958
rect 158872 535924 158888 535958
rect 158688 535908 158888 535924
rect 158946 535958 159146 536005
rect 158946 535924 158962 535958
rect 159130 535924 159146 535958
rect 158946 535908 159146 535924
rect 159204 535958 159404 536005
rect 159204 535924 159220 535958
rect 159388 535924 159404 535958
rect 159204 535908 159404 535924
rect 159462 535958 159662 536005
rect 159462 535924 159478 535958
rect 159646 535924 159662 535958
rect 159462 535908 159662 535924
rect 159720 535958 159920 536005
rect 159720 535924 159736 535958
rect 159904 535924 159920 535958
rect 159720 535908 159920 535924
rect 159978 535958 160178 536005
rect 159978 535924 159994 535958
rect 160162 535924 160178 535958
rect 159978 535908 160178 535924
rect 160236 535958 160436 536005
rect 160236 535924 160252 535958
rect 160420 535924 160436 535958
rect 160236 535908 160436 535924
rect 160494 535958 160694 536005
rect 160494 535924 160510 535958
rect 160678 535924 160694 535958
rect 160494 535908 160694 535924
rect 160878 535958 161078 536005
rect 160878 535924 160894 535958
rect 161062 535924 161078 535958
rect 160878 535908 161078 535924
rect 161136 535958 161336 536005
rect 161136 535924 161152 535958
rect 161320 535924 161336 535958
rect 161136 535908 161336 535924
rect 161394 535958 161594 536005
rect 161394 535924 161410 535958
rect 161578 535924 161594 535958
rect 161394 535908 161594 535924
rect 161776 535958 161976 536005
rect 161776 535924 161792 535958
rect 161960 535924 161976 535958
rect 161776 535908 161976 535924
rect 162034 535958 162234 536005
rect 162034 535924 162050 535958
rect 162218 535924 162234 535958
rect 162034 535908 162234 535924
rect 162414 535958 162614 536005
rect 162414 535924 162430 535958
rect 162598 535924 162614 535958
rect 162414 535908 162614 535924
rect 172287 530532 172405 530558
rect 172571 530532 172601 530558
rect 172657 530532 172687 530558
rect 172743 530532 172773 530558
rect 172829 530532 172859 530558
rect 172926 530532 172956 530558
rect 173115 530532 174061 530558
rect 174219 530532 174613 530558
rect 174963 530532 174993 530558
rect 175049 530532 175079 530558
rect 175135 530532 175165 530558
rect 175221 530532 175251 530558
rect 175318 530532 175348 530558
rect 175599 530532 175629 530558
rect 175807 530532 175837 530558
rect 175898 530532 175928 530558
rect 176047 530532 176077 530558
rect 176143 530532 176173 530558
rect 176252 530532 176282 530558
rect 176351 530532 176381 530558
rect 176483 530532 176513 530558
rect 176555 530532 176585 530558
rect 176721 530532 176751 530558
rect 176817 530532 176847 530558
rect 176912 530532 176942 530558
rect 177167 530532 177197 530558
rect 177251 530532 177281 530558
rect 177734 530532 177764 530558
rect 177829 530532 177929 530558
rect 178087 530532 178187 530558
rect 178241 530532 178271 530558
rect 178451 530532 178481 530558
rect 178539 530532 178569 530558
rect 178735 530532 178765 530558
rect 178821 530532 178851 530558
rect 178907 530532 178937 530558
rect 178993 530532 179023 530558
rect 179090 530532 179120 530558
rect 179280 530532 179310 530558
rect 179377 530532 179407 530558
rect 179463 530532 179493 530558
rect 179549 530532 179579 530558
rect 179635 530532 179665 530558
rect 180291 530532 180321 530558
rect 180400 530532 180430 530558
rect 180496 530532 180526 530558
rect 180621 530532 180651 530558
rect 180717 530532 180747 530558
rect 180885 530532 180915 530558
rect 181257 530532 181287 530558
rect 181425 530532 181455 530558
rect 181521 530532 181551 530558
rect 181646 530532 181676 530558
rect 181742 530532 181772 530558
rect 181851 530532 181881 530558
rect 182040 530532 182070 530558
rect 182137 530532 182167 530558
rect 182223 530532 182253 530558
rect 182309 530532 182339 530558
rect 182395 530532 182425 530558
rect 182683 530532 182893 530558
rect 183144 530532 183174 530558
rect 183241 530532 183271 530558
rect 183327 530532 183357 530558
rect 183413 530532 183443 530558
rect 183499 530532 183529 530558
rect 183695 530532 184641 530558
rect 184799 530532 185009 530558
rect 185260 530532 185290 530558
rect 185357 530532 185387 530558
rect 185443 530532 185473 530558
rect 185529 530532 185559 530558
rect 185615 530532 185645 530558
rect 185811 530532 186757 530558
rect 172287 530396 172405 530422
rect 172367 530394 172405 530396
rect 172367 530378 172433 530394
rect 172259 530338 172325 530354
rect 172259 530304 172275 530338
rect 172309 530304 172325 530338
rect 172367 530344 172383 530378
rect 172417 530344 172433 530378
rect 172367 530328 172433 530344
rect 172571 530375 172601 530448
rect 172657 530375 172687 530448
rect 172743 530375 172773 530448
rect 172829 530375 172859 530448
rect 172926 530380 172956 530448
rect 173115 530396 174061 530422
rect 174219 530396 174613 530422
rect 172571 530369 172859 530375
rect 172571 530364 172860 530369
rect 172571 530342 172635 530364
rect 172572 530330 172635 530342
rect 172669 530330 172703 530364
rect 172737 530330 172771 530364
rect 172805 530330 172860 530364
rect 172259 530288 172325 530304
rect 172287 530286 172325 530288
rect 172572 530320 172860 530330
rect 172287 530256 172405 530286
rect 172572 530282 172602 530320
rect 172658 530282 172688 530320
rect 172744 530282 172774 530320
rect 172830 530282 172860 530320
rect 172907 530364 172967 530380
rect 172907 530330 172917 530364
rect 172951 530330 172967 530364
rect 173607 530374 174061 530396
rect 172907 530314 172967 530330
rect 173115 530338 173565 530354
rect 172926 530282 172956 530314
rect 173115 530304 173387 530338
rect 173421 530304 173565 530338
rect 173607 530340 173751 530374
rect 173785 530340 174061 530374
rect 174437 530374 174613 530396
rect 173607 530324 174061 530340
rect 174219 530338 174395 530354
rect 173115 530282 173565 530304
rect 174219 530304 174235 530338
rect 174269 530304 174345 530338
rect 174379 530304 174395 530338
rect 174437 530340 174453 530374
rect 174487 530340 174563 530374
rect 174597 530340 174613 530374
rect 174963 530375 174993 530448
rect 175049 530375 175079 530448
rect 175135 530375 175165 530448
rect 175221 530375 175251 530448
rect 175318 530380 175348 530448
rect 175599 530380 175629 530402
rect 174963 530369 175251 530375
rect 174963 530364 175252 530369
rect 174963 530342 175027 530364
rect 174437 530324 174613 530340
rect 174964 530330 175027 530342
rect 175061 530330 175095 530364
rect 175129 530330 175163 530364
rect 175197 530330 175252 530364
rect 174219 530282 174395 530304
rect 174964 530320 175252 530330
rect 174964 530282 174994 530320
rect 175050 530282 175080 530320
rect 175136 530282 175166 530320
rect 175222 530282 175252 530320
rect 175299 530364 175359 530380
rect 175299 530330 175309 530364
rect 175343 530330 175359 530364
rect 175299 530314 175359 530330
rect 175599 530364 175658 530380
rect 175599 530330 175614 530364
rect 175648 530330 175658 530364
rect 175599 530314 175658 530330
rect 175318 530282 175348 530314
rect 175599 530282 175629 530314
rect 173115 530256 174061 530282
rect 174219 530256 174613 530282
rect 175807 530280 175837 530448
rect 175898 530388 175928 530448
rect 176047 530416 176077 530448
rect 175975 530400 176077 530416
rect 175879 530372 175933 530388
rect 175879 530338 175889 530372
rect 175923 530338 175933 530372
rect 175975 530366 175985 530400
rect 176019 530386 176077 530400
rect 176143 530390 176173 530460
rect 176252 530438 176282 530460
rect 176019 530366 176036 530386
rect 175975 530350 176036 530366
rect 175879 530322 175933 530338
rect 175802 530264 175856 530280
rect 175802 530230 175812 530264
rect 175846 530230 175856 530264
rect 175802 530214 175856 530230
rect 175814 530166 175844 530214
rect 175898 530166 175928 530322
rect 176006 530166 176036 530350
rect 176119 530374 176173 530390
rect 176119 530340 176129 530374
rect 176163 530342 176173 530374
rect 176215 530422 176282 530438
rect 176215 530388 176225 530422
rect 176259 530388 176282 530422
rect 176483 530426 176513 530448
rect 176459 530410 176513 530426
rect 176215 530372 176282 530388
rect 176351 530378 176381 530404
rect 176351 530362 176417 530378
rect 176163 530340 176185 530342
rect 176119 530330 176185 530340
rect 176119 530324 176206 530330
rect 176143 530312 176206 530324
rect 176156 530300 176206 530312
rect 176080 530248 176134 530264
rect 176080 530214 176090 530248
rect 176124 530214 176134 530248
rect 176080 530198 176134 530214
rect 176090 530166 176120 530198
rect 176176 530166 176206 530300
rect 176351 530328 176373 530362
rect 176407 530328 176417 530362
rect 176459 530376 176469 530410
rect 176503 530376 176513 530410
rect 176459 530360 176513 530376
rect 176351 530312 176417 530328
rect 176351 530295 176381 530312
rect 176275 530265 176381 530295
rect 176275 530250 176305 530265
rect 176472 530166 176502 530360
rect 176555 530290 176585 530448
rect 176721 530426 176751 530460
rect 176817 530426 176847 530460
rect 176708 530416 176774 530426
rect 176708 530382 176724 530416
rect 176758 530382 176774 530416
rect 176708 530372 176774 530382
rect 176816 530410 176870 530426
rect 176816 530376 176826 530410
rect 176860 530376 176870 530410
rect 176816 530360 176870 530376
rect 176816 530330 176847 530360
rect 176709 530300 176847 530330
rect 176912 530319 176942 530448
rect 177167 530359 177197 530448
rect 177251 530433 177281 530448
rect 177251 530403 177314 530433
rect 177284 530380 177314 530403
rect 177734 530380 177764 530402
rect 177829 530380 177929 530448
rect 177284 530364 177338 530380
rect 177167 530349 177242 530359
rect 176912 530303 177029 530319
rect 176544 530274 176599 530290
rect 176544 530240 176555 530274
rect 176589 530240 176599 530274
rect 176544 530224 176599 530240
rect 176569 530166 176599 530224
rect 176709 530166 176739 530300
rect 176912 530283 176985 530303
rect 176900 530269 176985 530283
rect 177019 530269 177029 530303
rect 176788 530248 176854 530258
rect 176788 530214 176804 530248
rect 176838 530214 176854 530248
rect 176788 530204 176854 530214
rect 176900 530253 177029 530269
rect 177167 530315 177192 530349
rect 177226 530315 177242 530349
rect 177167 530305 177242 530315
rect 177284 530330 177294 530364
rect 177328 530330 177338 530364
rect 177284 530314 177338 530330
rect 177733 530364 177787 530380
rect 177733 530330 177743 530364
rect 177777 530330 177787 530364
rect 177733 530314 177787 530330
rect 177829 530364 177983 530380
rect 177829 530330 177939 530364
rect 177973 530330 177983 530364
rect 177829 530314 177983 530330
rect 178087 530364 178187 530448
rect 178087 530330 178143 530364
rect 178177 530330 178187 530364
rect 176808 530166 176838 530204
rect 176900 530166 176930 530253
rect 177167 530216 177197 530305
rect 177284 530261 177314 530314
rect 177734 530282 177764 530314
rect 177251 530231 177314 530261
rect 177251 530216 177281 530231
rect 172287 530056 172405 530082
rect 172572 530056 172602 530082
rect 172658 530056 172688 530082
rect 172744 530056 172774 530082
rect 172830 530056 172860 530082
rect 172926 530056 172956 530082
rect 173115 530056 174061 530082
rect 174219 530056 174613 530082
rect 174964 530056 174994 530082
rect 175050 530056 175080 530082
rect 175136 530056 175166 530082
rect 175222 530056 175252 530082
rect 175318 530056 175348 530082
rect 175599 530056 175629 530082
rect 175814 530056 175844 530082
rect 175898 530056 175928 530082
rect 176006 530056 176036 530082
rect 176090 530056 176120 530082
rect 176176 530056 176206 530082
rect 176275 530056 176305 530082
rect 176472 530056 176502 530082
rect 176569 530056 176599 530082
rect 176709 530056 176739 530082
rect 176808 530056 176838 530082
rect 176900 530056 176930 530082
rect 177167 530062 177197 530088
rect 177251 530062 177281 530088
rect 177829 530166 177929 530314
rect 178087 530166 178187 530330
rect 178241 530380 178271 530448
rect 178241 530364 178301 530380
rect 178451 530367 178481 530428
rect 178539 530413 178569 530428
rect 178539 530389 178575 530413
rect 178545 530380 178575 530389
rect 178241 530330 178257 530364
rect 178291 530330 178301 530364
rect 178241 530314 178301 530330
rect 178447 530351 178501 530367
rect 178447 530317 178457 530351
rect 178491 530317 178501 530351
rect 178241 530166 178271 530314
rect 178447 530301 178501 530317
rect 178545 530364 178621 530380
rect 178545 530330 178577 530364
rect 178611 530330 178621 530364
rect 178735 530375 178765 530448
rect 178821 530375 178851 530448
rect 178907 530375 178937 530448
rect 178993 530375 179023 530448
rect 179090 530380 179120 530448
rect 179280 530380 179310 530448
rect 178735 530369 179023 530375
rect 178735 530364 179024 530369
rect 178735 530342 178799 530364
rect 178545 530314 178621 530330
rect 178736 530330 178799 530342
rect 178833 530330 178867 530364
rect 178901 530330 178935 530364
rect 178969 530330 179024 530364
rect 178736 530320 179024 530330
rect 178451 530240 178481 530301
rect 178545 530279 178575 530314
rect 178736 530282 178766 530320
rect 178822 530282 178852 530320
rect 178908 530282 178938 530320
rect 178994 530282 179024 530320
rect 179071 530364 179131 530380
rect 179071 530330 179081 530364
rect 179115 530330 179131 530364
rect 179071 530314 179131 530330
rect 179269 530364 179329 530380
rect 179377 530375 179407 530448
rect 179463 530375 179493 530448
rect 179549 530375 179579 530448
rect 179635 530375 179665 530448
rect 180291 530380 180321 530402
rect 180400 530380 180430 530448
rect 180496 530416 180526 530448
rect 180621 530416 180651 530448
rect 180496 530400 180579 530416
rect 179377 530369 179665 530375
rect 179269 530330 179285 530364
rect 179319 530330 179329 530364
rect 179269 530314 179329 530330
rect 179376 530364 179665 530369
rect 179376 530330 179431 530364
rect 179465 530330 179499 530364
rect 179533 530330 179567 530364
rect 179601 530342 179665 530364
rect 180288 530364 180342 530380
rect 179601 530330 179664 530342
rect 179376 530320 179664 530330
rect 179090 530282 179120 530314
rect 179280 530282 179310 530314
rect 179376 530282 179406 530320
rect 179462 530282 179492 530320
rect 179548 530282 179578 530320
rect 179634 530282 179664 530320
rect 180288 530330 180298 530364
rect 180332 530330 180342 530364
rect 180288 530314 180342 530330
rect 180384 530364 180438 530380
rect 180384 530330 180394 530364
rect 180428 530330 180438 530364
rect 180496 530366 180535 530400
rect 180569 530366 180579 530400
rect 180496 530350 180579 530366
rect 180621 530400 180675 530416
rect 180621 530366 180631 530400
rect 180665 530366 180675 530400
rect 180717 530410 180747 530448
rect 180717 530400 180843 530410
rect 180717 530380 180793 530400
rect 180621 530350 180675 530366
rect 180777 530366 180793 530380
rect 180827 530366 180843 530400
rect 180777 530356 180843 530366
rect 180384 530314 180438 530330
rect 180291 530282 180321 530314
rect 178539 530255 178575 530279
rect 178539 530240 178569 530255
rect 180400 530205 180430 530314
rect 180621 530250 180651 530350
rect 180503 530220 180651 530250
rect 180693 530287 180747 530303
rect 180693 530253 180703 530287
rect 180737 530253 180747 530287
rect 180693 530237 180747 530253
rect 180503 530205 180533 530220
rect 180717 530205 180747 530237
rect 180789 530205 180819 530356
rect 180885 530303 180915 530448
rect 180861 530287 180915 530303
rect 180861 530253 180871 530287
rect 180905 530253 180915 530287
rect 180861 530237 180915 530253
rect 180885 530205 180915 530237
rect 181257 530303 181287 530448
rect 181425 530410 181455 530448
rect 181521 530416 181551 530448
rect 181646 530416 181676 530448
rect 181329 530400 181455 530410
rect 181329 530366 181345 530400
rect 181379 530380 181455 530400
rect 181497 530400 181551 530416
rect 181379 530366 181395 530380
rect 181329 530356 181395 530366
rect 181497 530366 181507 530400
rect 181541 530366 181551 530400
rect 181257 530287 181311 530303
rect 181257 530253 181267 530287
rect 181301 530253 181311 530287
rect 181257 530237 181311 530253
rect 181257 530205 181287 530237
rect 181353 530205 181383 530356
rect 181497 530350 181551 530366
rect 181593 530400 181676 530416
rect 181593 530366 181603 530400
rect 181637 530366 181676 530400
rect 181742 530380 181772 530448
rect 181851 530380 181881 530402
rect 182040 530380 182070 530448
rect 181593 530350 181676 530366
rect 181734 530364 181788 530380
rect 181425 530287 181479 530303
rect 181425 530253 181435 530287
rect 181469 530253 181479 530287
rect 181425 530237 181479 530253
rect 181521 530250 181551 530350
rect 181734 530330 181744 530364
rect 181778 530330 181788 530364
rect 181734 530314 181788 530330
rect 181830 530364 181884 530380
rect 181830 530330 181840 530364
rect 181874 530330 181884 530364
rect 181830 530314 181884 530330
rect 182029 530364 182089 530380
rect 182137 530375 182167 530448
rect 182223 530375 182253 530448
rect 182309 530375 182339 530448
rect 182395 530375 182425 530448
rect 182683 530396 182893 530422
rect 182137 530369 182425 530375
rect 182029 530330 182045 530364
rect 182079 530330 182089 530364
rect 182029 530314 182089 530330
rect 182136 530364 182425 530369
rect 182136 530330 182191 530364
rect 182225 530330 182259 530364
rect 182293 530330 182327 530364
rect 182361 530342 182425 530364
rect 182809 530390 182893 530396
rect 182809 530374 182951 530390
rect 183144 530380 183174 530448
rect 182361 530330 182424 530342
rect 182136 530320 182424 530330
rect 181425 530205 181455 530237
rect 181521 530220 181669 530250
rect 181639 530205 181669 530220
rect 181742 530205 181772 530314
rect 181851 530282 181881 530314
rect 182040 530282 182070 530314
rect 182136 530282 182166 530320
rect 182222 530282 182252 530320
rect 182308 530282 182338 530320
rect 182394 530282 182424 530320
rect 182625 530338 182767 530354
rect 182625 530304 182641 530338
rect 182675 530304 182767 530338
rect 182809 530340 182901 530374
rect 182935 530340 182951 530374
rect 182809 530324 182951 530340
rect 183133 530364 183193 530380
rect 183241 530375 183271 530448
rect 183327 530375 183357 530448
rect 183413 530375 183443 530448
rect 183499 530375 183529 530448
rect 183695 530396 184641 530422
rect 184799 530396 185009 530422
rect 183241 530369 183529 530375
rect 183133 530330 183149 530364
rect 183183 530330 183193 530364
rect 183133 530314 183193 530330
rect 183240 530364 183529 530369
rect 183240 530330 183295 530364
rect 183329 530330 183363 530364
rect 183397 530330 183431 530364
rect 183465 530342 183529 530364
rect 184187 530374 184641 530396
rect 183465 530330 183528 530342
rect 183240 530320 183528 530330
rect 182625 530288 182767 530304
rect 182683 530282 182767 530288
rect 183144 530282 183174 530314
rect 183240 530282 183270 530320
rect 183326 530282 183356 530320
rect 183412 530282 183442 530320
rect 183498 530282 183528 530320
rect 183695 530338 184145 530354
rect 183695 530304 183967 530338
rect 184001 530304 184145 530338
rect 184187 530340 184331 530374
rect 184365 530340 184641 530374
rect 184925 530390 185009 530396
rect 184925 530374 185067 530390
rect 185260 530380 185290 530448
rect 184187 530324 184641 530340
rect 184741 530338 184883 530354
rect 183695 530282 184145 530304
rect 184741 530304 184757 530338
rect 184791 530304 184883 530338
rect 184925 530340 185017 530374
rect 185051 530340 185067 530374
rect 184925 530324 185067 530340
rect 185249 530364 185309 530380
rect 185357 530375 185387 530448
rect 185443 530375 185473 530448
rect 185529 530375 185559 530448
rect 185615 530375 185645 530448
rect 186949 530528 187045 530558
rect 186949 530494 186999 530528
rect 187033 530494 187045 530528
rect 186949 530460 187045 530494
rect 186949 530426 186999 530460
rect 187033 530426 187045 530460
rect 185811 530396 186757 530422
rect 185357 530369 185645 530375
rect 185249 530330 185265 530364
rect 185299 530330 185309 530364
rect 185249 530314 185309 530330
rect 185356 530364 185645 530369
rect 185356 530330 185411 530364
rect 185445 530330 185479 530364
rect 185513 530330 185547 530364
rect 185581 530342 185645 530364
rect 186303 530374 186757 530396
rect 185581 530330 185644 530342
rect 185356 530320 185644 530330
rect 184741 530288 184883 530304
rect 184799 530282 184883 530288
rect 185260 530282 185290 530314
rect 185356 530282 185386 530320
rect 185442 530282 185472 530320
rect 185528 530282 185558 530320
rect 185614 530282 185644 530320
rect 185811 530338 186261 530354
rect 185811 530304 186083 530338
rect 186117 530304 186261 530338
rect 186303 530340 186447 530374
rect 186481 530340 186757 530374
rect 186303 530324 186757 530340
rect 186949 530347 187045 530426
rect 185811 530282 186261 530304
rect 180400 530095 180430 530121
rect 180503 530095 180533 530121
rect 180717 530095 180747 530121
rect 180789 530095 180819 530121
rect 180885 530095 180915 530121
rect 181257 530095 181287 530121
rect 181353 530095 181383 530121
rect 181425 530095 181455 530121
rect 181639 530095 181669 530121
rect 181742 530095 181772 530121
rect 182683 530256 182893 530282
rect 183695 530256 184641 530282
rect 184799 530256 185009 530282
rect 185811 530256 186757 530282
rect 186949 530197 187045 530338
rect 186949 530163 186999 530197
rect 187033 530163 187045 530197
rect 186949 530129 187045 530163
rect 186949 530095 186999 530129
rect 187033 530095 187045 530129
rect 177734 530056 177764 530082
rect 177829 530056 177929 530082
rect 178087 530056 178187 530082
rect 178241 530056 178271 530082
rect 178451 530056 178481 530082
rect 178539 530056 178569 530082
rect 178736 530056 178766 530082
rect 178822 530056 178852 530082
rect 178908 530056 178938 530082
rect 178994 530056 179024 530082
rect 179090 530056 179120 530082
rect 179280 530056 179310 530082
rect 179376 530056 179406 530082
rect 179462 530056 179492 530082
rect 179548 530056 179578 530082
rect 179634 530056 179664 530082
rect 180291 530056 180321 530082
rect 181851 530056 181881 530082
rect 182040 530056 182070 530082
rect 182136 530056 182166 530082
rect 182222 530056 182252 530082
rect 182308 530056 182338 530082
rect 182394 530056 182424 530082
rect 182683 530056 182893 530082
rect 183144 530056 183174 530082
rect 183240 530056 183270 530082
rect 183326 530056 183356 530082
rect 183412 530056 183442 530082
rect 183498 530056 183528 530082
rect 183695 530056 184641 530082
rect 184799 530056 185009 530082
rect 185260 530056 185290 530082
rect 185356 530056 185386 530082
rect 185442 530056 185472 530082
rect 185528 530056 185558 530082
rect 185614 530056 185644 530082
rect 185811 530056 186757 530082
rect 186949 530056 187045 530095
rect 187087 530532 187183 530558
rect 187283 530532 187401 530558
rect 187087 530498 187099 530532
rect 187133 530498 187183 530532
rect 187087 530464 187183 530498
rect 187087 530430 187099 530464
rect 187133 530430 187183 530464
rect 187087 530347 187183 530430
rect 187283 530396 187401 530422
rect 187283 530394 187321 530396
rect 187087 530197 187183 530338
rect 187255 530378 187321 530394
rect 187255 530344 187271 530378
rect 187305 530344 187321 530378
rect 187255 530328 187321 530344
rect 187363 530338 187429 530354
rect 187363 530304 187379 530338
rect 187413 530304 187429 530338
rect 187363 530288 187429 530304
rect 187363 530286 187401 530288
rect 187283 530256 187401 530286
rect 187087 530163 187099 530197
rect 187133 530163 187183 530197
rect 187087 530129 187183 530163
rect 187087 530095 187099 530129
rect 187133 530095 187183 530129
rect 187087 530056 187183 530095
rect 187283 530056 187401 530082
rect 172287 529988 172405 530014
rect 172563 529988 173509 530014
rect 173667 529988 174613 530014
rect 174885 529988 174915 530014
rect 174969 529988 175069 530014
rect 175227 529988 175327 530014
rect 175392 529988 175422 530014
rect 172287 529784 172405 529814
rect 172563 529788 173509 529814
rect 173667 529788 174613 529814
rect 172287 529782 172325 529784
rect 172259 529766 172325 529782
rect 172259 529732 172275 529766
rect 172309 529732 172325 529766
rect 172563 529766 173013 529788
rect 172259 529716 172325 529732
rect 172367 529726 172433 529742
rect 172367 529692 172383 529726
rect 172417 529692 172433 529726
rect 172563 529732 172835 529766
rect 172869 529732 173013 529766
rect 173667 529766 174117 529788
rect 172563 529716 173013 529732
rect 173055 529730 173509 529746
rect 172367 529676 172433 529692
rect 173055 529696 173199 529730
rect 173233 529696 173509 529730
rect 173667 529732 173939 529766
rect 173973 529732 174117 529766
rect 174885 529756 174915 529904
rect 173667 529716 174117 529732
rect 174159 529730 174613 529746
rect 172367 529674 172405 529676
rect 173055 529674 173509 529696
rect 174159 529696 174303 529730
rect 174337 529696 174613 529730
rect 174159 529674 174613 529696
rect 174855 529740 174915 529756
rect 174855 529706 174865 529740
rect 174899 529706 174915 529740
rect 174855 529690 174915 529706
rect 172287 529648 172405 529674
rect 172563 529648 173509 529674
rect 173667 529648 174613 529674
rect 174885 529622 174915 529690
rect 174969 529740 175069 529904
rect 175227 529756 175327 529904
rect 175599 529982 175629 530008
rect 175683 529982 175713 530008
rect 175950 529988 175980 530014
rect 176042 529988 176072 530014
rect 176141 529988 176171 530014
rect 176281 529988 176311 530014
rect 176378 529988 176408 530014
rect 176575 529988 176605 530014
rect 176674 529988 176704 530014
rect 176760 529988 176790 530014
rect 176844 529988 176874 530014
rect 176952 529988 176982 530014
rect 177036 529988 177066 530014
rect 177251 529988 177281 530014
rect 178263 529988 178293 530014
rect 178451 529988 178481 530014
rect 178666 529988 178696 530014
rect 178750 529988 178780 530014
rect 178858 529988 178888 530014
rect 178942 529988 178972 530014
rect 179028 529988 179058 530014
rect 179127 529988 179157 530014
rect 179324 529988 179354 530014
rect 179421 529988 179451 530014
rect 179561 529988 179591 530014
rect 179660 529988 179690 530014
rect 179752 529988 179782 530014
rect 175599 529839 175629 529854
rect 175566 529809 175629 529839
rect 175392 529756 175422 529788
rect 175566 529756 175596 529809
rect 175683 529765 175713 529854
rect 175950 529817 175980 529904
rect 176042 529866 176072 529904
rect 174969 529706 174979 529740
rect 175013 529706 175069 529740
rect 174969 529622 175069 529706
rect 175173 529740 175327 529756
rect 175173 529706 175183 529740
rect 175217 529706 175327 529740
rect 175173 529690 175327 529706
rect 175369 529740 175423 529756
rect 175369 529706 175379 529740
rect 175413 529706 175423 529740
rect 175369 529690 175423 529706
rect 175542 529740 175596 529756
rect 175542 529706 175552 529740
rect 175586 529706 175596 529740
rect 175638 529755 175713 529765
rect 175638 529721 175654 529755
rect 175688 529721 175713 529755
rect 175851 529801 175980 529817
rect 176026 529856 176092 529866
rect 176026 529822 176042 529856
rect 176076 529822 176092 529856
rect 176026 529812 176092 529822
rect 175851 529767 175861 529801
rect 175895 529787 175980 529801
rect 175895 529767 175968 529787
rect 176141 529770 176171 529904
rect 176281 529846 176311 529904
rect 176281 529830 176336 529846
rect 176281 529796 176291 529830
rect 176325 529796 176336 529830
rect 176281 529780 176336 529796
rect 175851 529751 175968 529767
rect 175638 529711 175713 529721
rect 175542 529690 175596 529706
rect 175227 529622 175327 529690
rect 175392 529668 175422 529690
rect 175566 529667 175596 529690
rect 175566 529637 175629 529667
rect 175599 529622 175629 529637
rect 175683 529622 175713 529711
rect 175938 529622 175968 529751
rect 176033 529740 176171 529770
rect 176033 529710 176064 529740
rect 176010 529694 176064 529710
rect 176010 529660 176020 529694
rect 176054 529660 176064 529694
rect 176010 529644 176064 529660
rect 176106 529688 176172 529698
rect 176106 529654 176122 529688
rect 176156 529654 176172 529688
rect 176106 529644 176172 529654
rect 176033 529610 176063 529644
rect 176129 529610 176159 529644
rect 176295 529622 176325 529780
rect 176378 529710 176408 529904
rect 176575 529805 176605 529820
rect 176499 529775 176605 529805
rect 176499 529758 176529 529775
rect 176463 529742 176529 529758
rect 176367 529694 176421 529710
rect 176367 529660 176377 529694
rect 176411 529660 176421 529694
rect 176463 529708 176473 529742
rect 176507 529708 176529 529742
rect 176674 529770 176704 529904
rect 176760 529872 176790 529904
rect 176746 529856 176800 529872
rect 176746 529822 176756 529856
rect 176790 529822 176800 529856
rect 176746 529806 176800 529822
rect 176674 529758 176724 529770
rect 176674 529746 176737 529758
rect 176674 529740 176761 529746
rect 176695 529730 176761 529740
rect 176695 529728 176717 529730
rect 176463 529692 176529 529708
rect 176499 529666 176529 529692
rect 176598 529682 176665 529698
rect 176367 529644 176421 529660
rect 176367 529622 176397 529644
rect 176598 529648 176621 529682
rect 176655 529648 176665 529682
rect 176598 529632 176665 529648
rect 176707 529696 176717 529728
rect 176751 529696 176761 529730
rect 176707 529680 176761 529696
rect 176844 529720 176874 529904
rect 176952 529748 176982 529904
rect 177036 529856 177066 529904
rect 177024 529840 177078 529856
rect 177024 529806 177034 529840
rect 177068 529806 177078 529840
rect 177024 529790 177078 529806
rect 176947 529732 177001 529748
rect 176844 529704 176905 529720
rect 176844 529684 176861 529704
rect 176598 529610 176628 529632
rect 176707 529610 176737 529680
rect 176803 529670 176861 529684
rect 176895 529670 176905 529704
rect 176947 529698 176957 529732
rect 176991 529698 177001 529732
rect 176947 529682 177001 529698
rect 176803 529654 176905 529670
rect 176803 529622 176833 529654
rect 176952 529622 176982 529682
rect 177043 529622 177073 529790
rect 177669 529949 177699 529975
rect 177765 529949 177795 529975
rect 177837 529949 177867 529975
rect 178051 529949 178081 529975
rect 178154 529949 178184 529975
rect 177669 529833 177699 529865
rect 177669 529817 177723 529833
rect 177251 529756 177281 529788
rect 177222 529740 177281 529756
rect 177222 529706 177232 529740
rect 177266 529706 177281 529740
rect 177222 529690 177281 529706
rect 177251 529668 177281 529690
rect 177669 529783 177679 529817
rect 177713 529783 177723 529817
rect 177669 529767 177723 529783
rect 177669 529622 177699 529767
rect 177765 529714 177795 529865
rect 177837 529833 177867 529865
rect 178051 529850 178081 529865
rect 177837 529817 177891 529833
rect 177837 529783 177847 529817
rect 177881 529783 177891 529817
rect 177837 529767 177891 529783
rect 177933 529820 178081 529850
rect 177933 529720 177963 529820
rect 178154 529756 178184 529865
rect 178666 529856 178696 529904
rect 178654 529840 178708 529856
rect 178654 529806 178664 529840
rect 178698 529806 178708 529840
rect 178654 529790 178708 529806
rect 178263 529756 178293 529788
rect 178451 529756 178481 529788
rect 178146 529740 178200 529756
rect 177741 529704 177807 529714
rect 177741 529670 177757 529704
rect 177791 529690 177807 529704
rect 177909 529704 177963 529720
rect 177791 529670 177867 529690
rect 177741 529660 177867 529670
rect 177837 529622 177867 529660
rect 177909 529670 177919 529704
rect 177953 529670 177963 529704
rect 177909 529654 177963 529670
rect 178005 529704 178088 529720
rect 178005 529670 178015 529704
rect 178049 529670 178088 529704
rect 178146 529706 178156 529740
rect 178190 529706 178200 529740
rect 178146 529690 178200 529706
rect 178242 529740 178296 529756
rect 178242 529706 178252 529740
rect 178286 529706 178296 529740
rect 178242 529690 178296 529706
rect 178451 529740 178510 529756
rect 178451 529706 178466 529740
rect 178500 529706 178510 529740
rect 178451 529690 178510 529706
rect 178005 529654 178088 529670
rect 177933 529622 177963 529654
rect 178058 529622 178088 529654
rect 178154 529622 178184 529690
rect 178263 529668 178293 529690
rect 178451 529668 178481 529690
rect 178659 529622 178689 529790
rect 178750 529748 178780 529904
rect 178731 529732 178785 529748
rect 178731 529698 178741 529732
rect 178775 529698 178785 529732
rect 178858 529720 178888 529904
rect 178942 529872 178972 529904
rect 178932 529856 178986 529872
rect 178932 529822 178942 529856
rect 178976 529822 178986 529856
rect 178932 529806 178986 529822
rect 179028 529770 179058 529904
rect 180019 529982 180049 530008
rect 180103 529982 180133 530008
rect 180291 529982 180321 530008
rect 180375 529982 180405 530008
rect 180642 529988 180672 530014
rect 180734 529988 180764 530014
rect 180833 529988 180863 530014
rect 180973 529988 181003 530014
rect 181070 529988 181100 530014
rect 181267 529988 181297 530014
rect 181366 529988 181396 530014
rect 181452 529988 181482 530014
rect 181536 529988 181566 530014
rect 181644 529988 181674 530014
rect 181728 529988 181758 530014
rect 181943 529988 181973 530014
rect 182131 529988 182341 530014
rect 182702 529988 182732 530014
rect 182797 529988 182897 530014
rect 183055 529988 183155 530014
rect 183209 529988 183239 530014
rect 183419 529988 184365 530014
rect 184523 529988 185469 530014
rect 185627 529988 186573 530014
rect 186731 529988 187125 530014
rect 187283 529988 187401 530014
rect 179127 529805 179157 529820
rect 179127 529775 179233 529805
rect 179008 529758 179058 529770
rect 178995 529746 179058 529758
rect 178731 529682 178785 529698
rect 178827 529704 178888 529720
rect 178750 529622 178780 529682
rect 178827 529670 178837 529704
rect 178871 529684 178888 529704
rect 178971 529740 179058 529746
rect 179203 529758 179233 529775
rect 179203 529742 179269 529758
rect 178971 529730 179037 529740
rect 178971 529696 178981 529730
rect 179015 529728 179037 529730
rect 179015 529696 179025 529728
rect 179203 529708 179225 529742
rect 179259 529708 179269 529742
rect 179324 529710 179354 529904
rect 179421 529846 179451 529904
rect 179396 529830 179451 529846
rect 179396 529796 179407 529830
rect 179441 529796 179451 529830
rect 179396 529780 179451 529796
rect 178871 529670 178929 529684
rect 178971 529680 179025 529696
rect 178827 529654 178929 529670
rect 178899 529622 178929 529654
rect 178995 529610 179025 529680
rect 179067 529682 179134 529698
rect 179067 529648 179077 529682
rect 179111 529648 179134 529682
rect 179203 529692 179269 529708
rect 179311 529694 179365 529710
rect 179203 529666 179233 529692
rect 179067 529632 179134 529648
rect 179104 529610 179134 529632
rect 179311 529660 179321 529694
rect 179355 529660 179365 529694
rect 179311 529644 179365 529660
rect 179335 529622 179365 529644
rect 179407 529622 179437 529780
rect 179561 529770 179591 529904
rect 179660 529866 179690 529904
rect 179640 529856 179706 529866
rect 179640 529822 179656 529856
rect 179690 529822 179706 529856
rect 179640 529812 179706 529822
rect 179752 529817 179782 529904
rect 179752 529801 179881 529817
rect 179752 529787 179837 529801
rect 179561 529740 179699 529770
rect 179668 529710 179699 529740
rect 179764 529767 179837 529787
rect 179871 529767 179881 529801
rect 179764 529751 179881 529767
rect 180019 529765 180049 529854
rect 180103 529839 180133 529854
rect 180291 529839 180321 529854
rect 180103 529809 180166 529839
rect 180019 529755 180094 529765
rect 179560 529688 179626 529698
rect 179560 529654 179576 529688
rect 179610 529654 179626 529688
rect 179560 529644 179626 529654
rect 179668 529694 179722 529710
rect 179668 529660 179678 529694
rect 179712 529660 179722 529694
rect 179668 529644 179722 529660
rect 179573 529610 179603 529644
rect 179669 529610 179699 529644
rect 179764 529622 179794 529751
rect 180019 529721 180044 529755
rect 180078 529721 180094 529755
rect 180019 529711 180094 529721
rect 180136 529756 180166 529809
rect 180258 529809 180321 529839
rect 180258 529756 180288 529809
rect 180375 529765 180405 529854
rect 180642 529817 180672 529904
rect 180734 529866 180764 529904
rect 180136 529740 180190 529756
rect 180019 529622 180049 529711
rect 180136 529706 180146 529740
rect 180180 529706 180190 529740
rect 180136 529690 180190 529706
rect 180234 529740 180288 529756
rect 180234 529706 180244 529740
rect 180278 529706 180288 529740
rect 180330 529755 180405 529765
rect 180330 529721 180346 529755
rect 180380 529721 180405 529755
rect 180543 529801 180672 529817
rect 180718 529856 180784 529866
rect 180718 529822 180734 529856
rect 180768 529822 180784 529856
rect 180718 529812 180784 529822
rect 180543 529767 180553 529801
rect 180587 529787 180672 529801
rect 180587 529767 180660 529787
rect 180833 529770 180863 529904
rect 180973 529846 181003 529904
rect 180973 529830 181028 529846
rect 180973 529796 180983 529830
rect 181017 529796 181028 529830
rect 180973 529780 181028 529796
rect 180543 529751 180660 529767
rect 180330 529711 180405 529721
rect 180234 529690 180288 529706
rect 180136 529667 180166 529690
rect 180103 529637 180166 529667
rect 180258 529667 180288 529690
rect 180258 529637 180321 529667
rect 180103 529622 180133 529637
rect 180291 529622 180321 529637
rect 180375 529622 180405 529711
rect 180630 529622 180660 529751
rect 180725 529740 180863 529770
rect 180725 529710 180756 529740
rect 180702 529694 180756 529710
rect 180702 529660 180712 529694
rect 180746 529660 180756 529694
rect 180702 529644 180756 529660
rect 180798 529688 180864 529698
rect 180798 529654 180814 529688
rect 180848 529654 180864 529688
rect 180798 529644 180864 529654
rect 180725 529610 180755 529644
rect 180821 529610 180851 529644
rect 180987 529622 181017 529780
rect 181070 529710 181100 529904
rect 181267 529805 181297 529820
rect 181191 529775 181297 529805
rect 181191 529758 181221 529775
rect 181155 529742 181221 529758
rect 181059 529694 181113 529710
rect 181059 529660 181069 529694
rect 181103 529660 181113 529694
rect 181155 529708 181165 529742
rect 181199 529708 181221 529742
rect 181366 529770 181396 529904
rect 181452 529872 181482 529904
rect 181438 529856 181492 529872
rect 181438 529822 181448 529856
rect 181482 529822 181492 529856
rect 181438 529806 181492 529822
rect 181366 529758 181416 529770
rect 181366 529746 181429 529758
rect 181366 529740 181453 529746
rect 181387 529730 181453 529740
rect 181387 529728 181409 529730
rect 181155 529692 181221 529708
rect 181191 529666 181221 529692
rect 181290 529682 181357 529698
rect 181059 529644 181113 529660
rect 181059 529622 181089 529644
rect 181290 529648 181313 529682
rect 181347 529648 181357 529682
rect 181290 529632 181357 529648
rect 181399 529696 181409 529728
rect 181443 529696 181453 529730
rect 181399 529680 181453 529696
rect 181536 529720 181566 529904
rect 181644 529748 181674 529904
rect 181728 529856 181758 529904
rect 181716 529840 181770 529856
rect 181716 529806 181726 529840
rect 181760 529806 181770 529840
rect 181716 529790 181770 529806
rect 181639 529732 181693 529748
rect 181536 529704 181597 529720
rect 181536 529684 181553 529704
rect 181290 529610 181320 529632
rect 181399 529610 181429 529680
rect 181495 529670 181553 529684
rect 181587 529670 181597 529704
rect 181639 529698 181649 529732
rect 181683 529698 181693 529732
rect 181639 529682 181693 529698
rect 181495 529654 181597 529670
rect 181495 529622 181525 529654
rect 181644 529622 181674 529682
rect 181735 529622 181765 529790
rect 182131 529788 182341 529814
rect 181943 529756 181973 529788
rect 182131 529782 182215 529788
rect 181914 529740 181973 529756
rect 181914 529706 181924 529740
rect 181958 529706 181973 529740
rect 182073 529766 182215 529782
rect 182073 529732 182089 529766
rect 182123 529732 182215 529766
rect 182702 529756 182732 529788
rect 182797 529756 182897 529904
rect 182073 529716 182215 529732
rect 182257 529730 182399 529746
rect 181914 529690 181973 529706
rect 181943 529668 181973 529690
rect 182257 529696 182349 529730
rect 182383 529696 182399 529730
rect 182257 529680 182399 529696
rect 182701 529740 182755 529756
rect 182701 529706 182711 529740
rect 182745 529706 182755 529740
rect 182701 529690 182755 529706
rect 182797 529740 182951 529756
rect 182797 529706 182907 529740
rect 182941 529706 182951 529740
rect 182797 529690 182951 529706
rect 183055 529740 183155 529904
rect 183055 529706 183111 529740
rect 183145 529706 183155 529740
rect 182257 529674 182341 529680
rect 182131 529648 182341 529674
rect 182702 529668 182732 529690
rect 182797 529622 182897 529690
rect 183055 529622 183155 529706
rect 183209 529756 183239 529904
rect 183419 529788 184365 529814
rect 184523 529788 185469 529814
rect 185627 529788 186573 529814
rect 186731 529788 187125 529814
rect 183419 529766 183869 529788
rect 183209 529740 183269 529756
rect 183209 529706 183225 529740
rect 183259 529706 183269 529740
rect 183419 529732 183691 529766
rect 183725 529732 183869 529766
rect 184523 529766 184973 529788
rect 183419 529716 183869 529732
rect 183911 529730 184365 529746
rect 183209 529690 183269 529706
rect 183911 529696 184055 529730
rect 184089 529696 184365 529730
rect 184523 529732 184795 529766
rect 184829 529732 184973 529766
rect 185627 529766 186077 529788
rect 184523 529716 184973 529732
rect 185015 529730 185469 529746
rect 183209 529622 183239 529690
rect 183911 529674 184365 529696
rect 185015 529696 185159 529730
rect 185193 529696 185469 529730
rect 185627 529732 185899 529766
rect 185933 529732 186077 529766
rect 186731 529766 186907 529788
rect 187283 529784 187401 529814
rect 185627 529716 186077 529732
rect 186119 529730 186573 529746
rect 185015 529674 185469 529696
rect 186119 529696 186263 529730
rect 186297 529696 186573 529730
rect 186731 529732 186747 529766
rect 186781 529732 186857 529766
rect 186891 529732 186907 529766
rect 187363 529782 187401 529784
rect 187363 529766 187429 529782
rect 186731 529716 186907 529732
rect 186949 529730 187125 529746
rect 186119 529674 186573 529696
rect 186949 529696 186965 529730
rect 186999 529696 187075 529730
rect 187109 529696 187125 529730
rect 186949 529674 187125 529696
rect 187255 529726 187321 529742
rect 187255 529692 187271 529726
rect 187305 529692 187321 529726
rect 187363 529732 187379 529766
rect 187413 529732 187429 529766
rect 187363 529716 187429 529732
rect 187255 529676 187321 529692
rect 183419 529648 184365 529674
rect 184523 529648 185469 529674
rect 185627 529648 186573 529674
rect 186731 529648 187125 529674
rect 187283 529674 187321 529676
rect 187283 529648 187401 529674
rect 172287 529512 172405 529538
rect 172563 529512 173509 529538
rect 173667 529512 174613 529538
rect 174885 529512 174915 529538
rect 174969 529512 175069 529538
rect 175227 529512 175327 529538
rect 175392 529512 175422 529538
rect 175599 529512 175629 529538
rect 175683 529512 175713 529538
rect 175938 529512 175968 529538
rect 176033 529512 176063 529538
rect 176129 529512 176159 529538
rect 176295 529512 176325 529538
rect 176367 529512 176397 529538
rect 176499 529512 176529 529538
rect 176598 529512 176628 529538
rect 176707 529512 176737 529538
rect 176803 529512 176833 529538
rect 176952 529512 176982 529538
rect 177043 529512 177073 529538
rect 177251 529512 177281 529538
rect 177669 529512 177699 529538
rect 177837 529512 177867 529538
rect 177933 529512 177963 529538
rect 178058 529512 178088 529538
rect 178154 529512 178184 529538
rect 178263 529512 178293 529538
rect 178451 529512 178481 529538
rect 178659 529512 178689 529538
rect 178750 529512 178780 529538
rect 178899 529512 178929 529538
rect 178995 529512 179025 529538
rect 179104 529512 179134 529538
rect 179203 529512 179233 529538
rect 179335 529512 179365 529538
rect 179407 529512 179437 529538
rect 179573 529512 179603 529538
rect 179669 529512 179699 529538
rect 179764 529512 179794 529538
rect 180019 529512 180049 529538
rect 180103 529512 180133 529538
rect 180291 529512 180321 529538
rect 180375 529512 180405 529538
rect 180630 529512 180660 529538
rect 180725 529512 180755 529538
rect 180821 529512 180851 529538
rect 180987 529512 181017 529538
rect 181059 529512 181089 529538
rect 181191 529512 181221 529538
rect 181290 529512 181320 529538
rect 181399 529512 181429 529538
rect 181495 529512 181525 529538
rect 181644 529512 181674 529538
rect 181735 529512 181765 529538
rect 181943 529512 181973 529538
rect 182131 529512 182341 529538
rect 182702 529512 182732 529538
rect 182797 529512 182897 529538
rect 183055 529512 183155 529538
rect 183209 529512 183239 529538
rect 183419 529512 184365 529538
rect 184523 529512 185469 529538
rect 185627 529512 186573 529538
rect 186731 529512 187125 529538
rect 187283 529512 187401 529538
rect 172287 529444 172405 529470
rect 172563 529444 173509 529470
rect 173667 529444 174613 529470
rect 175185 529444 175215 529470
rect 175353 529444 175383 529470
rect 175449 529444 175479 529470
rect 175574 529444 175604 529470
rect 175670 529444 175700 529470
rect 175779 529444 175809 529470
rect 175985 529444 176015 529470
rect 176071 529444 176101 529470
rect 176157 529444 176187 529470
rect 176243 529444 176273 529470
rect 176329 529444 176359 529470
rect 176415 529444 176445 529470
rect 176501 529444 176531 529470
rect 176587 529444 176617 529470
rect 176672 529444 176702 529470
rect 176758 529444 176788 529470
rect 176844 529444 176874 529470
rect 176930 529444 176960 529470
rect 177016 529444 177046 529470
rect 177102 529444 177132 529470
rect 177188 529444 177218 529470
rect 177274 529444 177304 529470
rect 177360 529444 177390 529470
rect 177446 529444 177476 529470
rect 177532 529444 177562 529470
rect 177618 529444 177648 529470
rect 177807 529444 177837 529470
rect 177891 529444 177921 529470
rect 178146 529444 178176 529470
rect 178241 529444 178271 529470
rect 178337 529444 178367 529470
rect 178503 529444 178533 529470
rect 178575 529444 178605 529470
rect 178707 529444 178737 529470
rect 178806 529444 178836 529470
rect 178915 529444 178945 529470
rect 179011 529444 179041 529470
rect 179160 529444 179190 529470
rect 179251 529444 179281 529470
rect 179459 529444 179489 529470
rect 179739 529444 179769 529470
rect 179827 529444 179857 529470
rect 180107 529444 180501 529470
rect 180752 529444 180782 529470
rect 180838 529444 180868 529470
rect 180924 529444 180954 529470
rect 181010 529444 181040 529470
rect 181096 529444 181126 529470
rect 181182 529444 181212 529470
rect 181268 529444 181298 529470
rect 181354 529444 181384 529470
rect 181440 529444 181470 529470
rect 181526 529444 181556 529470
rect 181612 529444 181642 529470
rect 181698 529444 181728 529470
rect 181783 529444 181813 529470
rect 181869 529444 181899 529470
rect 181955 529444 181985 529470
rect 182041 529444 182071 529470
rect 182127 529444 182157 529470
rect 182213 529444 182243 529470
rect 182299 529444 182329 529470
rect 182385 529444 182415 529470
rect 182591 529444 182621 529470
rect 182679 529444 182709 529470
rect 182867 529444 183813 529470
rect 183971 529444 184917 529470
rect 185259 529444 186205 529470
rect 186363 529444 186941 529470
rect 187283 529444 187401 529470
rect 172287 529308 172405 529334
rect 172563 529308 173509 529334
rect 173667 529308 174613 529334
rect 172367 529306 172405 529308
rect 172367 529290 172433 529306
rect 172259 529250 172325 529266
rect 172259 529216 172275 529250
rect 172309 529216 172325 529250
rect 172367 529256 172383 529290
rect 172417 529256 172433 529290
rect 173055 529286 173509 529308
rect 172367 529240 172433 529256
rect 172563 529250 173013 529266
rect 172259 529200 172325 529216
rect 172287 529198 172325 529200
rect 172563 529216 172835 529250
rect 172869 529216 173013 529250
rect 173055 529252 173199 529286
rect 173233 529252 173509 529286
rect 174159 529286 174613 529308
rect 173055 529236 173509 529252
rect 173667 529250 174117 529266
rect 172287 529168 172405 529198
rect 172563 529194 173013 529216
rect 173667 529216 173939 529250
rect 173973 529216 174117 529250
rect 174159 529252 174303 529286
rect 174337 529252 174613 529286
rect 174159 529236 174613 529252
rect 173667 529194 174117 529216
rect 175185 529215 175215 529360
rect 175353 529322 175383 529360
rect 175449 529328 175479 529360
rect 175574 529328 175604 529360
rect 175257 529312 175383 529322
rect 175257 529278 175273 529312
rect 175307 529292 175383 529312
rect 175425 529312 175479 529328
rect 175307 529278 175323 529292
rect 175257 529268 175323 529278
rect 175425 529278 175435 529312
rect 175469 529278 175479 529312
rect 175185 529199 175239 529215
rect 172563 529168 173509 529194
rect 173667 529168 174613 529194
rect 175185 529165 175195 529199
rect 175229 529165 175239 529199
rect 175185 529149 175239 529165
rect 175185 529117 175215 529149
rect 175281 529117 175311 529268
rect 175425 529262 175479 529278
rect 175521 529312 175604 529328
rect 175521 529278 175531 529312
rect 175565 529278 175604 529312
rect 175670 529292 175700 529360
rect 175779 529292 175809 529314
rect 175985 529301 176015 529360
rect 176071 529301 176101 529360
rect 176157 529301 176187 529360
rect 176243 529301 176273 529360
rect 176329 529301 176359 529360
rect 176415 529301 176445 529360
rect 176501 529301 176531 529360
rect 176587 529301 176617 529360
rect 176672 529301 176702 529360
rect 176758 529301 176788 529360
rect 176844 529301 176874 529360
rect 176930 529301 176960 529360
rect 177016 529301 177046 529360
rect 177102 529301 177132 529360
rect 177188 529301 177218 529360
rect 177274 529301 177304 529360
rect 175521 529262 175604 529278
rect 175662 529276 175716 529292
rect 175353 529199 175407 529215
rect 175353 529165 175363 529199
rect 175397 529165 175407 529199
rect 175353 529149 175407 529165
rect 175449 529162 175479 529262
rect 175662 529242 175672 529276
rect 175706 529242 175716 529276
rect 175662 529226 175716 529242
rect 175758 529276 175812 529292
rect 175758 529242 175768 529276
rect 175802 529242 175812 529276
rect 175758 529226 175812 529242
rect 175985 529276 177304 529301
rect 175985 529242 176210 529276
rect 176244 529242 176278 529276
rect 176312 529242 176346 529276
rect 176380 529242 176414 529276
rect 176448 529242 176482 529276
rect 176516 529242 176550 529276
rect 176584 529242 176618 529276
rect 176652 529242 176686 529276
rect 176720 529242 176754 529276
rect 176788 529242 176822 529276
rect 176856 529242 176890 529276
rect 176924 529242 176958 529276
rect 176992 529242 177026 529276
rect 177060 529242 177094 529276
rect 177128 529242 177162 529276
rect 177196 529242 177230 529276
rect 177264 529242 177304 529276
rect 175985 529226 177304 529242
rect 175353 529117 175383 529149
rect 175449 529132 175597 529162
rect 175567 529117 175597 529132
rect 175670 529117 175700 529226
rect 175779 529194 175809 529226
rect 175985 529194 176015 529226
rect 176071 529194 176101 529226
rect 176157 529194 176187 529226
rect 176243 529194 176273 529226
rect 176329 529194 176359 529226
rect 176415 529194 176445 529226
rect 176501 529194 176531 529226
rect 176587 529194 176617 529226
rect 176672 529194 176702 529226
rect 176758 529194 176788 529226
rect 176844 529194 176874 529226
rect 176930 529194 176960 529226
rect 177016 529194 177046 529226
rect 177102 529194 177132 529226
rect 177188 529194 177218 529226
rect 177274 529194 177304 529226
rect 177360 529311 177390 529360
rect 177446 529311 177476 529360
rect 177532 529311 177562 529360
rect 177618 529311 177648 529360
rect 177807 529345 177837 529360
rect 177774 529315 177837 529345
rect 177360 529276 177707 529311
rect 177774 529292 177804 529315
rect 177360 529242 177657 529276
rect 177691 529242 177707 529276
rect 177360 529209 177707 529242
rect 177750 529276 177804 529292
rect 177750 529242 177760 529276
rect 177794 529242 177804 529276
rect 177891 529271 177921 529360
rect 177750 529226 177804 529242
rect 177360 529194 177390 529209
rect 177446 529194 177476 529209
rect 177532 529194 177562 529209
rect 177618 529194 177648 529209
rect 175185 529007 175215 529033
rect 175281 529007 175311 529033
rect 175353 529007 175383 529033
rect 175567 529007 175597 529033
rect 175670 529007 175700 529033
rect 177774 529173 177804 529226
rect 177846 529261 177921 529271
rect 177846 529227 177862 529261
rect 177896 529227 177921 529261
rect 178146 529231 178176 529360
rect 178241 529338 178271 529372
rect 178337 529338 178367 529372
rect 178218 529322 178272 529338
rect 178218 529288 178228 529322
rect 178262 529288 178272 529322
rect 178218 529272 178272 529288
rect 178314 529328 178380 529338
rect 178314 529294 178330 529328
rect 178364 529294 178380 529328
rect 178314 529284 178380 529294
rect 177846 529217 177921 529227
rect 177774 529143 177837 529173
rect 177807 529128 177837 529143
rect 177891 529128 177921 529217
rect 178059 529215 178176 529231
rect 178059 529181 178069 529215
rect 178103 529195 178176 529215
rect 178241 529242 178272 529272
rect 178241 529212 178379 529242
rect 178103 529181 178188 529195
rect 178059 529165 178188 529181
rect 178158 529078 178188 529165
rect 178234 529160 178300 529170
rect 178234 529126 178250 529160
rect 178284 529126 178300 529160
rect 178234 529116 178300 529126
rect 178250 529078 178280 529116
rect 178349 529078 178379 529212
rect 178503 529202 178533 529360
rect 178575 529338 178605 529360
rect 178575 529322 178629 529338
rect 178575 529288 178585 529322
rect 178619 529288 178629 529322
rect 178806 529350 178836 529372
rect 178806 529334 178873 529350
rect 178707 529290 178737 529316
rect 178575 529272 178629 529288
rect 178671 529274 178737 529290
rect 178806 529300 178829 529334
rect 178863 529300 178873 529334
rect 178806 529284 178873 529300
rect 178915 529302 178945 529372
rect 179011 529328 179041 529360
rect 179011 529312 179113 529328
rect 178915 529286 178969 529302
rect 179011 529298 179069 529312
rect 178489 529186 178544 529202
rect 178489 529152 178499 529186
rect 178533 529152 178544 529186
rect 178489 529136 178544 529152
rect 178489 529078 178519 529136
rect 178586 529078 178616 529272
rect 178671 529240 178681 529274
rect 178715 529240 178737 529274
rect 178915 529254 178925 529286
rect 178903 529252 178925 529254
rect 178959 529252 178969 529286
rect 178903 529242 178969 529252
rect 178671 529224 178737 529240
rect 178707 529207 178737 529224
rect 178882 529236 178969 529242
rect 179052 529278 179069 529298
rect 179103 529278 179113 529312
rect 179160 529300 179190 529360
rect 179052 529262 179113 529278
rect 179155 529284 179209 529300
rect 178882 529224 178945 529236
rect 178882 529212 178932 529224
rect 178707 529177 178813 529207
rect 178783 529162 178813 529177
rect 172287 528968 172405 528994
rect 172563 528968 173509 528994
rect 173667 528968 174613 528994
rect 175779 528968 175809 528994
rect 175985 528968 176015 528994
rect 176071 528968 176101 528994
rect 176157 528968 176187 528994
rect 176243 528968 176273 528994
rect 176329 528968 176359 528994
rect 176415 528968 176445 528994
rect 176501 528968 176531 528994
rect 176587 528968 176617 528994
rect 176672 528968 176702 528994
rect 176758 528968 176788 528994
rect 176844 528968 176874 528994
rect 176930 528968 176960 528994
rect 177016 528968 177046 528994
rect 177102 528968 177132 528994
rect 177188 528968 177218 528994
rect 177274 528968 177304 528994
rect 177360 528968 177390 528994
rect 177446 528968 177476 528994
rect 177532 528968 177562 528994
rect 177618 528968 177648 528994
rect 177807 528974 177837 529000
rect 177891 528974 177921 529000
rect 178882 529078 178912 529212
rect 178954 529160 179008 529176
rect 178954 529126 178964 529160
rect 178998 529126 179008 529160
rect 178954 529110 179008 529126
rect 178968 529078 178998 529110
rect 179052 529078 179082 529262
rect 179155 529250 179165 529284
rect 179199 529250 179209 529284
rect 179155 529234 179209 529250
rect 179160 529078 179190 529234
rect 179251 529192 179281 529360
rect 179739 529325 179769 529340
rect 179459 529292 179489 529314
rect 179733 529301 179769 529325
rect 179733 529292 179763 529301
rect 179430 529276 179489 529292
rect 179430 529242 179440 529276
rect 179474 529242 179489 529276
rect 179430 529226 179489 529242
rect 179687 529276 179763 529292
rect 179827 529279 179857 529340
rect 180107 529308 180501 529334
rect 180752 529311 180782 529360
rect 180838 529311 180868 529360
rect 180924 529311 180954 529360
rect 181010 529311 181040 529360
rect 180325 529286 180501 529308
rect 179687 529242 179697 529276
rect 179731 529242 179763 529276
rect 179687 529226 179763 529242
rect 179459 529194 179489 529226
rect 179232 529176 179286 529192
rect 179232 529142 179242 529176
rect 179276 529142 179286 529176
rect 179232 529126 179286 529142
rect 179244 529078 179274 529126
rect 179733 529191 179763 529226
rect 179807 529263 179861 529279
rect 179807 529229 179817 529263
rect 179851 529229 179861 529263
rect 179807 529213 179861 529229
rect 180107 529250 180283 529266
rect 180107 529216 180123 529250
rect 180157 529216 180233 529250
rect 180267 529216 180283 529250
rect 180325 529252 180341 529286
rect 180375 529252 180451 529286
rect 180485 529252 180501 529286
rect 180325 529236 180501 529252
rect 180693 529276 181040 529311
rect 180693 529242 180709 529276
rect 180743 529242 181040 529276
rect 179733 529167 179769 529191
rect 179739 529152 179769 529167
rect 179827 529152 179857 529213
rect 180107 529194 180283 529216
rect 180693 529209 181040 529242
rect 180752 529194 180782 529209
rect 180838 529194 180868 529209
rect 180924 529194 180954 529209
rect 181010 529194 181040 529209
rect 181096 529301 181126 529360
rect 181182 529301 181212 529360
rect 181268 529301 181298 529360
rect 181354 529301 181384 529360
rect 181440 529301 181470 529360
rect 181526 529301 181556 529360
rect 181612 529301 181642 529360
rect 181698 529301 181728 529360
rect 181783 529301 181813 529360
rect 181869 529301 181899 529360
rect 181955 529301 181985 529360
rect 182041 529301 182071 529360
rect 182127 529301 182157 529360
rect 182213 529301 182243 529360
rect 182299 529301 182329 529360
rect 182385 529301 182415 529360
rect 181096 529276 182415 529301
rect 182591 529279 182621 529340
rect 182679 529325 182709 529340
rect 182679 529301 182715 529325
rect 182867 529308 183813 529334
rect 183971 529308 184917 529334
rect 185259 529308 186205 529334
rect 186363 529308 186941 529334
rect 182685 529292 182715 529301
rect 181096 529242 181136 529276
rect 181170 529242 181204 529276
rect 181238 529242 181272 529276
rect 181306 529242 181340 529276
rect 181374 529242 181408 529276
rect 181442 529242 181476 529276
rect 181510 529242 181544 529276
rect 181578 529242 181612 529276
rect 181646 529242 181680 529276
rect 181714 529242 181748 529276
rect 181782 529242 181816 529276
rect 181850 529242 181884 529276
rect 181918 529242 181952 529276
rect 181986 529242 182020 529276
rect 182054 529242 182088 529276
rect 182122 529242 182156 529276
rect 182190 529242 182415 529276
rect 181096 529226 182415 529242
rect 181096 529194 181126 529226
rect 181182 529194 181212 529226
rect 181268 529194 181298 529226
rect 181354 529194 181384 529226
rect 181440 529194 181470 529226
rect 181526 529194 181556 529226
rect 181612 529194 181642 529226
rect 181698 529194 181728 529226
rect 181783 529194 181813 529226
rect 181869 529194 181899 529226
rect 181955 529194 181985 529226
rect 182041 529194 182071 529226
rect 182127 529194 182157 529226
rect 182213 529194 182243 529226
rect 182299 529194 182329 529226
rect 182385 529194 182415 529226
rect 182587 529263 182641 529279
rect 182587 529229 182597 529263
rect 182631 529229 182641 529263
rect 182587 529213 182641 529229
rect 182685 529276 182761 529292
rect 182685 529242 182717 529276
rect 182751 529242 182761 529276
rect 183359 529286 183813 529308
rect 182685 529226 182761 529242
rect 182867 529250 183317 529266
rect 180107 529168 180501 529194
rect 182591 529152 182621 529213
rect 182685 529191 182715 529226
rect 182679 529167 182715 529191
rect 182867 529216 183139 529250
rect 183173 529216 183317 529250
rect 183359 529252 183503 529286
rect 183537 529252 183813 529286
rect 184463 529286 184917 529308
rect 183359 529236 183813 529252
rect 183971 529250 184421 529266
rect 182867 529194 183317 529216
rect 183971 529216 184243 529250
rect 184277 529216 184421 529250
rect 184463 529252 184607 529286
rect 184641 529252 184917 529286
rect 185751 529286 186205 529308
rect 184463 529236 184917 529252
rect 185259 529250 185709 529266
rect 183971 529194 184421 529216
rect 185259 529216 185531 529250
rect 185565 529216 185709 529250
rect 185751 529252 185895 529286
rect 185929 529252 186205 529286
rect 186669 529286 186941 529308
rect 187283 529308 187401 529334
rect 187283 529306 187321 529308
rect 185751 529236 186205 529252
rect 186363 529250 186627 529266
rect 185259 529194 185709 529216
rect 186363 529216 186379 529250
rect 186413 529216 186478 529250
rect 186512 529216 186577 529250
rect 186611 529216 186627 529250
rect 186669 529252 186685 529286
rect 186719 529252 186788 529286
rect 186822 529252 186891 529286
rect 186925 529252 186941 529286
rect 186669 529236 186941 529252
rect 187255 529290 187321 529306
rect 187255 529256 187271 529290
rect 187305 529256 187321 529290
rect 187255 529240 187321 529256
rect 187363 529250 187429 529266
rect 186363 529194 186627 529216
rect 187363 529216 187379 529250
rect 187413 529216 187429 529250
rect 187363 529200 187429 529216
rect 187363 529198 187401 529200
rect 182867 529168 183813 529194
rect 183971 529168 184917 529194
rect 182679 529152 182709 529167
rect 185259 529168 186205 529194
rect 186363 529168 186941 529194
rect 187283 529168 187401 529198
rect 178158 528968 178188 528994
rect 178250 528968 178280 528994
rect 178349 528968 178379 528994
rect 178489 528968 178519 528994
rect 178586 528968 178616 528994
rect 178783 528968 178813 528994
rect 178882 528968 178912 528994
rect 178968 528968 178998 528994
rect 179052 528968 179082 528994
rect 179160 528968 179190 528994
rect 179244 528968 179274 528994
rect 179459 528968 179489 528994
rect 179739 528968 179769 528994
rect 179827 528968 179857 528994
rect 180107 528968 180501 528994
rect 180752 528968 180782 528994
rect 180838 528968 180868 528994
rect 180924 528968 180954 528994
rect 181010 528968 181040 528994
rect 181096 528968 181126 528994
rect 181182 528968 181212 528994
rect 181268 528968 181298 528994
rect 181354 528968 181384 528994
rect 181440 528968 181470 528994
rect 181526 528968 181556 528994
rect 181612 528968 181642 528994
rect 181698 528968 181728 528994
rect 181783 528968 181813 528994
rect 181869 528968 181899 528994
rect 181955 528968 181985 528994
rect 182041 528968 182071 528994
rect 182127 528968 182157 528994
rect 182213 528968 182243 528994
rect 182299 528968 182329 528994
rect 182385 528968 182415 528994
rect 182591 528968 182621 528994
rect 182679 528968 182709 528994
rect 182867 528968 183813 528994
rect 183971 528968 184917 528994
rect 185259 528968 186205 528994
rect 186363 528968 186941 528994
rect 187283 528968 187401 528994
rect 172287 528900 172405 528926
rect 172563 528900 173509 528926
rect 173667 528900 174613 528926
rect 174771 528900 175717 528926
rect 175967 528900 175997 528926
rect 176055 528900 176085 528926
rect 176243 528900 176273 528926
rect 176331 528900 176361 528926
rect 177159 528900 177189 528926
rect 177550 528900 177580 528926
rect 177645 528900 177745 528926
rect 177903 528900 178003 528926
rect 178057 528900 178087 528926
rect 178452 528900 178482 528926
rect 178538 528900 178568 528926
rect 178624 528900 178654 528926
rect 178710 528900 178740 528926
rect 178796 528900 178826 528926
rect 178882 528900 178912 528926
rect 178968 528900 178998 528926
rect 179054 528900 179084 528926
rect 179140 528900 179170 528926
rect 179226 528900 179256 528926
rect 179312 528900 179342 528926
rect 179398 528900 179428 528926
rect 179483 528900 179513 528926
rect 179569 528900 179599 528926
rect 179655 528900 179685 528926
rect 179741 528900 179771 528926
rect 179827 528900 179857 528926
rect 179913 528900 179943 528926
rect 179999 528900 180029 528926
rect 180085 528900 180115 528926
rect 180291 528900 180321 528926
rect 180379 528900 180409 528926
rect 176565 528861 176595 528887
rect 176661 528861 176691 528887
rect 176733 528861 176763 528887
rect 176947 528861 176977 528887
rect 177050 528861 177080 528887
rect 176565 528745 176595 528777
rect 175967 528727 175997 528742
rect 172287 528696 172405 528726
rect 172563 528700 173509 528726
rect 173667 528700 174613 528726
rect 174771 528700 175717 528726
rect 175961 528703 175997 528727
rect 172287 528694 172325 528696
rect 172259 528678 172325 528694
rect 172259 528644 172275 528678
rect 172309 528644 172325 528678
rect 172563 528678 173013 528700
rect 172259 528628 172325 528644
rect 172367 528638 172433 528654
rect 172367 528604 172383 528638
rect 172417 528604 172433 528638
rect 172563 528644 172835 528678
rect 172869 528644 173013 528678
rect 173667 528678 174117 528700
rect 172563 528628 173013 528644
rect 173055 528642 173509 528658
rect 172367 528588 172433 528604
rect 173055 528608 173199 528642
rect 173233 528608 173509 528642
rect 173667 528644 173939 528678
rect 173973 528644 174117 528678
rect 174771 528678 175221 528700
rect 173667 528628 174117 528644
rect 174159 528642 174613 528658
rect 172367 528586 172405 528588
rect 173055 528586 173509 528608
rect 174159 528608 174303 528642
rect 174337 528608 174613 528642
rect 174771 528644 175043 528678
rect 175077 528644 175221 528678
rect 175961 528668 175991 528703
rect 176055 528681 176085 528742
rect 176243 528727 176273 528742
rect 176237 528703 176273 528727
rect 174771 528628 175221 528644
rect 175263 528642 175717 528658
rect 174159 528586 174613 528608
rect 175263 528608 175407 528642
rect 175441 528608 175717 528642
rect 175263 528586 175717 528608
rect 175915 528652 175991 528668
rect 175915 528618 175925 528652
rect 175959 528618 175991 528652
rect 175915 528602 175991 528618
rect 176035 528665 176089 528681
rect 176237 528668 176267 528703
rect 176331 528681 176361 528742
rect 176565 528729 176619 528745
rect 176565 528695 176575 528729
rect 176609 528695 176619 528729
rect 176035 528631 176045 528665
rect 176079 528631 176089 528665
rect 176035 528615 176089 528631
rect 176191 528652 176267 528668
rect 176191 528618 176201 528652
rect 176235 528618 176267 528652
rect 172287 528560 172405 528586
rect 172563 528560 173509 528586
rect 173667 528560 174613 528586
rect 174771 528560 175717 528586
rect 175961 528593 175991 528602
rect 175961 528569 175997 528593
rect 175967 528554 175997 528569
rect 176055 528554 176085 528615
rect 176191 528602 176267 528618
rect 176311 528665 176365 528681
rect 176311 528631 176321 528665
rect 176355 528631 176365 528665
rect 176311 528615 176365 528631
rect 176565 528679 176619 528695
rect 176237 528593 176267 528602
rect 176237 528569 176273 528593
rect 176243 528554 176273 528569
rect 176331 528554 176361 528615
rect 176565 528534 176595 528679
rect 176661 528626 176691 528777
rect 176733 528745 176763 528777
rect 176947 528762 176977 528777
rect 176733 528729 176787 528745
rect 176733 528695 176743 528729
rect 176777 528695 176787 528729
rect 176733 528679 176787 528695
rect 176829 528732 176977 528762
rect 176829 528632 176859 528732
rect 177050 528668 177080 528777
rect 177159 528668 177189 528700
rect 177550 528668 177580 528700
rect 177645 528668 177745 528816
rect 177042 528652 177096 528668
rect 176637 528616 176703 528626
rect 176637 528582 176653 528616
rect 176687 528602 176703 528616
rect 176805 528616 176859 528632
rect 176687 528582 176763 528602
rect 176637 528572 176763 528582
rect 176733 528534 176763 528572
rect 176805 528582 176815 528616
rect 176849 528582 176859 528616
rect 176805 528566 176859 528582
rect 176901 528616 176984 528632
rect 176901 528582 176911 528616
rect 176945 528582 176984 528616
rect 177042 528618 177052 528652
rect 177086 528618 177096 528652
rect 177042 528602 177096 528618
rect 177138 528652 177192 528668
rect 177138 528618 177148 528652
rect 177182 528618 177192 528652
rect 177138 528602 177192 528618
rect 177549 528652 177603 528668
rect 177549 528618 177559 528652
rect 177593 528618 177603 528652
rect 177549 528602 177603 528618
rect 177645 528652 177799 528668
rect 177645 528618 177755 528652
rect 177789 528618 177799 528652
rect 177645 528602 177799 528618
rect 177903 528652 178003 528816
rect 177903 528618 177959 528652
rect 177993 528618 178003 528652
rect 176901 528566 176984 528582
rect 176829 528534 176859 528566
rect 176954 528534 176984 528566
rect 177050 528534 177080 528602
rect 177159 528580 177189 528602
rect 177550 528580 177580 528602
rect 177645 528534 177745 528602
rect 177903 528534 178003 528618
rect 178057 528668 178087 528816
rect 180567 528894 180597 528920
rect 180651 528894 180681 528920
rect 180918 528900 180948 528926
rect 181010 528900 181040 528926
rect 181109 528900 181139 528926
rect 181249 528900 181279 528926
rect 181346 528900 181376 528926
rect 181543 528900 181573 528926
rect 181642 528900 181672 528926
rect 181728 528900 181758 528926
rect 181812 528900 181842 528926
rect 181920 528900 181950 528926
rect 182004 528900 182034 528926
rect 182219 528900 182249 528926
rect 182683 528900 183629 528926
rect 183787 528900 184733 528926
rect 184891 528900 185837 528926
rect 185995 528900 186941 528926
rect 187283 528900 187401 528926
rect 180567 528751 180597 528766
rect 180291 528727 180321 528742
rect 180285 528703 180321 528727
rect 178452 528685 178482 528700
rect 178538 528685 178568 528700
rect 178624 528685 178654 528700
rect 178710 528685 178740 528700
rect 178057 528652 178117 528668
rect 178057 528618 178073 528652
rect 178107 528618 178117 528652
rect 178057 528602 178117 528618
rect 178393 528652 178740 528685
rect 178393 528618 178409 528652
rect 178443 528618 178740 528652
rect 178057 528534 178087 528602
rect 178393 528583 178740 528618
rect 178452 528534 178482 528583
rect 178538 528534 178568 528583
rect 178624 528534 178654 528583
rect 178710 528534 178740 528583
rect 178796 528668 178826 528700
rect 178882 528668 178912 528700
rect 178968 528668 178998 528700
rect 179054 528668 179084 528700
rect 179140 528668 179170 528700
rect 179226 528668 179256 528700
rect 179312 528668 179342 528700
rect 179398 528668 179428 528700
rect 179483 528668 179513 528700
rect 179569 528668 179599 528700
rect 179655 528668 179685 528700
rect 179741 528668 179771 528700
rect 179827 528668 179857 528700
rect 179913 528668 179943 528700
rect 179999 528668 180029 528700
rect 180085 528668 180115 528700
rect 180285 528668 180315 528703
rect 180379 528681 180409 528742
rect 180534 528721 180597 528751
rect 178796 528652 180115 528668
rect 178796 528618 178836 528652
rect 178870 528618 178904 528652
rect 178938 528618 178972 528652
rect 179006 528618 179040 528652
rect 179074 528618 179108 528652
rect 179142 528618 179176 528652
rect 179210 528618 179244 528652
rect 179278 528618 179312 528652
rect 179346 528618 179380 528652
rect 179414 528618 179448 528652
rect 179482 528618 179516 528652
rect 179550 528618 179584 528652
rect 179618 528618 179652 528652
rect 179686 528618 179720 528652
rect 179754 528618 179788 528652
rect 179822 528618 179856 528652
rect 179890 528618 180115 528652
rect 178796 528593 180115 528618
rect 180239 528652 180315 528668
rect 180239 528618 180249 528652
rect 180283 528618 180315 528652
rect 180239 528602 180315 528618
rect 180359 528665 180413 528681
rect 180534 528668 180564 528721
rect 180651 528677 180681 528766
rect 180918 528729 180948 528816
rect 181010 528778 181040 528816
rect 180359 528631 180369 528665
rect 180403 528631 180413 528665
rect 180359 528615 180413 528631
rect 180510 528652 180564 528668
rect 180510 528618 180520 528652
rect 180554 528618 180564 528652
rect 180606 528667 180681 528677
rect 180606 528633 180622 528667
rect 180656 528633 180681 528667
rect 180819 528713 180948 528729
rect 180994 528768 181060 528778
rect 180994 528734 181010 528768
rect 181044 528734 181060 528768
rect 180994 528724 181060 528734
rect 180819 528679 180829 528713
rect 180863 528699 180948 528713
rect 180863 528679 180936 528699
rect 181109 528682 181139 528816
rect 181249 528758 181279 528816
rect 181249 528742 181304 528758
rect 181249 528708 181259 528742
rect 181293 528708 181304 528742
rect 181249 528692 181304 528708
rect 180819 528663 180936 528679
rect 180606 528623 180681 528633
rect 178796 528534 178826 528593
rect 178882 528534 178912 528593
rect 178968 528534 178998 528593
rect 179054 528534 179084 528593
rect 179140 528534 179170 528593
rect 179226 528534 179256 528593
rect 179312 528534 179342 528593
rect 179398 528534 179428 528593
rect 179483 528534 179513 528593
rect 179569 528534 179599 528593
rect 179655 528534 179685 528593
rect 179741 528534 179771 528593
rect 179827 528534 179857 528593
rect 179913 528534 179943 528593
rect 179999 528534 180029 528593
rect 180085 528534 180115 528593
rect 180285 528593 180315 528602
rect 180285 528569 180321 528593
rect 180291 528554 180321 528569
rect 180379 528554 180409 528615
rect 180510 528602 180564 528618
rect 180534 528579 180564 528602
rect 180534 528549 180597 528579
rect 180567 528534 180597 528549
rect 180651 528534 180681 528623
rect 180906 528534 180936 528663
rect 181001 528652 181139 528682
rect 181001 528622 181032 528652
rect 180978 528606 181032 528622
rect 180978 528572 180988 528606
rect 181022 528572 181032 528606
rect 180978 528556 181032 528572
rect 181074 528600 181140 528610
rect 181074 528566 181090 528600
rect 181124 528566 181140 528600
rect 181074 528556 181140 528566
rect 181001 528522 181031 528556
rect 181097 528522 181127 528556
rect 181263 528534 181293 528692
rect 181346 528622 181376 528816
rect 181543 528717 181573 528732
rect 181467 528687 181573 528717
rect 181467 528670 181497 528687
rect 181431 528654 181497 528670
rect 181335 528606 181389 528622
rect 181335 528572 181345 528606
rect 181379 528572 181389 528606
rect 181431 528620 181441 528654
rect 181475 528620 181497 528654
rect 181642 528682 181672 528816
rect 181728 528784 181758 528816
rect 181714 528768 181768 528784
rect 181714 528734 181724 528768
rect 181758 528734 181768 528768
rect 181714 528718 181768 528734
rect 181642 528670 181692 528682
rect 181642 528658 181705 528670
rect 181642 528652 181729 528658
rect 181663 528642 181729 528652
rect 181663 528640 181685 528642
rect 181431 528604 181497 528620
rect 181467 528578 181497 528604
rect 181566 528594 181633 528610
rect 181335 528556 181389 528572
rect 181335 528534 181365 528556
rect 181566 528560 181589 528594
rect 181623 528560 181633 528594
rect 181566 528544 181633 528560
rect 181675 528608 181685 528640
rect 181719 528608 181729 528642
rect 181675 528592 181729 528608
rect 181812 528632 181842 528816
rect 181920 528660 181950 528816
rect 182004 528768 182034 528816
rect 181992 528752 182046 528768
rect 181992 528718 182002 528752
rect 182036 528718 182046 528752
rect 181992 528702 182046 528718
rect 181915 528644 181969 528660
rect 181812 528616 181873 528632
rect 181812 528596 181829 528616
rect 181566 528522 181596 528544
rect 181675 528522 181705 528592
rect 181771 528582 181829 528596
rect 181863 528582 181873 528616
rect 181915 528610 181925 528644
rect 181959 528610 181969 528644
rect 181915 528594 181969 528610
rect 181771 528566 181873 528582
rect 181771 528534 181801 528566
rect 181920 528534 181950 528594
rect 182011 528534 182041 528702
rect 182683 528700 183629 528726
rect 183787 528700 184733 528726
rect 184891 528700 185837 528726
rect 185995 528700 186941 528726
rect 182219 528668 182249 528700
rect 182190 528652 182249 528668
rect 182190 528618 182200 528652
rect 182234 528618 182249 528652
rect 182683 528678 183133 528700
rect 182683 528644 182955 528678
rect 182989 528644 183133 528678
rect 183787 528678 184237 528700
rect 182683 528628 183133 528644
rect 183175 528642 183629 528658
rect 182190 528602 182249 528618
rect 182219 528580 182249 528602
rect 183175 528608 183319 528642
rect 183353 528608 183629 528642
rect 183787 528644 184059 528678
rect 184093 528644 184237 528678
rect 184891 528678 185341 528700
rect 183787 528628 184237 528644
rect 184279 528642 184733 528658
rect 183175 528586 183629 528608
rect 184279 528608 184423 528642
rect 184457 528608 184733 528642
rect 184891 528644 185163 528678
rect 185197 528644 185341 528678
rect 185995 528678 186445 528700
rect 187283 528696 187401 528726
rect 184891 528628 185341 528644
rect 185383 528642 185837 528658
rect 184279 528586 184733 528608
rect 185383 528608 185527 528642
rect 185561 528608 185837 528642
rect 185995 528644 186267 528678
rect 186301 528644 186445 528678
rect 187363 528694 187401 528696
rect 187363 528678 187429 528694
rect 185995 528628 186445 528644
rect 186487 528642 186941 528658
rect 185383 528586 185837 528608
rect 186487 528608 186631 528642
rect 186665 528608 186941 528642
rect 186487 528586 186941 528608
rect 187255 528638 187321 528654
rect 187255 528604 187271 528638
rect 187305 528604 187321 528638
rect 187363 528644 187379 528678
rect 187413 528644 187429 528678
rect 187363 528628 187429 528644
rect 187255 528588 187321 528604
rect 182683 528560 183629 528586
rect 183787 528560 184733 528586
rect 184891 528560 185837 528586
rect 185995 528560 186941 528586
rect 187283 528586 187321 528588
rect 187283 528560 187401 528586
rect 172287 528424 172405 528450
rect 172563 528424 173509 528450
rect 173667 528424 174613 528450
rect 174771 528424 175717 528450
rect 175967 528424 175997 528450
rect 176055 528424 176085 528450
rect 176243 528424 176273 528450
rect 176331 528424 176361 528450
rect 176565 528424 176595 528450
rect 176733 528424 176763 528450
rect 176829 528424 176859 528450
rect 176954 528424 176984 528450
rect 177050 528424 177080 528450
rect 177159 528424 177189 528450
rect 177550 528424 177580 528450
rect 177645 528424 177745 528450
rect 177903 528424 178003 528450
rect 178057 528424 178087 528450
rect 178452 528424 178482 528450
rect 178538 528424 178568 528450
rect 178624 528424 178654 528450
rect 178710 528424 178740 528450
rect 178796 528424 178826 528450
rect 178882 528424 178912 528450
rect 178968 528424 178998 528450
rect 179054 528424 179084 528450
rect 179140 528424 179170 528450
rect 179226 528424 179256 528450
rect 179312 528424 179342 528450
rect 179398 528424 179428 528450
rect 179483 528424 179513 528450
rect 179569 528424 179599 528450
rect 179655 528424 179685 528450
rect 179741 528424 179771 528450
rect 179827 528424 179857 528450
rect 179913 528424 179943 528450
rect 179999 528424 180029 528450
rect 180085 528424 180115 528450
rect 180291 528424 180321 528450
rect 180379 528424 180409 528450
rect 180567 528424 180597 528450
rect 180651 528424 180681 528450
rect 180906 528424 180936 528450
rect 181001 528424 181031 528450
rect 181097 528424 181127 528450
rect 181263 528424 181293 528450
rect 181335 528424 181365 528450
rect 181467 528424 181497 528450
rect 181566 528424 181596 528450
rect 181675 528424 181705 528450
rect 181771 528424 181801 528450
rect 181920 528424 181950 528450
rect 182011 528424 182041 528450
rect 182219 528424 182249 528450
rect 182683 528424 183629 528450
rect 183787 528424 184733 528450
rect 184891 528424 185837 528450
rect 185995 528424 186941 528450
rect 187283 528424 187401 528450
rect 172287 528356 172405 528382
rect 172563 528356 173509 528382
rect 173667 528356 174613 528382
rect 174955 528356 175901 528382
rect 176151 528356 176181 528382
rect 176235 528356 176265 528382
rect 176490 528356 176520 528382
rect 176585 528356 176615 528382
rect 176681 528356 176711 528382
rect 176847 528356 176877 528382
rect 176919 528356 176949 528382
rect 177051 528356 177081 528382
rect 177150 528356 177180 528382
rect 177259 528356 177289 528382
rect 177355 528356 177385 528382
rect 177504 528356 177534 528382
rect 177595 528356 177625 528382
rect 177803 528356 177833 528382
rect 177991 528356 178021 528382
rect 178079 528356 178109 528382
rect 178267 528356 178845 528382
rect 179003 528356 179033 528382
rect 179112 528356 179142 528382
rect 179208 528356 179238 528382
rect 179333 528356 179363 528382
rect 179429 528356 179459 528382
rect 179597 528356 179627 528382
rect 180107 528356 180685 528382
rect 181027 528356 181057 528382
rect 181136 528356 181166 528382
rect 181232 528356 181262 528382
rect 181357 528356 181387 528382
rect 181453 528356 181483 528382
rect 181621 528356 181651 528382
rect 181855 528356 182801 528382
rect 182959 528356 183905 528382
rect 184063 528356 185009 528382
rect 185259 528356 186205 528382
rect 186363 528356 186941 528382
rect 187283 528356 187401 528382
rect 172287 528220 172405 528246
rect 172563 528220 173509 528246
rect 173667 528220 174613 528246
rect 176151 528257 176181 528272
rect 174955 528220 175901 528246
rect 172367 528218 172405 528220
rect 172367 528202 172433 528218
rect 172259 528162 172325 528178
rect 172259 528128 172275 528162
rect 172309 528128 172325 528162
rect 172367 528168 172383 528202
rect 172417 528168 172433 528202
rect 173055 528198 173509 528220
rect 172367 528152 172433 528168
rect 172563 528162 173013 528178
rect 172259 528112 172325 528128
rect 172287 528110 172325 528112
rect 172563 528128 172835 528162
rect 172869 528128 173013 528162
rect 173055 528164 173199 528198
rect 173233 528164 173509 528198
rect 174159 528198 174613 528220
rect 173055 528148 173509 528164
rect 173667 528162 174117 528178
rect 172287 528080 172405 528110
rect 172563 528106 173013 528128
rect 173667 528128 173939 528162
rect 173973 528128 174117 528162
rect 174159 528164 174303 528198
rect 174337 528164 174613 528198
rect 175447 528198 175901 528220
rect 176118 528227 176181 528257
rect 176118 528204 176148 528227
rect 174159 528148 174613 528164
rect 174955 528162 175405 528178
rect 173667 528106 174117 528128
rect 174955 528128 175227 528162
rect 175261 528128 175405 528162
rect 175447 528164 175591 528198
rect 175625 528164 175901 528198
rect 175447 528148 175901 528164
rect 176094 528188 176148 528204
rect 176094 528154 176104 528188
rect 176138 528154 176148 528188
rect 176235 528183 176265 528272
rect 176094 528138 176148 528154
rect 174955 528106 175405 528128
rect 172563 528080 173509 528106
rect 173667 528080 174613 528106
rect 174955 528080 175901 528106
rect 176118 528085 176148 528138
rect 176190 528173 176265 528183
rect 176190 528139 176206 528173
rect 176240 528139 176265 528173
rect 176490 528143 176520 528272
rect 176585 528250 176615 528284
rect 176681 528250 176711 528284
rect 176562 528234 176616 528250
rect 176562 528200 176572 528234
rect 176606 528200 176616 528234
rect 176562 528184 176616 528200
rect 176658 528240 176724 528250
rect 176658 528206 176674 528240
rect 176708 528206 176724 528240
rect 176658 528196 176724 528206
rect 176190 528129 176265 528139
rect 176118 528055 176181 528085
rect 176151 528040 176181 528055
rect 176235 528040 176265 528129
rect 176403 528127 176520 528143
rect 176403 528093 176413 528127
rect 176447 528107 176520 528127
rect 176585 528154 176616 528184
rect 176585 528124 176723 528154
rect 176447 528093 176532 528107
rect 176403 528077 176532 528093
rect 176502 527990 176532 528077
rect 176578 528072 176644 528082
rect 176578 528038 176594 528072
rect 176628 528038 176644 528072
rect 176578 528028 176644 528038
rect 176594 527990 176624 528028
rect 176693 527990 176723 528124
rect 176847 528114 176877 528272
rect 176919 528250 176949 528272
rect 176919 528234 176973 528250
rect 176919 528200 176929 528234
rect 176963 528200 176973 528234
rect 177150 528262 177180 528284
rect 177150 528246 177217 528262
rect 177051 528202 177081 528228
rect 176919 528184 176973 528200
rect 177015 528186 177081 528202
rect 177150 528212 177173 528246
rect 177207 528212 177217 528246
rect 177150 528196 177217 528212
rect 177259 528214 177289 528284
rect 177355 528240 177385 528272
rect 177355 528224 177457 528240
rect 177259 528198 177313 528214
rect 177355 528210 177413 528224
rect 176833 528098 176888 528114
rect 176833 528064 176843 528098
rect 176877 528064 176888 528098
rect 176833 528048 176888 528064
rect 176833 527990 176863 528048
rect 176930 527990 176960 528184
rect 177015 528152 177025 528186
rect 177059 528152 177081 528186
rect 177259 528166 177269 528198
rect 177247 528164 177269 528166
rect 177303 528164 177313 528198
rect 177247 528154 177313 528164
rect 177015 528136 177081 528152
rect 177051 528119 177081 528136
rect 177226 528148 177313 528154
rect 177396 528190 177413 528210
rect 177447 528190 177457 528224
rect 177504 528212 177534 528272
rect 177396 528174 177457 528190
rect 177499 528196 177553 528212
rect 177226 528136 177289 528148
rect 177226 528124 177276 528136
rect 177051 528089 177157 528119
rect 177127 528074 177157 528089
rect 172287 527880 172405 527906
rect 172563 527880 173509 527906
rect 173667 527880 174613 527906
rect 174955 527880 175901 527906
rect 176151 527886 176181 527912
rect 176235 527886 176265 527912
rect 177226 527990 177256 528124
rect 177298 528072 177352 528088
rect 177298 528038 177308 528072
rect 177342 528038 177352 528072
rect 177298 528022 177352 528038
rect 177312 527990 177342 528022
rect 177396 527990 177426 528174
rect 177499 528162 177509 528196
rect 177543 528162 177553 528196
rect 177499 528146 177553 528162
rect 177504 527990 177534 528146
rect 177595 528104 177625 528272
rect 177803 528204 177833 528226
rect 177774 528188 177833 528204
rect 177991 528191 178021 528252
rect 178079 528237 178109 528252
rect 178079 528213 178115 528237
rect 178267 528220 178845 528246
rect 178085 528204 178115 528213
rect 177774 528154 177784 528188
rect 177818 528154 177833 528188
rect 177774 528138 177833 528154
rect 177803 528106 177833 528138
rect 177987 528175 178041 528191
rect 177987 528141 177997 528175
rect 178031 528141 178041 528175
rect 177987 528125 178041 528141
rect 178085 528188 178161 528204
rect 178085 528154 178117 528188
rect 178151 528154 178161 528188
rect 178573 528198 178845 528220
rect 179003 528204 179033 528226
rect 179112 528204 179142 528272
rect 179208 528240 179238 528272
rect 179333 528240 179363 528272
rect 179208 528224 179291 528240
rect 178085 528138 178161 528154
rect 178267 528162 178531 528178
rect 177576 528088 177630 528104
rect 177576 528054 177586 528088
rect 177620 528054 177630 528088
rect 177576 528038 177630 528054
rect 177588 527990 177618 528038
rect 177991 528064 178021 528125
rect 178085 528103 178115 528138
rect 178079 528079 178115 528103
rect 178267 528128 178283 528162
rect 178317 528128 178382 528162
rect 178416 528128 178481 528162
rect 178515 528128 178531 528162
rect 178573 528164 178589 528198
rect 178623 528164 178692 528198
rect 178726 528164 178795 528198
rect 178829 528164 178845 528198
rect 178573 528148 178845 528164
rect 179000 528188 179054 528204
rect 179000 528154 179010 528188
rect 179044 528154 179054 528188
rect 179000 528138 179054 528154
rect 179096 528188 179150 528204
rect 179096 528154 179106 528188
rect 179140 528154 179150 528188
rect 179208 528190 179247 528224
rect 179281 528190 179291 528224
rect 179208 528174 179291 528190
rect 179333 528224 179387 528240
rect 179333 528190 179343 528224
rect 179377 528190 179387 528224
rect 179429 528234 179459 528272
rect 179429 528224 179555 528234
rect 179429 528204 179505 528224
rect 179333 528174 179387 528190
rect 179489 528190 179505 528204
rect 179539 528190 179555 528224
rect 179489 528180 179555 528190
rect 179096 528138 179150 528154
rect 178267 528106 178531 528128
rect 179003 528106 179033 528138
rect 178267 528080 178845 528106
rect 178079 528064 178109 528079
rect 179112 528029 179142 528138
rect 179333 528074 179363 528174
rect 179215 528044 179363 528074
rect 179405 528111 179459 528127
rect 179405 528077 179415 528111
rect 179449 528077 179459 528111
rect 179405 528061 179459 528077
rect 179215 528029 179245 528044
rect 179429 528029 179459 528061
rect 179501 528029 179531 528180
rect 179597 528127 179627 528272
rect 180107 528220 180685 528246
rect 180413 528198 180685 528220
rect 181027 528204 181057 528226
rect 181136 528204 181166 528272
rect 181232 528240 181262 528272
rect 181357 528240 181387 528272
rect 181232 528224 181315 528240
rect 179573 528111 179627 528127
rect 179573 528077 179583 528111
rect 179617 528077 179627 528111
rect 180107 528162 180371 528178
rect 180107 528128 180123 528162
rect 180157 528128 180222 528162
rect 180256 528128 180321 528162
rect 180355 528128 180371 528162
rect 180413 528164 180429 528198
rect 180463 528164 180532 528198
rect 180566 528164 180635 528198
rect 180669 528164 180685 528198
rect 180413 528148 180685 528164
rect 181024 528188 181078 528204
rect 181024 528154 181034 528188
rect 181068 528154 181078 528188
rect 181024 528138 181078 528154
rect 181120 528188 181174 528204
rect 181120 528154 181130 528188
rect 181164 528154 181174 528188
rect 181232 528190 181271 528224
rect 181305 528190 181315 528224
rect 181232 528174 181315 528190
rect 181357 528224 181411 528240
rect 181357 528190 181367 528224
rect 181401 528190 181411 528224
rect 181453 528234 181483 528272
rect 181453 528224 181579 528234
rect 181453 528204 181529 528224
rect 181357 528174 181411 528190
rect 181513 528190 181529 528204
rect 181563 528190 181579 528224
rect 181513 528180 181579 528190
rect 181120 528138 181174 528154
rect 180107 528106 180371 528128
rect 181027 528106 181057 528138
rect 179573 528061 179627 528077
rect 179597 528029 179627 528061
rect 180107 528080 180685 528106
rect 179112 527919 179142 527945
rect 179215 527919 179245 527945
rect 179429 527919 179459 527945
rect 179501 527919 179531 527945
rect 179597 527919 179627 527945
rect 181136 528029 181166 528138
rect 181357 528074 181387 528174
rect 181239 528044 181387 528074
rect 181429 528111 181483 528127
rect 181429 528077 181439 528111
rect 181473 528077 181483 528111
rect 181429 528061 181483 528077
rect 181239 528029 181269 528044
rect 181453 528029 181483 528061
rect 181525 528029 181555 528180
rect 181621 528127 181651 528272
rect 181855 528220 182801 528246
rect 182959 528220 183905 528246
rect 184063 528220 185009 528246
rect 185259 528220 186205 528246
rect 186363 528220 186941 528246
rect 182347 528198 182801 528220
rect 181597 528111 181651 528127
rect 181597 528077 181607 528111
rect 181641 528077 181651 528111
rect 181855 528162 182305 528178
rect 181855 528128 182127 528162
rect 182161 528128 182305 528162
rect 182347 528164 182491 528198
rect 182525 528164 182801 528198
rect 183451 528198 183905 528220
rect 182347 528148 182801 528164
rect 182959 528162 183409 528178
rect 181855 528106 182305 528128
rect 182959 528128 183231 528162
rect 183265 528128 183409 528162
rect 183451 528164 183595 528198
rect 183629 528164 183905 528198
rect 184555 528198 185009 528220
rect 183451 528148 183905 528164
rect 184063 528162 184513 528178
rect 182959 528106 183409 528128
rect 184063 528128 184335 528162
rect 184369 528128 184513 528162
rect 184555 528164 184699 528198
rect 184733 528164 185009 528198
rect 185751 528198 186205 528220
rect 184555 528148 185009 528164
rect 185259 528162 185709 528178
rect 184063 528106 184513 528128
rect 185259 528128 185531 528162
rect 185565 528128 185709 528162
rect 185751 528164 185895 528198
rect 185929 528164 186205 528198
rect 186669 528198 186941 528220
rect 187283 528220 187401 528246
rect 187283 528218 187321 528220
rect 185751 528148 186205 528164
rect 186363 528162 186627 528178
rect 185259 528106 185709 528128
rect 186363 528128 186379 528162
rect 186413 528128 186478 528162
rect 186512 528128 186577 528162
rect 186611 528128 186627 528162
rect 186669 528164 186685 528198
rect 186719 528164 186788 528198
rect 186822 528164 186891 528198
rect 186925 528164 186941 528198
rect 186669 528148 186941 528164
rect 187255 528202 187321 528218
rect 187255 528168 187271 528202
rect 187305 528168 187321 528202
rect 187255 528152 187321 528168
rect 187363 528162 187429 528178
rect 186363 528106 186627 528128
rect 187363 528128 187379 528162
rect 187413 528128 187429 528162
rect 187363 528112 187429 528128
rect 187363 528110 187401 528112
rect 181855 528080 182801 528106
rect 182959 528080 183905 528106
rect 184063 528080 185009 528106
rect 181597 528061 181651 528077
rect 181621 528029 181651 528061
rect 181136 527919 181166 527945
rect 181239 527919 181269 527945
rect 181453 527919 181483 527945
rect 181525 527919 181555 527945
rect 181621 527919 181651 527945
rect 185259 528080 186205 528106
rect 186363 528080 186941 528106
rect 187283 528080 187401 528110
rect 176502 527880 176532 527906
rect 176594 527880 176624 527906
rect 176693 527880 176723 527906
rect 176833 527880 176863 527906
rect 176930 527880 176960 527906
rect 177127 527880 177157 527906
rect 177226 527880 177256 527906
rect 177312 527880 177342 527906
rect 177396 527880 177426 527906
rect 177504 527880 177534 527906
rect 177588 527880 177618 527906
rect 177803 527880 177833 527906
rect 177991 527880 178021 527906
rect 178079 527880 178109 527906
rect 178267 527880 178845 527906
rect 179003 527880 179033 527906
rect 180107 527880 180685 527906
rect 181027 527880 181057 527906
rect 181855 527880 182801 527906
rect 182959 527880 183905 527906
rect 184063 527880 185009 527906
rect 185259 527880 186205 527906
rect 186363 527880 186941 527906
rect 187283 527880 187401 527906
rect 172287 527812 172405 527838
rect 172563 527812 173509 527838
rect 173667 527812 174613 527838
rect 174771 527812 175717 527838
rect 175875 527812 176269 527838
rect 176446 527812 176476 527838
rect 176541 527812 176641 527838
rect 176799 527812 176899 527838
rect 176953 527812 176983 527838
rect 177163 527812 177281 527838
rect 177531 527812 178477 527838
rect 178635 527812 178845 527838
rect 179022 527812 179052 527838
rect 179117 527812 179217 527838
rect 179375 527812 179475 527838
rect 179529 527812 179559 527838
rect 179739 527812 180685 527838
rect 180843 527812 181789 527838
rect 181947 527812 182341 527838
rect 182683 527812 183629 527838
rect 183787 527812 184733 527838
rect 184891 527812 185837 527838
rect 185995 527812 186941 527838
rect 187283 527812 187401 527838
rect 172287 527608 172405 527638
rect 172563 527612 173509 527638
rect 173667 527612 174613 527638
rect 174771 527612 175717 527638
rect 175875 527612 176269 527638
rect 172287 527606 172325 527608
rect 172259 527590 172325 527606
rect 172259 527556 172275 527590
rect 172309 527556 172325 527590
rect 172563 527590 173013 527612
rect 172259 527540 172325 527556
rect 172367 527550 172433 527566
rect 172367 527516 172383 527550
rect 172417 527516 172433 527550
rect 172563 527556 172835 527590
rect 172869 527556 173013 527590
rect 173667 527590 174117 527612
rect 172563 527540 173013 527556
rect 173055 527554 173509 527570
rect 172367 527500 172433 527516
rect 173055 527520 173199 527554
rect 173233 527520 173509 527554
rect 173667 527556 173939 527590
rect 173973 527556 174117 527590
rect 174771 527590 175221 527612
rect 173667 527540 174117 527556
rect 174159 527554 174613 527570
rect 172367 527498 172405 527500
rect 173055 527498 173509 527520
rect 174159 527520 174303 527554
rect 174337 527520 174613 527554
rect 174771 527556 175043 527590
rect 175077 527556 175221 527590
rect 175875 527590 176051 527612
rect 174771 527540 175221 527556
rect 175263 527554 175717 527570
rect 174159 527498 174613 527520
rect 175263 527520 175407 527554
rect 175441 527520 175717 527554
rect 175875 527556 175891 527590
rect 175925 527556 176001 527590
rect 176035 527556 176051 527590
rect 176446 527580 176476 527612
rect 176541 527580 176641 527728
rect 175875 527540 176051 527556
rect 176093 527554 176269 527570
rect 175263 527498 175717 527520
rect 176093 527520 176109 527554
rect 176143 527520 176219 527554
rect 176253 527520 176269 527554
rect 176093 527498 176269 527520
rect 176445 527564 176499 527580
rect 176445 527530 176455 527564
rect 176489 527530 176499 527564
rect 176445 527514 176499 527530
rect 176541 527564 176695 527580
rect 176541 527530 176651 527564
rect 176685 527530 176695 527564
rect 176541 527514 176695 527530
rect 176799 527564 176899 527728
rect 176799 527530 176855 527564
rect 176889 527530 176899 527564
rect 172287 527472 172405 527498
rect 172563 527472 173509 527498
rect 173667 527472 174613 527498
rect 174771 527472 175717 527498
rect 175875 527472 176269 527498
rect 176446 527492 176476 527514
rect 176541 527446 176641 527514
rect 176799 527446 176899 527530
rect 176953 527580 176983 527728
rect 177163 527608 177281 527638
rect 177531 527612 178477 527638
rect 178635 527612 178845 527638
rect 177163 527606 177201 527608
rect 177135 527590 177201 527606
rect 176953 527564 177013 527580
rect 176953 527530 176969 527564
rect 177003 527530 177013 527564
rect 177135 527556 177151 527590
rect 177185 527556 177201 527590
rect 177531 527590 177981 527612
rect 178635 527606 178719 527612
rect 177135 527540 177201 527556
rect 177243 527550 177309 527566
rect 176953 527514 177013 527530
rect 177243 527516 177259 527550
rect 177293 527516 177309 527550
rect 177531 527556 177803 527590
rect 177837 527556 177981 527590
rect 178577 527590 178719 527606
rect 177531 527540 177981 527556
rect 178023 527554 178477 527570
rect 176953 527446 176983 527514
rect 177243 527500 177309 527516
rect 178023 527520 178167 527554
rect 178201 527520 178477 527554
rect 178577 527556 178593 527590
rect 178627 527556 178719 527590
rect 179022 527580 179052 527612
rect 179117 527580 179217 527728
rect 178577 527540 178719 527556
rect 178761 527554 178903 527570
rect 177243 527498 177281 527500
rect 178023 527498 178477 527520
rect 178761 527520 178853 527554
rect 178887 527520 178903 527554
rect 178761 527504 178903 527520
rect 179021 527564 179075 527580
rect 179021 527530 179031 527564
rect 179065 527530 179075 527564
rect 179021 527514 179075 527530
rect 179117 527564 179271 527580
rect 179117 527530 179227 527564
rect 179261 527530 179271 527564
rect 179117 527514 179271 527530
rect 179375 527564 179475 527728
rect 179375 527530 179431 527564
rect 179465 527530 179475 527564
rect 178761 527498 178845 527504
rect 177163 527472 177281 527498
rect 177531 527472 178477 527498
rect 178635 527472 178845 527498
rect 179022 527492 179052 527514
rect 179117 527446 179217 527514
rect 179375 527446 179475 527530
rect 179529 527580 179559 527728
rect 179739 527612 180685 527638
rect 180843 527612 181789 527638
rect 181947 527612 182341 527638
rect 182683 527612 183629 527638
rect 183787 527612 184733 527638
rect 184891 527612 185837 527638
rect 185995 527612 186941 527638
rect 179739 527590 180189 527612
rect 179529 527564 179589 527580
rect 179529 527530 179545 527564
rect 179579 527530 179589 527564
rect 179739 527556 180011 527590
rect 180045 527556 180189 527590
rect 180843 527590 181293 527612
rect 179739 527540 180189 527556
rect 180231 527554 180685 527570
rect 179529 527514 179589 527530
rect 180231 527520 180375 527554
rect 180409 527520 180685 527554
rect 180843 527556 181115 527590
rect 181149 527556 181293 527590
rect 181947 527590 182123 527612
rect 180843 527540 181293 527556
rect 181335 527554 181789 527570
rect 179529 527446 179559 527514
rect 180231 527498 180685 527520
rect 181335 527520 181479 527554
rect 181513 527520 181789 527554
rect 181947 527556 181963 527590
rect 181997 527556 182073 527590
rect 182107 527556 182123 527590
rect 182683 527590 183133 527612
rect 181947 527540 182123 527556
rect 182165 527554 182341 527570
rect 181335 527498 181789 527520
rect 182165 527520 182181 527554
rect 182215 527520 182291 527554
rect 182325 527520 182341 527554
rect 182683 527556 182955 527590
rect 182989 527556 183133 527590
rect 183787 527590 184237 527612
rect 182683 527540 183133 527556
rect 183175 527554 183629 527570
rect 182165 527498 182341 527520
rect 183175 527520 183319 527554
rect 183353 527520 183629 527554
rect 183787 527556 184059 527590
rect 184093 527556 184237 527590
rect 184891 527590 185341 527612
rect 183787 527540 184237 527556
rect 184279 527554 184733 527570
rect 183175 527498 183629 527520
rect 184279 527520 184423 527554
rect 184457 527520 184733 527554
rect 184891 527556 185163 527590
rect 185197 527556 185341 527590
rect 185995 527590 186445 527612
rect 187283 527608 187401 527638
rect 184891 527540 185341 527556
rect 185383 527554 185837 527570
rect 184279 527498 184733 527520
rect 185383 527520 185527 527554
rect 185561 527520 185837 527554
rect 185995 527556 186267 527590
rect 186301 527556 186445 527590
rect 187363 527606 187401 527608
rect 187363 527590 187429 527606
rect 185995 527540 186445 527556
rect 186487 527554 186941 527570
rect 185383 527498 185837 527520
rect 186487 527520 186631 527554
rect 186665 527520 186941 527554
rect 186487 527498 186941 527520
rect 187255 527550 187321 527566
rect 187255 527516 187271 527550
rect 187305 527516 187321 527550
rect 187363 527556 187379 527590
rect 187413 527556 187429 527590
rect 187363 527540 187429 527556
rect 187255 527500 187321 527516
rect 179739 527472 180685 527498
rect 180843 527472 181789 527498
rect 181947 527472 182341 527498
rect 182683 527472 183629 527498
rect 183787 527472 184733 527498
rect 184891 527472 185837 527498
rect 185995 527472 186941 527498
rect 187283 527498 187321 527500
rect 187283 527472 187401 527498
rect 172287 527336 172405 527362
rect 172563 527336 173509 527362
rect 173667 527336 174613 527362
rect 174771 527336 175717 527362
rect 175875 527336 176269 527362
rect 176446 527336 176476 527362
rect 176541 527336 176641 527362
rect 176799 527336 176899 527362
rect 176953 527336 176983 527362
rect 177163 527336 177281 527362
rect 177531 527336 178477 527362
rect 178635 527336 178845 527362
rect 179022 527336 179052 527362
rect 179117 527336 179217 527362
rect 179375 527336 179475 527362
rect 179529 527336 179559 527362
rect 179739 527336 180685 527362
rect 180843 527336 181789 527362
rect 181947 527336 182341 527362
rect 182683 527336 183629 527362
rect 183787 527336 184733 527362
rect 184891 527336 185837 527362
rect 185995 527336 186941 527362
rect 187283 527336 187401 527362
rect 172287 527268 172405 527294
rect 172563 527268 173509 527294
rect 173667 527268 174613 527294
rect 174955 527268 175901 527294
rect 176059 527268 177005 527294
rect 177163 527268 178109 527294
rect 178267 527268 179213 527294
rect 179371 527268 179765 527294
rect 180107 527268 181053 527294
rect 181211 527268 182157 527294
rect 182315 527268 183261 527294
rect 183419 527268 184365 527294
rect 184523 527268 184917 527294
rect 185259 527268 186205 527294
rect 186363 527268 186941 527294
rect 187283 527268 187401 527294
rect 172287 527132 172405 527158
rect 172563 527132 173509 527158
rect 173667 527132 174613 527158
rect 174955 527132 175901 527158
rect 176059 527132 177005 527158
rect 177163 527132 178109 527158
rect 178267 527132 179213 527158
rect 179371 527132 179765 527158
rect 180107 527132 181053 527158
rect 181211 527132 182157 527158
rect 182315 527132 183261 527158
rect 183419 527132 184365 527158
rect 184523 527132 184917 527158
rect 185259 527132 186205 527158
rect 186363 527132 186941 527158
rect 172367 527130 172405 527132
rect 172367 527114 172433 527130
rect 172259 527074 172325 527090
rect 172259 527040 172275 527074
rect 172309 527040 172325 527074
rect 172367 527080 172383 527114
rect 172417 527080 172433 527114
rect 173055 527110 173509 527132
rect 172367 527064 172433 527080
rect 172563 527074 173013 527090
rect 172259 527024 172325 527040
rect 172287 527022 172325 527024
rect 172563 527040 172835 527074
rect 172869 527040 173013 527074
rect 173055 527076 173199 527110
rect 173233 527076 173509 527110
rect 174159 527110 174613 527132
rect 173055 527060 173509 527076
rect 173667 527074 174117 527090
rect 172287 526992 172405 527022
rect 172563 527018 173013 527040
rect 173667 527040 173939 527074
rect 173973 527040 174117 527074
rect 174159 527076 174303 527110
rect 174337 527076 174613 527110
rect 175447 527110 175901 527132
rect 174159 527060 174613 527076
rect 174955 527074 175405 527090
rect 173667 527018 174117 527040
rect 174955 527040 175227 527074
rect 175261 527040 175405 527074
rect 175447 527076 175591 527110
rect 175625 527076 175901 527110
rect 176551 527110 177005 527132
rect 175447 527060 175901 527076
rect 176059 527074 176509 527090
rect 174955 527018 175405 527040
rect 176059 527040 176331 527074
rect 176365 527040 176509 527074
rect 176551 527076 176695 527110
rect 176729 527076 177005 527110
rect 177655 527110 178109 527132
rect 176551 527060 177005 527076
rect 177163 527074 177613 527090
rect 176059 527018 176509 527040
rect 177163 527040 177435 527074
rect 177469 527040 177613 527074
rect 177655 527076 177799 527110
rect 177833 527076 178109 527110
rect 178759 527110 179213 527132
rect 177655 527060 178109 527076
rect 178267 527074 178717 527090
rect 177163 527018 177613 527040
rect 178267 527040 178539 527074
rect 178573 527040 178717 527074
rect 178759 527076 178903 527110
rect 178937 527076 179213 527110
rect 179589 527110 179765 527132
rect 178759 527060 179213 527076
rect 179371 527074 179547 527090
rect 178267 527018 178717 527040
rect 179371 527040 179387 527074
rect 179421 527040 179497 527074
rect 179531 527040 179547 527074
rect 179589 527076 179605 527110
rect 179639 527076 179715 527110
rect 179749 527076 179765 527110
rect 180599 527110 181053 527132
rect 179589 527060 179765 527076
rect 180107 527074 180557 527090
rect 179371 527018 179547 527040
rect 180107 527040 180379 527074
rect 180413 527040 180557 527074
rect 180599 527076 180743 527110
rect 180777 527076 181053 527110
rect 181703 527110 182157 527132
rect 180599 527060 181053 527076
rect 181211 527074 181661 527090
rect 180107 527018 180557 527040
rect 181211 527040 181483 527074
rect 181517 527040 181661 527074
rect 181703 527076 181847 527110
rect 181881 527076 182157 527110
rect 182807 527110 183261 527132
rect 181703 527060 182157 527076
rect 182315 527074 182765 527090
rect 181211 527018 181661 527040
rect 182315 527040 182587 527074
rect 182621 527040 182765 527074
rect 182807 527076 182951 527110
rect 182985 527076 183261 527110
rect 183911 527110 184365 527132
rect 182807 527060 183261 527076
rect 183419 527074 183869 527090
rect 182315 527018 182765 527040
rect 183419 527040 183691 527074
rect 183725 527040 183869 527074
rect 183911 527076 184055 527110
rect 184089 527076 184365 527110
rect 184741 527110 184917 527132
rect 183911 527060 184365 527076
rect 184523 527074 184699 527090
rect 183419 527018 183869 527040
rect 184523 527040 184539 527074
rect 184573 527040 184649 527074
rect 184683 527040 184699 527074
rect 184741 527076 184757 527110
rect 184791 527076 184867 527110
rect 184901 527076 184917 527110
rect 185751 527110 186205 527132
rect 184741 527060 184917 527076
rect 185259 527074 185709 527090
rect 184523 527018 184699 527040
rect 185259 527040 185531 527074
rect 185565 527040 185709 527074
rect 185751 527076 185895 527110
rect 185929 527076 186205 527110
rect 186669 527110 186941 527132
rect 187283 527132 187401 527158
rect 187283 527130 187321 527132
rect 185751 527060 186205 527076
rect 186363 527074 186627 527090
rect 185259 527018 185709 527040
rect 186363 527040 186379 527074
rect 186413 527040 186478 527074
rect 186512 527040 186577 527074
rect 186611 527040 186627 527074
rect 186669 527076 186685 527110
rect 186719 527076 186788 527110
rect 186822 527076 186891 527110
rect 186925 527076 186941 527110
rect 186669 527060 186941 527076
rect 187255 527114 187321 527130
rect 187255 527080 187271 527114
rect 187305 527080 187321 527114
rect 187255 527064 187321 527080
rect 187363 527074 187429 527090
rect 186363 527018 186627 527040
rect 187363 527040 187379 527074
rect 187413 527040 187429 527074
rect 187363 527024 187429 527040
rect 187363 527022 187401 527024
rect 172563 526992 173509 527018
rect 173667 526992 174613 527018
rect 174955 526992 175901 527018
rect 176059 526992 177005 527018
rect 177163 526992 178109 527018
rect 178267 526992 179213 527018
rect 179371 526992 179765 527018
rect 180107 526992 181053 527018
rect 181211 526992 182157 527018
rect 182315 526992 183261 527018
rect 183419 526992 184365 527018
rect 184523 526992 184917 527018
rect 185259 526992 186205 527018
rect 186363 526992 186941 527018
rect 187283 526992 187401 527022
rect 172287 526792 172405 526818
rect 172563 526792 173509 526818
rect 173667 526792 174613 526818
rect 174955 526792 175901 526818
rect 176059 526792 177005 526818
rect 177163 526792 178109 526818
rect 178267 526792 179213 526818
rect 179371 526792 179765 526818
rect 180107 526792 181053 526818
rect 181211 526792 182157 526818
rect 182315 526792 183261 526818
rect 183419 526792 184365 526818
rect 184523 526792 184917 526818
rect 185259 526792 186205 526818
rect 186363 526792 186941 526818
rect 187283 526792 187401 526818
rect 172287 526724 172405 526750
rect 172563 526724 173509 526750
rect 173667 526724 174613 526750
rect 174771 526724 175717 526750
rect 175875 526724 176821 526750
rect 176979 526724 177189 526750
rect 177531 526724 178477 526750
rect 178635 526724 179581 526750
rect 179739 526724 180685 526750
rect 180843 526724 181789 526750
rect 181947 526724 182341 526750
rect 182683 526724 183629 526750
rect 183787 526724 184733 526750
rect 184891 526724 185837 526750
rect 185995 526724 186941 526750
rect 187283 526724 187401 526750
rect 172287 526520 172405 526550
rect 172563 526524 173509 526550
rect 173667 526524 174613 526550
rect 174771 526524 175717 526550
rect 175875 526524 176821 526550
rect 176979 526524 177189 526550
rect 177531 526524 178477 526550
rect 178635 526524 179581 526550
rect 179739 526524 180685 526550
rect 180843 526524 181789 526550
rect 181947 526524 182341 526550
rect 182683 526524 183629 526550
rect 183787 526524 184733 526550
rect 184891 526524 185837 526550
rect 185995 526524 186941 526550
rect 172287 526518 172325 526520
rect 172259 526502 172325 526518
rect 172259 526468 172275 526502
rect 172309 526468 172325 526502
rect 172563 526502 173013 526524
rect 172259 526452 172325 526468
rect 172367 526462 172433 526478
rect 172367 526428 172383 526462
rect 172417 526428 172433 526462
rect 172563 526468 172835 526502
rect 172869 526468 173013 526502
rect 173667 526502 174117 526524
rect 172563 526452 173013 526468
rect 173055 526466 173509 526482
rect 172367 526412 172433 526428
rect 173055 526432 173199 526466
rect 173233 526432 173509 526466
rect 173667 526468 173939 526502
rect 173973 526468 174117 526502
rect 174771 526502 175221 526524
rect 173667 526452 174117 526468
rect 174159 526466 174613 526482
rect 172367 526410 172405 526412
rect 173055 526410 173509 526432
rect 174159 526432 174303 526466
rect 174337 526432 174613 526466
rect 174771 526468 175043 526502
rect 175077 526468 175221 526502
rect 175875 526502 176325 526524
rect 176979 526518 177063 526524
rect 174771 526452 175221 526468
rect 175263 526466 175717 526482
rect 174159 526410 174613 526432
rect 175263 526432 175407 526466
rect 175441 526432 175717 526466
rect 175875 526468 176147 526502
rect 176181 526468 176325 526502
rect 176921 526502 177063 526518
rect 175875 526452 176325 526468
rect 176367 526466 176821 526482
rect 175263 526410 175717 526432
rect 176367 526432 176511 526466
rect 176545 526432 176821 526466
rect 176921 526468 176937 526502
rect 176971 526468 177063 526502
rect 177531 526502 177981 526524
rect 176921 526452 177063 526468
rect 177105 526466 177247 526482
rect 176367 526410 176821 526432
rect 177105 526432 177197 526466
rect 177231 526432 177247 526466
rect 177531 526468 177803 526502
rect 177837 526468 177981 526502
rect 178635 526502 179085 526524
rect 177531 526452 177981 526468
rect 178023 526466 178477 526482
rect 177105 526416 177247 526432
rect 178023 526432 178167 526466
rect 178201 526432 178477 526466
rect 178635 526468 178907 526502
rect 178941 526468 179085 526502
rect 179739 526502 180189 526524
rect 178635 526452 179085 526468
rect 179127 526466 179581 526482
rect 177105 526410 177189 526416
rect 178023 526410 178477 526432
rect 179127 526432 179271 526466
rect 179305 526432 179581 526466
rect 179739 526468 180011 526502
rect 180045 526468 180189 526502
rect 180843 526502 181293 526524
rect 179739 526452 180189 526468
rect 180231 526466 180685 526482
rect 179127 526410 179581 526432
rect 180231 526432 180375 526466
rect 180409 526432 180685 526466
rect 180843 526468 181115 526502
rect 181149 526468 181293 526502
rect 181947 526502 182123 526524
rect 180843 526452 181293 526468
rect 181335 526466 181789 526482
rect 180231 526410 180685 526432
rect 181335 526432 181479 526466
rect 181513 526432 181789 526466
rect 181947 526468 181963 526502
rect 181997 526468 182073 526502
rect 182107 526468 182123 526502
rect 182683 526502 183133 526524
rect 181947 526452 182123 526468
rect 182165 526466 182341 526482
rect 181335 526410 181789 526432
rect 182165 526432 182181 526466
rect 182215 526432 182291 526466
rect 182325 526432 182341 526466
rect 182683 526468 182955 526502
rect 182989 526468 183133 526502
rect 183787 526502 184237 526524
rect 182683 526452 183133 526468
rect 183175 526466 183629 526482
rect 182165 526410 182341 526432
rect 183175 526432 183319 526466
rect 183353 526432 183629 526466
rect 183787 526468 184059 526502
rect 184093 526468 184237 526502
rect 184891 526502 185341 526524
rect 183787 526452 184237 526468
rect 184279 526466 184733 526482
rect 183175 526410 183629 526432
rect 184279 526432 184423 526466
rect 184457 526432 184733 526466
rect 184891 526468 185163 526502
rect 185197 526468 185341 526502
rect 185995 526502 186445 526524
rect 187283 526520 187401 526550
rect 184891 526452 185341 526468
rect 185383 526466 185837 526482
rect 184279 526410 184733 526432
rect 185383 526432 185527 526466
rect 185561 526432 185837 526466
rect 185995 526468 186267 526502
rect 186301 526468 186445 526502
rect 187363 526518 187401 526520
rect 187363 526502 187429 526518
rect 185995 526452 186445 526468
rect 186487 526466 186941 526482
rect 185383 526410 185837 526432
rect 186487 526432 186631 526466
rect 186665 526432 186941 526466
rect 186487 526410 186941 526432
rect 187255 526462 187321 526478
rect 187255 526428 187271 526462
rect 187305 526428 187321 526462
rect 187363 526468 187379 526502
rect 187413 526468 187429 526502
rect 187363 526452 187429 526468
rect 187255 526412 187321 526428
rect 172287 526384 172405 526410
rect 172563 526384 173509 526410
rect 173667 526384 174613 526410
rect 174771 526384 175717 526410
rect 175875 526384 176821 526410
rect 176979 526384 177189 526410
rect 177531 526384 178477 526410
rect 178635 526384 179581 526410
rect 179739 526384 180685 526410
rect 180843 526384 181789 526410
rect 181947 526384 182341 526410
rect 182683 526384 183629 526410
rect 183787 526384 184733 526410
rect 184891 526384 185837 526410
rect 185995 526384 186941 526410
rect 187283 526410 187321 526412
rect 187283 526384 187401 526410
rect 172287 526248 172405 526274
rect 172563 526248 173509 526274
rect 173667 526248 174613 526274
rect 174771 526248 175717 526274
rect 175875 526248 176821 526274
rect 176979 526248 177189 526274
rect 177531 526248 178477 526274
rect 178635 526248 179581 526274
rect 179739 526248 180685 526274
rect 180843 526248 181789 526274
rect 181947 526248 182341 526274
rect 182683 526248 183629 526274
rect 183787 526248 184733 526274
rect 184891 526248 185837 526274
rect 185995 526248 186941 526274
rect 187283 526248 187401 526274
rect 172287 526180 172405 526206
rect 172563 526180 173509 526206
rect 173667 526180 174613 526206
rect 174955 526180 175901 526206
rect 176059 526180 177005 526206
rect 177163 526180 178109 526206
rect 178267 526180 179213 526206
rect 179371 526180 179765 526206
rect 180107 526180 181053 526206
rect 181211 526180 182157 526206
rect 182315 526180 183261 526206
rect 183419 526180 184365 526206
rect 184523 526180 184917 526206
rect 185259 526180 186205 526206
rect 186363 526180 186941 526206
rect 187283 526180 187401 526206
rect 172287 526044 172405 526070
rect 172563 526044 173509 526070
rect 173667 526044 174613 526070
rect 174955 526044 175901 526070
rect 176059 526044 177005 526070
rect 177163 526044 178109 526070
rect 178267 526044 179213 526070
rect 179371 526044 179765 526070
rect 180107 526044 181053 526070
rect 181211 526044 182157 526070
rect 182315 526044 183261 526070
rect 183419 526044 184365 526070
rect 184523 526044 184917 526070
rect 185259 526044 186205 526070
rect 186363 526044 186941 526070
rect 172367 526042 172405 526044
rect 172367 526026 172433 526042
rect 172259 525986 172325 526002
rect 172259 525952 172275 525986
rect 172309 525952 172325 525986
rect 172367 525992 172383 526026
rect 172417 525992 172433 526026
rect 173055 526022 173509 526044
rect 172367 525976 172433 525992
rect 172563 525986 173013 526002
rect 172259 525936 172325 525952
rect 172287 525934 172325 525936
rect 172563 525952 172835 525986
rect 172869 525952 173013 525986
rect 173055 525988 173199 526022
rect 173233 525988 173509 526022
rect 174159 526022 174613 526044
rect 173055 525972 173509 525988
rect 173667 525986 174117 526002
rect 172287 525904 172405 525934
rect 172563 525930 173013 525952
rect 173667 525952 173939 525986
rect 173973 525952 174117 525986
rect 174159 525988 174303 526022
rect 174337 525988 174613 526022
rect 175447 526022 175901 526044
rect 174159 525972 174613 525988
rect 174955 525986 175405 526002
rect 173667 525930 174117 525952
rect 174955 525952 175227 525986
rect 175261 525952 175405 525986
rect 175447 525988 175591 526022
rect 175625 525988 175901 526022
rect 176551 526022 177005 526044
rect 175447 525972 175901 525988
rect 176059 525986 176509 526002
rect 174955 525930 175405 525952
rect 176059 525952 176331 525986
rect 176365 525952 176509 525986
rect 176551 525988 176695 526022
rect 176729 525988 177005 526022
rect 177655 526022 178109 526044
rect 176551 525972 177005 525988
rect 177163 525986 177613 526002
rect 176059 525930 176509 525952
rect 177163 525952 177435 525986
rect 177469 525952 177613 525986
rect 177655 525988 177799 526022
rect 177833 525988 178109 526022
rect 178759 526022 179213 526044
rect 177655 525972 178109 525988
rect 178267 525986 178717 526002
rect 177163 525930 177613 525952
rect 178267 525952 178539 525986
rect 178573 525952 178717 525986
rect 178759 525988 178903 526022
rect 178937 525988 179213 526022
rect 179589 526022 179765 526044
rect 178759 525972 179213 525988
rect 179371 525986 179547 526002
rect 178267 525930 178717 525952
rect 179371 525952 179387 525986
rect 179421 525952 179497 525986
rect 179531 525952 179547 525986
rect 179589 525988 179605 526022
rect 179639 525988 179715 526022
rect 179749 525988 179765 526022
rect 180599 526022 181053 526044
rect 179589 525972 179765 525988
rect 180107 525986 180557 526002
rect 179371 525930 179547 525952
rect 180107 525952 180379 525986
rect 180413 525952 180557 525986
rect 180599 525988 180743 526022
rect 180777 525988 181053 526022
rect 181703 526022 182157 526044
rect 180599 525972 181053 525988
rect 181211 525986 181661 526002
rect 180107 525930 180557 525952
rect 181211 525952 181483 525986
rect 181517 525952 181661 525986
rect 181703 525988 181847 526022
rect 181881 525988 182157 526022
rect 182807 526022 183261 526044
rect 181703 525972 182157 525988
rect 182315 525986 182765 526002
rect 181211 525930 181661 525952
rect 182315 525952 182587 525986
rect 182621 525952 182765 525986
rect 182807 525988 182951 526022
rect 182985 525988 183261 526022
rect 183911 526022 184365 526044
rect 182807 525972 183261 525988
rect 183419 525986 183869 526002
rect 182315 525930 182765 525952
rect 183419 525952 183691 525986
rect 183725 525952 183869 525986
rect 183911 525988 184055 526022
rect 184089 525988 184365 526022
rect 184741 526022 184917 526044
rect 183911 525972 184365 525988
rect 184523 525986 184699 526002
rect 183419 525930 183869 525952
rect 184523 525952 184539 525986
rect 184573 525952 184649 525986
rect 184683 525952 184699 525986
rect 184741 525988 184757 526022
rect 184791 525988 184867 526022
rect 184901 525988 184917 526022
rect 185751 526022 186205 526044
rect 184741 525972 184917 525988
rect 185259 525986 185709 526002
rect 184523 525930 184699 525952
rect 185259 525952 185531 525986
rect 185565 525952 185709 525986
rect 185751 525988 185895 526022
rect 185929 525988 186205 526022
rect 186669 526022 186941 526044
rect 187283 526044 187401 526070
rect 187283 526042 187321 526044
rect 185751 525972 186205 525988
rect 186363 525986 186627 526002
rect 185259 525930 185709 525952
rect 186363 525952 186379 525986
rect 186413 525952 186478 525986
rect 186512 525952 186577 525986
rect 186611 525952 186627 525986
rect 186669 525988 186685 526022
rect 186719 525988 186788 526022
rect 186822 525988 186891 526022
rect 186925 525988 186941 526022
rect 186669 525972 186941 525988
rect 187255 526026 187321 526042
rect 187255 525992 187271 526026
rect 187305 525992 187321 526026
rect 187255 525976 187321 525992
rect 187363 525986 187429 526002
rect 186363 525930 186627 525952
rect 187363 525952 187379 525986
rect 187413 525952 187429 525986
rect 187363 525936 187429 525952
rect 187363 525934 187401 525936
rect 172563 525904 173509 525930
rect 173667 525904 174613 525930
rect 174955 525904 175901 525930
rect 176059 525904 177005 525930
rect 177163 525904 178109 525930
rect 178267 525904 179213 525930
rect 179371 525904 179765 525930
rect 180107 525904 181053 525930
rect 181211 525904 182157 525930
rect 182315 525904 183261 525930
rect 183419 525904 184365 525930
rect 184523 525904 184917 525930
rect 185259 525904 186205 525930
rect 186363 525904 186941 525930
rect 187283 525904 187401 525934
rect 172287 525704 172405 525730
rect 172563 525704 173509 525730
rect 173667 525704 174613 525730
rect 174955 525704 175901 525730
rect 176059 525704 177005 525730
rect 177163 525704 178109 525730
rect 178267 525704 179213 525730
rect 179371 525704 179765 525730
rect 180107 525704 181053 525730
rect 181211 525704 182157 525730
rect 182315 525704 183261 525730
rect 183419 525704 184365 525730
rect 184523 525704 184917 525730
rect 185259 525704 186205 525730
rect 186363 525704 186941 525730
rect 187283 525704 187401 525730
rect 172287 525636 172405 525662
rect 172563 525636 173509 525662
rect 173667 525636 174613 525662
rect 174771 525636 175717 525662
rect 175875 525636 176821 525662
rect 176979 525636 177189 525662
rect 177531 525636 178477 525662
rect 178635 525636 179581 525662
rect 179739 525636 180685 525662
rect 180843 525636 181789 525662
rect 181947 525636 182341 525662
rect 182683 525636 183629 525662
rect 183787 525636 184733 525662
rect 184891 525636 185837 525662
rect 185995 525636 186941 525662
rect 187283 525636 187401 525662
rect 172287 525432 172405 525462
rect 172563 525436 173509 525462
rect 173667 525436 174613 525462
rect 174771 525436 175717 525462
rect 175875 525436 176821 525462
rect 176979 525436 177189 525462
rect 177531 525436 178477 525462
rect 178635 525436 179581 525462
rect 179739 525436 180685 525462
rect 180843 525436 181789 525462
rect 181947 525436 182341 525462
rect 182683 525436 183629 525462
rect 183787 525436 184733 525462
rect 184891 525436 185837 525462
rect 185995 525436 186941 525462
rect 172287 525430 172325 525432
rect 172259 525414 172325 525430
rect 172259 525380 172275 525414
rect 172309 525380 172325 525414
rect 172563 525414 173013 525436
rect 172259 525364 172325 525380
rect 172367 525374 172433 525390
rect 172367 525340 172383 525374
rect 172417 525340 172433 525374
rect 172563 525380 172835 525414
rect 172869 525380 173013 525414
rect 173667 525414 174117 525436
rect 172563 525364 173013 525380
rect 173055 525378 173509 525394
rect 172367 525324 172433 525340
rect 173055 525344 173199 525378
rect 173233 525344 173509 525378
rect 173667 525380 173939 525414
rect 173973 525380 174117 525414
rect 174771 525414 175221 525436
rect 173667 525364 174117 525380
rect 174159 525378 174613 525394
rect 172367 525322 172405 525324
rect 173055 525322 173509 525344
rect 174159 525344 174303 525378
rect 174337 525344 174613 525378
rect 174771 525380 175043 525414
rect 175077 525380 175221 525414
rect 175875 525414 176325 525436
rect 176979 525430 177063 525436
rect 174771 525364 175221 525380
rect 175263 525378 175717 525394
rect 174159 525322 174613 525344
rect 175263 525344 175407 525378
rect 175441 525344 175717 525378
rect 175875 525380 176147 525414
rect 176181 525380 176325 525414
rect 176921 525414 177063 525430
rect 175875 525364 176325 525380
rect 176367 525378 176821 525394
rect 175263 525322 175717 525344
rect 176367 525344 176511 525378
rect 176545 525344 176821 525378
rect 176921 525380 176937 525414
rect 176971 525380 177063 525414
rect 177531 525414 177981 525436
rect 176921 525364 177063 525380
rect 177105 525378 177247 525394
rect 176367 525322 176821 525344
rect 177105 525344 177197 525378
rect 177231 525344 177247 525378
rect 177531 525380 177803 525414
rect 177837 525380 177981 525414
rect 178635 525414 179085 525436
rect 177531 525364 177981 525380
rect 178023 525378 178477 525394
rect 177105 525328 177247 525344
rect 178023 525344 178167 525378
rect 178201 525344 178477 525378
rect 178635 525380 178907 525414
rect 178941 525380 179085 525414
rect 179739 525414 180189 525436
rect 178635 525364 179085 525380
rect 179127 525378 179581 525394
rect 177105 525322 177189 525328
rect 178023 525322 178477 525344
rect 179127 525344 179271 525378
rect 179305 525344 179581 525378
rect 179739 525380 180011 525414
rect 180045 525380 180189 525414
rect 180843 525414 181293 525436
rect 179739 525364 180189 525380
rect 180231 525378 180685 525394
rect 179127 525322 179581 525344
rect 180231 525344 180375 525378
rect 180409 525344 180685 525378
rect 180843 525380 181115 525414
rect 181149 525380 181293 525414
rect 181947 525414 182123 525436
rect 180843 525364 181293 525380
rect 181335 525378 181789 525394
rect 180231 525322 180685 525344
rect 181335 525344 181479 525378
rect 181513 525344 181789 525378
rect 181947 525380 181963 525414
rect 181997 525380 182073 525414
rect 182107 525380 182123 525414
rect 182683 525414 183133 525436
rect 181947 525364 182123 525380
rect 182165 525378 182341 525394
rect 181335 525322 181789 525344
rect 182165 525344 182181 525378
rect 182215 525344 182291 525378
rect 182325 525344 182341 525378
rect 182683 525380 182955 525414
rect 182989 525380 183133 525414
rect 183787 525414 184237 525436
rect 182683 525364 183133 525380
rect 183175 525378 183629 525394
rect 182165 525322 182341 525344
rect 183175 525344 183319 525378
rect 183353 525344 183629 525378
rect 183787 525380 184059 525414
rect 184093 525380 184237 525414
rect 184891 525414 185341 525436
rect 183787 525364 184237 525380
rect 184279 525378 184733 525394
rect 183175 525322 183629 525344
rect 184279 525344 184423 525378
rect 184457 525344 184733 525378
rect 184891 525380 185163 525414
rect 185197 525380 185341 525414
rect 185995 525414 186445 525436
rect 187283 525432 187401 525462
rect 184891 525364 185341 525380
rect 185383 525378 185837 525394
rect 184279 525322 184733 525344
rect 185383 525344 185527 525378
rect 185561 525344 185837 525378
rect 185995 525380 186267 525414
rect 186301 525380 186445 525414
rect 187363 525430 187401 525432
rect 187363 525414 187429 525430
rect 185995 525364 186445 525380
rect 186487 525378 186941 525394
rect 185383 525322 185837 525344
rect 186487 525344 186631 525378
rect 186665 525344 186941 525378
rect 186487 525322 186941 525344
rect 187255 525374 187321 525390
rect 187255 525340 187271 525374
rect 187305 525340 187321 525374
rect 187363 525380 187379 525414
rect 187413 525380 187429 525414
rect 187363 525364 187429 525380
rect 187255 525324 187321 525340
rect 172287 525296 172405 525322
rect 172563 525296 173509 525322
rect 173667 525296 174613 525322
rect 174771 525296 175717 525322
rect 175875 525296 176821 525322
rect 176979 525296 177189 525322
rect 177531 525296 178477 525322
rect 178635 525296 179581 525322
rect 179739 525296 180685 525322
rect 180843 525296 181789 525322
rect 181947 525296 182341 525322
rect 182683 525296 183629 525322
rect 183787 525296 184733 525322
rect 184891 525296 185837 525322
rect 185995 525296 186941 525322
rect 187283 525322 187321 525324
rect 187283 525296 187401 525322
rect 172287 525160 172405 525186
rect 172563 525160 173509 525186
rect 173667 525160 174613 525186
rect 174771 525160 175717 525186
rect 175875 525160 176821 525186
rect 176979 525160 177189 525186
rect 177531 525160 178477 525186
rect 178635 525160 179581 525186
rect 179739 525160 180685 525186
rect 180843 525160 181789 525186
rect 181947 525160 182341 525186
rect 182683 525160 183629 525186
rect 183787 525160 184733 525186
rect 184891 525160 185837 525186
rect 185995 525160 186941 525186
rect 187283 525160 187401 525186
rect 172287 525092 172405 525118
rect 172563 525092 173509 525118
rect 173667 525092 174613 525118
rect 174955 525092 175901 525118
rect 176059 525092 177005 525118
rect 177163 525092 178109 525118
rect 178267 525092 179213 525118
rect 179371 525092 179765 525118
rect 180107 525092 181053 525118
rect 181211 525092 182157 525118
rect 182315 525092 183261 525118
rect 183419 525092 184365 525118
rect 184523 525092 184917 525118
rect 185259 525092 186205 525118
rect 186363 525092 186941 525118
rect 187283 525092 187401 525118
rect 172287 524956 172405 524982
rect 172563 524956 173509 524982
rect 173667 524956 174613 524982
rect 174955 524956 175901 524982
rect 176059 524956 177005 524982
rect 177163 524956 178109 524982
rect 178267 524956 179213 524982
rect 179371 524956 179765 524982
rect 180107 524956 181053 524982
rect 181211 524956 182157 524982
rect 182315 524956 183261 524982
rect 183419 524956 184365 524982
rect 184523 524956 184917 524982
rect 185259 524956 186205 524982
rect 186363 524956 186941 524982
rect 172367 524954 172405 524956
rect 172367 524938 172433 524954
rect 172259 524898 172325 524914
rect 172259 524864 172275 524898
rect 172309 524864 172325 524898
rect 172367 524904 172383 524938
rect 172417 524904 172433 524938
rect 173055 524934 173509 524956
rect 172367 524888 172433 524904
rect 172563 524898 173013 524914
rect 172259 524848 172325 524864
rect 172287 524846 172325 524848
rect 172563 524864 172835 524898
rect 172869 524864 173013 524898
rect 173055 524900 173199 524934
rect 173233 524900 173509 524934
rect 174159 524934 174613 524956
rect 173055 524884 173509 524900
rect 173667 524898 174117 524914
rect 172287 524816 172405 524846
rect 172563 524842 173013 524864
rect 173667 524864 173939 524898
rect 173973 524864 174117 524898
rect 174159 524900 174303 524934
rect 174337 524900 174613 524934
rect 175447 524934 175901 524956
rect 174159 524884 174613 524900
rect 174955 524898 175405 524914
rect 173667 524842 174117 524864
rect 174955 524864 175227 524898
rect 175261 524864 175405 524898
rect 175447 524900 175591 524934
rect 175625 524900 175901 524934
rect 176551 524934 177005 524956
rect 175447 524884 175901 524900
rect 176059 524898 176509 524914
rect 174955 524842 175405 524864
rect 176059 524864 176331 524898
rect 176365 524864 176509 524898
rect 176551 524900 176695 524934
rect 176729 524900 177005 524934
rect 177655 524934 178109 524956
rect 176551 524884 177005 524900
rect 177163 524898 177613 524914
rect 176059 524842 176509 524864
rect 177163 524864 177435 524898
rect 177469 524864 177613 524898
rect 177655 524900 177799 524934
rect 177833 524900 178109 524934
rect 178759 524934 179213 524956
rect 177655 524884 178109 524900
rect 178267 524898 178717 524914
rect 177163 524842 177613 524864
rect 178267 524864 178539 524898
rect 178573 524864 178717 524898
rect 178759 524900 178903 524934
rect 178937 524900 179213 524934
rect 179589 524934 179765 524956
rect 178759 524884 179213 524900
rect 179371 524898 179547 524914
rect 178267 524842 178717 524864
rect 179371 524864 179387 524898
rect 179421 524864 179497 524898
rect 179531 524864 179547 524898
rect 179589 524900 179605 524934
rect 179639 524900 179715 524934
rect 179749 524900 179765 524934
rect 180599 524934 181053 524956
rect 179589 524884 179765 524900
rect 180107 524898 180557 524914
rect 179371 524842 179547 524864
rect 180107 524864 180379 524898
rect 180413 524864 180557 524898
rect 180599 524900 180743 524934
rect 180777 524900 181053 524934
rect 181703 524934 182157 524956
rect 180599 524884 181053 524900
rect 181211 524898 181661 524914
rect 180107 524842 180557 524864
rect 181211 524864 181483 524898
rect 181517 524864 181661 524898
rect 181703 524900 181847 524934
rect 181881 524900 182157 524934
rect 182807 524934 183261 524956
rect 181703 524884 182157 524900
rect 182315 524898 182765 524914
rect 181211 524842 181661 524864
rect 182315 524864 182587 524898
rect 182621 524864 182765 524898
rect 182807 524900 182951 524934
rect 182985 524900 183261 524934
rect 183911 524934 184365 524956
rect 182807 524884 183261 524900
rect 183419 524898 183869 524914
rect 182315 524842 182765 524864
rect 183419 524864 183691 524898
rect 183725 524864 183869 524898
rect 183911 524900 184055 524934
rect 184089 524900 184365 524934
rect 184741 524934 184917 524956
rect 183911 524884 184365 524900
rect 184523 524898 184699 524914
rect 183419 524842 183869 524864
rect 184523 524864 184539 524898
rect 184573 524864 184649 524898
rect 184683 524864 184699 524898
rect 184741 524900 184757 524934
rect 184791 524900 184867 524934
rect 184901 524900 184917 524934
rect 185751 524934 186205 524956
rect 184741 524884 184917 524900
rect 185259 524898 185709 524914
rect 184523 524842 184699 524864
rect 185259 524864 185531 524898
rect 185565 524864 185709 524898
rect 185751 524900 185895 524934
rect 185929 524900 186205 524934
rect 186669 524934 186941 524956
rect 187283 524956 187401 524982
rect 187283 524954 187321 524956
rect 185751 524884 186205 524900
rect 186363 524898 186627 524914
rect 185259 524842 185709 524864
rect 186363 524864 186379 524898
rect 186413 524864 186478 524898
rect 186512 524864 186577 524898
rect 186611 524864 186627 524898
rect 186669 524900 186685 524934
rect 186719 524900 186788 524934
rect 186822 524900 186891 524934
rect 186925 524900 186941 524934
rect 186669 524884 186941 524900
rect 187255 524938 187321 524954
rect 187255 524904 187271 524938
rect 187305 524904 187321 524938
rect 187255 524888 187321 524904
rect 187363 524898 187429 524914
rect 186363 524842 186627 524864
rect 187363 524864 187379 524898
rect 187413 524864 187429 524898
rect 187363 524848 187429 524864
rect 187363 524846 187401 524848
rect 172563 524816 173509 524842
rect 173667 524816 174613 524842
rect 174955 524816 175901 524842
rect 176059 524816 177005 524842
rect 177163 524816 178109 524842
rect 178267 524816 179213 524842
rect 179371 524816 179765 524842
rect 180107 524816 181053 524842
rect 181211 524816 182157 524842
rect 182315 524816 183261 524842
rect 183419 524816 184365 524842
rect 184523 524816 184917 524842
rect 185259 524816 186205 524842
rect 186363 524816 186941 524842
rect 187283 524816 187401 524846
rect 172287 524616 172405 524642
rect 172563 524616 173509 524642
rect 173667 524616 174613 524642
rect 174955 524616 175901 524642
rect 176059 524616 177005 524642
rect 177163 524616 178109 524642
rect 178267 524616 179213 524642
rect 179371 524616 179765 524642
rect 180107 524616 181053 524642
rect 181211 524616 182157 524642
rect 182315 524616 183261 524642
rect 183419 524616 184365 524642
rect 184523 524616 184917 524642
rect 185259 524616 186205 524642
rect 186363 524616 186941 524642
rect 187283 524616 187401 524642
rect 172287 524548 172405 524574
rect 172563 524548 173509 524574
rect 173667 524548 174613 524574
rect 174771 524548 175717 524574
rect 175875 524548 176821 524574
rect 176979 524548 177189 524574
rect 177531 524548 178477 524574
rect 178635 524548 179581 524574
rect 179739 524548 180685 524574
rect 180843 524548 181789 524574
rect 181947 524548 182341 524574
rect 182683 524548 183629 524574
rect 183787 524548 184733 524574
rect 184891 524548 185837 524574
rect 185995 524548 186941 524574
rect 187283 524548 187401 524574
rect 172287 524344 172405 524374
rect 172563 524348 173509 524374
rect 173667 524348 174613 524374
rect 174771 524348 175717 524374
rect 175875 524348 176821 524374
rect 176979 524348 177189 524374
rect 177531 524348 178477 524374
rect 178635 524348 179581 524374
rect 179739 524348 180685 524374
rect 180843 524348 181789 524374
rect 181947 524348 182341 524374
rect 182683 524348 183629 524374
rect 183787 524348 184733 524374
rect 184891 524348 185837 524374
rect 185995 524348 186941 524374
rect 172287 524342 172325 524344
rect 172259 524326 172325 524342
rect 172259 524292 172275 524326
rect 172309 524292 172325 524326
rect 172563 524326 173013 524348
rect 172259 524276 172325 524292
rect 172367 524286 172433 524302
rect 172367 524252 172383 524286
rect 172417 524252 172433 524286
rect 172563 524292 172835 524326
rect 172869 524292 173013 524326
rect 173667 524326 174117 524348
rect 172563 524276 173013 524292
rect 173055 524290 173509 524306
rect 172367 524236 172433 524252
rect 173055 524256 173199 524290
rect 173233 524256 173509 524290
rect 173667 524292 173939 524326
rect 173973 524292 174117 524326
rect 174771 524326 175221 524348
rect 173667 524276 174117 524292
rect 174159 524290 174613 524306
rect 172367 524234 172405 524236
rect 173055 524234 173509 524256
rect 174159 524256 174303 524290
rect 174337 524256 174613 524290
rect 174771 524292 175043 524326
rect 175077 524292 175221 524326
rect 175875 524326 176325 524348
rect 176979 524342 177063 524348
rect 174771 524276 175221 524292
rect 175263 524290 175717 524306
rect 174159 524234 174613 524256
rect 175263 524256 175407 524290
rect 175441 524256 175717 524290
rect 175875 524292 176147 524326
rect 176181 524292 176325 524326
rect 176921 524326 177063 524342
rect 175875 524276 176325 524292
rect 176367 524290 176821 524306
rect 175263 524234 175717 524256
rect 176367 524256 176511 524290
rect 176545 524256 176821 524290
rect 176921 524292 176937 524326
rect 176971 524292 177063 524326
rect 177531 524326 177981 524348
rect 176921 524276 177063 524292
rect 177105 524290 177247 524306
rect 176367 524234 176821 524256
rect 177105 524256 177197 524290
rect 177231 524256 177247 524290
rect 177531 524292 177803 524326
rect 177837 524292 177981 524326
rect 178635 524326 179085 524348
rect 177531 524276 177981 524292
rect 178023 524290 178477 524306
rect 177105 524240 177247 524256
rect 178023 524256 178167 524290
rect 178201 524256 178477 524290
rect 178635 524292 178907 524326
rect 178941 524292 179085 524326
rect 179739 524326 180189 524348
rect 178635 524276 179085 524292
rect 179127 524290 179581 524306
rect 177105 524234 177189 524240
rect 178023 524234 178477 524256
rect 179127 524256 179271 524290
rect 179305 524256 179581 524290
rect 179739 524292 180011 524326
rect 180045 524292 180189 524326
rect 180843 524326 181293 524348
rect 179739 524276 180189 524292
rect 180231 524290 180685 524306
rect 179127 524234 179581 524256
rect 180231 524256 180375 524290
rect 180409 524256 180685 524290
rect 180843 524292 181115 524326
rect 181149 524292 181293 524326
rect 181947 524326 182123 524348
rect 180843 524276 181293 524292
rect 181335 524290 181789 524306
rect 180231 524234 180685 524256
rect 181335 524256 181479 524290
rect 181513 524256 181789 524290
rect 181947 524292 181963 524326
rect 181997 524292 182073 524326
rect 182107 524292 182123 524326
rect 182683 524326 183133 524348
rect 181947 524276 182123 524292
rect 182165 524290 182341 524306
rect 181335 524234 181789 524256
rect 182165 524256 182181 524290
rect 182215 524256 182291 524290
rect 182325 524256 182341 524290
rect 182683 524292 182955 524326
rect 182989 524292 183133 524326
rect 183787 524326 184237 524348
rect 182683 524276 183133 524292
rect 183175 524290 183629 524306
rect 182165 524234 182341 524256
rect 183175 524256 183319 524290
rect 183353 524256 183629 524290
rect 183787 524292 184059 524326
rect 184093 524292 184237 524326
rect 184891 524326 185341 524348
rect 183787 524276 184237 524292
rect 184279 524290 184733 524306
rect 183175 524234 183629 524256
rect 184279 524256 184423 524290
rect 184457 524256 184733 524290
rect 184891 524292 185163 524326
rect 185197 524292 185341 524326
rect 185995 524326 186445 524348
rect 187283 524344 187401 524374
rect 184891 524276 185341 524292
rect 185383 524290 185837 524306
rect 184279 524234 184733 524256
rect 185383 524256 185527 524290
rect 185561 524256 185837 524290
rect 185995 524292 186267 524326
rect 186301 524292 186445 524326
rect 187363 524342 187401 524344
rect 187363 524326 187429 524342
rect 185995 524276 186445 524292
rect 186487 524290 186941 524306
rect 185383 524234 185837 524256
rect 186487 524256 186631 524290
rect 186665 524256 186941 524290
rect 186487 524234 186941 524256
rect 187255 524286 187321 524302
rect 187255 524252 187271 524286
rect 187305 524252 187321 524286
rect 187363 524292 187379 524326
rect 187413 524292 187429 524326
rect 187363 524276 187429 524292
rect 187255 524236 187321 524252
rect 172287 524208 172405 524234
rect 172563 524208 173509 524234
rect 173667 524208 174613 524234
rect 174771 524208 175717 524234
rect 175875 524208 176821 524234
rect 176979 524208 177189 524234
rect 177531 524208 178477 524234
rect 178635 524208 179581 524234
rect 179739 524208 180685 524234
rect 180843 524208 181789 524234
rect 181947 524208 182341 524234
rect 182683 524208 183629 524234
rect 183787 524208 184733 524234
rect 184891 524208 185837 524234
rect 185995 524208 186941 524234
rect 187283 524234 187321 524236
rect 187283 524208 187401 524234
rect 172287 524072 172405 524098
rect 172563 524072 173509 524098
rect 173667 524072 174613 524098
rect 174771 524072 175717 524098
rect 175875 524072 176821 524098
rect 176979 524072 177189 524098
rect 177531 524072 178477 524098
rect 178635 524072 179581 524098
rect 179739 524072 180685 524098
rect 180843 524072 181789 524098
rect 181947 524072 182341 524098
rect 182683 524072 183629 524098
rect 183787 524072 184733 524098
rect 184891 524072 185837 524098
rect 185995 524072 186941 524098
rect 187283 524072 187401 524098
rect 172287 524004 172405 524030
rect 172563 524004 173509 524030
rect 173667 524004 174613 524030
rect 174955 524004 175901 524030
rect 176059 524004 177005 524030
rect 177163 524004 178109 524030
rect 178267 524004 179213 524030
rect 179371 524004 179765 524030
rect 180107 524004 181053 524030
rect 181211 524004 182157 524030
rect 182315 524004 183261 524030
rect 183419 524004 184365 524030
rect 184523 524004 184917 524030
rect 185259 524004 186205 524030
rect 186363 524004 186941 524030
rect 187283 524004 187401 524030
rect 172287 523868 172405 523894
rect 172563 523868 173509 523894
rect 173667 523868 174613 523894
rect 174955 523868 175901 523894
rect 176059 523868 177005 523894
rect 177163 523868 178109 523894
rect 178267 523868 179213 523894
rect 179371 523868 179765 523894
rect 180107 523868 181053 523894
rect 181211 523868 182157 523894
rect 182315 523868 183261 523894
rect 183419 523868 184365 523894
rect 184523 523868 184917 523894
rect 185259 523868 186205 523894
rect 186363 523868 186941 523894
rect 172367 523866 172405 523868
rect 172367 523850 172433 523866
rect 172259 523810 172325 523826
rect 172259 523776 172275 523810
rect 172309 523776 172325 523810
rect 172367 523816 172383 523850
rect 172417 523816 172433 523850
rect 173055 523846 173509 523868
rect 172367 523800 172433 523816
rect 172563 523810 173013 523826
rect 172259 523760 172325 523776
rect 172287 523758 172325 523760
rect 172563 523776 172835 523810
rect 172869 523776 173013 523810
rect 173055 523812 173199 523846
rect 173233 523812 173509 523846
rect 174159 523846 174613 523868
rect 173055 523796 173509 523812
rect 173667 523810 174117 523826
rect 172287 523728 172405 523758
rect 172563 523754 173013 523776
rect 173667 523776 173939 523810
rect 173973 523776 174117 523810
rect 174159 523812 174303 523846
rect 174337 523812 174613 523846
rect 175447 523846 175901 523868
rect 174159 523796 174613 523812
rect 174955 523810 175405 523826
rect 173667 523754 174117 523776
rect 174955 523776 175227 523810
rect 175261 523776 175405 523810
rect 175447 523812 175591 523846
rect 175625 523812 175901 523846
rect 176551 523846 177005 523868
rect 175447 523796 175901 523812
rect 176059 523810 176509 523826
rect 174955 523754 175405 523776
rect 176059 523776 176331 523810
rect 176365 523776 176509 523810
rect 176551 523812 176695 523846
rect 176729 523812 177005 523846
rect 177655 523846 178109 523868
rect 176551 523796 177005 523812
rect 177163 523810 177613 523826
rect 176059 523754 176509 523776
rect 177163 523776 177435 523810
rect 177469 523776 177613 523810
rect 177655 523812 177799 523846
rect 177833 523812 178109 523846
rect 178759 523846 179213 523868
rect 177655 523796 178109 523812
rect 178267 523810 178717 523826
rect 177163 523754 177613 523776
rect 178267 523776 178539 523810
rect 178573 523776 178717 523810
rect 178759 523812 178903 523846
rect 178937 523812 179213 523846
rect 179589 523846 179765 523868
rect 178759 523796 179213 523812
rect 179371 523810 179547 523826
rect 178267 523754 178717 523776
rect 179371 523776 179387 523810
rect 179421 523776 179497 523810
rect 179531 523776 179547 523810
rect 179589 523812 179605 523846
rect 179639 523812 179715 523846
rect 179749 523812 179765 523846
rect 180599 523846 181053 523868
rect 179589 523796 179765 523812
rect 180107 523810 180557 523826
rect 179371 523754 179547 523776
rect 180107 523776 180379 523810
rect 180413 523776 180557 523810
rect 180599 523812 180743 523846
rect 180777 523812 181053 523846
rect 181703 523846 182157 523868
rect 180599 523796 181053 523812
rect 181211 523810 181661 523826
rect 180107 523754 180557 523776
rect 181211 523776 181483 523810
rect 181517 523776 181661 523810
rect 181703 523812 181847 523846
rect 181881 523812 182157 523846
rect 182807 523846 183261 523868
rect 181703 523796 182157 523812
rect 182315 523810 182765 523826
rect 181211 523754 181661 523776
rect 182315 523776 182587 523810
rect 182621 523776 182765 523810
rect 182807 523812 182951 523846
rect 182985 523812 183261 523846
rect 183911 523846 184365 523868
rect 182807 523796 183261 523812
rect 183419 523810 183869 523826
rect 182315 523754 182765 523776
rect 183419 523776 183691 523810
rect 183725 523776 183869 523810
rect 183911 523812 184055 523846
rect 184089 523812 184365 523846
rect 184741 523846 184917 523868
rect 183911 523796 184365 523812
rect 184523 523810 184699 523826
rect 183419 523754 183869 523776
rect 184523 523776 184539 523810
rect 184573 523776 184649 523810
rect 184683 523776 184699 523810
rect 184741 523812 184757 523846
rect 184791 523812 184867 523846
rect 184901 523812 184917 523846
rect 185751 523846 186205 523868
rect 184741 523796 184917 523812
rect 185259 523810 185709 523826
rect 184523 523754 184699 523776
rect 185259 523776 185531 523810
rect 185565 523776 185709 523810
rect 185751 523812 185895 523846
rect 185929 523812 186205 523846
rect 186669 523846 186941 523868
rect 187283 523868 187401 523894
rect 187283 523866 187321 523868
rect 185751 523796 186205 523812
rect 186363 523810 186627 523826
rect 185259 523754 185709 523776
rect 186363 523776 186379 523810
rect 186413 523776 186478 523810
rect 186512 523776 186577 523810
rect 186611 523776 186627 523810
rect 186669 523812 186685 523846
rect 186719 523812 186788 523846
rect 186822 523812 186891 523846
rect 186925 523812 186941 523846
rect 186669 523796 186941 523812
rect 187255 523850 187321 523866
rect 187255 523816 187271 523850
rect 187305 523816 187321 523850
rect 187255 523800 187321 523816
rect 187363 523810 187429 523826
rect 186363 523754 186627 523776
rect 187363 523776 187379 523810
rect 187413 523776 187429 523810
rect 187363 523760 187429 523776
rect 187363 523758 187401 523760
rect 172563 523728 173509 523754
rect 173667 523728 174613 523754
rect 174955 523728 175901 523754
rect 176059 523728 177005 523754
rect 177163 523728 178109 523754
rect 178267 523728 179213 523754
rect 179371 523728 179765 523754
rect 180107 523728 181053 523754
rect 181211 523728 182157 523754
rect 182315 523728 183261 523754
rect 183419 523728 184365 523754
rect 184523 523728 184917 523754
rect 185259 523728 186205 523754
rect 186363 523728 186941 523754
rect 187283 523728 187401 523758
rect 172287 523528 172405 523554
rect 172563 523528 173509 523554
rect 173667 523528 174613 523554
rect 174955 523528 175901 523554
rect 176059 523528 177005 523554
rect 177163 523528 178109 523554
rect 178267 523528 179213 523554
rect 179371 523528 179765 523554
rect 180107 523528 181053 523554
rect 181211 523528 182157 523554
rect 182315 523528 183261 523554
rect 183419 523528 184365 523554
rect 184523 523528 184917 523554
rect 185259 523528 186205 523554
rect 186363 523528 186941 523554
rect 187283 523528 187401 523554
rect 172287 523460 172405 523486
rect 172563 523460 173509 523486
rect 173667 523460 174613 523486
rect 174771 523460 175717 523486
rect 175875 523460 176821 523486
rect 176979 523460 177189 523486
rect 177531 523460 178477 523486
rect 178635 523460 179581 523486
rect 179739 523460 180685 523486
rect 180843 523460 181789 523486
rect 181947 523460 182341 523486
rect 182683 523460 183629 523486
rect 183787 523460 184733 523486
rect 184891 523460 185837 523486
rect 185995 523460 186941 523486
rect 187283 523460 187401 523486
rect 172287 523256 172405 523286
rect 172563 523260 173509 523286
rect 173667 523260 174613 523286
rect 174771 523260 175717 523286
rect 175875 523260 176821 523286
rect 176979 523260 177189 523286
rect 177531 523260 178477 523286
rect 178635 523260 179581 523286
rect 179739 523260 180685 523286
rect 180843 523260 181789 523286
rect 181947 523260 182341 523286
rect 182683 523260 183629 523286
rect 183787 523260 184733 523286
rect 184891 523260 185837 523286
rect 185995 523260 186941 523286
rect 172287 523254 172325 523256
rect 172259 523238 172325 523254
rect 172259 523204 172275 523238
rect 172309 523204 172325 523238
rect 172563 523238 173013 523260
rect 172259 523188 172325 523204
rect 172367 523198 172433 523214
rect 172367 523164 172383 523198
rect 172417 523164 172433 523198
rect 172563 523204 172835 523238
rect 172869 523204 173013 523238
rect 173667 523238 174117 523260
rect 172563 523188 173013 523204
rect 173055 523202 173509 523218
rect 172367 523148 172433 523164
rect 173055 523168 173199 523202
rect 173233 523168 173509 523202
rect 173667 523204 173939 523238
rect 173973 523204 174117 523238
rect 174771 523238 175221 523260
rect 173667 523188 174117 523204
rect 174159 523202 174613 523218
rect 172367 523146 172405 523148
rect 173055 523146 173509 523168
rect 174159 523168 174303 523202
rect 174337 523168 174613 523202
rect 174771 523204 175043 523238
rect 175077 523204 175221 523238
rect 175875 523238 176325 523260
rect 176979 523254 177063 523260
rect 174771 523188 175221 523204
rect 175263 523202 175717 523218
rect 174159 523146 174613 523168
rect 175263 523168 175407 523202
rect 175441 523168 175717 523202
rect 175875 523204 176147 523238
rect 176181 523204 176325 523238
rect 176921 523238 177063 523254
rect 175875 523188 176325 523204
rect 176367 523202 176821 523218
rect 175263 523146 175717 523168
rect 176367 523168 176511 523202
rect 176545 523168 176821 523202
rect 176921 523204 176937 523238
rect 176971 523204 177063 523238
rect 177531 523238 177981 523260
rect 176921 523188 177063 523204
rect 177105 523202 177247 523218
rect 176367 523146 176821 523168
rect 177105 523168 177197 523202
rect 177231 523168 177247 523202
rect 177531 523204 177803 523238
rect 177837 523204 177981 523238
rect 178635 523238 179085 523260
rect 177531 523188 177981 523204
rect 178023 523202 178477 523218
rect 177105 523152 177247 523168
rect 178023 523168 178167 523202
rect 178201 523168 178477 523202
rect 178635 523204 178907 523238
rect 178941 523204 179085 523238
rect 179739 523238 180189 523260
rect 178635 523188 179085 523204
rect 179127 523202 179581 523218
rect 177105 523146 177189 523152
rect 178023 523146 178477 523168
rect 179127 523168 179271 523202
rect 179305 523168 179581 523202
rect 179739 523204 180011 523238
rect 180045 523204 180189 523238
rect 180843 523238 181293 523260
rect 179739 523188 180189 523204
rect 180231 523202 180685 523218
rect 179127 523146 179581 523168
rect 180231 523168 180375 523202
rect 180409 523168 180685 523202
rect 180843 523204 181115 523238
rect 181149 523204 181293 523238
rect 181947 523238 182123 523260
rect 180843 523188 181293 523204
rect 181335 523202 181789 523218
rect 180231 523146 180685 523168
rect 181335 523168 181479 523202
rect 181513 523168 181789 523202
rect 181947 523204 181963 523238
rect 181997 523204 182073 523238
rect 182107 523204 182123 523238
rect 182683 523238 183133 523260
rect 181947 523188 182123 523204
rect 182165 523202 182341 523218
rect 181335 523146 181789 523168
rect 182165 523168 182181 523202
rect 182215 523168 182291 523202
rect 182325 523168 182341 523202
rect 182683 523204 182955 523238
rect 182989 523204 183133 523238
rect 183787 523238 184237 523260
rect 182683 523188 183133 523204
rect 183175 523202 183629 523218
rect 182165 523146 182341 523168
rect 183175 523168 183319 523202
rect 183353 523168 183629 523202
rect 183787 523204 184059 523238
rect 184093 523204 184237 523238
rect 184891 523238 185341 523260
rect 183787 523188 184237 523204
rect 184279 523202 184733 523218
rect 183175 523146 183629 523168
rect 184279 523168 184423 523202
rect 184457 523168 184733 523202
rect 184891 523204 185163 523238
rect 185197 523204 185341 523238
rect 185995 523238 186445 523260
rect 187283 523256 187401 523286
rect 184891 523188 185341 523204
rect 185383 523202 185837 523218
rect 184279 523146 184733 523168
rect 185383 523168 185527 523202
rect 185561 523168 185837 523202
rect 185995 523204 186267 523238
rect 186301 523204 186445 523238
rect 187363 523254 187401 523256
rect 187363 523238 187429 523254
rect 185995 523188 186445 523204
rect 186487 523202 186941 523218
rect 185383 523146 185837 523168
rect 186487 523168 186631 523202
rect 186665 523168 186941 523202
rect 186487 523146 186941 523168
rect 187255 523198 187321 523214
rect 187255 523164 187271 523198
rect 187305 523164 187321 523198
rect 187363 523204 187379 523238
rect 187413 523204 187429 523238
rect 187363 523188 187429 523204
rect 187255 523148 187321 523164
rect 172287 523120 172405 523146
rect 172563 523120 173509 523146
rect 173667 523120 174613 523146
rect 174771 523120 175717 523146
rect 175875 523120 176821 523146
rect 176979 523120 177189 523146
rect 177531 523120 178477 523146
rect 178635 523120 179581 523146
rect 179739 523120 180685 523146
rect 180843 523120 181789 523146
rect 181947 523120 182341 523146
rect 182683 523120 183629 523146
rect 183787 523120 184733 523146
rect 184891 523120 185837 523146
rect 185995 523120 186941 523146
rect 187283 523146 187321 523148
rect 187283 523120 187401 523146
rect 172287 522984 172405 523010
rect 172563 522984 173509 523010
rect 173667 522984 174613 523010
rect 174771 522984 175717 523010
rect 175875 522984 176821 523010
rect 176979 522984 177189 523010
rect 177531 522984 178477 523010
rect 178635 522984 179581 523010
rect 179739 522984 180685 523010
rect 180843 522984 181789 523010
rect 181947 522984 182341 523010
rect 182683 522984 183629 523010
rect 183787 522984 184733 523010
rect 184891 522984 185837 523010
rect 185995 522984 186941 523010
rect 187283 522984 187401 523010
rect 172287 522916 172405 522942
rect 172563 522916 173509 522942
rect 173667 522916 174613 522942
rect 174955 522916 175901 522942
rect 176059 522916 177005 522942
rect 177163 522916 178109 522942
rect 178267 522916 179213 522942
rect 179371 522916 179765 522942
rect 180107 522916 181053 522942
rect 181211 522916 182157 522942
rect 182315 522916 183261 522942
rect 183419 522916 184365 522942
rect 184523 522916 184917 522942
rect 185259 522916 186205 522942
rect 186363 522916 186941 522942
rect 187283 522916 187401 522942
rect 172287 522780 172405 522806
rect 172563 522780 173509 522806
rect 173667 522780 174613 522806
rect 174955 522780 175901 522806
rect 176059 522780 177005 522806
rect 177163 522780 178109 522806
rect 178267 522780 179213 522806
rect 179371 522780 179765 522806
rect 180107 522780 181053 522806
rect 181211 522780 182157 522806
rect 182315 522780 183261 522806
rect 183419 522780 184365 522806
rect 184523 522780 184917 522806
rect 185259 522780 186205 522806
rect 186363 522780 186941 522806
rect 172367 522778 172405 522780
rect 172367 522762 172433 522778
rect 172259 522722 172325 522738
rect 172259 522688 172275 522722
rect 172309 522688 172325 522722
rect 172367 522728 172383 522762
rect 172417 522728 172433 522762
rect 173055 522758 173509 522780
rect 172367 522712 172433 522728
rect 172563 522722 173013 522738
rect 172259 522672 172325 522688
rect 172287 522670 172325 522672
rect 172563 522688 172835 522722
rect 172869 522688 173013 522722
rect 173055 522724 173199 522758
rect 173233 522724 173509 522758
rect 174159 522758 174613 522780
rect 173055 522708 173509 522724
rect 173667 522722 174117 522738
rect 172287 522640 172405 522670
rect 172563 522666 173013 522688
rect 173667 522688 173939 522722
rect 173973 522688 174117 522722
rect 174159 522724 174303 522758
rect 174337 522724 174613 522758
rect 175447 522758 175901 522780
rect 174159 522708 174613 522724
rect 174955 522722 175405 522738
rect 173667 522666 174117 522688
rect 174955 522688 175227 522722
rect 175261 522688 175405 522722
rect 175447 522724 175591 522758
rect 175625 522724 175901 522758
rect 176551 522758 177005 522780
rect 175447 522708 175901 522724
rect 176059 522722 176509 522738
rect 174955 522666 175405 522688
rect 176059 522688 176331 522722
rect 176365 522688 176509 522722
rect 176551 522724 176695 522758
rect 176729 522724 177005 522758
rect 177655 522758 178109 522780
rect 176551 522708 177005 522724
rect 177163 522722 177613 522738
rect 176059 522666 176509 522688
rect 177163 522688 177435 522722
rect 177469 522688 177613 522722
rect 177655 522724 177799 522758
rect 177833 522724 178109 522758
rect 178759 522758 179213 522780
rect 177655 522708 178109 522724
rect 178267 522722 178717 522738
rect 177163 522666 177613 522688
rect 178267 522688 178539 522722
rect 178573 522688 178717 522722
rect 178759 522724 178903 522758
rect 178937 522724 179213 522758
rect 179589 522758 179765 522780
rect 178759 522708 179213 522724
rect 179371 522722 179547 522738
rect 178267 522666 178717 522688
rect 179371 522688 179387 522722
rect 179421 522688 179497 522722
rect 179531 522688 179547 522722
rect 179589 522724 179605 522758
rect 179639 522724 179715 522758
rect 179749 522724 179765 522758
rect 180599 522758 181053 522780
rect 179589 522708 179765 522724
rect 180107 522722 180557 522738
rect 179371 522666 179547 522688
rect 180107 522688 180379 522722
rect 180413 522688 180557 522722
rect 180599 522724 180743 522758
rect 180777 522724 181053 522758
rect 181703 522758 182157 522780
rect 180599 522708 181053 522724
rect 181211 522722 181661 522738
rect 180107 522666 180557 522688
rect 181211 522688 181483 522722
rect 181517 522688 181661 522722
rect 181703 522724 181847 522758
rect 181881 522724 182157 522758
rect 182807 522758 183261 522780
rect 181703 522708 182157 522724
rect 182315 522722 182765 522738
rect 181211 522666 181661 522688
rect 182315 522688 182587 522722
rect 182621 522688 182765 522722
rect 182807 522724 182951 522758
rect 182985 522724 183261 522758
rect 183911 522758 184365 522780
rect 182807 522708 183261 522724
rect 183419 522722 183869 522738
rect 182315 522666 182765 522688
rect 183419 522688 183691 522722
rect 183725 522688 183869 522722
rect 183911 522724 184055 522758
rect 184089 522724 184365 522758
rect 184741 522758 184917 522780
rect 183911 522708 184365 522724
rect 184523 522722 184699 522738
rect 183419 522666 183869 522688
rect 184523 522688 184539 522722
rect 184573 522688 184649 522722
rect 184683 522688 184699 522722
rect 184741 522724 184757 522758
rect 184791 522724 184867 522758
rect 184901 522724 184917 522758
rect 185751 522758 186205 522780
rect 184741 522708 184917 522724
rect 185259 522722 185709 522738
rect 184523 522666 184699 522688
rect 185259 522688 185531 522722
rect 185565 522688 185709 522722
rect 185751 522724 185895 522758
rect 185929 522724 186205 522758
rect 186669 522758 186941 522780
rect 187283 522780 187401 522806
rect 187283 522778 187321 522780
rect 185751 522708 186205 522724
rect 186363 522722 186627 522738
rect 185259 522666 185709 522688
rect 186363 522688 186379 522722
rect 186413 522688 186478 522722
rect 186512 522688 186577 522722
rect 186611 522688 186627 522722
rect 186669 522724 186685 522758
rect 186719 522724 186788 522758
rect 186822 522724 186891 522758
rect 186925 522724 186941 522758
rect 186669 522708 186941 522724
rect 187255 522762 187321 522778
rect 187255 522728 187271 522762
rect 187305 522728 187321 522762
rect 187255 522712 187321 522728
rect 187363 522722 187429 522738
rect 186363 522666 186627 522688
rect 187363 522688 187379 522722
rect 187413 522688 187429 522722
rect 187363 522672 187429 522688
rect 187363 522670 187401 522672
rect 172563 522640 173509 522666
rect 173667 522640 174613 522666
rect 174955 522640 175901 522666
rect 176059 522640 177005 522666
rect 177163 522640 178109 522666
rect 178267 522640 179213 522666
rect 179371 522640 179765 522666
rect 180107 522640 181053 522666
rect 181211 522640 182157 522666
rect 182315 522640 183261 522666
rect 183419 522640 184365 522666
rect 184523 522640 184917 522666
rect 185259 522640 186205 522666
rect 186363 522640 186941 522666
rect 187283 522640 187401 522670
rect 172287 522440 172405 522466
rect 172563 522440 173509 522466
rect 173667 522440 174613 522466
rect 174955 522440 175901 522466
rect 176059 522440 177005 522466
rect 177163 522440 178109 522466
rect 178267 522440 179213 522466
rect 179371 522440 179765 522466
rect 180107 522440 181053 522466
rect 181211 522440 182157 522466
rect 182315 522440 183261 522466
rect 183419 522440 184365 522466
rect 184523 522440 184917 522466
rect 185259 522440 186205 522466
rect 186363 522440 186941 522466
rect 187283 522440 187401 522466
rect 172287 522372 172405 522398
rect 172563 522372 173509 522398
rect 173667 522372 174613 522398
rect 174771 522372 175717 522398
rect 175875 522372 176821 522398
rect 176979 522372 177189 522398
rect 177531 522372 178477 522398
rect 178635 522372 179581 522398
rect 179739 522372 180685 522398
rect 180843 522372 181789 522398
rect 181947 522372 182341 522398
rect 182683 522372 183629 522398
rect 183787 522372 184733 522398
rect 184891 522372 185837 522398
rect 185995 522372 186941 522398
rect 187283 522372 187401 522398
rect 172287 522168 172405 522198
rect 172563 522172 173509 522198
rect 173667 522172 174613 522198
rect 174771 522172 175717 522198
rect 175875 522172 176821 522198
rect 176979 522172 177189 522198
rect 177531 522172 178477 522198
rect 178635 522172 179581 522198
rect 179739 522172 180685 522198
rect 180843 522172 181789 522198
rect 181947 522172 182341 522198
rect 182683 522172 183629 522198
rect 183787 522172 184733 522198
rect 184891 522172 185837 522198
rect 185995 522172 186941 522198
rect 172287 522166 172325 522168
rect 172259 522150 172325 522166
rect 172259 522116 172275 522150
rect 172309 522116 172325 522150
rect 172563 522150 173013 522172
rect 172259 522100 172325 522116
rect 172367 522110 172433 522126
rect 172367 522076 172383 522110
rect 172417 522076 172433 522110
rect 172563 522116 172835 522150
rect 172869 522116 173013 522150
rect 173667 522150 174117 522172
rect 172563 522100 173013 522116
rect 173055 522114 173509 522130
rect 172367 522060 172433 522076
rect 173055 522080 173199 522114
rect 173233 522080 173509 522114
rect 173667 522116 173939 522150
rect 173973 522116 174117 522150
rect 174771 522150 175221 522172
rect 173667 522100 174117 522116
rect 174159 522114 174613 522130
rect 172367 522058 172405 522060
rect 173055 522058 173509 522080
rect 174159 522080 174303 522114
rect 174337 522080 174613 522114
rect 174771 522116 175043 522150
rect 175077 522116 175221 522150
rect 175875 522150 176325 522172
rect 176979 522166 177063 522172
rect 174771 522100 175221 522116
rect 175263 522114 175717 522130
rect 174159 522058 174613 522080
rect 175263 522080 175407 522114
rect 175441 522080 175717 522114
rect 175875 522116 176147 522150
rect 176181 522116 176325 522150
rect 176921 522150 177063 522166
rect 175875 522100 176325 522116
rect 176367 522114 176821 522130
rect 175263 522058 175717 522080
rect 176367 522080 176511 522114
rect 176545 522080 176821 522114
rect 176921 522116 176937 522150
rect 176971 522116 177063 522150
rect 177531 522150 177981 522172
rect 176921 522100 177063 522116
rect 177105 522114 177247 522130
rect 176367 522058 176821 522080
rect 177105 522080 177197 522114
rect 177231 522080 177247 522114
rect 177531 522116 177803 522150
rect 177837 522116 177981 522150
rect 178635 522150 179085 522172
rect 177531 522100 177981 522116
rect 178023 522114 178477 522130
rect 177105 522064 177247 522080
rect 178023 522080 178167 522114
rect 178201 522080 178477 522114
rect 178635 522116 178907 522150
rect 178941 522116 179085 522150
rect 179739 522150 180189 522172
rect 178635 522100 179085 522116
rect 179127 522114 179581 522130
rect 177105 522058 177189 522064
rect 178023 522058 178477 522080
rect 179127 522080 179271 522114
rect 179305 522080 179581 522114
rect 179739 522116 180011 522150
rect 180045 522116 180189 522150
rect 180843 522150 181293 522172
rect 179739 522100 180189 522116
rect 180231 522114 180685 522130
rect 179127 522058 179581 522080
rect 180231 522080 180375 522114
rect 180409 522080 180685 522114
rect 180843 522116 181115 522150
rect 181149 522116 181293 522150
rect 181947 522150 182123 522172
rect 180843 522100 181293 522116
rect 181335 522114 181789 522130
rect 180231 522058 180685 522080
rect 181335 522080 181479 522114
rect 181513 522080 181789 522114
rect 181947 522116 181963 522150
rect 181997 522116 182073 522150
rect 182107 522116 182123 522150
rect 182683 522150 183133 522172
rect 181947 522100 182123 522116
rect 182165 522114 182341 522130
rect 181335 522058 181789 522080
rect 182165 522080 182181 522114
rect 182215 522080 182291 522114
rect 182325 522080 182341 522114
rect 182683 522116 182955 522150
rect 182989 522116 183133 522150
rect 183787 522150 184237 522172
rect 182683 522100 183133 522116
rect 183175 522114 183629 522130
rect 182165 522058 182341 522080
rect 183175 522080 183319 522114
rect 183353 522080 183629 522114
rect 183787 522116 184059 522150
rect 184093 522116 184237 522150
rect 184891 522150 185341 522172
rect 183787 522100 184237 522116
rect 184279 522114 184733 522130
rect 183175 522058 183629 522080
rect 184279 522080 184423 522114
rect 184457 522080 184733 522114
rect 184891 522116 185163 522150
rect 185197 522116 185341 522150
rect 185995 522150 186445 522172
rect 187283 522168 187401 522198
rect 184891 522100 185341 522116
rect 185383 522114 185837 522130
rect 184279 522058 184733 522080
rect 185383 522080 185527 522114
rect 185561 522080 185837 522114
rect 185995 522116 186267 522150
rect 186301 522116 186445 522150
rect 187363 522166 187401 522168
rect 187363 522150 187429 522166
rect 185995 522100 186445 522116
rect 186487 522114 186941 522130
rect 185383 522058 185837 522080
rect 186487 522080 186631 522114
rect 186665 522080 186941 522114
rect 186487 522058 186941 522080
rect 187255 522110 187321 522126
rect 187255 522076 187271 522110
rect 187305 522076 187321 522110
rect 187363 522116 187379 522150
rect 187413 522116 187429 522150
rect 187363 522100 187429 522116
rect 187255 522060 187321 522076
rect 172287 522032 172405 522058
rect 172563 522032 173509 522058
rect 173667 522032 174613 522058
rect 174771 522032 175717 522058
rect 175875 522032 176821 522058
rect 176979 522032 177189 522058
rect 177531 522032 178477 522058
rect 178635 522032 179581 522058
rect 179739 522032 180685 522058
rect 180843 522032 181789 522058
rect 181947 522032 182341 522058
rect 182683 522032 183629 522058
rect 183787 522032 184733 522058
rect 184891 522032 185837 522058
rect 185995 522032 186941 522058
rect 187283 522058 187321 522060
rect 187283 522032 187401 522058
rect 172287 521896 172405 521922
rect 172563 521896 173509 521922
rect 173667 521896 174613 521922
rect 174771 521896 175717 521922
rect 175875 521896 176821 521922
rect 176979 521896 177189 521922
rect 177531 521896 178477 521922
rect 178635 521896 179581 521922
rect 179739 521896 180685 521922
rect 180843 521896 181789 521922
rect 181947 521896 182341 521922
rect 182683 521896 183629 521922
rect 183787 521896 184733 521922
rect 184891 521896 185837 521922
rect 185995 521896 186941 521922
rect 187283 521896 187401 521922
rect 172287 521828 172405 521854
rect 172563 521828 173509 521854
rect 173667 521828 174613 521854
rect 174955 521828 175901 521854
rect 176059 521828 177005 521854
rect 177163 521828 178109 521854
rect 178267 521828 179213 521854
rect 179371 521828 179765 521854
rect 180107 521828 181053 521854
rect 181211 521828 182157 521854
rect 182315 521828 183261 521854
rect 183419 521828 184365 521854
rect 184523 521828 184917 521854
rect 185259 521828 186205 521854
rect 186363 521828 186941 521854
rect 187283 521828 187401 521854
rect 172287 521692 172405 521718
rect 172563 521692 173509 521718
rect 173667 521692 174613 521718
rect 174955 521692 175901 521718
rect 176059 521692 177005 521718
rect 177163 521692 178109 521718
rect 178267 521692 179213 521718
rect 179371 521692 179765 521718
rect 180107 521692 181053 521718
rect 181211 521692 182157 521718
rect 182315 521692 183261 521718
rect 183419 521692 184365 521718
rect 184523 521692 184917 521718
rect 185259 521692 186205 521718
rect 186363 521692 186941 521718
rect 172367 521690 172405 521692
rect 172367 521674 172433 521690
rect 172259 521634 172325 521650
rect 172259 521600 172275 521634
rect 172309 521600 172325 521634
rect 172367 521640 172383 521674
rect 172417 521640 172433 521674
rect 173055 521670 173509 521692
rect 172367 521624 172433 521640
rect 172563 521634 173013 521650
rect 172259 521584 172325 521600
rect 172287 521582 172325 521584
rect 172563 521600 172835 521634
rect 172869 521600 173013 521634
rect 173055 521636 173199 521670
rect 173233 521636 173509 521670
rect 174159 521670 174613 521692
rect 173055 521620 173509 521636
rect 173667 521634 174117 521650
rect 172287 521552 172405 521582
rect 172563 521578 173013 521600
rect 173667 521600 173939 521634
rect 173973 521600 174117 521634
rect 174159 521636 174303 521670
rect 174337 521636 174613 521670
rect 175447 521670 175901 521692
rect 174159 521620 174613 521636
rect 174955 521634 175405 521650
rect 173667 521578 174117 521600
rect 174955 521600 175227 521634
rect 175261 521600 175405 521634
rect 175447 521636 175591 521670
rect 175625 521636 175901 521670
rect 176551 521670 177005 521692
rect 175447 521620 175901 521636
rect 176059 521634 176509 521650
rect 174955 521578 175405 521600
rect 176059 521600 176331 521634
rect 176365 521600 176509 521634
rect 176551 521636 176695 521670
rect 176729 521636 177005 521670
rect 177655 521670 178109 521692
rect 176551 521620 177005 521636
rect 177163 521634 177613 521650
rect 176059 521578 176509 521600
rect 177163 521600 177435 521634
rect 177469 521600 177613 521634
rect 177655 521636 177799 521670
rect 177833 521636 178109 521670
rect 178759 521670 179213 521692
rect 177655 521620 178109 521636
rect 178267 521634 178717 521650
rect 177163 521578 177613 521600
rect 178267 521600 178539 521634
rect 178573 521600 178717 521634
rect 178759 521636 178903 521670
rect 178937 521636 179213 521670
rect 179589 521670 179765 521692
rect 178759 521620 179213 521636
rect 179371 521634 179547 521650
rect 178267 521578 178717 521600
rect 179371 521600 179387 521634
rect 179421 521600 179497 521634
rect 179531 521600 179547 521634
rect 179589 521636 179605 521670
rect 179639 521636 179715 521670
rect 179749 521636 179765 521670
rect 180599 521670 181053 521692
rect 179589 521620 179765 521636
rect 180107 521634 180557 521650
rect 179371 521578 179547 521600
rect 180107 521600 180379 521634
rect 180413 521600 180557 521634
rect 180599 521636 180743 521670
rect 180777 521636 181053 521670
rect 181703 521670 182157 521692
rect 180599 521620 181053 521636
rect 181211 521634 181661 521650
rect 180107 521578 180557 521600
rect 181211 521600 181483 521634
rect 181517 521600 181661 521634
rect 181703 521636 181847 521670
rect 181881 521636 182157 521670
rect 182807 521670 183261 521692
rect 181703 521620 182157 521636
rect 182315 521634 182765 521650
rect 181211 521578 181661 521600
rect 182315 521600 182587 521634
rect 182621 521600 182765 521634
rect 182807 521636 182951 521670
rect 182985 521636 183261 521670
rect 183911 521670 184365 521692
rect 182807 521620 183261 521636
rect 183419 521634 183869 521650
rect 182315 521578 182765 521600
rect 183419 521600 183691 521634
rect 183725 521600 183869 521634
rect 183911 521636 184055 521670
rect 184089 521636 184365 521670
rect 184741 521670 184917 521692
rect 183911 521620 184365 521636
rect 184523 521634 184699 521650
rect 183419 521578 183869 521600
rect 184523 521600 184539 521634
rect 184573 521600 184649 521634
rect 184683 521600 184699 521634
rect 184741 521636 184757 521670
rect 184791 521636 184867 521670
rect 184901 521636 184917 521670
rect 185751 521670 186205 521692
rect 184741 521620 184917 521636
rect 185259 521634 185709 521650
rect 184523 521578 184699 521600
rect 185259 521600 185531 521634
rect 185565 521600 185709 521634
rect 185751 521636 185895 521670
rect 185929 521636 186205 521670
rect 186669 521670 186941 521692
rect 187283 521692 187401 521718
rect 187283 521690 187321 521692
rect 185751 521620 186205 521636
rect 186363 521634 186627 521650
rect 185259 521578 185709 521600
rect 186363 521600 186379 521634
rect 186413 521600 186478 521634
rect 186512 521600 186577 521634
rect 186611 521600 186627 521634
rect 186669 521636 186685 521670
rect 186719 521636 186788 521670
rect 186822 521636 186891 521670
rect 186925 521636 186941 521670
rect 186669 521620 186941 521636
rect 187255 521674 187321 521690
rect 187255 521640 187271 521674
rect 187305 521640 187321 521674
rect 187255 521624 187321 521640
rect 187363 521634 187429 521650
rect 186363 521578 186627 521600
rect 187363 521600 187379 521634
rect 187413 521600 187429 521634
rect 187363 521584 187429 521600
rect 187363 521582 187401 521584
rect 172563 521552 173509 521578
rect 173667 521552 174613 521578
rect 174955 521552 175901 521578
rect 176059 521552 177005 521578
rect 177163 521552 178109 521578
rect 178267 521552 179213 521578
rect 179371 521552 179765 521578
rect 180107 521552 181053 521578
rect 181211 521552 182157 521578
rect 182315 521552 183261 521578
rect 183419 521552 184365 521578
rect 184523 521552 184917 521578
rect 185259 521552 186205 521578
rect 186363 521552 186941 521578
rect 187283 521552 187401 521582
rect 172287 521352 172405 521378
rect 172563 521352 173509 521378
rect 173667 521352 174613 521378
rect 174955 521352 175901 521378
rect 176059 521352 177005 521378
rect 177163 521352 178109 521378
rect 178267 521352 179213 521378
rect 179371 521352 179765 521378
rect 180107 521352 181053 521378
rect 181211 521352 182157 521378
rect 182315 521352 183261 521378
rect 183419 521352 184365 521378
rect 184523 521352 184917 521378
rect 185259 521352 186205 521378
rect 186363 521352 186941 521378
rect 187283 521352 187401 521378
rect 172287 521284 172405 521310
rect 172563 521284 173509 521310
rect 173667 521284 174613 521310
rect 174771 521284 175717 521310
rect 175875 521284 176821 521310
rect 176979 521284 177189 521310
rect 177531 521284 178477 521310
rect 178635 521284 179581 521310
rect 179739 521284 180685 521310
rect 180843 521284 181789 521310
rect 181947 521284 182341 521310
rect 182683 521284 183629 521310
rect 183787 521284 184733 521310
rect 184891 521284 185837 521310
rect 185995 521284 186941 521310
rect 187283 521284 187401 521310
rect 172287 521080 172405 521110
rect 172563 521084 173509 521110
rect 173667 521084 174613 521110
rect 174771 521084 175717 521110
rect 175875 521084 176821 521110
rect 176979 521084 177189 521110
rect 177531 521084 178477 521110
rect 178635 521084 179581 521110
rect 179739 521084 180685 521110
rect 180843 521084 181789 521110
rect 181947 521084 182341 521110
rect 182683 521084 183629 521110
rect 183787 521084 184733 521110
rect 184891 521084 185837 521110
rect 185995 521084 186941 521110
rect 172287 521078 172325 521080
rect 172259 521062 172325 521078
rect 172259 521028 172275 521062
rect 172309 521028 172325 521062
rect 172563 521062 173013 521084
rect 172259 521012 172325 521028
rect 172367 521022 172433 521038
rect 172367 520988 172383 521022
rect 172417 520988 172433 521022
rect 172563 521028 172835 521062
rect 172869 521028 173013 521062
rect 173667 521062 174117 521084
rect 172563 521012 173013 521028
rect 173055 521026 173509 521042
rect 172367 520972 172433 520988
rect 173055 520992 173199 521026
rect 173233 520992 173509 521026
rect 173667 521028 173939 521062
rect 173973 521028 174117 521062
rect 174771 521062 175221 521084
rect 173667 521012 174117 521028
rect 174159 521026 174613 521042
rect 172367 520970 172405 520972
rect 173055 520970 173509 520992
rect 174159 520992 174303 521026
rect 174337 520992 174613 521026
rect 174771 521028 175043 521062
rect 175077 521028 175221 521062
rect 175875 521062 176325 521084
rect 176979 521078 177063 521084
rect 174771 521012 175221 521028
rect 175263 521026 175717 521042
rect 174159 520970 174613 520992
rect 175263 520992 175407 521026
rect 175441 520992 175717 521026
rect 175875 521028 176147 521062
rect 176181 521028 176325 521062
rect 176921 521062 177063 521078
rect 175875 521012 176325 521028
rect 176367 521026 176821 521042
rect 175263 520970 175717 520992
rect 176367 520992 176511 521026
rect 176545 520992 176821 521026
rect 176921 521028 176937 521062
rect 176971 521028 177063 521062
rect 177531 521062 177981 521084
rect 176921 521012 177063 521028
rect 177105 521026 177247 521042
rect 176367 520970 176821 520992
rect 177105 520992 177197 521026
rect 177231 520992 177247 521026
rect 177531 521028 177803 521062
rect 177837 521028 177981 521062
rect 178635 521062 179085 521084
rect 177531 521012 177981 521028
rect 178023 521026 178477 521042
rect 177105 520976 177247 520992
rect 178023 520992 178167 521026
rect 178201 520992 178477 521026
rect 178635 521028 178907 521062
rect 178941 521028 179085 521062
rect 179739 521062 180189 521084
rect 178635 521012 179085 521028
rect 179127 521026 179581 521042
rect 177105 520970 177189 520976
rect 178023 520970 178477 520992
rect 179127 520992 179271 521026
rect 179305 520992 179581 521026
rect 179739 521028 180011 521062
rect 180045 521028 180189 521062
rect 180843 521062 181293 521084
rect 179739 521012 180189 521028
rect 180231 521026 180685 521042
rect 179127 520970 179581 520992
rect 180231 520992 180375 521026
rect 180409 520992 180685 521026
rect 180843 521028 181115 521062
rect 181149 521028 181293 521062
rect 181947 521062 182123 521084
rect 180843 521012 181293 521028
rect 181335 521026 181789 521042
rect 180231 520970 180685 520992
rect 181335 520992 181479 521026
rect 181513 520992 181789 521026
rect 181947 521028 181963 521062
rect 181997 521028 182073 521062
rect 182107 521028 182123 521062
rect 182683 521062 183133 521084
rect 181947 521012 182123 521028
rect 182165 521026 182341 521042
rect 181335 520970 181789 520992
rect 182165 520992 182181 521026
rect 182215 520992 182291 521026
rect 182325 520992 182341 521026
rect 182683 521028 182955 521062
rect 182989 521028 183133 521062
rect 183787 521062 184237 521084
rect 182683 521012 183133 521028
rect 183175 521026 183629 521042
rect 182165 520970 182341 520992
rect 183175 520992 183319 521026
rect 183353 520992 183629 521026
rect 183787 521028 184059 521062
rect 184093 521028 184237 521062
rect 184891 521062 185341 521084
rect 183787 521012 184237 521028
rect 184279 521026 184733 521042
rect 183175 520970 183629 520992
rect 184279 520992 184423 521026
rect 184457 520992 184733 521026
rect 184891 521028 185163 521062
rect 185197 521028 185341 521062
rect 185995 521062 186445 521084
rect 187283 521080 187401 521110
rect 184891 521012 185341 521028
rect 185383 521026 185837 521042
rect 184279 520970 184733 520992
rect 185383 520992 185527 521026
rect 185561 520992 185837 521026
rect 185995 521028 186267 521062
rect 186301 521028 186445 521062
rect 187363 521078 187401 521080
rect 187363 521062 187429 521078
rect 185995 521012 186445 521028
rect 186487 521026 186941 521042
rect 185383 520970 185837 520992
rect 186487 520992 186631 521026
rect 186665 520992 186941 521026
rect 186487 520970 186941 520992
rect 187255 521022 187321 521038
rect 187255 520988 187271 521022
rect 187305 520988 187321 521022
rect 187363 521028 187379 521062
rect 187413 521028 187429 521062
rect 187363 521012 187429 521028
rect 187255 520972 187321 520988
rect 172287 520944 172405 520970
rect 172563 520944 173509 520970
rect 173667 520944 174613 520970
rect 174771 520944 175717 520970
rect 175875 520944 176821 520970
rect 176979 520944 177189 520970
rect 177531 520944 178477 520970
rect 178635 520944 179581 520970
rect 179739 520944 180685 520970
rect 180843 520944 181789 520970
rect 181947 520944 182341 520970
rect 182683 520944 183629 520970
rect 183787 520944 184733 520970
rect 184891 520944 185837 520970
rect 185995 520944 186941 520970
rect 187283 520970 187321 520972
rect 187283 520944 187401 520970
rect 172287 520808 172405 520834
rect 172563 520808 173509 520834
rect 173667 520808 174613 520834
rect 174771 520808 175717 520834
rect 175875 520808 176821 520834
rect 176979 520808 177189 520834
rect 177531 520808 178477 520834
rect 178635 520808 179581 520834
rect 179739 520808 180685 520834
rect 180843 520808 181789 520834
rect 181947 520808 182341 520834
rect 182683 520808 183629 520834
rect 183787 520808 184733 520834
rect 184891 520808 185837 520834
rect 185995 520808 186941 520834
rect 187283 520808 187401 520834
rect 172287 520740 172405 520766
rect 172563 520740 173509 520766
rect 173667 520740 174613 520766
rect 174955 520740 175901 520766
rect 176059 520740 177005 520766
rect 177163 520740 178109 520766
rect 178267 520740 179213 520766
rect 179371 520740 179765 520766
rect 180107 520740 181053 520766
rect 181211 520740 182157 520766
rect 182315 520740 183261 520766
rect 183419 520740 184365 520766
rect 184523 520740 184917 520766
rect 185259 520740 186205 520766
rect 186363 520740 186941 520766
rect 187283 520740 187401 520766
rect 172287 520604 172405 520630
rect 172563 520604 173509 520630
rect 173667 520604 174613 520630
rect 174955 520604 175901 520630
rect 176059 520604 177005 520630
rect 177163 520604 178109 520630
rect 178267 520604 179213 520630
rect 179371 520604 179765 520630
rect 180107 520604 181053 520630
rect 181211 520604 182157 520630
rect 182315 520604 183261 520630
rect 183419 520604 184365 520630
rect 184523 520604 184917 520630
rect 185259 520604 186205 520630
rect 186363 520604 186941 520630
rect 172367 520602 172405 520604
rect 172367 520586 172433 520602
rect 172259 520546 172325 520562
rect 172259 520512 172275 520546
rect 172309 520512 172325 520546
rect 172367 520552 172383 520586
rect 172417 520552 172433 520586
rect 173055 520582 173509 520604
rect 172367 520536 172433 520552
rect 172563 520546 173013 520562
rect 172259 520496 172325 520512
rect 172287 520494 172325 520496
rect 172563 520512 172835 520546
rect 172869 520512 173013 520546
rect 173055 520548 173199 520582
rect 173233 520548 173509 520582
rect 174159 520582 174613 520604
rect 173055 520532 173509 520548
rect 173667 520546 174117 520562
rect 172287 520464 172405 520494
rect 172563 520490 173013 520512
rect 173667 520512 173939 520546
rect 173973 520512 174117 520546
rect 174159 520548 174303 520582
rect 174337 520548 174613 520582
rect 175447 520582 175901 520604
rect 174159 520532 174613 520548
rect 174955 520546 175405 520562
rect 173667 520490 174117 520512
rect 174955 520512 175227 520546
rect 175261 520512 175405 520546
rect 175447 520548 175591 520582
rect 175625 520548 175901 520582
rect 176551 520582 177005 520604
rect 175447 520532 175901 520548
rect 176059 520546 176509 520562
rect 174955 520490 175405 520512
rect 176059 520512 176331 520546
rect 176365 520512 176509 520546
rect 176551 520548 176695 520582
rect 176729 520548 177005 520582
rect 177655 520582 178109 520604
rect 176551 520532 177005 520548
rect 177163 520546 177613 520562
rect 176059 520490 176509 520512
rect 177163 520512 177435 520546
rect 177469 520512 177613 520546
rect 177655 520548 177799 520582
rect 177833 520548 178109 520582
rect 178759 520582 179213 520604
rect 177655 520532 178109 520548
rect 178267 520546 178717 520562
rect 177163 520490 177613 520512
rect 178267 520512 178539 520546
rect 178573 520512 178717 520546
rect 178759 520548 178903 520582
rect 178937 520548 179213 520582
rect 179589 520582 179765 520604
rect 178759 520532 179213 520548
rect 179371 520546 179547 520562
rect 178267 520490 178717 520512
rect 179371 520512 179387 520546
rect 179421 520512 179497 520546
rect 179531 520512 179547 520546
rect 179589 520548 179605 520582
rect 179639 520548 179715 520582
rect 179749 520548 179765 520582
rect 180599 520582 181053 520604
rect 179589 520532 179765 520548
rect 180107 520546 180557 520562
rect 179371 520490 179547 520512
rect 180107 520512 180379 520546
rect 180413 520512 180557 520546
rect 180599 520548 180743 520582
rect 180777 520548 181053 520582
rect 181703 520582 182157 520604
rect 180599 520532 181053 520548
rect 181211 520546 181661 520562
rect 180107 520490 180557 520512
rect 181211 520512 181483 520546
rect 181517 520512 181661 520546
rect 181703 520548 181847 520582
rect 181881 520548 182157 520582
rect 182807 520582 183261 520604
rect 181703 520532 182157 520548
rect 182315 520546 182765 520562
rect 181211 520490 181661 520512
rect 182315 520512 182587 520546
rect 182621 520512 182765 520546
rect 182807 520548 182951 520582
rect 182985 520548 183261 520582
rect 183911 520582 184365 520604
rect 182807 520532 183261 520548
rect 183419 520546 183869 520562
rect 182315 520490 182765 520512
rect 183419 520512 183691 520546
rect 183725 520512 183869 520546
rect 183911 520548 184055 520582
rect 184089 520548 184365 520582
rect 184741 520582 184917 520604
rect 183911 520532 184365 520548
rect 184523 520546 184699 520562
rect 183419 520490 183869 520512
rect 184523 520512 184539 520546
rect 184573 520512 184649 520546
rect 184683 520512 184699 520546
rect 184741 520548 184757 520582
rect 184791 520548 184867 520582
rect 184901 520548 184917 520582
rect 185751 520582 186205 520604
rect 184741 520532 184917 520548
rect 185259 520546 185709 520562
rect 184523 520490 184699 520512
rect 185259 520512 185531 520546
rect 185565 520512 185709 520546
rect 185751 520548 185895 520582
rect 185929 520548 186205 520582
rect 186669 520582 186941 520604
rect 187283 520604 187401 520630
rect 187283 520602 187321 520604
rect 185751 520532 186205 520548
rect 186363 520546 186627 520562
rect 185259 520490 185709 520512
rect 186363 520512 186379 520546
rect 186413 520512 186478 520546
rect 186512 520512 186577 520546
rect 186611 520512 186627 520546
rect 186669 520548 186685 520582
rect 186719 520548 186788 520582
rect 186822 520548 186891 520582
rect 186925 520548 186941 520582
rect 186669 520532 186941 520548
rect 187255 520586 187321 520602
rect 187255 520552 187271 520586
rect 187305 520552 187321 520586
rect 187255 520536 187321 520552
rect 187363 520546 187429 520562
rect 186363 520490 186627 520512
rect 187363 520512 187379 520546
rect 187413 520512 187429 520546
rect 187363 520496 187429 520512
rect 187363 520494 187401 520496
rect 172563 520464 173509 520490
rect 173667 520464 174613 520490
rect 174955 520464 175901 520490
rect 176059 520464 177005 520490
rect 177163 520464 178109 520490
rect 178267 520464 179213 520490
rect 179371 520464 179765 520490
rect 180107 520464 181053 520490
rect 181211 520464 182157 520490
rect 182315 520464 183261 520490
rect 183419 520464 184365 520490
rect 184523 520464 184917 520490
rect 185259 520464 186205 520490
rect 186363 520464 186941 520490
rect 187283 520464 187401 520494
rect 172287 520264 172405 520290
rect 172563 520264 173509 520290
rect 173667 520264 174613 520290
rect 174955 520264 175901 520290
rect 176059 520264 177005 520290
rect 177163 520264 178109 520290
rect 178267 520264 179213 520290
rect 179371 520264 179765 520290
rect 180107 520264 181053 520290
rect 181211 520264 182157 520290
rect 182315 520264 183261 520290
rect 183419 520264 184365 520290
rect 184523 520264 184917 520290
rect 185259 520264 186205 520290
rect 186363 520264 186941 520290
rect 187283 520264 187401 520290
rect 172287 520196 172405 520222
rect 172563 520196 173509 520222
rect 173667 520196 174613 520222
rect 174771 520196 175717 520222
rect 175875 520196 176821 520222
rect 176979 520196 177189 520222
rect 177531 520196 178477 520222
rect 178635 520196 179581 520222
rect 179739 520196 180685 520222
rect 180843 520196 181789 520222
rect 181947 520196 182341 520222
rect 182683 520196 183629 520222
rect 183787 520196 184733 520222
rect 184891 520196 185837 520222
rect 185995 520196 186941 520222
rect 187283 520196 187401 520222
rect 172287 519992 172405 520022
rect 172563 519996 173509 520022
rect 173667 519996 174613 520022
rect 174771 519996 175717 520022
rect 175875 519996 176821 520022
rect 176979 519996 177189 520022
rect 177531 519996 178477 520022
rect 178635 519996 179581 520022
rect 179739 519996 180685 520022
rect 180843 519996 181789 520022
rect 181947 519996 182341 520022
rect 182683 519996 183629 520022
rect 183787 519996 184733 520022
rect 184891 519996 185837 520022
rect 185995 519996 186941 520022
rect 172287 519990 172325 519992
rect 172259 519974 172325 519990
rect 172259 519940 172275 519974
rect 172309 519940 172325 519974
rect 172563 519974 173013 519996
rect 172259 519924 172325 519940
rect 172367 519934 172433 519950
rect 172367 519900 172383 519934
rect 172417 519900 172433 519934
rect 172563 519940 172835 519974
rect 172869 519940 173013 519974
rect 173667 519974 174117 519996
rect 172563 519924 173013 519940
rect 173055 519938 173509 519954
rect 172367 519884 172433 519900
rect 173055 519904 173199 519938
rect 173233 519904 173509 519938
rect 173667 519940 173939 519974
rect 173973 519940 174117 519974
rect 174771 519974 175221 519996
rect 173667 519924 174117 519940
rect 174159 519938 174613 519954
rect 172367 519882 172405 519884
rect 173055 519882 173509 519904
rect 174159 519904 174303 519938
rect 174337 519904 174613 519938
rect 174771 519940 175043 519974
rect 175077 519940 175221 519974
rect 175875 519974 176325 519996
rect 176979 519990 177063 519996
rect 174771 519924 175221 519940
rect 175263 519938 175717 519954
rect 174159 519882 174613 519904
rect 175263 519904 175407 519938
rect 175441 519904 175717 519938
rect 175875 519940 176147 519974
rect 176181 519940 176325 519974
rect 176921 519974 177063 519990
rect 175875 519924 176325 519940
rect 176367 519938 176821 519954
rect 175263 519882 175717 519904
rect 176367 519904 176511 519938
rect 176545 519904 176821 519938
rect 176921 519940 176937 519974
rect 176971 519940 177063 519974
rect 177531 519974 177981 519996
rect 176921 519924 177063 519940
rect 177105 519938 177247 519954
rect 176367 519882 176821 519904
rect 177105 519904 177197 519938
rect 177231 519904 177247 519938
rect 177531 519940 177803 519974
rect 177837 519940 177981 519974
rect 178635 519974 179085 519996
rect 177531 519924 177981 519940
rect 178023 519938 178477 519954
rect 177105 519888 177247 519904
rect 178023 519904 178167 519938
rect 178201 519904 178477 519938
rect 178635 519940 178907 519974
rect 178941 519940 179085 519974
rect 179739 519974 180189 519996
rect 178635 519924 179085 519940
rect 179127 519938 179581 519954
rect 177105 519882 177189 519888
rect 178023 519882 178477 519904
rect 179127 519904 179271 519938
rect 179305 519904 179581 519938
rect 179739 519940 180011 519974
rect 180045 519940 180189 519974
rect 180843 519974 181293 519996
rect 179739 519924 180189 519940
rect 180231 519938 180685 519954
rect 179127 519882 179581 519904
rect 180231 519904 180375 519938
rect 180409 519904 180685 519938
rect 180843 519940 181115 519974
rect 181149 519940 181293 519974
rect 181947 519974 182123 519996
rect 180843 519924 181293 519940
rect 181335 519938 181789 519954
rect 180231 519882 180685 519904
rect 181335 519904 181479 519938
rect 181513 519904 181789 519938
rect 181947 519940 181963 519974
rect 181997 519940 182073 519974
rect 182107 519940 182123 519974
rect 182683 519974 183133 519996
rect 181947 519924 182123 519940
rect 182165 519938 182341 519954
rect 181335 519882 181789 519904
rect 182165 519904 182181 519938
rect 182215 519904 182291 519938
rect 182325 519904 182341 519938
rect 182683 519940 182955 519974
rect 182989 519940 183133 519974
rect 183787 519974 184237 519996
rect 182683 519924 183133 519940
rect 183175 519938 183629 519954
rect 182165 519882 182341 519904
rect 183175 519904 183319 519938
rect 183353 519904 183629 519938
rect 183787 519940 184059 519974
rect 184093 519940 184237 519974
rect 184891 519974 185341 519996
rect 183787 519924 184237 519940
rect 184279 519938 184733 519954
rect 183175 519882 183629 519904
rect 184279 519904 184423 519938
rect 184457 519904 184733 519938
rect 184891 519940 185163 519974
rect 185197 519940 185341 519974
rect 185995 519974 186445 519996
rect 187283 519992 187401 520022
rect 184891 519924 185341 519940
rect 185383 519938 185837 519954
rect 184279 519882 184733 519904
rect 185383 519904 185527 519938
rect 185561 519904 185837 519938
rect 185995 519940 186267 519974
rect 186301 519940 186445 519974
rect 187363 519990 187401 519992
rect 187363 519974 187429 519990
rect 185995 519924 186445 519940
rect 186487 519938 186941 519954
rect 185383 519882 185837 519904
rect 186487 519904 186631 519938
rect 186665 519904 186941 519938
rect 186487 519882 186941 519904
rect 187255 519934 187321 519950
rect 187255 519900 187271 519934
rect 187305 519900 187321 519934
rect 187363 519940 187379 519974
rect 187413 519940 187429 519974
rect 187363 519924 187429 519940
rect 187255 519884 187321 519900
rect 172287 519856 172405 519882
rect 172563 519856 173509 519882
rect 173667 519856 174613 519882
rect 174771 519856 175717 519882
rect 175875 519856 176821 519882
rect 176979 519856 177189 519882
rect 177531 519856 178477 519882
rect 178635 519856 179581 519882
rect 179739 519856 180685 519882
rect 180843 519856 181789 519882
rect 181947 519856 182341 519882
rect 182683 519856 183629 519882
rect 183787 519856 184733 519882
rect 184891 519856 185837 519882
rect 185995 519856 186941 519882
rect 187283 519882 187321 519884
rect 187283 519856 187401 519882
rect 172287 519720 172405 519746
rect 172563 519720 173509 519746
rect 173667 519720 174613 519746
rect 174771 519720 175717 519746
rect 175875 519720 176821 519746
rect 176979 519720 177189 519746
rect 177531 519720 178477 519746
rect 178635 519720 179581 519746
rect 179739 519720 180685 519746
rect 180843 519720 181789 519746
rect 181947 519720 182341 519746
rect 182683 519720 183629 519746
rect 183787 519720 184733 519746
rect 184891 519720 185837 519746
rect 185995 519720 186941 519746
rect 187283 519720 187401 519746
rect 172287 519652 172405 519678
rect 172563 519652 173509 519678
rect 173667 519652 174613 519678
rect 174955 519652 175901 519678
rect 176059 519652 177005 519678
rect 177163 519652 178109 519678
rect 178267 519652 179213 519678
rect 179371 519652 179765 519678
rect 180107 519652 181053 519678
rect 181211 519652 182157 519678
rect 182315 519652 183261 519678
rect 183419 519652 184365 519678
rect 184523 519652 184917 519678
rect 185259 519652 186205 519678
rect 186363 519652 186941 519678
rect 187283 519652 187401 519678
rect 172287 519516 172405 519542
rect 172563 519516 173509 519542
rect 173667 519516 174613 519542
rect 174955 519516 175901 519542
rect 176059 519516 177005 519542
rect 177163 519516 178109 519542
rect 178267 519516 179213 519542
rect 179371 519516 179765 519542
rect 180107 519516 181053 519542
rect 181211 519516 182157 519542
rect 182315 519516 183261 519542
rect 183419 519516 184365 519542
rect 184523 519516 184917 519542
rect 185259 519516 186205 519542
rect 186363 519516 186941 519542
rect 172367 519514 172405 519516
rect 172367 519498 172433 519514
rect 172259 519458 172325 519474
rect 172259 519424 172275 519458
rect 172309 519424 172325 519458
rect 172367 519464 172383 519498
rect 172417 519464 172433 519498
rect 173055 519494 173509 519516
rect 172367 519448 172433 519464
rect 172563 519458 173013 519474
rect 172259 519408 172325 519424
rect 172287 519406 172325 519408
rect 172563 519424 172835 519458
rect 172869 519424 173013 519458
rect 173055 519460 173199 519494
rect 173233 519460 173509 519494
rect 174159 519494 174613 519516
rect 173055 519444 173509 519460
rect 173667 519458 174117 519474
rect 172287 519376 172405 519406
rect 172563 519402 173013 519424
rect 173667 519424 173939 519458
rect 173973 519424 174117 519458
rect 174159 519460 174303 519494
rect 174337 519460 174613 519494
rect 175447 519494 175901 519516
rect 174159 519444 174613 519460
rect 174955 519458 175405 519474
rect 173667 519402 174117 519424
rect 174955 519424 175227 519458
rect 175261 519424 175405 519458
rect 175447 519460 175591 519494
rect 175625 519460 175901 519494
rect 176551 519494 177005 519516
rect 175447 519444 175901 519460
rect 176059 519458 176509 519474
rect 174955 519402 175405 519424
rect 176059 519424 176331 519458
rect 176365 519424 176509 519458
rect 176551 519460 176695 519494
rect 176729 519460 177005 519494
rect 177655 519494 178109 519516
rect 176551 519444 177005 519460
rect 177163 519458 177613 519474
rect 176059 519402 176509 519424
rect 177163 519424 177435 519458
rect 177469 519424 177613 519458
rect 177655 519460 177799 519494
rect 177833 519460 178109 519494
rect 178759 519494 179213 519516
rect 177655 519444 178109 519460
rect 178267 519458 178717 519474
rect 177163 519402 177613 519424
rect 178267 519424 178539 519458
rect 178573 519424 178717 519458
rect 178759 519460 178903 519494
rect 178937 519460 179213 519494
rect 179589 519494 179765 519516
rect 178759 519444 179213 519460
rect 179371 519458 179547 519474
rect 178267 519402 178717 519424
rect 179371 519424 179387 519458
rect 179421 519424 179497 519458
rect 179531 519424 179547 519458
rect 179589 519460 179605 519494
rect 179639 519460 179715 519494
rect 179749 519460 179765 519494
rect 180599 519494 181053 519516
rect 179589 519444 179765 519460
rect 180107 519458 180557 519474
rect 179371 519402 179547 519424
rect 180107 519424 180379 519458
rect 180413 519424 180557 519458
rect 180599 519460 180743 519494
rect 180777 519460 181053 519494
rect 181703 519494 182157 519516
rect 180599 519444 181053 519460
rect 181211 519458 181661 519474
rect 180107 519402 180557 519424
rect 181211 519424 181483 519458
rect 181517 519424 181661 519458
rect 181703 519460 181847 519494
rect 181881 519460 182157 519494
rect 182807 519494 183261 519516
rect 181703 519444 182157 519460
rect 182315 519458 182765 519474
rect 181211 519402 181661 519424
rect 182315 519424 182587 519458
rect 182621 519424 182765 519458
rect 182807 519460 182951 519494
rect 182985 519460 183261 519494
rect 183911 519494 184365 519516
rect 182807 519444 183261 519460
rect 183419 519458 183869 519474
rect 182315 519402 182765 519424
rect 183419 519424 183691 519458
rect 183725 519424 183869 519458
rect 183911 519460 184055 519494
rect 184089 519460 184365 519494
rect 184741 519494 184917 519516
rect 183911 519444 184365 519460
rect 184523 519458 184699 519474
rect 183419 519402 183869 519424
rect 184523 519424 184539 519458
rect 184573 519424 184649 519458
rect 184683 519424 184699 519458
rect 184741 519460 184757 519494
rect 184791 519460 184867 519494
rect 184901 519460 184917 519494
rect 185751 519494 186205 519516
rect 184741 519444 184917 519460
rect 185259 519458 185709 519474
rect 184523 519402 184699 519424
rect 185259 519424 185531 519458
rect 185565 519424 185709 519458
rect 185751 519460 185895 519494
rect 185929 519460 186205 519494
rect 186669 519494 186941 519516
rect 187283 519516 187401 519542
rect 187283 519514 187321 519516
rect 185751 519444 186205 519460
rect 186363 519458 186627 519474
rect 185259 519402 185709 519424
rect 186363 519424 186379 519458
rect 186413 519424 186478 519458
rect 186512 519424 186577 519458
rect 186611 519424 186627 519458
rect 186669 519460 186685 519494
rect 186719 519460 186788 519494
rect 186822 519460 186891 519494
rect 186925 519460 186941 519494
rect 186669 519444 186941 519460
rect 187255 519498 187321 519514
rect 187255 519464 187271 519498
rect 187305 519464 187321 519498
rect 187255 519448 187321 519464
rect 187363 519458 187429 519474
rect 186363 519402 186627 519424
rect 187363 519424 187379 519458
rect 187413 519424 187429 519458
rect 187363 519408 187429 519424
rect 187363 519406 187401 519408
rect 172563 519376 173509 519402
rect 173667 519376 174613 519402
rect 174955 519376 175901 519402
rect 176059 519376 177005 519402
rect 177163 519376 178109 519402
rect 178267 519376 179213 519402
rect 179371 519376 179765 519402
rect 180107 519376 181053 519402
rect 181211 519376 182157 519402
rect 182315 519376 183261 519402
rect 183419 519376 184365 519402
rect 184523 519376 184917 519402
rect 185259 519376 186205 519402
rect 186363 519376 186941 519402
rect 187283 519376 187401 519406
rect 172287 519176 172405 519202
rect 172563 519176 173509 519202
rect 173667 519176 174613 519202
rect 174955 519176 175901 519202
rect 176059 519176 177005 519202
rect 177163 519176 178109 519202
rect 178267 519176 179213 519202
rect 179371 519176 179765 519202
rect 180107 519176 181053 519202
rect 181211 519176 182157 519202
rect 182315 519176 183261 519202
rect 183419 519176 184365 519202
rect 184523 519176 184917 519202
rect 185259 519176 186205 519202
rect 186363 519176 186941 519202
rect 187283 519176 187401 519202
rect 172287 519108 172405 519134
rect 172563 519108 173509 519134
rect 173667 519108 174613 519134
rect 174771 519108 175717 519134
rect 175875 519108 176821 519134
rect 176979 519108 177189 519134
rect 177531 519108 178477 519134
rect 178635 519108 179581 519134
rect 179739 519108 180685 519134
rect 180843 519108 181789 519134
rect 181947 519108 182341 519134
rect 182683 519108 183629 519134
rect 183787 519108 184733 519134
rect 184891 519108 185837 519134
rect 185995 519108 186941 519134
rect 187283 519108 187401 519134
rect 172287 518904 172405 518934
rect 172563 518908 173509 518934
rect 173667 518908 174613 518934
rect 174771 518908 175717 518934
rect 175875 518908 176821 518934
rect 176979 518908 177189 518934
rect 177531 518908 178477 518934
rect 178635 518908 179581 518934
rect 179739 518908 180685 518934
rect 180843 518908 181789 518934
rect 181947 518908 182341 518934
rect 182683 518908 183629 518934
rect 183787 518908 184733 518934
rect 184891 518908 185837 518934
rect 185995 518908 186941 518934
rect 172287 518902 172325 518904
rect 172259 518886 172325 518902
rect 172259 518852 172275 518886
rect 172309 518852 172325 518886
rect 172563 518886 173013 518908
rect 172259 518836 172325 518852
rect 172367 518846 172433 518862
rect 172367 518812 172383 518846
rect 172417 518812 172433 518846
rect 172563 518852 172835 518886
rect 172869 518852 173013 518886
rect 173667 518886 174117 518908
rect 172563 518836 173013 518852
rect 173055 518850 173509 518866
rect 172367 518796 172433 518812
rect 173055 518816 173199 518850
rect 173233 518816 173509 518850
rect 173667 518852 173939 518886
rect 173973 518852 174117 518886
rect 174771 518886 175221 518908
rect 173667 518836 174117 518852
rect 174159 518850 174613 518866
rect 172367 518794 172405 518796
rect 173055 518794 173509 518816
rect 174159 518816 174303 518850
rect 174337 518816 174613 518850
rect 174771 518852 175043 518886
rect 175077 518852 175221 518886
rect 175875 518886 176325 518908
rect 176979 518902 177063 518908
rect 174771 518836 175221 518852
rect 175263 518850 175717 518866
rect 174159 518794 174613 518816
rect 175263 518816 175407 518850
rect 175441 518816 175717 518850
rect 175875 518852 176147 518886
rect 176181 518852 176325 518886
rect 176921 518886 177063 518902
rect 175875 518836 176325 518852
rect 176367 518850 176821 518866
rect 175263 518794 175717 518816
rect 176367 518816 176511 518850
rect 176545 518816 176821 518850
rect 176921 518852 176937 518886
rect 176971 518852 177063 518886
rect 177531 518886 177981 518908
rect 176921 518836 177063 518852
rect 177105 518850 177247 518866
rect 176367 518794 176821 518816
rect 177105 518816 177197 518850
rect 177231 518816 177247 518850
rect 177531 518852 177803 518886
rect 177837 518852 177981 518886
rect 178635 518886 179085 518908
rect 177531 518836 177981 518852
rect 178023 518850 178477 518866
rect 177105 518800 177247 518816
rect 178023 518816 178167 518850
rect 178201 518816 178477 518850
rect 178635 518852 178907 518886
rect 178941 518852 179085 518886
rect 179739 518886 180189 518908
rect 178635 518836 179085 518852
rect 179127 518850 179581 518866
rect 177105 518794 177189 518800
rect 178023 518794 178477 518816
rect 179127 518816 179271 518850
rect 179305 518816 179581 518850
rect 179739 518852 180011 518886
rect 180045 518852 180189 518886
rect 180843 518886 181293 518908
rect 179739 518836 180189 518852
rect 180231 518850 180685 518866
rect 179127 518794 179581 518816
rect 180231 518816 180375 518850
rect 180409 518816 180685 518850
rect 180843 518852 181115 518886
rect 181149 518852 181293 518886
rect 181947 518886 182123 518908
rect 180843 518836 181293 518852
rect 181335 518850 181789 518866
rect 180231 518794 180685 518816
rect 181335 518816 181479 518850
rect 181513 518816 181789 518850
rect 181947 518852 181963 518886
rect 181997 518852 182073 518886
rect 182107 518852 182123 518886
rect 182683 518886 183133 518908
rect 181947 518836 182123 518852
rect 182165 518850 182341 518866
rect 181335 518794 181789 518816
rect 182165 518816 182181 518850
rect 182215 518816 182291 518850
rect 182325 518816 182341 518850
rect 182683 518852 182955 518886
rect 182989 518852 183133 518886
rect 183787 518886 184237 518908
rect 182683 518836 183133 518852
rect 183175 518850 183629 518866
rect 182165 518794 182341 518816
rect 183175 518816 183319 518850
rect 183353 518816 183629 518850
rect 183787 518852 184059 518886
rect 184093 518852 184237 518886
rect 184891 518886 185341 518908
rect 183787 518836 184237 518852
rect 184279 518850 184733 518866
rect 183175 518794 183629 518816
rect 184279 518816 184423 518850
rect 184457 518816 184733 518850
rect 184891 518852 185163 518886
rect 185197 518852 185341 518886
rect 185995 518886 186445 518908
rect 187283 518904 187401 518934
rect 184891 518836 185341 518852
rect 185383 518850 185837 518866
rect 184279 518794 184733 518816
rect 185383 518816 185527 518850
rect 185561 518816 185837 518850
rect 185995 518852 186267 518886
rect 186301 518852 186445 518886
rect 187363 518902 187401 518904
rect 187363 518886 187429 518902
rect 185995 518836 186445 518852
rect 186487 518850 186941 518866
rect 185383 518794 185837 518816
rect 186487 518816 186631 518850
rect 186665 518816 186941 518850
rect 186487 518794 186941 518816
rect 187255 518846 187321 518862
rect 187255 518812 187271 518846
rect 187305 518812 187321 518846
rect 187363 518852 187379 518886
rect 187413 518852 187429 518886
rect 187363 518836 187429 518852
rect 187255 518796 187321 518812
rect 172287 518768 172405 518794
rect 172563 518768 173509 518794
rect 173667 518768 174613 518794
rect 174771 518768 175717 518794
rect 175875 518768 176821 518794
rect 176979 518768 177189 518794
rect 177531 518768 178477 518794
rect 178635 518768 179581 518794
rect 179739 518768 180685 518794
rect 180843 518768 181789 518794
rect 181947 518768 182341 518794
rect 182683 518768 183629 518794
rect 183787 518768 184733 518794
rect 184891 518768 185837 518794
rect 185995 518768 186941 518794
rect 187283 518794 187321 518796
rect 187283 518768 187401 518794
rect 172287 518632 172405 518658
rect 172563 518632 173509 518658
rect 173667 518632 174613 518658
rect 174771 518632 175717 518658
rect 175875 518632 176821 518658
rect 176979 518632 177189 518658
rect 177531 518632 178477 518658
rect 178635 518632 179581 518658
rect 179739 518632 180685 518658
rect 180843 518632 181789 518658
rect 181947 518632 182341 518658
rect 182683 518632 183629 518658
rect 183787 518632 184733 518658
rect 184891 518632 185837 518658
rect 185995 518632 186941 518658
rect 187283 518632 187401 518658
rect 172287 518564 172405 518590
rect 172563 518564 173509 518590
rect 173667 518564 174613 518590
rect 174955 518564 175901 518590
rect 176059 518564 177005 518590
rect 177163 518564 178109 518590
rect 178267 518564 179213 518590
rect 179371 518564 179765 518590
rect 180107 518564 181053 518590
rect 181211 518564 182157 518590
rect 182315 518564 183261 518590
rect 183419 518564 184365 518590
rect 184523 518564 184917 518590
rect 185259 518564 186205 518590
rect 186363 518564 186941 518590
rect 187283 518564 187401 518590
rect 172287 518428 172405 518454
rect 172563 518428 173509 518454
rect 173667 518428 174613 518454
rect 174955 518428 175901 518454
rect 176059 518428 177005 518454
rect 177163 518428 178109 518454
rect 178267 518428 179213 518454
rect 179371 518428 179765 518454
rect 180107 518428 181053 518454
rect 181211 518428 182157 518454
rect 182315 518428 183261 518454
rect 183419 518428 184365 518454
rect 184523 518428 184917 518454
rect 185259 518428 186205 518454
rect 186363 518428 186941 518454
rect 172367 518426 172405 518428
rect 172367 518410 172433 518426
rect 172259 518370 172325 518386
rect 172259 518336 172275 518370
rect 172309 518336 172325 518370
rect 172367 518376 172383 518410
rect 172417 518376 172433 518410
rect 173055 518406 173509 518428
rect 172367 518360 172433 518376
rect 172563 518370 173013 518386
rect 172259 518320 172325 518336
rect 172287 518318 172325 518320
rect 172563 518336 172835 518370
rect 172869 518336 173013 518370
rect 173055 518372 173199 518406
rect 173233 518372 173509 518406
rect 174159 518406 174613 518428
rect 173055 518356 173509 518372
rect 173667 518370 174117 518386
rect 172287 518288 172405 518318
rect 172563 518314 173013 518336
rect 173667 518336 173939 518370
rect 173973 518336 174117 518370
rect 174159 518372 174303 518406
rect 174337 518372 174613 518406
rect 175447 518406 175901 518428
rect 174159 518356 174613 518372
rect 174955 518370 175405 518386
rect 173667 518314 174117 518336
rect 174955 518336 175227 518370
rect 175261 518336 175405 518370
rect 175447 518372 175591 518406
rect 175625 518372 175901 518406
rect 176551 518406 177005 518428
rect 175447 518356 175901 518372
rect 176059 518370 176509 518386
rect 174955 518314 175405 518336
rect 176059 518336 176331 518370
rect 176365 518336 176509 518370
rect 176551 518372 176695 518406
rect 176729 518372 177005 518406
rect 177655 518406 178109 518428
rect 176551 518356 177005 518372
rect 177163 518370 177613 518386
rect 176059 518314 176509 518336
rect 177163 518336 177435 518370
rect 177469 518336 177613 518370
rect 177655 518372 177799 518406
rect 177833 518372 178109 518406
rect 178759 518406 179213 518428
rect 177655 518356 178109 518372
rect 178267 518370 178717 518386
rect 177163 518314 177613 518336
rect 178267 518336 178539 518370
rect 178573 518336 178717 518370
rect 178759 518372 178903 518406
rect 178937 518372 179213 518406
rect 179589 518406 179765 518428
rect 178759 518356 179213 518372
rect 179371 518370 179547 518386
rect 178267 518314 178717 518336
rect 179371 518336 179387 518370
rect 179421 518336 179497 518370
rect 179531 518336 179547 518370
rect 179589 518372 179605 518406
rect 179639 518372 179715 518406
rect 179749 518372 179765 518406
rect 180599 518406 181053 518428
rect 179589 518356 179765 518372
rect 180107 518370 180557 518386
rect 179371 518314 179547 518336
rect 180107 518336 180379 518370
rect 180413 518336 180557 518370
rect 180599 518372 180743 518406
rect 180777 518372 181053 518406
rect 181703 518406 182157 518428
rect 180599 518356 181053 518372
rect 181211 518370 181661 518386
rect 180107 518314 180557 518336
rect 181211 518336 181483 518370
rect 181517 518336 181661 518370
rect 181703 518372 181847 518406
rect 181881 518372 182157 518406
rect 182807 518406 183261 518428
rect 181703 518356 182157 518372
rect 182315 518370 182765 518386
rect 181211 518314 181661 518336
rect 182315 518336 182587 518370
rect 182621 518336 182765 518370
rect 182807 518372 182951 518406
rect 182985 518372 183261 518406
rect 183911 518406 184365 518428
rect 182807 518356 183261 518372
rect 183419 518370 183869 518386
rect 182315 518314 182765 518336
rect 183419 518336 183691 518370
rect 183725 518336 183869 518370
rect 183911 518372 184055 518406
rect 184089 518372 184365 518406
rect 184741 518406 184917 518428
rect 183911 518356 184365 518372
rect 184523 518370 184699 518386
rect 183419 518314 183869 518336
rect 184523 518336 184539 518370
rect 184573 518336 184649 518370
rect 184683 518336 184699 518370
rect 184741 518372 184757 518406
rect 184791 518372 184867 518406
rect 184901 518372 184917 518406
rect 185751 518406 186205 518428
rect 184741 518356 184917 518372
rect 185259 518370 185709 518386
rect 184523 518314 184699 518336
rect 185259 518336 185531 518370
rect 185565 518336 185709 518370
rect 185751 518372 185895 518406
rect 185929 518372 186205 518406
rect 186669 518406 186941 518428
rect 187283 518428 187401 518454
rect 187283 518426 187321 518428
rect 185751 518356 186205 518372
rect 186363 518370 186627 518386
rect 185259 518314 185709 518336
rect 186363 518336 186379 518370
rect 186413 518336 186478 518370
rect 186512 518336 186577 518370
rect 186611 518336 186627 518370
rect 186669 518372 186685 518406
rect 186719 518372 186788 518406
rect 186822 518372 186891 518406
rect 186925 518372 186941 518406
rect 186669 518356 186941 518372
rect 187255 518410 187321 518426
rect 187255 518376 187271 518410
rect 187305 518376 187321 518410
rect 187255 518360 187321 518376
rect 187363 518370 187429 518386
rect 186363 518314 186627 518336
rect 187363 518336 187379 518370
rect 187413 518336 187429 518370
rect 187363 518320 187429 518336
rect 187363 518318 187401 518320
rect 172563 518288 173509 518314
rect 173667 518288 174613 518314
rect 174955 518288 175901 518314
rect 176059 518288 177005 518314
rect 177163 518288 178109 518314
rect 178267 518288 179213 518314
rect 179371 518288 179765 518314
rect 180107 518288 181053 518314
rect 181211 518288 182157 518314
rect 182315 518288 183261 518314
rect 183419 518288 184365 518314
rect 184523 518288 184917 518314
rect 185259 518288 186205 518314
rect 186363 518288 186941 518314
rect 187283 518288 187401 518318
rect 172287 518088 172405 518114
rect 172563 518088 173509 518114
rect 173667 518088 174613 518114
rect 174955 518088 175901 518114
rect 176059 518088 177005 518114
rect 177163 518088 178109 518114
rect 178267 518088 179213 518114
rect 179371 518088 179765 518114
rect 180107 518088 181053 518114
rect 181211 518088 182157 518114
rect 182315 518088 183261 518114
rect 183419 518088 184365 518114
rect 184523 518088 184917 518114
rect 185259 518088 186205 518114
rect 186363 518088 186941 518114
rect 187283 518088 187401 518114
rect 172287 518020 172405 518046
rect 172563 518020 173509 518046
rect 173667 518020 174613 518046
rect 174771 518020 175717 518046
rect 175875 518020 176821 518046
rect 176979 518020 177189 518046
rect 177531 518020 178477 518046
rect 178635 518020 179581 518046
rect 179739 518020 180685 518046
rect 180843 518020 181789 518046
rect 181947 518020 182341 518046
rect 182683 518020 183629 518046
rect 183787 518020 184733 518046
rect 184891 518020 185837 518046
rect 185995 518020 186941 518046
rect 187283 518020 187401 518046
rect 172287 517816 172405 517846
rect 172563 517820 173509 517846
rect 173667 517820 174613 517846
rect 174771 517820 175717 517846
rect 175875 517820 176821 517846
rect 176979 517820 177189 517846
rect 177531 517820 178477 517846
rect 178635 517820 179581 517846
rect 179739 517820 180685 517846
rect 180843 517820 181789 517846
rect 181947 517820 182341 517846
rect 182683 517820 183629 517846
rect 183787 517820 184733 517846
rect 184891 517820 185837 517846
rect 185995 517820 186941 517846
rect 172287 517814 172325 517816
rect 172259 517798 172325 517814
rect 172259 517764 172275 517798
rect 172309 517764 172325 517798
rect 172563 517798 173013 517820
rect 172259 517748 172325 517764
rect 172367 517758 172433 517774
rect 172367 517724 172383 517758
rect 172417 517724 172433 517758
rect 172563 517764 172835 517798
rect 172869 517764 173013 517798
rect 173667 517798 174117 517820
rect 172563 517748 173013 517764
rect 173055 517762 173509 517778
rect 172367 517708 172433 517724
rect 173055 517728 173199 517762
rect 173233 517728 173509 517762
rect 173667 517764 173939 517798
rect 173973 517764 174117 517798
rect 174771 517798 175221 517820
rect 173667 517748 174117 517764
rect 174159 517762 174613 517778
rect 172367 517706 172405 517708
rect 173055 517706 173509 517728
rect 174159 517728 174303 517762
rect 174337 517728 174613 517762
rect 174771 517764 175043 517798
rect 175077 517764 175221 517798
rect 175875 517798 176325 517820
rect 176979 517814 177063 517820
rect 174771 517748 175221 517764
rect 175263 517762 175717 517778
rect 174159 517706 174613 517728
rect 175263 517728 175407 517762
rect 175441 517728 175717 517762
rect 175875 517764 176147 517798
rect 176181 517764 176325 517798
rect 176921 517798 177063 517814
rect 175875 517748 176325 517764
rect 176367 517762 176821 517778
rect 175263 517706 175717 517728
rect 176367 517728 176511 517762
rect 176545 517728 176821 517762
rect 176921 517764 176937 517798
rect 176971 517764 177063 517798
rect 177531 517798 177981 517820
rect 176921 517748 177063 517764
rect 177105 517762 177247 517778
rect 176367 517706 176821 517728
rect 177105 517728 177197 517762
rect 177231 517728 177247 517762
rect 177531 517764 177803 517798
rect 177837 517764 177981 517798
rect 178635 517798 179085 517820
rect 177531 517748 177981 517764
rect 178023 517762 178477 517778
rect 177105 517712 177247 517728
rect 178023 517728 178167 517762
rect 178201 517728 178477 517762
rect 178635 517764 178907 517798
rect 178941 517764 179085 517798
rect 179739 517798 180189 517820
rect 178635 517748 179085 517764
rect 179127 517762 179581 517778
rect 177105 517706 177189 517712
rect 178023 517706 178477 517728
rect 179127 517728 179271 517762
rect 179305 517728 179581 517762
rect 179739 517764 180011 517798
rect 180045 517764 180189 517798
rect 180843 517798 181293 517820
rect 179739 517748 180189 517764
rect 180231 517762 180685 517778
rect 179127 517706 179581 517728
rect 180231 517728 180375 517762
rect 180409 517728 180685 517762
rect 180843 517764 181115 517798
rect 181149 517764 181293 517798
rect 181947 517798 182123 517820
rect 180843 517748 181293 517764
rect 181335 517762 181789 517778
rect 180231 517706 180685 517728
rect 181335 517728 181479 517762
rect 181513 517728 181789 517762
rect 181947 517764 181963 517798
rect 181997 517764 182073 517798
rect 182107 517764 182123 517798
rect 182683 517798 183133 517820
rect 181947 517748 182123 517764
rect 182165 517762 182341 517778
rect 181335 517706 181789 517728
rect 182165 517728 182181 517762
rect 182215 517728 182291 517762
rect 182325 517728 182341 517762
rect 182683 517764 182955 517798
rect 182989 517764 183133 517798
rect 183787 517798 184237 517820
rect 182683 517748 183133 517764
rect 183175 517762 183629 517778
rect 182165 517706 182341 517728
rect 183175 517728 183319 517762
rect 183353 517728 183629 517762
rect 183787 517764 184059 517798
rect 184093 517764 184237 517798
rect 184891 517798 185341 517820
rect 183787 517748 184237 517764
rect 184279 517762 184733 517778
rect 183175 517706 183629 517728
rect 184279 517728 184423 517762
rect 184457 517728 184733 517762
rect 184891 517764 185163 517798
rect 185197 517764 185341 517798
rect 185995 517798 186445 517820
rect 187283 517816 187401 517846
rect 184891 517748 185341 517764
rect 185383 517762 185837 517778
rect 184279 517706 184733 517728
rect 185383 517728 185527 517762
rect 185561 517728 185837 517762
rect 185995 517764 186267 517798
rect 186301 517764 186445 517798
rect 187363 517814 187401 517816
rect 187363 517798 187429 517814
rect 185995 517748 186445 517764
rect 186487 517762 186941 517778
rect 185383 517706 185837 517728
rect 186487 517728 186631 517762
rect 186665 517728 186941 517762
rect 186487 517706 186941 517728
rect 187255 517758 187321 517774
rect 187255 517724 187271 517758
rect 187305 517724 187321 517758
rect 187363 517764 187379 517798
rect 187413 517764 187429 517798
rect 187363 517748 187429 517764
rect 187255 517708 187321 517724
rect 172287 517680 172405 517706
rect 172563 517680 173509 517706
rect 173667 517680 174613 517706
rect 174771 517680 175717 517706
rect 175875 517680 176821 517706
rect 176979 517680 177189 517706
rect 177531 517680 178477 517706
rect 178635 517680 179581 517706
rect 179739 517680 180685 517706
rect 180843 517680 181789 517706
rect 181947 517680 182341 517706
rect 182683 517680 183629 517706
rect 183787 517680 184733 517706
rect 184891 517680 185837 517706
rect 185995 517680 186941 517706
rect 187283 517706 187321 517708
rect 187283 517680 187401 517706
rect 172287 517544 172405 517570
rect 172563 517544 173509 517570
rect 173667 517544 174613 517570
rect 174771 517544 175717 517570
rect 175875 517544 176821 517570
rect 176979 517544 177189 517570
rect 177531 517544 178477 517570
rect 178635 517544 179581 517570
rect 179739 517544 180685 517570
rect 180843 517544 181789 517570
rect 181947 517544 182341 517570
rect 182683 517544 183629 517570
rect 183787 517544 184733 517570
rect 184891 517544 185837 517570
rect 185995 517544 186941 517570
rect 187283 517544 187401 517570
rect 172287 517476 172405 517502
rect 172563 517476 173509 517502
rect 173667 517476 174613 517502
rect 174955 517476 175901 517502
rect 176059 517476 177005 517502
rect 177163 517476 178109 517502
rect 178267 517476 179213 517502
rect 179371 517476 179765 517502
rect 180107 517476 181053 517502
rect 181211 517476 182157 517502
rect 182315 517476 183261 517502
rect 183419 517476 184365 517502
rect 184523 517476 184917 517502
rect 185259 517476 186205 517502
rect 186363 517476 186941 517502
rect 187283 517476 187401 517502
rect 172287 517340 172405 517366
rect 172563 517340 173509 517366
rect 173667 517340 174613 517366
rect 174955 517340 175901 517366
rect 176059 517340 177005 517366
rect 177163 517340 178109 517366
rect 178267 517340 179213 517366
rect 179371 517340 179765 517366
rect 180107 517340 181053 517366
rect 181211 517340 182157 517366
rect 182315 517340 183261 517366
rect 183419 517340 184365 517366
rect 184523 517340 184917 517366
rect 185259 517340 186205 517366
rect 186363 517340 186941 517366
rect 172367 517338 172405 517340
rect 172367 517322 172433 517338
rect 172259 517282 172325 517298
rect 172259 517248 172275 517282
rect 172309 517248 172325 517282
rect 172367 517288 172383 517322
rect 172417 517288 172433 517322
rect 173055 517318 173509 517340
rect 172367 517272 172433 517288
rect 172563 517282 173013 517298
rect 172259 517232 172325 517248
rect 172287 517230 172325 517232
rect 172563 517248 172835 517282
rect 172869 517248 173013 517282
rect 173055 517284 173199 517318
rect 173233 517284 173509 517318
rect 174159 517318 174613 517340
rect 173055 517268 173509 517284
rect 173667 517282 174117 517298
rect 172287 517200 172405 517230
rect 172563 517226 173013 517248
rect 173667 517248 173939 517282
rect 173973 517248 174117 517282
rect 174159 517284 174303 517318
rect 174337 517284 174613 517318
rect 175447 517318 175901 517340
rect 174159 517268 174613 517284
rect 174955 517282 175405 517298
rect 173667 517226 174117 517248
rect 174955 517248 175227 517282
rect 175261 517248 175405 517282
rect 175447 517284 175591 517318
rect 175625 517284 175901 517318
rect 176551 517318 177005 517340
rect 175447 517268 175901 517284
rect 176059 517282 176509 517298
rect 174955 517226 175405 517248
rect 176059 517248 176331 517282
rect 176365 517248 176509 517282
rect 176551 517284 176695 517318
rect 176729 517284 177005 517318
rect 177655 517318 178109 517340
rect 176551 517268 177005 517284
rect 177163 517282 177613 517298
rect 176059 517226 176509 517248
rect 177163 517248 177435 517282
rect 177469 517248 177613 517282
rect 177655 517284 177799 517318
rect 177833 517284 178109 517318
rect 178759 517318 179213 517340
rect 177655 517268 178109 517284
rect 178267 517282 178717 517298
rect 177163 517226 177613 517248
rect 178267 517248 178539 517282
rect 178573 517248 178717 517282
rect 178759 517284 178903 517318
rect 178937 517284 179213 517318
rect 179589 517318 179765 517340
rect 178759 517268 179213 517284
rect 179371 517282 179547 517298
rect 178267 517226 178717 517248
rect 179371 517248 179387 517282
rect 179421 517248 179497 517282
rect 179531 517248 179547 517282
rect 179589 517284 179605 517318
rect 179639 517284 179715 517318
rect 179749 517284 179765 517318
rect 180599 517318 181053 517340
rect 179589 517268 179765 517284
rect 180107 517282 180557 517298
rect 179371 517226 179547 517248
rect 180107 517248 180379 517282
rect 180413 517248 180557 517282
rect 180599 517284 180743 517318
rect 180777 517284 181053 517318
rect 181703 517318 182157 517340
rect 180599 517268 181053 517284
rect 181211 517282 181661 517298
rect 180107 517226 180557 517248
rect 181211 517248 181483 517282
rect 181517 517248 181661 517282
rect 181703 517284 181847 517318
rect 181881 517284 182157 517318
rect 182807 517318 183261 517340
rect 181703 517268 182157 517284
rect 182315 517282 182765 517298
rect 181211 517226 181661 517248
rect 182315 517248 182587 517282
rect 182621 517248 182765 517282
rect 182807 517284 182951 517318
rect 182985 517284 183261 517318
rect 183911 517318 184365 517340
rect 182807 517268 183261 517284
rect 183419 517282 183869 517298
rect 182315 517226 182765 517248
rect 183419 517248 183691 517282
rect 183725 517248 183869 517282
rect 183911 517284 184055 517318
rect 184089 517284 184365 517318
rect 184741 517318 184917 517340
rect 183911 517268 184365 517284
rect 184523 517282 184699 517298
rect 183419 517226 183869 517248
rect 184523 517248 184539 517282
rect 184573 517248 184649 517282
rect 184683 517248 184699 517282
rect 184741 517284 184757 517318
rect 184791 517284 184867 517318
rect 184901 517284 184917 517318
rect 185751 517318 186205 517340
rect 184741 517268 184917 517284
rect 185259 517282 185709 517298
rect 184523 517226 184699 517248
rect 185259 517248 185531 517282
rect 185565 517248 185709 517282
rect 185751 517284 185895 517318
rect 185929 517284 186205 517318
rect 186669 517318 186941 517340
rect 187283 517340 187401 517366
rect 187283 517338 187321 517340
rect 185751 517268 186205 517284
rect 186363 517282 186627 517298
rect 185259 517226 185709 517248
rect 186363 517248 186379 517282
rect 186413 517248 186478 517282
rect 186512 517248 186577 517282
rect 186611 517248 186627 517282
rect 186669 517284 186685 517318
rect 186719 517284 186788 517318
rect 186822 517284 186891 517318
rect 186925 517284 186941 517318
rect 186669 517268 186941 517284
rect 187255 517322 187321 517338
rect 187255 517288 187271 517322
rect 187305 517288 187321 517322
rect 187255 517272 187321 517288
rect 187363 517282 187429 517298
rect 186363 517226 186627 517248
rect 187363 517248 187379 517282
rect 187413 517248 187429 517282
rect 187363 517232 187429 517248
rect 187363 517230 187401 517232
rect 172563 517200 173509 517226
rect 173667 517200 174613 517226
rect 174955 517200 175901 517226
rect 176059 517200 177005 517226
rect 177163 517200 178109 517226
rect 178267 517200 179213 517226
rect 179371 517200 179765 517226
rect 180107 517200 181053 517226
rect 181211 517200 182157 517226
rect 182315 517200 183261 517226
rect 183419 517200 184365 517226
rect 184523 517200 184917 517226
rect 185259 517200 186205 517226
rect 186363 517200 186941 517226
rect 187283 517200 187401 517230
rect 172287 517000 172405 517026
rect 172563 517000 173509 517026
rect 173667 517000 174613 517026
rect 174955 517000 175901 517026
rect 176059 517000 177005 517026
rect 177163 517000 178109 517026
rect 178267 517000 179213 517026
rect 179371 517000 179765 517026
rect 180107 517000 181053 517026
rect 181211 517000 182157 517026
rect 182315 517000 183261 517026
rect 183419 517000 184365 517026
rect 184523 517000 184917 517026
rect 185259 517000 186205 517026
rect 186363 517000 186941 517026
rect 187283 517000 187401 517026
rect 172287 516932 172405 516958
rect 172563 516932 173509 516958
rect 173667 516932 174613 516958
rect 174771 516932 175717 516958
rect 175875 516932 176821 516958
rect 176979 516932 177189 516958
rect 177531 516932 178477 516958
rect 178635 516932 179581 516958
rect 179739 516932 180685 516958
rect 180843 516932 181789 516958
rect 181947 516932 182341 516958
rect 182683 516932 183629 516958
rect 183787 516932 184733 516958
rect 184891 516932 185837 516958
rect 185995 516932 186941 516958
rect 187283 516932 187401 516958
rect 172287 516728 172405 516758
rect 172563 516732 173509 516758
rect 173667 516732 174613 516758
rect 174771 516732 175717 516758
rect 175875 516732 176821 516758
rect 176979 516732 177189 516758
rect 177531 516732 178477 516758
rect 178635 516732 179581 516758
rect 179739 516732 180685 516758
rect 180843 516732 181789 516758
rect 181947 516732 182341 516758
rect 182683 516732 183629 516758
rect 183787 516732 184733 516758
rect 184891 516732 185837 516758
rect 185995 516732 186941 516758
rect 172287 516726 172325 516728
rect 172259 516710 172325 516726
rect 172259 516676 172275 516710
rect 172309 516676 172325 516710
rect 172563 516710 173013 516732
rect 172259 516660 172325 516676
rect 172367 516670 172433 516686
rect 172367 516636 172383 516670
rect 172417 516636 172433 516670
rect 172563 516676 172835 516710
rect 172869 516676 173013 516710
rect 173667 516710 174117 516732
rect 172563 516660 173013 516676
rect 173055 516674 173509 516690
rect 172367 516620 172433 516636
rect 173055 516640 173199 516674
rect 173233 516640 173509 516674
rect 173667 516676 173939 516710
rect 173973 516676 174117 516710
rect 174771 516710 175221 516732
rect 173667 516660 174117 516676
rect 174159 516674 174613 516690
rect 172367 516618 172405 516620
rect 173055 516618 173509 516640
rect 174159 516640 174303 516674
rect 174337 516640 174613 516674
rect 174771 516676 175043 516710
rect 175077 516676 175221 516710
rect 175875 516710 176325 516732
rect 176979 516726 177063 516732
rect 174771 516660 175221 516676
rect 175263 516674 175717 516690
rect 174159 516618 174613 516640
rect 175263 516640 175407 516674
rect 175441 516640 175717 516674
rect 175875 516676 176147 516710
rect 176181 516676 176325 516710
rect 176921 516710 177063 516726
rect 175875 516660 176325 516676
rect 176367 516674 176821 516690
rect 175263 516618 175717 516640
rect 176367 516640 176511 516674
rect 176545 516640 176821 516674
rect 176921 516676 176937 516710
rect 176971 516676 177063 516710
rect 177531 516710 177981 516732
rect 176921 516660 177063 516676
rect 177105 516674 177247 516690
rect 176367 516618 176821 516640
rect 177105 516640 177197 516674
rect 177231 516640 177247 516674
rect 177531 516676 177803 516710
rect 177837 516676 177981 516710
rect 178635 516710 179085 516732
rect 177531 516660 177981 516676
rect 178023 516674 178477 516690
rect 177105 516624 177247 516640
rect 178023 516640 178167 516674
rect 178201 516640 178477 516674
rect 178635 516676 178907 516710
rect 178941 516676 179085 516710
rect 179739 516710 180189 516732
rect 178635 516660 179085 516676
rect 179127 516674 179581 516690
rect 177105 516618 177189 516624
rect 178023 516618 178477 516640
rect 179127 516640 179271 516674
rect 179305 516640 179581 516674
rect 179739 516676 180011 516710
rect 180045 516676 180189 516710
rect 180843 516710 181293 516732
rect 179739 516660 180189 516676
rect 180231 516674 180685 516690
rect 179127 516618 179581 516640
rect 180231 516640 180375 516674
rect 180409 516640 180685 516674
rect 180843 516676 181115 516710
rect 181149 516676 181293 516710
rect 181947 516710 182123 516732
rect 180843 516660 181293 516676
rect 181335 516674 181789 516690
rect 180231 516618 180685 516640
rect 181335 516640 181479 516674
rect 181513 516640 181789 516674
rect 181947 516676 181963 516710
rect 181997 516676 182073 516710
rect 182107 516676 182123 516710
rect 182683 516710 183133 516732
rect 181947 516660 182123 516676
rect 182165 516674 182341 516690
rect 181335 516618 181789 516640
rect 182165 516640 182181 516674
rect 182215 516640 182291 516674
rect 182325 516640 182341 516674
rect 182683 516676 182955 516710
rect 182989 516676 183133 516710
rect 183787 516710 184237 516732
rect 182683 516660 183133 516676
rect 183175 516674 183629 516690
rect 182165 516618 182341 516640
rect 183175 516640 183319 516674
rect 183353 516640 183629 516674
rect 183787 516676 184059 516710
rect 184093 516676 184237 516710
rect 184891 516710 185341 516732
rect 183787 516660 184237 516676
rect 184279 516674 184733 516690
rect 183175 516618 183629 516640
rect 184279 516640 184423 516674
rect 184457 516640 184733 516674
rect 184891 516676 185163 516710
rect 185197 516676 185341 516710
rect 185995 516710 186445 516732
rect 187283 516728 187401 516758
rect 184891 516660 185341 516676
rect 185383 516674 185837 516690
rect 184279 516618 184733 516640
rect 185383 516640 185527 516674
rect 185561 516640 185837 516674
rect 185995 516676 186267 516710
rect 186301 516676 186445 516710
rect 187363 516726 187401 516728
rect 187363 516710 187429 516726
rect 185995 516660 186445 516676
rect 186487 516674 186941 516690
rect 185383 516618 185837 516640
rect 186487 516640 186631 516674
rect 186665 516640 186941 516674
rect 186487 516618 186941 516640
rect 187255 516670 187321 516686
rect 187255 516636 187271 516670
rect 187305 516636 187321 516670
rect 187363 516676 187379 516710
rect 187413 516676 187429 516710
rect 187363 516660 187429 516676
rect 187255 516620 187321 516636
rect 172287 516592 172405 516618
rect 172563 516592 173509 516618
rect 173667 516592 174613 516618
rect 174771 516592 175717 516618
rect 175875 516592 176821 516618
rect 176979 516592 177189 516618
rect 177531 516592 178477 516618
rect 178635 516592 179581 516618
rect 179739 516592 180685 516618
rect 180843 516592 181789 516618
rect 181947 516592 182341 516618
rect 182683 516592 183629 516618
rect 183787 516592 184733 516618
rect 184891 516592 185837 516618
rect 185995 516592 186941 516618
rect 187283 516618 187321 516620
rect 187283 516592 187401 516618
rect 172287 516456 172405 516482
rect 172563 516456 173509 516482
rect 173667 516456 174613 516482
rect 174771 516456 175717 516482
rect 175875 516456 176821 516482
rect 176979 516456 177189 516482
rect 177531 516456 178477 516482
rect 178635 516456 179581 516482
rect 179739 516456 180685 516482
rect 180843 516456 181789 516482
rect 181947 516456 182341 516482
rect 182683 516456 183629 516482
rect 183787 516456 184733 516482
rect 184891 516456 185837 516482
rect 185995 516456 186941 516482
rect 187283 516456 187401 516482
rect 172287 516388 172405 516414
rect 172563 516388 173509 516414
rect 173667 516388 174613 516414
rect 174955 516388 175901 516414
rect 176059 516388 177005 516414
rect 177163 516388 178109 516414
rect 178267 516388 179213 516414
rect 179371 516388 179765 516414
rect 180107 516388 181053 516414
rect 181211 516388 182157 516414
rect 182315 516388 183261 516414
rect 183419 516388 184365 516414
rect 184523 516388 184917 516414
rect 185259 516388 186205 516414
rect 186363 516388 186941 516414
rect 187283 516388 187401 516414
rect 172287 516252 172405 516278
rect 172563 516252 173509 516278
rect 173667 516252 174613 516278
rect 174955 516252 175901 516278
rect 176059 516252 177005 516278
rect 177163 516252 178109 516278
rect 178267 516252 179213 516278
rect 179371 516252 179765 516278
rect 180107 516252 181053 516278
rect 181211 516252 182157 516278
rect 182315 516252 183261 516278
rect 183419 516252 184365 516278
rect 184523 516252 184917 516278
rect 185259 516252 186205 516278
rect 186363 516252 186941 516278
rect 172367 516250 172405 516252
rect 172367 516234 172433 516250
rect 172259 516194 172325 516210
rect 172259 516160 172275 516194
rect 172309 516160 172325 516194
rect 172367 516200 172383 516234
rect 172417 516200 172433 516234
rect 173055 516230 173509 516252
rect 172367 516184 172433 516200
rect 172563 516194 173013 516210
rect 172259 516144 172325 516160
rect 172287 516142 172325 516144
rect 172563 516160 172835 516194
rect 172869 516160 173013 516194
rect 173055 516196 173199 516230
rect 173233 516196 173509 516230
rect 174159 516230 174613 516252
rect 173055 516180 173509 516196
rect 173667 516194 174117 516210
rect 172287 516112 172405 516142
rect 172563 516138 173013 516160
rect 173667 516160 173939 516194
rect 173973 516160 174117 516194
rect 174159 516196 174303 516230
rect 174337 516196 174613 516230
rect 175447 516230 175901 516252
rect 174159 516180 174613 516196
rect 174955 516194 175405 516210
rect 173667 516138 174117 516160
rect 174955 516160 175227 516194
rect 175261 516160 175405 516194
rect 175447 516196 175591 516230
rect 175625 516196 175901 516230
rect 176551 516230 177005 516252
rect 175447 516180 175901 516196
rect 176059 516194 176509 516210
rect 174955 516138 175405 516160
rect 176059 516160 176331 516194
rect 176365 516160 176509 516194
rect 176551 516196 176695 516230
rect 176729 516196 177005 516230
rect 177655 516230 178109 516252
rect 176551 516180 177005 516196
rect 177163 516194 177613 516210
rect 176059 516138 176509 516160
rect 177163 516160 177435 516194
rect 177469 516160 177613 516194
rect 177655 516196 177799 516230
rect 177833 516196 178109 516230
rect 178759 516230 179213 516252
rect 177655 516180 178109 516196
rect 178267 516194 178717 516210
rect 177163 516138 177613 516160
rect 178267 516160 178539 516194
rect 178573 516160 178717 516194
rect 178759 516196 178903 516230
rect 178937 516196 179213 516230
rect 179589 516230 179765 516252
rect 178759 516180 179213 516196
rect 179371 516194 179547 516210
rect 178267 516138 178717 516160
rect 179371 516160 179387 516194
rect 179421 516160 179497 516194
rect 179531 516160 179547 516194
rect 179589 516196 179605 516230
rect 179639 516196 179715 516230
rect 179749 516196 179765 516230
rect 180599 516230 181053 516252
rect 179589 516180 179765 516196
rect 180107 516194 180557 516210
rect 179371 516138 179547 516160
rect 180107 516160 180379 516194
rect 180413 516160 180557 516194
rect 180599 516196 180743 516230
rect 180777 516196 181053 516230
rect 181703 516230 182157 516252
rect 180599 516180 181053 516196
rect 181211 516194 181661 516210
rect 180107 516138 180557 516160
rect 181211 516160 181483 516194
rect 181517 516160 181661 516194
rect 181703 516196 181847 516230
rect 181881 516196 182157 516230
rect 182807 516230 183261 516252
rect 181703 516180 182157 516196
rect 182315 516194 182765 516210
rect 181211 516138 181661 516160
rect 182315 516160 182587 516194
rect 182621 516160 182765 516194
rect 182807 516196 182951 516230
rect 182985 516196 183261 516230
rect 183911 516230 184365 516252
rect 182807 516180 183261 516196
rect 183419 516194 183869 516210
rect 182315 516138 182765 516160
rect 183419 516160 183691 516194
rect 183725 516160 183869 516194
rect 183911 516196 184055 516230
rect 184089 516196 184365 516230
rect 184741 516230 184917 516252
rect 183911 516180 184365 516196
rect 184523 516194 184699 516210
rect 183419 516138 183869 516160
rect 184523 516160 184539 516194
rect 184573 516160 184649 516194
rect 184683 516160 184699 516194
rect 184741 516196 184757 516230
rect 184791 516196 184867 516230
rect 184901 516196 184917 516230
rect 185751 516230 186205 516252
rect 184741 516180 184917 516196
rect 185259 516194 185709 516210
rect 184523 516138 184699 516160
rect 185259 516160 185531 516194
rect 185565 516160 185709 516194
rect 185751 516196 185895 516230
rect 185929 516196 186205 516230
rect 186669 516230 186941 516252
rect 187283 516252 187401 516278
rect 187283 516250 187321 516252
rect 185751 516180 186205 516196
rect 186363 516194 186627 516210
rect 185259 516138 185709 516160
rect 186363 516160 186379 516194
rect 186413 516160 186478 516194
rect 186512 516160 186577 516194
rect 186611 516160 186627 516194
rect 186669 516196 186685 516230
rect 186719 516196 186788 516230
rect 186822 516196 186891 516230
rect 186925 516196 186941 516230
rect 186669 516180 186941 516196
rect 187255 516234 187321 516250
rect 187255 516200 187271 516234
rect 187305 516200 187321 516234
rect 187255 516184 187321 516200
rect 187363 516194 187429 516210
rect 186363 516138 186627 516160
rect 187363 516160 187379 516194
rect 187413 516160 187429 516194
rect 187363 516144 187429 516160
rect 187363 516142 187401 516144
rect 172563 516112 173509 516138
rect 173667 516112 174613 516138
rect 174955 516112 175901 516138
rect 176059 516112 177005 516138
rect 177163 516112 178109 516138
rect 178267 516112 179213 516138
rect 179371 516112 179765 516138
rect 180107 516112 181053 516138
rect 181211 516112 182157 516138
rect 182315 516112 183261 516138
rect 183419 516112 184365 516138
rect 184523 516112 184917 516138
rect 185259 516112 186205 516138
rect 186363 516112 186941 516138
rect 187283 516112 187401 516142
rect 172287 515912 172405 515938
rect 172563 515912 173509 515938
rect 173667 515912 174613 515938
rect 174955 515912 175901 515938
rect 176059 515912 177005 515938
rect 177163 515912 178109 515938
rect 178267 515912 179213 515938
rect 179371 515912 179765 515938
rect 180107 515912 181053 515938
rect 181211 515912 182157 515938
rect 182315 515912 183261 515938
rect 183419 515912 184365 515938
rect 184523 515912 184917 515938
rect 185259 515912 186205 515938
rect 186363 515912 186941 515938
rect 187283 515912 187401 515938
rect 172287 515844 172405 515870
rect 172563 515844 173141 515870
rect 173484 515844 173514 515870
rect 173580 515844 173610 515870
rect 173666 515844 173696 515870
rect 173752 515844 173782 515870
rect 173838 515844 173868 515870
rect 174035 515844 174613 515870
rect 174955 515844 175901 515870
rect 176059 515844 177005 515870
rect 177163 515844 177281 515870
rect 177531 515844 178477 515870
rect 178635 515844 179581 515870
rect 179739 515844 179857 515870
rect 180107 515844 181053 515870
rect 181211 515844 181789 515870
rect 182131 515844 182161 515870
rect 182219 515844 182249 515870
rect 182683 515844 183629 515870
rect 183787 515844 184733 515870
rect 184891 515844 185009 515870
rect 185259 515844 186205 515870
rect 186456 515844 186486 515870
rect 186552 515844 186582 515870
rect 186638 515844 186668 515870
rect 186724 515844 186754 515870
rect 186810 515844 186840 515870
rect 187007 515844 187125 515870
rect 187283 515844 187401 515870
rect 172287 515640 172405 515670
rect 172563 515644 173141 515670
rect 174035 515644 174613 515670
rect 174955 515644 175901 515670
rect 176059 515644 177005 515670
rect 172287 515638 172325 515640
rect 172259 515622 172325 515638
rect 172259 515588 172275 515622
rect 172309 515588 172325 515622
rect 172563 515622 172827 515644
rect 172259 515572 172325 515588
rect 172367 515582 172433 515598
rect 172367 515548 172383 515582
rect 172417 515548 172433 515582
rect 172563 515588 172579 515622
rect 172613 515588 172678 515622
rect 172712 515588 172777 515622
rect 172811 515588 172827 515622
rect 173484 515612 173514 515644
rect 172563 515572 172827 515588
rect 172869 515586 173141 515602
rect 172367 515532 172433 515548
rect 172869 515552 172885 515586
rect 172919 515552 172988 515586
rect 173022 515552 173091 515586
rect 173125 515552 173141 515586
rect 172367 515530 172405 515532
rect 172869 515530 173141 515552
rect 173473 515596 173533 515612
rect 173473 515562 173489 515596
rect 173523 515562 173533 515596
rect 173473 515546 173533 515562
rect 173580 515606 173610 515644
rect 173666 515606 173696 515644
rect 173752 515606 173782 515644
rect 173838 515606 173868 515644
rect 173580 515596 173868 515606
rect 173580 515562 173635 515596
rect 173669 515562 173703 515596
rect 173737 515562 173771 515596
rect 173805 515584 173868 515596
rect 174035 515622 174299 515644
rect 174035 515588 174051 515622
rect 174085 515588 174150 515622
rect 174184 515588 174249 515622
rect 174283 515588 174299 515622
rect 174955 515622 175405 515644
rect 173805 515562 173869 515584
rect 174035 515572 174299 515588
rect 174341 515586 174613 515602
rect 173580 515557 173869 515562
rect 173581 515551 173869 515557
rect 172287 515504 172405 515530
rect 172563 515504 173141 515530
rect 173484 515478 173514 515546
rect 173581 515478 173611 515551
rect 173667 515478 173697 515551
rect 173753 515478 173783 515551
rect 173839 515478 173869 515551
rect 174341 515552 174357 515586
rect 174391 515552 174460 515586
rect 174494 515552 174563 515586
rect 174597 515552 174613 515586
rect 174955 515588 175227 515622
rect 175261 515588 175405 515622
rect 176059 515622 176509 515644
rect 177163 515640 177281 515670
rect 177531 515644 178477 515670
rect 178635 515644 179581 515670
rect 177163 515638 177201 515640
rect 174955 515572 175405 515588
rect 175447 515586 175901 515602
rect 174341 515530 174613 515552
rect 175447 515552 175591 515586
rect 175625 515552 175901 515586
rect 176059 515588 176331 515622
rect 176365 515588 176509 515622
rect 177135 515622 177201 515638
rect 176059 515572 176509 515588
rect 176551 515586 177005 515602
rect 175447 515530 175901 515552
rect 176551 515552 176695 515586
rect 176729 515552 177005 515586
rect 177135 515588 177151 515622
rect 177185 515588 177201 515622
rect 177531 515622 177981 515644
rect 177135 515572 177201 515588
rect 177243 515582 177309 515598
rect 176551 515530 177005 515552
rect 177243 515548 177259 515582
rect 177293 515548 177309 515582
rect 177531 515588 177803 515622
rect 177837 515588 177981 515622
rect 178635 515622 179085 515644
rect 179739 515640 179857 515670
rect 180107 515644 181053 515670
rect 181211 515644 181789 515670
rect 179739 515638 179777 515640
rect 177531 515572 177981 515588
rect 178023 515586 178477 515602
rect 177243 515532 177309 515548
rect 178023 515552 178167 515586
rect 178201 515552 178477 515586
rect 178635 515588 178907 515622
rect 178941 515588 179085 515622
rect 179711 515622 179777 515638
rect 178635 515572 179085 515588
rect 179127 515586 179581 515602
rect 177243 515530 177281 515532
rect 178023 515530 178477 515552
rect 179127 515552 179271 515586
rect 179305 515552 179581 515586
rect 179711 515588 179727 515622
rect 179761 515588 179777 515622
rect 180107 515622 180557 515644
rect 179711 515572 179777 515588
rect 179819 515582 179885 515598
rect 179127 515530 179581 515552
rect 179819 515548 179835 515582
rect 179869 515548 179885 515582
rect 180107 515588 180379 515622
rect 180413 515588 180557 515622
rect 181211 515622 181475 515644
rect 182131 515625 182161 515686
rect 182219 515671 182249 515686
rect 182219 515647 182255 515671
rect 180107 515572 180557 515588
rect 180599 515586 181053 515602
rect 179819 515532 179885 515548
rect 180599 515552 180743 515586
rect 180777 515552 181053 515586
rect 181211 515588 181227 515622
rect 181261 515588 181326 515622
rect 181360 515588 181425 515622
rect 181459 515588 181475 515622
rect 182129 515609 182183 515625
rect 181211 515572 181475 515588
rect 181517 515586 181789 515602
rect 179819 515530 179857 515532
rect 180599 515530 181053 515552
rect 181517 515552 181533 515586
rect 181567 515552 181636 515586
rect 181670 515552 181739 515586
rect 181773 515552 181789 515586
rect 182129 515575 182139 515609
rect 182173 515575 182183 515609
rect 182129 515559 182183 515575
rect 182225 515612 182255 515647
rect 182683 515644 183629 515670
rect 183787 515644 184733 515670
rect 182683 515622 183133 515644
rect 182225 515596 182301 515612
rect 182225 515562 182257 515596
rect 182291 515562 182301 515596
rect 182683 515588 182955 515622
rect 182989 515588 183133 515622
rect 183787 515622 184237 515644
rect 184891 515640 185009 515670
rect 185259 515644 186205 515670
rect 184891 515638 184929 515640
rect 182683 515572 183133 515588
rect 183175 515586 183629 515602
rect 181517 515530 181789 515552
rect 174035 515504 174613 515530
rect 174955 515504 175901 515530
rect 176059 515504 177005 515530
rect 177163 515504 177281 515530
rect 177531 515504 178477 515530
rect 178635 515504 179581 515530
rect 179739 515504 179857 515530
rect 180107 515504 181053 515530
rect 181211 515504 181789 515530
rect 182131 515498 182161 515559
rect 182225 515546 182301 515562
rect 183175 515552 183319 515586
rect 183353 515552 183629 515586
rect 183787 515588 184059 515622
rect 184093 515588 184237 515622
rect 184863 515622 184929 515638
rect 183787 515572 184237 515588
rect 184279 515586 184733 515602
rect 182225 515537 182255 515546
rect 182219 515513 182255 515537
rect 183175 515530 183629 515552
rect 184279 515552 184423 515586
rect 184457 515552 184733 515586
rect 184863 515588 184879 515622
rect 184913 515588 184929 515622
rect 185259 515622 185709 515644
rect 184863 515572 184929 515588
rect 184971 515582 185037 515598
rect 184279 515530 184733 515552
rect 184971 515548 184987 515582
rect 185021 515548 185037 515582
rect 185259 515588 185531 515622
rect 185565 515588 185709 515622
rect 186456 515612 186486 515644
rect 185259 515572 185709 515588
rect 185751 515586 186205 515602
rect 184971 515532 185037 515548
rect 185751 515552 185895 515586
rect 185929 515552 186205 515586
rect 184971 515530 185009 515532
rect 185751 515530 186205 515552
rect 186445 515596 186505 515612
rect 186445 515562 186461 515596
rect 186495 515562 186505 515596
rect 186445 515546 186505 515562
rect 186552 515606 186582 515644
rect 186638 515606 186668 515644
rect 186724 515606 186754 515644
rect 186810 515606 186840 515644
rect 187007 515640 187125 515670
rect 187283 515640 187401 515670
rect 187007 515638 187045 515640
rect 186552 515596 186840 515606
rect 186552 515562 186607 515596
rect 186641 515562 186675 515596
rect 186709 515562 186743 515596
rect 186777 515584 186840 515596
rect 186979 515622 187045 515638
rect 186979 515588 186995 515622
rect 187029 515588 187045 515622
rect 187363 515638 187401 515640
rect 187363 515622 187429 515638
rect 186777 515562 186841 515584
rect 186979 515572 187045 515588
rect 187087 515582 187153 515598
rect 186552 515557 186841 515562
rect 186553 515551 186841 515557
rect 182219 515498 182249 515513
rect 182683 515504 183629 515530
rect 183787 515504 184733 515530
rect 184891 515504 185009 515530
rect 185259 515504 186205 515530
rect 186456 515478 186486 515546
rect 186553 515478 186583 515551
rect 186639 515478 186669 515551
rect 186725 515478 186755 515551
rect 186811 515478 186841 515551
rect 187087 515548 187103 515582
rect 187137 515548 187153 515582
rect 187087 515532 187153 515548
rect 187255 515582 187321 515598
rect 187255 515548 187271 515582
rect 187305 515548 187321 515582
rect 187363 515588 187379 515622
rect 187413 515588 187429 515622
rect 187363 515572 187429 515588
rect 187255 515532 187321 515548
rect 187087 515530 187125 515532
rect 187007 515504 187125 515530
rect 187283 515530 187321 515532
rect 187283 515504 187401 515530
rect 172287 515368 172405 515394
rect 172563 515368 173141 515394
rect 173484 515368 173514 515394
rect 173581 515368 173611 515394
rect 173667 515368 173697 515394
rect 173753 515368 173783 515394
rect 173839 515368 173869 515394
rect 174035 515368 174613 515394
rect 174955 515368 175901 515394
rect 176059 515368 177005 515394
rect 177163 515368 177281 515394
rect 177531 515368 178477 515394
rect 178635 515368 179581 515394
rect 179739 515368 179857 515394
rect 180107 515368 181053 515394
rect 181211 515368 181789 515394
rect 182131 515368 182161 515394
rect 182219 515368 182249 515394
rect 182683 515368 183629 515394
rect 183787 515368 184733 515394
rect 184891 515368 185009 515394
rect 185259 515368 186205 515394
rect 186456 515368 186486 515394
rect 186553 515368 186583 515394
rect 186639 515368 186669 515394
rect 186725 515368 186755 515394
rect 186811 515368 186841 515394
rect 187007 515368 187125 515394
rect 187283 515368 187401 515394
<< polycont >>
rect 164728 541085 164762 541119
rect 165031 541092 165065 541126
rect 165223 541092 165257 541126
rect 165415 541092 165449 541126
rect 165607 541092 165641 541126
rect 165799 541092 165833 541126
rect 165991 541092 166025 541126
rect 166408 541085 166442 541119
rect 166208 540285 166242 540319
rect 164728 539975 164762 540009
rect 164935 539982 164969 540016
rect 165127 539982 165161 540016
rect 165319 539982 165353 540016
rect 165511 539982 165545 540016
rect 165703 539982 165737 540016
rect 165895 539982 165929 540016
rect 166208 539975 166242 540009
rect 166408 539975 166442 540009
rect 168528 541085 168562 541119
rect 168831 541092 168865 541126
rect 169023 541092 169057 541126
rect 169215 541092 169249 541126
rect 169407 541092 169441 541126
rect 169599 541092 169633 541126
rect 169791 541092 169825 541126
rect 170208 541085 170242 541119
rect 170008 540285 170042 540319
rect 168528 539975 168562 540009
rect 168735 539982 168769 540016
rect 168927 539982 168961 540016
rect 169119 539982 169153 540016
rect 169311 539982 169345 540016
rect 169503 539982 169537 540016
rect 169695 539982 169729 540016
rect 170008 539975 170042 540009
rect 170208 539975 170242 540009
rect 172228 541085 172262 541119
rect 172531 541092 172565 541126
rect 172723 541092 172757 541126
rect 172915 541092 172949 541126
rect 173107 541092 173141 541126
rect 173299 541092 173333 541126
rect 173491 541092 173525 541126
rect 173908 541085 173942 541119
rect 173708 540285 173742 540319
rect 172228 539975 172262 540009
rect 172435 539982 172469 540016
rect 172627 539982 172661 540016
rect 172819 539982 172853 540016
rect 173011 539982 173045 540016
rect 173203 539982 173237 540016
rect 173395 539982 173429 540016
rect 173708 539975 173742 540009
rect 173908 539975 173942 540009
rect 175728 541085 175762 541119
rect 176031 541092 176065 541126
rect 176223 541092 176257 541126
rect 176415 541092 176449 541126
rect 176607 541092 176641 541126
rect 176799 541092 176833 541126
rect 176991 541092 177025 541126
rect 177408 541085 177442 541119
rect 177208 540285 177242 540319
rect 175728 539975 175762 540009
rect 175935 539982 175969 540016
rect 176127 539982 176161 540016
rect 176319 539982 176353 540016
rect 176511 539982 176545 540016
rect 176703 539982 176737 540016
rect 176895 539982 176929 540016
rect 177208 539975 177242 540009
rect 177408 539975 177442 540009
rect 179328 541085 179362 541119
rect 179631 541092 179665 541126
rect 179823 541092 179857 541126
rect 180015 541092 180049 541126
rect 180207 541092 180241 541126
rect 180399 541092 180433 541126
rect 180591 541092 180625 541126
rect 181008 541085 181042 541119
rect 180808 540285 180842 540319
rect 179328 539975 179362 540009
rect 179535 539982 179569 540016
rect 179727 539982 179761 540016
rect 179919 539982 179953 540016
rect 180111 539982 180145 540016
rect 180303 539982 180337 540016
rect 180495 539982 180529 540016
rect 180808 539975 180842 540009
rect 181008 539975 181042 540009
rect 182628 541085 182662 541119
rect 182931 541092 182965 541126
rect 183123 541092 183157 541126
rect 183315 541092 183349 541126
rect 183507 541092 183541 541126
rect 183699 541092 183733 541126
rect 183891 541092 183925 541126
rect 184308 541085 184342 541119
rect 184108 540285 184142 540319
rect 182628 539975 182662 540009
rect 182835 539982 182869 540016
rect 183027 539982 183061 540016
rect 183219 539982 183253 540016
rect 183411 539982 183445 540016
rect 183603 539982 183637 540016
rect 183795 539982 183829 540016
rect 184108 539975 184142 540009
rect 184308 539975 184342 540009
rect 185928 541085 185962 541119
rect 186231 541092 186265 541126
rect 186423 541092 186457 541126
rect 186615 541092 186649 541126
rect 186807 541092 186841 541126
rect 186999 541092 187033 541126
rect 187191 541092 187225 541126
rect 187608 541085 187642 541119
rect 187408 540285 187442 540319
rect 185928 539975 185962 540009
rect 186135 539982 186169 540016
rect 186327 539982 186361 540016
rect 186519 539982 186553 540016
rect 186711 539982 186745 540016
rect 186903 539982 186937 540016
rect 187095 539982 187129 540016
rect 187408 539975 187442 540009
rect 187608 539975 187642 540009
rect 189228 541085 189262 541119
rect 189531 541092 189565 541126
rect 189723 541092 189757 541126
rect 189915 541092 189949 541126
rect 190107 541092 190141 541126
rect 190299 541092 190333 541126
rect 190491 541092 190525 541126
rect 190908 541085 190942 541119
rect 190708 540285 190742 540319
rect 189228 539975 189262 540009
rect 189435 539982 189469 540016
rect 189627 539982 189661 540016
rect 189819 539982 189853 540016
rect 190011 539982 190045 540016
rect 190203 539982 190237 540016
rect 190395 539982 190429 540016
rect 190708 539975 190742 540009
rect 190908 539975 190942 540009
rect 158726 538435 158894 538469
rect 159102 538435 159270 538469
rect 159360 538435 159528 538469
rect 159618 538435 159786 538469
rect 159876 538435 160044 538469
rect 160134 538435 160302 538469
rect 160392 538435 160560 538469
rect 160650 538435 160818 538469
rect 160908 538435 161076 538469
rect 161166 538435 161334 538469
rect 161546 538435 161714 538469
rect 161946 538435 162114 538469
rect 162326 538435 162494 538469
rect 158726 538125 158894 538159
rect 159102 538125 159270 538159
rect 159360 538125 159528 538159
rect 159618 538125 159786 538159
rect 159876 538125 160044 538159
rect 160134 538125 160302 538159
rect 160392 538125 160560 538159
rect 160650 538125 160818 538159
rect 160908 538125 161076 538159
rect 161166 538125 161334 538159
rect 161546 538125 161714 538159
rect 161946 538125 162114 538159
rect 162326 538125 162494 538159
rect 164712 539572 164746 539606
rect 165035 539579 165069 539613
rect 165227 539579 165261 539613
rect 165419 539579 165453 539613
rect 165611 539579 165645 539613
rect 165803 539579 165837 539613
rect 165995 539579 166029 539613
rect 166212 539572 166246 539606
rect 166412 539572 166446 539606
rect 166212 538844 166246 538878
rect 164712 538444 164746 538478
rect 164939 538451 164973 538485
rect 165131 538451 165165 538485
rect 165323 538451 165357 538485
rect 165515 538451 165549 538485
rect 165707 538451 165741 538485
rect 165899 538451 165933 538485
rect 166412 538444 166446 538478
rect 168512 539572 168546 539606
rect 168835 539579 168869 539613
rect 169027 539579 169061 539613
rect 169219 539579 169253 539613
rect 169411 539579 169445 539613
rect 169603 539579 169637 539613
rect 169795 539579 169829 539613
rect 170012 539572 170046 539606
rect 170212 539572 170246 539606
rect 170012 538844 170046 538878
rect 168512 538444 168546 538478
rect 168739 538451 168773 538485
rect 168931 538451 168965 538485
rect 169123 538451 169157 538485
rect 169315 538451 169349 538485
rect 169507 538451 169541 538485
rect 169699 538451 169733 538485
rect 170212 538444 170246 538478
rect 172212 539572 172246 539606
rect 172535 539579 172569 539613
rect 172727 539579 172761 539613
rect 172919 539579 172953 539613
rect 173111 539579 173145 539613
rect 173303 539579 173337 539613
rect 173495 539579 173529 539613
rect 173712 539572 173746 539606
rect 173912 539572 173946 539606
rect 173712 538844 173746 538878
rect 172212 538444 172246 538478
rect 172439 538451 172473 538485
rect 172631 538451 172665 538485
rect 172823 538451 172857 538485
rect 173015 538451 173049 538485
rect 173207 538451 173241 538485
rect 173399 538451 173433 538485
rect 173912 538444 173946 538478
rect 175712 539572 175746 539606
rect 176035 539579 176069 539613
rect 176227 539579 176261 539613
rect 176419 539579 176453 539613
rect 176611 539579 176645 539613
rect 176803 539579 176837 539613
rect 176995 539579 177029 539613
rect 177212 539572 177246 539606
rect 177412 539572 177446 539606
rect 177212 538844 177246 538878
rect 175712 538444 175746 538478
rect 175939 538451 175973 538485
rect 176131 538451 176165 538485
rect 176323 538451 176357 538485
rect 176515 538451 176549 538485
rect 176707 538451 176741 538485
rect 176899 538451 176933 538485
rect 177412 538444 177446 538478
rect 179312 539572 179346 539606
rect 179635 539579 179669 539613
rect 179827 539579 179861 539613
rect 180019 539579 180053 539613
rect 180211 539579 180245 539613
rect 180403 539579 180437 539613
rect 180595 539579 180629 539613
rect 180812 539572 180846 539606
rect 181012 539572 181046 539606
rect 180812 538844 180846 538878
rect 179312 538444 179346 538478
rect 179539 538451 179573 538485
rect 179731 538451 179765 538485
rect 179923 538451 179957 538485
rect 180115 538451 180149 538485
rect 180307 538451 180341 538485
rect 180499 538451 180533 538485
rect 181012 538444 181046 538478
rect 182612 539572 182646 539606
rect 182935 539579 182969 539613
rect 183127 539579 183161 539613
rect 183319 539579 183353 539613
rect 183511 539579 183545 539613
rect 183703 539579 183737 539613
rect 183895 539579 183929 539613
rect 184112 539572 184146 539606
rect 184312 539572 184346 539606
rect 184112 538844 184146 538878
rect 182612 538444 182646 538478
rect 182839 538451 182873 538485
rect 183031 538451 183065 538485
rect 183223 538451 183257 538485
rect 183415 538451 183449 538485
rect 183607 538451 183641 538485
rect 183799 538451 183833 538485
rect 184312 538444 184346 538478
rect 185912 539572 185946 539606
rect 186235 539579 186269 539613
rect 186427 539579 186461 539613
rect 186619 539579 186653 539613
rect 186811 539579 186845 539613
rect 187003 539579 187037 539613
rect 187195 539579 187229 539613
rect 187412 539572 187446 539606
rect 187612 539572 187646 539606
rect 187412 538844 187446 538878
rect 185912 538444 185946 538478
rect 186139 538451 186173 538485
rect 186331 538451 186365 538485
rect 186523 538451 186557 538485
rect 186715 538451 186749 538485
rect 186907 538451 186941 538485
rect 187099 538451 187133 538485
rect 187612 538444 187646 538478
rect 189212 539572 189246 539606
rect 189535 539579 189569 539613
rect 189727 539579 189761 539613
rect 189919 539579 189953 539613
rect 190111 539579 190145 539613
rect 190303 539579 190337 539613
rect 190495 539579 190529 539613
rect 190712 539572 190746 539606
rect 190912 539572 190946 539606
rect 190712 538844 190746 538878
rect 189212 538444 189246 538478
rect 189439 538451 189473 538485
rect 189631 538451 189665 538485
rect 189823 538451 189857 538485
rect 190015 538451 190049 538485
rect 190207 538451 190241 538485
rect 190399 538451 190433 538485
rect 190912 538444 190946 538478
rect 161302 537672 161336 537706
rect 161506 537672 161540 537706
rect 161698 537672 161732 537706
rect 161906 537672 161940 537706
rect 162098 537672 162132 537706
rect 162322 537672 162356 537706
rect 161302 536944 161336 536978
rect 161602 536944 161636 536978
rect 162002 536944 162036 536978
rect 162322 536944 162356 536978
rect 157810 536652 157978 536686
rect 158188 536652 158356 536686
rect 158446 536652 158614 536686
rect 158704 536652 158872 536686
rect 158962 536652 159130 536686
rect 159220 536652 159388 536686
rect 159478 536652 159646 536686
rect 159736 536652 159904 536686
rect 159994 536652 160162 536686
rect 160252 536652 160420 536686
rect 160510 536652 160678 536686
rect 160894 536652 161062 536686
rect 161152 536652 161320 536686
rect 161410 536652 161578 536686
rect 161792 536652 161960 536686
rect 162050 536652 162218 536686
rect 162430 536652 162598 536686
rect 157810 535924 157978 535958
rect 158188 535924 158356 535958
rect 158446 535924 158614 535958
rect 158704 535924 158872 535958
rect 158962 535924 159130 535958
rect 159220 535924 159388 535958
rect 159478 535924 159646 535958
rect 159736 535924 159904 535958
rect 159994 535924 160162 535958
rect 160252 535924 160420 535958
rect 160510 535924 160678 535958
rect 160894 535924 161062 535958
rect 161152 535924 161320 535958
rect 161410 535924 161578 535958
rect 161792 535924 161960 535958
rect 162050 535924 162218 535958
rect 162430 535924 162598 535958
rect 172275 530304 172309 530338
rect 172383 530344 172417 530378
rect 172635 530330 172669 530364
rect 172703 530330 172737 530364
rect 172771 530330 172805 530364
rect 172917 530330 172951 530364
rect 173387 530304 173421 530338
rect 173751 530340 173785 530374
rect 174235 530304 174269 530338
rect 174345 530304 174379 530338
rect 174453 530340 174487 530374
rect 174563 530340 174597 530374
rect 175027 530330 175061 530364
rect 175095 530330 175129 530364
rect 175163 530330 175197 530364
rect 175309 530330 175343 530364
rect 175614 530330 175648 530364
rect 175889 530338 175923 530372
rect 175985 530366 176019 530400
rect 175812 530230 175846 530264
rect 176129 530340 176163 530374
rect 176225 530388 176259 530422
rect 176090 530214 176124 530248
rect 176373 530328 176407 530362
rect 176469 530376 176503 530410
rect 176724 530382 176758 530416
rect 176826 530376 176860 530410
rect 176555 530240 176589 530274
rect 176985 530269 177019 530303
rect 176804 530214 176838 530248
rect 177192 530315 177226 530349
rect 177294 530330 177328 530364
rect 177743 530330 177777 530364
rect 177939 530330 177973 530364
rect 178143 530330 178177 530364
rect 178257 530330 178291 530364
rect 178457 530317 178491 530351
rect 178577 530330 178611 530364
rect 178799 530330 178833 530364
rect 178867 530330 178901 530364
rect 178935 530330 178969 530364
rect 179081 530330 179115 530364
rect 179285 530330 179319 530364
rect 179431 530330 179465 530364
rect 179499 530330 179533 530364
rect 179567 530330 179601 530364
rect 180298 530330 180332 530364
rect 180394 530330 180428 530364
rect 180535 530366 180569 530400
rect 180631 530366 180665 530400
rect 180793 530366 180827 530400
rect 180703 530253 180737 530287
rect 180871 530253 180905 530287
rect 181345 530366 181379 530400
rect 181507 530366 181541 530400
rect 181267 530253 181301 530287
rect 181603 530366 181637 530400
rect 181435 530253 181469 530287
rect 181744 530330 181778 530364
rect 181840 530330 181874 530364
rect 182045 530330 182079 530364
rect 182191 530330 182225 530364
rect 182259 530330 182293 530364
rect 182327 530330 182361 530364
rect 182641 530304 182675 530338
rect 182901 530340 182935 530374
rect 183149 530330 183183 530364
rect 183295 530330 183329 530364
rect 183363 530330 183397 530364
rect 183431 530330 183465 530364
rect 183967 530304 184001 530338
rect 184331 530340 184365 530374
rect 184757 530304 184791 530338
rect 185017 530340 185051 530374
rect 186999 530494 187033 530528
rect 186999 530426 187033 530460
rect 185265 530330 185299 530364
rect 185411 530330 185445 530364
rect 185479 530330 185513 530364
rect 185547 530330 185581 530364
rect 186083 530304 186117 530338
rect 186447 530340 186481 530374
rect 186999 530163 187033 530197
rect 186999 530095 187033 530129
rect 187099 530498 187133 530532
rect 187099 530430 187133 530464
rect 187271 530344 187305 530378
rect 187379 530304 187413 530338
rect 187099 530163 187133 530197
rect 187099 530095 187133 530129
rect 172275 529732 172309 529766
rect 172383 529692 172417 529726
rect 172835 529732 172869 529766
rect 173199 529696 173233 529730
rect 173939 529732 173973 529766
rect 174303 529696 174337 529730
rect 174865 529706 174899 529740
rect 174979 529706 175013 529740
rect 175183 529706 175217 529740
rect 175379 529706 175413 529740
rect 175552 529706 175586 529740
rect 175654 529721 175688 529755
rect 176042 529822 176076 529856
rect 175861 529767 175895 529801
rect 176291 529796 176325 529830
rect 176020 529660 176054 529694
rect 176122 529654 176156 529688
rect 176377 529660 176411 529694
rect 176473 529708 176507 529742
rect 176756 529822 176790 529856
rect 176621 529648 176655 529682
rect 176717 529696 176751 529730
rect 177034 529806 177068 529840
rect 176861 529670 176895 529704
rect 176957 529698 176991 529732
rect 177232 529706 177266 529740
rect 177679 529783 177713 529817
rect 177847 529783 177881 529817
rect 178664 529806 178698 529840
rect 177757 529670 177791 529704
rect 177919 529670 177953 529704
rect 178015 529670 178049 529704
rect 178156 529706 178190 529740
rect 178252 529706 178286 529740
rect 178466 529706 178500 529740
rect 178741 529698 178775 529732
rect 178942 529822 178976 529856
rect 178837 529670 178871 529704
rect 178981 529696 179015 529730
rect 179225 529708 179259 529742
rect 179407 529796 179441 529830
rect 179077 529648 179111 529682
rect 179321 529660 179355 529694
rect 179656 529822 179690 529856
rect 179837 529767 179871 529801
rect 179576 529654 179610 529688
rect 179678 529660 179712 529694
rect 180044 529721 180078 529755
rect 180146 529706 180180 529740
rect 180244 529706 180278 529740
rect 180346 529721 180380 529755
rect 180734 529822 180768 529856
rect 180553 529767 180587 529801
rect 180983 529796 181017 529830
rect 180712 529660 180746 529694
rect 180814 529654 180848 529688
rect 181069 529660 181103 529694
rect 181165 529708 181199 529742
rect 181448 529822 181482 529856
rect 181313 529648 181347 529682
rect 181409 529696 181443 529730
rect 181726 529806 181760 529840
rect 181553 529670 181587 529704
rect 181649 529698 181683 529732
rect 181924 529706 181958 529740
rect 182089 529732 182123 529766
rect 182349 529696 182383 529730
rect 182711 529706 182745 529740
rect 182907 529706 182941 529740
rect 183111 529706 183145 529740
rect 183225 529706 183259 529740
rect 183691 529732 183725 529766
rect 184055 529696 184089 529730
rect 184795 529732 184829 529766
rect 185159 529696 185193 529730
rect 185899 529732 185933 529766
rect 186263 529696 186297 529730
rect 186747 529732 186781 529766
rect 186857 529732 186891 529766
rect 186965 529696 186999 529730
rect 187075 529696 187109 529730
rect 187271 529692 187305 529726
rect 187379 529732 187413 529766
rect 172275 529216 172309 529250
rect 172383 529256 172417 529290
rect 172835 529216 172869 529250
rect 173199 529252 173233 529286
rect 173939 529216 173973 529250
rect 174303 529252 174337 529286
rect 175273 529278 175307 529312
rect 175435 529278 175469 529312
rect 175195 529165 175229 529199
rect 175531 529278 175565 529312
rect 175363 529165 175397 529199
rect 175672 529242 175706 529276
rect 175768 529242 175802 529276
rect 176210 529242 176244 529276
rect 176278 529242 176312 529276
rect 176346 529242 176380 529276
rect 176414 529242 176448 529276
rect 176482 529242 176516 529276
rect 176550 529242 176584 529276
rect 176618 529242 176652 529276
rect 176686 529242 176720 529276
rect 176754 529242 176788 529276
rect 176822 529242 176856 529276
rect 176890 529242 176924 529276
rect 176958 529242 176992 529276
rect 177026 529242 177060 529276
rect 177094 529242 177128 529276
rect 177162 529242 177196 529276
rect 177230 529242 177264 529276
rect 177657 529242 177691 529276
rect 177760 529242 177794 529276
rect 177862 529227 177896 529261
rect 178228 529288 178262 529322
rect 178330 529294 178364 529328
rect 178069 529181 178103 529215
rect 178250 529126 178284 529160
rect 178585 529288 178619 529322
rect 178829 529300 178863 529334
rect 178499 529152 178533 529186
rect 178681 529240 178715 529274
rect 178925 529252 178959 529286
rect 179069 529278 179103 529312
rect 178964 529126 178998 529160
rect 179165 529250 179199 529284
rect 179440 529242 179474 529276
rect 179697 529242 179731 529276
rect 179242 529142 179276 529176
rect 179817 529229 179851 529263
rect 180123 529216 180157 529250
rect 180233 529216 180267 529250
rect 180341 529252 180375 529286
rect 180451 529252 180485 529286
rect 180709 529242 180743 529276
rect 181136 529242 181170 529276
rect 181204 529242 181238 529276
rect 181272 529242 181306 529276
rect 181340 529242 181374 529276
rect 181408 529242 181442 529276
rect 181476 529242 181510 529276
rect 181544 529242 181578 529276
rect 181612 529242 181646 529276
rect 181680 529242 181714 529276
rect 181748 529242 181782 529276
rect 181816 529242 181850 529276
rect 181884 529242 181918 529276
rect 181952 529242 181986 529276
rect 182020 529242 182054 529276
rect 182088 529242 182122 529276
rect 182156 529242 182190 529276
rect 182597 529229 182631 529263
rect 182717 529242 182751 529276
rect 183139 529216 183173 529250
rect 183503 529252 183537 529286
rect 184243 529216 184277 529250
rect 184607 529252 184641 529286
rect 185531 529216 185565 529250
rect 185895 529252 185929 529286
rect 186379 529216 186413 529250
rect 186478 529216 186512 529250
rect 186577 529216 186611 529250
rect 186685 529252 186719 529286
rect 186788 529252 186822 529286
rect 186891 529252 186925 529286
rect 187271 529256 187305 529290
rect 187379 529216 187413 529250
rect 172275 528644 172309 528678
rect 172383 528604 172417 528638
rect 172835 528644 172869 528678
rect 173199 528608 173233 528642
rect 173939 528644 173973 528678
rect 174303 528608 174337 528642
rect 175043 528644 175077 528678
rect 175407 528608 175441 528642
rect 175925 528618 175959 528652
rect 176575 528695 176609 528729
rect 176045 528631 176079 528665
rect 176201 528618 176235 528652
rect 176321 528631 176355 528665
rect 176743 528695 176777 528729
rect 176653 528582 176687 528616
rect 176815 528582 176849 528616
rect 176911 528582 176945 528616
rect 177052 528618 177086 528652
rect 177148 528618 177182 528652
rect 177559 528618 177593 528652
rect 177755 528618 177789 528652
rect 177959 528618 177993 528652
rect 178073 528618 178107 528652
rect 178409 528618 178443 528652
rect 178836 528618 178870 528652
rect 178904 528618 178938 528652
rect 178972 528618 179006 528652
rect 179040 528618 179074 528652
rect 179108 528618 179142 528652
rect 179176 528618 179210 528652
rect 179244 528618 179278 528652
rect 179312 528618 179346 528652
rect 179380 528618 179414 528652
rect 179448 528618 179482 528652
rect 179516 528618 179550 528652
rect 179584 528618 179618 528652
rect 179652 528618 179686 528652
rect 179720 528618 179754 528652
rect 179788 528618 179822 528652
rect 179856 528618 179890 528652
rect 180249 528618 180283 528652
rect 180369 528631 180403 528665
rect 180520 528618 180554 528652
rect 180622 528633 180656 528667
rect 181010 528734 181044 528768
rect 180829 528679 180863 528713
rect 181259 528708 181293 528742
rect 180988 528572 181022 528606
rect 181090 528566 181124 528600
rect 181345 528572 181379 528606
rect 181441 528620 181475 528654
rect 181724 528734 181758 528768
rect 181589 528560 181623 528594
rect 181685 528608 181719 528642
rect 182002 528718 182036 528752
rect 181829 528582 181863 528616
rect 181925 528610 181959 528644
rect 182200 528618 182234 528652
rect 182955 528644 182989 528678
rect 183319 528608 183353 528642
rect 184059 528644 184093 528678
rect 184423 528608 184457 528642
rect 185163 528644 185197 528678
rect 185527 528608 185561 528642
rect 186267 528644 186301 528678
rect 186631 528608 186665 528642
rect 187271 528604 187305 528638
rect 187379 528644 187413 528678
rect 172275 528128 172309 528162
rect 172383 528168 172417 528202
rect 172835 528128 172869 528162
rect 173199 528164 173233 528198
rect 173939 528128 173973 528162
rect 174303 528164 174337 528198
rect 175227 528128 175261 528162
rect 175591 528164 175625 528198
rect 176104 528154 176138 528188
rect 176206 528139 176240 528173
rect 176572 528200 176606 528234
rect 176674 528206 176708 528240
rect 176413 528093 176447 528127
rect 176594 528038 176628 528072
rect 176929 528200 176963 528234
rect 177173 528212 177207 528246
rect 176843 528064 176877 528098
rect 177025 528152 177059 528186
rect 177269 528164 177303 528198
rect 177413 528190 177447 528224
rect 177308 528038 177342 528072
rect 177509 528162 177543 528196
rect 177784 528154 177818 528188
rect 177997 528141 178031 528175
rect 178117 528154 178151 528188
rect 177586 528054 177620 528088
rect 178283 528128 178317 528162
rect 178382 528128 178416 528162
rect 178481 528128 178515 528162
rect 178589 528164 178623 528198
rect 178692 528164 178726 528198
rect 178795 528164 178829 528198
rect 179010 528154 179044 528188
rect 179106 528154 179140 528188
rect 179247 528190 179281 528224
rect 179343 528190 179377 528224
rect 179505 528190 179539 528224
rect 179415 528077 179449 528111
rect 179583 528077 179617 528111
rect 180123 528128 180157 528162
rect 180222 528128 180256 528162
rect 180321 528128 180355 528162
rect 180429 528164 180463 528198
rect 180532 528164 180566 528198
rect 180635 528164 180669 528198
rect 181034 528154 181068 528188
rect 181130 528154 181164 528188
rect 181271 528190 181305 528224
rect 181367 528190 181401 528224
rect 181529 528190 181563 528224
rect 181439 528077 181473 528111
rect 181607 528077 181641 528111
rect 182127 528128 182161 528162
rect 182491 528164 182525 528198
rect 183231 528128 183265 528162
rect 183595 528164 183629 528198
rect 184335 528128 184369 528162
rect 184699 528164 184733 528198
rect 185531 528128 185565 528162
rect 185895 528164 185929 528198
rect 186379 528128 186413 528162
rect 186478 528128 186512 528162
rect 186577 528128 186611 528162
rect 186685 528164 186719 528198
rect 186788 528164 186822 528198
rect 186891 528164 186925 528198
rect 187271 528168 187305 528202
rect 187379 528128 187413 528162
rect 172275 527556 172309 527590
rect 172383 527516 172417 527550
rect 172835 527556 172869 527590
rect 173199 527520 173233 527554
rect 173939 527556 173973 527590
rect 174303 527520 174337 527554
rect 175043 527556 175077 527590
rect 175407 527520 175441 527554
rect 175891 527556 175925 527590
rect 176001 527556 176035 527590
rect 176109 527520 176143 527554
rect 176219 527520 176253 527554
rect 176455 527530 176489 527564
rect 176651 527530 176685 527564
rect 176855 527530 176889 527564
rect 176969 527530 177003 527564
rect 177151 527556 177185 527590
rect 177259 527516 177293 527550
rect 177803 527556 177837 527590
rect 178167 527520 178201 527554
rect 178593 527556 178627 527590
rect 178853 527520 178887 527554
rect 179031 527530 179065 527564
rect 179227 527530 179261 527564
rect 179431 527530 179465 527564
rect 179545 527530 179579 527564
rect 180011 527556 180045 527590
rect 180375 527520 180409 527554
rect 181115 527556 181149 527590
rect 181479 527520 181513 527554
rect 181963 527556 181997 527590
rect 182073 527556 182107 527590
rect 182181 527520 182215 527554
rect 182291 527520 182325 527554
rect 182955 527556 182989 527590
rect 183319 527520 183353 527554
rect 184059 527556 184093 527590
rect 184423 527520 184457 527554
rect 185163 527556 185197 527590
rect 185527 527520 185561 527554
rect 186267 527556 186301 527590
rect 186631 527520 186665 527554
rect 187271 527516 187305 527550
rect 187379 527556 187413 527590
rect 172275 527040 172309 527074
rect 172383 527080 172417 527114
rect 172835 527040 172869 527074
rect 173199 527076 173233 527110
rect 173939 527040 173973 527074
rect 174303 527076 174337 527110
rect 175227 527040 175261 527074
rect 175591 527076 175625 527110
rect 176331 527040 176365 527074
rect 176695 527076 176729 527110
rect 177435 527040 177469 527074
rect 177799 527076 177833 527110
rect 178539 527040 178573 527074
rect 178903 527076 178937 527110
rect 179387 527040 179421 527074
rect 179497 527040 179531 527074
rect 179605 527076 179639 527110
rect 179715 527076 179749 527110
rect 180379 527040 180413 527074
rect 180743 527076 180777 527110
rect 181483 527040 181517 527074
rect 181847 527076 181881 527110
rect 182587 527040 182621 527074
rect 182951 527076 182985 527110
rect 183691 527040 183725 527074
rect 184055 527076 184089 527110
rect 184539 527040 184573 527074
rect 184649 527040 184683 527074
rect 184757 527076 184791 527110
rect 184867 527076 184901 527110
rect 185531 527040 185565 527074
rect 185895 527076 185929 527110
rect 186379 527040 186413 527074
rect 186478 527040 186512 527074
rect 186577 527040 186611 527074
rect 186685 527076 186719 527110
rect 186788 527076 186822 527110
rect 186891 527076 186925 527110
rect 187271 527080 187305 527114
rect 187379 527040 187413 527074
rect 172275 526468 172309 526502
rect 172383 526428 172417 526462
rect 172835 526468 172869 526502
rect 173199 526432 173233 526466
rect 173939 526468 173973 526502
rect 174303 526432 174337 526466
rect 175043 526468 175077 526502
rect 175407 526432 175441 526466
rect 176147 526468 176181 526502
rect 176511 526432 176545 526466
rect 176937 526468 176971 526502
rect 177197 526432 177231 526466
rect 177803 526468 177837 526502
rect 178167 526432 178201 526466
rect 178907 526468 178941 526502
rect 179271 526432 179305 526466
rect 180011 526468 180045 526502
rect 180375 526432 180409 526466
rect 181115 526468 181149 526502
rect 181479 526432 181513 526466
rect 181963 526468 181997 526502
rect 182073 526468 182107 526502
rect 182181 526432 182215 526466
rect 182291 526432 182325 526466
rect 182955 526468 182989 526502
rect 183319 526432 183353 526466
rect 184059 526468 184093 526502
rect 184423 526432 184457 526466
rect 185163 526468 185197 526502
rect 185527 526432 185561 526466
rect 186267 526468 186301 526502
rect 186631 526432 186665 526466
rect 187271 526428 187305 526462
rect 187379 526468 187413 526502
rect 172275 525952 172309 525986
rect 172383 525992 172417 526026
rect 172835 525952 172869 525986
rect 173199 525988 173233 526022
rect 173939 525952 173973 525986
rect 174303 525988 174337 526022
rect 175227 525952 175261 525986
rect 175591 525988 175625 526022
rect 176331 525952 176365 525986
rect 176695 525988 176729 526022
rect 177435 525952 177469 525986
rect 177799 525988 177833 526022
rect 178539 525952 178573 525986
rect 178903 525988 178937 526022
rect 179387 525952 179421 525986
rect 179497 525952 179531 525986
rect 179605 525988 179639 526022
rect 179715 525988 179749 526022
rect 180379 525952 180413 525986
rect 180743 525988 180777 526022
rect 181483 525952 181517 525986
rect 181847 525988 181881 526022
rect 182587 525952 182621 525986
rect 182951 525988 182985 526022
rect 183691 525952 183725 525986
rect 184055 525988 184089 526022
rect 184539 525952 184573 525986
rect 184649 525952 184683 525986
rect 184757 525988 184791 526022
rect 184867 525988 184901 526022
rect 185531 525952 185565 525986
rect 185895 525988 185929 526022
rect 186379 525952 186413 525986
rect 186478 525952 186512 525986
rect 186577 525952 186611 525986
rect 186685 525988 186719 526022
rect 186788 525988 186822 526022
rect 186891 525988 186925 526022
rect 187271 525992 187305 526026
rect 187379 525952 187413 525986
rect 172275 525380 172309 525414
rect 172383 525340 172417 525374
rect 172835 525380 172869 525414
rect 173199 525344 173233 525378
rect 173939 525380 173973 525414
rect 174303 525344 174337 525378
rect 175043 525380 175077 525414
rect 175407 525344 175441 525378
rect 176147 525380 176181 525414
rect 176511 525344 176545 525378
rect 176937 525380 176971 525414
rect 177197 525344 177231 525378
rect 177803 525380 177837 525414
rect 178167 525344 178201 525378
rect 178907 525380 178941 525414
rect 179271 525344 179305 525378
rect 180011 525380 180045 525414
rect 180375 525344 180409 525378
rect 181115 525380 181149 525414
rect 181479 525344 181513 525378
rect 181963 525380 181997 525414
rect 182073 525380 182107 525414
rect 182181 525344 182215 525378
rect 182291 525344 182325 525378
rect 182955 525380 182989 525414
rect 183319 525344 183353 525378
rect 184059 525380 184093 525414
rect 184423 525344 184457 525378
rect 185163 525380 185197 525414
rect 185527 525344 185561 525378
rect 186267 525380 186301 525414
rect 186631 525344 186665 525378
rect 187271 525340 187305 525374
rect 187379 525380 187413 525414
rect 172275 524864 172309 524898
rect 172383 524904 172417 524938
rect 172835 524864 172869 524898
rect 173199 524900 173233 524934
rect 173939 524864 173973 524898
rect 174303 524900 174337 524934
rect 175227 524864 175261 524898
rect 175591 524900 175625 524934
rect 176331 524864 176365 524898
rect 176695 524900 176729 524934
rect 177435 524864 177469 524898
rect 177799 524900 177833 524934
rect 178539 524864 178573 524898
rect 178903 524900 178937 524934
rect 179387 524864 179421 524898
rect 179497 524864 179531 524898
rect 179605 524900 179639 524934
rect 179715 524900 179749 524934
rect 180379 524864 180413 524898
rect 180743 524900 180777 524934
rect 181483 524864 181517 524898
rect 181847 524900 181881 524934
rect 182587 524864 182621 524898
rect 182951 524900 182985 524934
rect 183691 524864 183725 524898
rect 184055 524900 184089 524934
rect 184539 524864 184573 524898
rect 184649 524864 184683 524898
rect 184757 524900 184791 524934
rect 184867 524900 184901 524934
rect 185531 524864 185565 524898
rect 185895 524900 185929 524934
rect 186379 524864 186413 524898
rect 186478 524864 186512 524898
rect 186577 524864 186611 524898
rect 186685 524900 186719 524934
rect 186788 524900 186822 524934
rect 186891 524900 186925 524934
rect 187271 524904 187305 524938
rect 187379 524864 187413 524898
rect 172275 524292 172309 524326
rect 172383 524252 172417 524286
rect 172835 524292 172869 524326
rect 173199 524256 173233 524290
rect 173939 524292 173973 524326
rect 174303 524256 174337 524290
rect 175043 524292 175077 524326
rect 175407 524256 175441 524290
rect 176147 524292 176181 524326
rect 176511 524256 176545 524290
rect 176937 524292 176971 524326
rect 177197 524256 177231 524290
rect 177803 524292 177837 524326
rect 178167 524256 178201 524290
rect 178907 524292 178941 524326
rect 179271 524256 179305 524290
rect 180011 524292 180045 524326
rect 180375 524256 180409 524290
rect 181115 524292 181149 524326
rect 181479 524256 181513 524290
rect 181963 524292 181997 524326
rect 182073 524292 182107 524326
rect 182181 524256 182215 524290
rect 182291 524256 182325 524290
rect 182955 524292 182989 524326
rect 183319 524256 183353 524290
rect 184059 524292 184093 524326
rect 184423 524256 184457 524290
rect 185163 524292 185197 524326
rect 185527 524256 185561 524290
rect 186267 524292 186301 524326
rect 186631 524256 186665 524290
rect 187271 524252 187305 524286
rect 187379 524292 187413 524326
rect 172275 523776 172309 523810
rect 172383 523816 172417 523850
rect 172835 523776 172869 523810
rect 173199 523812 173233 523846
rect 173939 523776 173973 523810
rect 174303 523812 174337 523846
rect 175227 523776 175261 523810
rect 175591 523812 175625 523846
rect 176331 523776 176365 523810
rect 176695 523812 176729 523846
rect 177435 523776 177469 523810
rect 177799 523812 177833 523846
rect 178539 523776 178573 523810
rect 178903 523812 178937 523846
rect 179387 523776 179421 523810
rect 179497 523776 179531 523810
rect 179605 523812 179639 523846
rect 179715 523812 179749 523846
rect 180379 523776 180413 523810
rect 180743 523812 180777 523846
rect 181483 523776 181517 523810
rect 181847 523812 181881 523846
rect 182587 523776 182621 523810
rect 182951 523812 182985 523846
rect 183691 523776 183725 523810
rect 184055 523812 184089 523846
rect 184539 523776 184573 523810
rect 184649 523776 184683 523810
rect 184757 523812 184791 523846
rect 184867 523812 184901 523846
rect 185531 523776 185565 523810
rect 185895 523812 185929 523846
rect 186379 523776 186413 523810
rect 186478 523776 186512 523810
rect 186577 523776 186611 523810
rect 186685 523812 186719 523846
rect 186788 523812 186822 523846
rect 186891 523812 186925 523846
rect 187271 523816 187305 523850
rect 187379 523776 187413 523810
rect 172275 523204 172309 523238
rect 172383 523164 172417 523198
rect 172835 523204 172869 523238
rect 173199 523168 173233 523202
rect 173939 523204 173973 523238
rect 174303 523168 174337 523202
rect 175043 523204 175077 523238
rect 175407 523168 175441 523202
rect 176147 523204 176181 523238
rect 176511 523168 176545 523202
rect 176937 523204 176971 523238
rect 177197 523168 177231 523202
rect 177803 523204 177837 523238
rect 178167 523168 178201 523202
rect 178907 523204 178941 523238
rect 179271 523168 179305 523202
rect 180011 523204 180045 523238
rect 180375 523168 180409 523202
rect 181115 523204 181149 523238
rect 181479 523168 181513 523202
rect 181963 523204 181997 523238
rect 182073 523204 182107 523238
rect 182181 523168 182215 523202
rect 182291 523168 182325 523202
rect 182955 523204 182989 523238
rect 183319 523168 183353 523202
rect 184059 523204 184093 523238
rect 184423 523168 184457 523202
rect 185163 523204 185197 523238
rect 185527 523168 185561 523202
rect 186267 523204 186301 523238
rect 186631 523168 186665 523202
rect 187271 523164 187305 523198
rect 187379 523204 187413 523238
rect 172275 522688 172309 522722
rect 172383 522728 172417 522762
rect 172835 522688 172869 522722
rect 173199 522724 173233 522758
rect 173939 522688 173973 522722
rect 174303 522724 174337 522758
rect 175227 522688 175261 522722
rect 175591 522724 175625 522758
rect 176331 522688 176365 522722
rect 176695 522724 176729 522758
rect 177435 522688 177469 522722
rect 177799 522724 177833 522758
rect 178539 522688 178573 522722
rect 178903 522724 178937 522758
rect 179387 522688 179421 522722
rect 179497 522688 179531 522722
rect 179605 522724 179639 522758
rect 179715 522724 179749 522758
rect 180379 522688 180413 522722
rect 180743 522724 180777 522758
rect 181483 522688 181517 522722
rect 181847 522724 181881 522758
rect 182587 522688 182621 522722
rect 182951 522724 182985 522758
rect 183691 522688 183725 522722
rect 184055 522724 184089 522758
rect 184539 522688 184573 522722
rect 184649 522688 184683 522722
rect 184757 522724 184791 522758
rect 184867 522724 184901 522758
rect 185531 522688 185565 522722
rect 185895 522724 185929 522758
rect 186379 522688 186413 522722
rect 186478 522688 186512 522722
rect 186577 522688 186611 522722
rect 186685 522724 186719 522758
rect 186788 522724 186822 522758
rect 186891 522724 186925 522758
rect 187271 522728 187305 522762
rect 187379 522688 187413 522722
rect 172275 522116 172309 522150
rect 172383 522076 172417 522110
rect 172835 522116 172869 522150
rect 173199 522080 173233 522114
rect 173939 522116 173973 522150
rect 174303 522080 174337 522114
rect 175043 522116 175077 522150
rect 175407 522080 175441 522114
rect 176147 522116 176181 522150
rect 176511 522080 176545 522114
rect 176937 522116 176971 522150
rect 177197 522080 177231 522114
rect 177803 522116 177837 522150
rect 178167 522080 178201 522114
rect 178907 522116 178941 522150
rect 179271 522080 179305 522114
rect 180011 522116 180045 522150
rect 180375 522080 180409 522114
rect 181115 522116 181149 522150
rect 181479 522080 181513 522114
rect 181963 522116 181997 522150
rect 182073 522116 182107 522150
rect 182181 522080 182215 522114
rect 182291 522080 182325 522114
rect 182955 522116 182989 522150
rect 183319 522080 183353 522114
rect 184059 522116 184093 522150
rect 184423 522080 184457 522114
rect 185163 522116 185197 522150
rect 185527 522080 185561 522114
rect 186267 522116 186301 522150
rect 186631 522080 186665 522114
rect 187271 522076 187305 522110
rect 187379 522116 187413 522150
rect 172275 521600 172309 521634
rect 172383 521640 172417 521674
rect 172835 521600 172869 521634
rect 173199 521636 173233 521670
rect 173939 521600 173973 521634
rect 174303 521636 174337 521670
rect 175227 521600 175261 521634
rect 175591 521636 175625 521670
rect 176331 521600 176365 521634
rect 176695 521636 176729 521670
rect 177435 521600 177469 521634
rect 177799 521636 177833 521670
rect 178539 521600 178573 521634
rect 178903 521636 178937 521670
rect 179387 521600 179421 521634
rect 179497 521600 179531 521634
rect 179605 521636 179639 521670
rect 179715 521636 179749 521670
rect 180379 521600 180413 521634
rect 180743 521636 180777 521670
rect 181483 521600 181517 521634
rect 181847 521636 181881 521670
rect 182587 521600 182621 521634
rect 182951 521636 182985 521670
rect 183691 521600 183725 521634
rect 184055 521636 184089 521670
rect 184539 521600 184573 521634
rect 184649 521600 184683 521634
rect 184757 521636 184791 521670
rect 184867 521636 184901 521670
rect 185531 521600 185565 521634
rect 185895 521636 185929 521670
rect 186379 521600 186413 521634
rect 186478 521600 186512 521634
rect 186577 521600 186611 521634
rect 186685 521636 186719 521670
rect 186788 521636 186822 521670
rect 186891 521636 186925 521670
rect 187271 521640 187305 521674
rect 187379 521600 187413 521634
rect 172275 521028 172309 521062
rect 172383 520988 172417 521022
rect 172835 521028 172869 521062
rect 173199 520992 173233 521026
rect 173939 521028 173973 521062
rect 174303 520992 174337 521026
rect 175043 521028 175077 521062
rect 175407 520992 175441 521026
rect 176147 521028 176181 521062
rect 176511 520992 176545 521026
rect 176937 521028 176971 521062
rect 177197 520992 177231 521026
rect 177803 521028 177837 521062
rect 178167 520992 178201 521026
rect 178907 521028 178941 521062
rect 179271 520992 179305 521026
rect 180011 521028 180045 521062
rect 180375 520992 180409 521026
rect 181115 521028 181149 521062
rect 181479 520992 181513 521026
rect 181963 521028 181997 521062
rect 182073 521028 182107 521062
rect 182181 520992 182215 521026
rect 182291 520992 182325 521026
rect 182955 521028 182989 521062
rect 183319 520992 183353 521026
rect 184059 521028 184093 521062
rect 184423 520992 184457 521026
rect 185163 521028 185197 521062
rect 185527 520992 185561 521026
rect 186267 521028 186301 521062
rect 186631 520992 186665 521026
rect 187271 520988 187305 521022
rect 187379 521028 187413 521062
rect 172275 520512 172309 520546
rect 172383 520552 172417 520586
rect 172835 520512 172869 520546
rect 173199 520548 173233 520582
rect 173939 520512 173973 520546
rect 174303 520548 174337 520582
rect 175227 520512 175261 520546
rect 175591 520548 175625 520582
rect 176331 520512 176365 520546
rect 176695 520548 176729 520582
rect 177435 520512 177469 520546
rect 177799 520548 177833 520582
rect 178539 520512 178573 520546
rect 178903 520548 178937 520582
rect 179387 520512 179421 520546
rect 179497 520512 179531 520546
rect 179605 520548 179639 520582
rect 179715 520548 179749 520582
rect 180379 520512 180413 520546
rect 180743 520548 180777 520582
rect 181483 520512 181517 520546
rect 181847 520548 181881 520582
rect 182587 520512 182621 520546
rect 182951 520548 182985 520582
rect 183691 520512 183725 520546
rect 184055 520548 184089 520582
rect 184539 520512 184573 520546
rect 184649 520512 184683 520546
rect 184757 520548 184791 520582
rect 184867 520548 184901 520582
rect 185531 520512 185565 520546
rect 185895 520548 185929 520582
rect 186379 520512 186413 520546
rect 186478 520512 186512 520546
rect 186577 520512 186611 520546
rect 186685 520548 186719 520582
rect 186788 520548 186822 520582
rect 186891 520548 186925 520582
rect 187271 520552 187305 520586
rect 187379 520512 187413 520546
rect 172275 519940 172309 519974
rect 172383 519900 172417 519934
rect 172835 519940 172869 519974
rect 173199 519904 173233 519938
rect 173939 519940 173973 519974
rect 174303 519904 174337 519938
rect 175043 519940 175077 519974
rect 175407 519904 175441 519938
rect 176147 519940 176181 519974
rect 176511 519904 176545 519938
rect 176937 519940 176971 519974
rect 177197 519904 177231 519938
rect 177803 519940 177837 519974
rect 178167 519904 178201 519938
rect 178907 519940 178941 519974
rect 179271 519904 179305 519938
rect 180011 519940 180045 519974
rect 180375 519904 180409 519938
rect 181115 519940 181149 519974
rect 181479 519904 181513 519938
rect 181963 519940 181997 519974
rect 182073 519940 182107 519974
rect 182181 519904 182215 519938
rect 182291 519904 182325 519938
rect 182955 519940 182989 519974
rect 183319 519904 183353 519938
rect 184059 519940 184093 519974
rect 184423 519904 184457 519938
rect 185163 519940 185197 519974
rect 185527 519904 185561 519938
rect 186267 519940 186301 519974
rect 186631 519904 186665 519938
rect 187271 519900 187305 519934
rect 187379 519940 187413 519974
rect 172275 519424 172309 519458
rect 172383 519464 172417 519498
rect 172835 519424 172869 519458
rect 173199 519460 173233 519494
rect 173939 519424 173973 519458
rect 174303 519460 174337 519494
rect 175227 519424 175261 519458
rect 175591 519460 175625 519494
rect 176331 519424 176365 519458
rect 176695 519460 176729 519494
rect 177435 519424 177469 519458
rect 177799 519460 177833 519494
rect 178539 519424 178573 519458
rect 178903 519460 178937 519494
rect 179387 519424 179421 519458
rect 179497 519424 179531 519458
rect 179605 519460 179639 519494
rect 179715 519460 179749 519494
rect 180379 519424 180413 519458
rect 180743 519460 180777 519494
rect 181483 519424 181517 519458
rect 181847 519460 181881 519494
rect 182587 519424 182621 519458
rect 182951 519460 182985 519494
rect 183691 519424 183725 519458
rect 184055 519460 184089 519494
rect 184539 519424 184573 519458
rect 184649 519424 184683 519458
rect 184757 519460 184791 519494
rect 184867 519460 184901 519494
rect 185531 519424 185565 519458
rect 185895 519460 185929 519494
rect 186379 519424 186413 519458
rect 186478 519424 186512 519458
rect 186577 519424 186611 519458
rect 186685 519460 186719 519494
rect 186788 519460 186822 519494
rect 186891 519460 186925 519494
rect 187271 519464 187305 519498
rect 187379 519424 187413 519458
rect 172275 518852 172309 518886
rect 172383 518812 172417 518846
rect 172835 518852 172869 518886
rect 173199 518816 173233 518850
rect 173939 518852 173973 518886
rect 174303 518816 174337 518850
rect 175043 518852 175077 518886
rect 175407 518816 175441 518850
rect 176147 518852 176181 518886
rect 176511 518816 176545 518850
rect 176937 518852 176971 518886
rect 177197 518816 177231 518850
rect 177803 518852 177837 518886
rect 178167 518816 178201 518850
rect 178907 518852 178941 518886
rect 179271 518816 179305 518850
rect 180011 518852 180045 518886
rect 180375 518816 180409 518850
rect 181115 518852 181149 518886
rect 181479 518816 181513 518850
rect 181963 518852 181997 518886
rect 182073 518852 182107 518886
rect 182181 518816 182215 518850
rect 182291 518816 182325 518850
rect 182955 518852 182989 518886
rect 183319 518816 183353 518850
rect 184059 518852 184093 518886
rect 184423 518816 184457 518850
rect 185163 518852 185197 518886
rect 185527 518816 185561 518850
rect 186267 518852 186301 518886
rect 186631 518816 186665 518850
rect 187271 518812 187305 518846
rect 187379 518852 187413 518886
rect 172275 518336 172309 518370
rect 172383 518376 172417 518410
rect 172835 518336 172869 518370
rect 173199 518372 173233 518406
rect 173939 518336 173973 518370
rect 174303 518372 174337 518406
rect 175227 518336 175261 518370
rect 175591 518372 175625 518406
rect 176331 518336 176365 518370
rect 176695 518372 176729 518406
rect 177435 518336 177469 518370
rect 177799 518372 177833 518406
rect 178539 518336 178573 518370
rect 178903 518372 178937 518406
rect 179387 518336 179421 518370
rect 179497 518336 179531 518370
rect 179605 518372 179639 518406
rect 179715 518372 179749 518406
rect 180379 518336 180413 518370
rect 180743 518372 180777 518406
rect 181483 518336 181517 518370
rect 181847 518372 181881 518406
rect 182587 518336 182621 518370
rect 182951 518372 182985 518406
rect 183691 518336 183725 518370
rect 184055 518372 184089 518406
rect 184539 518336 184573 518370
rect 184649 518336 184683 518370
rect 184757 518372 184791 518406
rect 184867 518372 184901 518406
rect 185531 518336 185565 518370
rect 185895 518372 185929 518406
rect 186379 518336 186413 518370
rect 186478 518336 186512 518370
rect 186577 518336 186611 518370
rect 186685 518372 186719 518406
rect 186788 518372 186822 518406
rect 186891 518372 186925 518406
rect 187271 518376 187305 518410
rect 187379 518336 187413 518370
rect 172275 517764 172309 517798
rect 172383 517724 172417 517758
rect 172835 517764 172869 517798
rect 173199 517728 173233 517762
rect 173939 517764 173973 517798
rect 174303 517728 174337 517762
rect 175043 517764 175077 517798
rect 175407 517728 175441 517762
rect 176147 517764 176181 517798
rect 176511 517728 176545 517762
rect 176937 517764 176971 517798
rect 177197 517728 177231 517762
rect 177803 517764 177837 517798
rect 178167 517728 178201 517762
rect 178907 517764 178941 517798
rect 179271 517728 179305 517762
rect 180011 517764 180045 517798
rect 180375 517728 180409 517762
rect 181115 517764 181149 517798
rect 181479 517728 181513 517762
rect 181963 517764 181997 517798
rect 182073 517764 182107 517798
rect 182181 517728 182215 517762
rect 182291 517728 182325 517762
rect 182955 517764 182989 517798
rect 183319 517728 183353 517762
rect 184059 517764 184093 517798
rect 184423 517728 184457 517762
rect 185163 517764 185197 517798
rect 185527 517728 185561 517762
rect 186267 517764 186301 517798
rect 186631 517728 186665 517762
rect 187271 517724 187305 517758
rect 187379 517764 187413 517798
rect 172275 517248 172309 517282
rect 172383 517288 172417 517322
rect 172835 517248 172869 517282
rect 173199 517284 173233 517318
rect 173939 517248 173973 517282
rect 174303 517284 174337 517318
rect 175227 517248 175261 517282
rect 175591 517284 175625 517318
rect 176331 517248 176365 517282
rect 176695 517284 176729 517318
rect 177435 517248 177469 517282
rect 177799 517284 177833 517318
rect 178539 517248 178573 517282
rect 178903 517284 178937 517318
rect 179387 517248 179421 517282
rect 179497 517248 179531 517282
rect 179605 517284 179639 517318
rect 179715 517284 179749 517318
rect 180379 517248 180413 517282
rect 180743 517284 180777 517318
rect 181483 517248 181517 517282
rect 181847 517284 181881 517318
rect 182587 517248 182621 517282
rect 182951 517284 182985 517318
rect 183691 517248 183725 517282
rect 184055 517284 184089 517318
rect 184539 517248 184573 517282
rect 184649 517248 184683 517282
rect 184757 517284 184791 517318
rect 184867 517284 184901 517318
rect 185531 517248 185565 517282
rect 185895 517284 185929 517318
rect 186379 517248 186413 517282
rect 186478 517248 186512 517282
rect 186577 517248 186611 517282
rect 186685 517284 186719 517318
rect 186788 517284 186822 517318
rect 186891 517284 186925 517318
rect 187271 517288 187305 517322
rect 187379 517248 187413 517282
rect 172275 516676 172309 516710
rect 172383 516636 172417 516670
rect 172835 516676 172869 516710
rect 173199 516640 173233 516674
rect 173939 516676 173973 516710
rect 174303 516640 174337 516674
rect 175043 516676 175077 516710
rect 175407 516640 175441 516674
rect 176147 516676 176181 516710
rect 176511 516640 176545 516674
rect 176937 516676 176971 516710
rect 177197 516640 177231 516674
rect 177803 516676 177837 516710
rect 178167 516640 178201 516674
rect 178907 516676 178941 516710
rect 179271 516640 179305 516674
rect 180011 516676 180045 516710
rect 180375 516640 180409 516674
rect 181115 516676 181149 516710
rect 181479 516640 181513 516674
rect 181963 516676 181997 516710
rect 182073 516676 182107 516710
rect 182181 516640 182215 516674
rect 182291 516640 182325 516674
rect 182955 516676 182989 516710
rect 183319 516640 183353 516674
rect 184059 516676 184093 516710
rect 184423 516640 184457 516674
rect 185163 516676 185197 516710
rect 185527 516640 185561 516674
rect 186267 516676 186301 516710
rect 186631 516640 186665 516674
rect 187271 516636 187305 516670
rect 187379 516676 187413 516710
rect 172275 516160 172309 516194
rect 172383 516200 172417 516234
rect 172835 516160 172869 516194
rect 173199 516196 173233 516230
rect 173939 516160 173973 516194
rect 174303 516196 174337 516230
rect 175227 516160 175261 516194
rect 175591 516196 175625 516230
rect 176331 516160 176365 516194
rect 176695 516196 176729 516230
rect 177435 516160 177469 516194
rect 177799 516196 177833 516230
rect 178539 516160 178573 516194
rect 178903 516196 178937 516230
rect 179387 516160 179421 516194
rect 179497 516160 179531 516194
rect 179605 516196 179639 516230
rect 179715 516196 179749 516230
rect 180379 516160 180413 516194
rect 180743 516196 180777 516230
rect 181483 516160 181517 516194
rect 181847 516196 181881 516230
rect 182587 516160 182621 516194
rect 182951 516196 182985 516230
rect 183691 516160 183725 516194
rect 184055 516196 184089 516230
rect 184539 516160 184573 516194
rect 184649 516160 184683 516194
rect 184757 516196 184791 516230
rect 184867 516196 184901 516230
rect 185531 516160 185565 516194
rect 185895 516196 185929 516230
rect 186379 516160 186413 516194
rect 186478 516160 186512 516194
rect 186577 516160 186611 516194
rect 186685 516196 186719 516230
rect 186788 516196 186822 516230
rect 186891 516196 186925 516230
rect 187271 516200 187305 516234
rect 187379 516160 187413 516194
rect 172275 515588 172309 515622
rect 172383 515548 172417 515582
rect 172579 515588 172613 515622
rect 172678 515588 172712 515622
rect 172777 515588 172811 515622
rect 172885 515552 172919 515586
rect 172988 515552 173022 515586
rect 173091 515552 173125 515586
rect 173489 515562 173523 515596
rect 173635 515562 173669 515596
rect 173703 515562 173737 515596
rect 173771 515562 173805 515596
rect 174051 515588 174085 515622
rect 174150 515588 174184 515622
rect 174249 515588 174283 515622
rect 174357 515552 174391 515586
rect 174460 515552 174494 515586
rect 174563 515552 174597 515586
rect 175227 515588 175261 515622
rect 175591 515552 175625 515586
rect 176331 515588 176365 515622
rect 176695 515552 176729 515586
rect 177151 515588 177185 515622
rect 177259 515548 177293 515582
rect 177803 515588 177837 515622
rect 178167 515552 178201 515586
rect 178907 515588 178941 515622
rect 179271 515552 179305 515586
rect 179727 515588 179761 515622
rect 179835 515548 179869 515582
rect 180379 515588 180413 515622
rect 180743 515552 180777 515586
rect 181227 515588 181261 515622
rect 181326 515588 181360 515622
rect 181425 515588 181459 515622
rect 181533 515552 181567 515586
rect 181636 515552 181670 515586
rect 181739 515552 181773 515586
rect 182139 515575 182173 515609
rect 182257 515562 182291 515596
rect 182955 515588 182989 515622
rect 183319 515552 183353 515586
rect 184059 515588 184093 515622
rect 184423 515552 184457 515586
rect 184879 515588 184913 515622
rect 184987 515548 185021 515582
rect 185531 515588 185565 515622
rect 185895 515552 185929 515586
rect 186461 515562 186495 515596
rect 186607 515562 186641 515596
rect 186675 515562 186709 515596
rect 186743 515562 186777 515596
rect 186995 515588 187029 515622
rect 187103 515548 187137 515582
rect 187271 515548 187305 515582
rect 187379 515588 187413 515622
<< xpolycontact >>
rect 164316 537517 164386 537949
rect 164316 536001 164386 536433
rect 164634 537517 164704 537949
rect 164634 536001 164704 536433
rect 164952 537517 165022 537949
rect 164952 536001 165022 536433
rect 165270 537517 165340 537949
rect 165270 536001 165340 536433
rect 165588 537517 165658 537949
rect 165588 536001 165658 536433
rect 165906 537517 165976 537949
rect 165906 536001 165976 536433
rect 166224 537517 166294 537949
rect 166224 536001 166294 536433
rect 166542 537517 166612 537949
rect 166542 536001 166612 536433
rect 168088 537517 168158 537949
rect 168088 536001 168158 536433
rect 168406 537517 168476 537949
rect 168406 536001 168476 536433
rect 168724 537517 168794 537949
rect 168724 536001 168794 536433
rect 169042 537517 169112 537949
rect 169042 536001 169112 536433
rect 171824 537517 171894 537949
rect 171824 536001 171894 536433
rect 172142 537517 172212 537949
rect 172142 536001 172212 536433
rect 175342 537517 175412 537949
rect 175342 536001 175412 536433
rect 178942 537517 179012 537949
rect 178942 536561 179012 536993
rect 182242 537517 182312 537949
rect 182242 536841 182312 537273
rect 185542 537517 185612 537949
rect 185542 536981 185612 537413
rect 188842 537517 188912 537949
rect 188842 536885 188912 537317
rect 164286 535177 164356 535609
rect 164286 533661 164356 534093
rect 164604 535177 164674 535609
rect 164604 533661 164674 534093
rect 164922 535177 164992 535609
rect 164922 533661 164992 534093
rect 165240 535177 165310 535609
rect 165240 533661 165310 534093
rect 165558 535177 165628 535609
rect 165558 533661 165628 534093
rect 165876 535177 165946 535609
rect 165876 533661 165946 534093
rect 166194 535177 166264 535609
rect 166194 533661 166264 534093
rect 166512 535177 166582 535609
rect 166512 533661 166582 534093
<< ppolyres >>
rect 188842 537317 188912 537517
<< xpolyres >>
rect 164316 536433 164386 537517
rect 164634 536433 164704 537517
rect 164952 536433 165022 537517
rect 165270 536433 165340 537517
rect 165588 536433 165658 537517
rect 165906 536433 165976 537517
rect 166224 536433 166294 537517
rect 166542 536433 166612 537517
rect 168088 536433 168158 537517
rect 168406 536433 168476 537517
rect 168724 536433 168794 537517
rect 169042 536433 169112 537517
rect 171824 536433 171894 537517
rect 172142 536433 172212 537517
rect 175342 536433 175412 537517
rect 178942 536993 179012 537517
rect 182242 537273 182312 537517
rect 185542 537413 185612 537517
rect 164286 534093 164356 535177
rect 164604 534093 164674 535177
rect 164922 534093 164992 535177
rect 165240 534093 165310 535177
rect 165558 534093 165628 535177
rect 165876 534093 165946 535177
rect 166194 534093 166264 535177
rect 166512 534093 166582 535177
<< rmp >>
rect 186949 530338 187045 530347
rect 187087 530338 187183 530347
<< locali >>
rect 164518 541255 166648 541275
rect 164518 541245 164618 541255
rect 164518 539865 164538 541245
rect 164578 541215 164618 541245
rect 166538 541235 166648 541255
rect 166538 541215 166578 541235
rect 164578 541185 166578 541215
rect 164578 539915 164598 541185
rect 164712 541085 164728 541119
rect 164762 541085 164778 541119
rect 165015 541092 165031 541126
rect 165065 541092 165081 541126
rect 165207 541092 165223 541126
rect 165257 541092 165273 541126
rect 165399 541092 165415 541126
rect 165449 541092 165465 541126
rect 165591 541092 165607 541126
rect 165641 541092 165657 541126
rect 165783 541092 165799 541126
rect 165833 541092 165849 541126
rect 165975 541092 165991 541126
rect 166025 541092 166041 541126
rect 166392 541085 166408 541119
rect 166442 541085 166458 541119
rect 164684 541035 164718 541051
rect 164684 540043 164718 540059
rect 164772 541035 164806 541051
rect 164772 540043 164806 540059
rect 164887 541042 164921 541058
rect 164887 540050 164921 540066
rect 164983 541042 165017 541058
rect 164983 540050 165017 540066
rect 165079 541042 165113 541058
rect 165079 540050 165113 540066
rect 165175 541042 165209 541058
rect 165175 540050 165209 540066
rect 165271 541042 165305 541058
rect 165271 540050 165305 540066
rect 165367 541042 165401 541058
rect 165367 540050 165401 540066
rect 165463 541042 165497 541058
rect 165463 540050 165497 540066
rect 165559 541042 165593 541058
rect 165559 540050 165593 540066
rect 165655 541042 165689 541058
rect 165655 540050 165689 540066
rect 165751 541042 165785 541058
rect 165751 540050 165785 540066
rect 165847 541042 165881 541058
rect 165847 540050 165881 540066
rect 165943 541042 165977 541058
rect 165943 540050 165977 540066
rect 166039 541042 166073 541058
rect 166364 541035 166398 541051
rect 166192 540285 166208 540319
rect 166242 540285 166258 540319
rect 166039 540050 166073 540066
rect 166164 540235 166198 540251
rect 166164 540043 166198 540059
rect 166252 540235 166286 540251
rect 166252 540043 166286 540059
rect 166364 540043 166398 540059
rect 166452 541035 166486 541051
rect 166452 540043 166486 540059
rect 166558 540215 166578 541185
rect 166618 540215 166648 541235
rect 166558 540085 166568 540215
rect 166628 540085 166648 540215
rect 164712 539975 164728 540009
rect 164762 539975 164778 540009
rect 164919 539982 164935 540016
rect 164969 539982 164985 540016
rect 165111 539982 165127 540016
rect 165161 539982 165177 540016
rect 165303 539982 165319 540016
rect 165353 539982 165369 540016
rect 165495 539982 165511 540016
rect 165545 539982 165561 540016
rect 165687 539982 165703 540016
rect 165737 539982 165753 540016
rect 165879 539982 165895 540016
rect 165929 539982 165945 540016
rect 166192 539975 166208 540009
rect 166242 539975 166258 540009
rect 166392 539975 166408 540009
rect 166442 539975 166458 540009
rect 166558 539915 166578 540085
rect 164578 539895 166578 539915
rect 164578 539865 164618 539895
rect 164518 539855 164618 539865
rect 166538 539855 166578 539895
rect 166618 539855 166648 540085
rect 164518 539825 166648 539855
rect 168318 541255 170448 541275
rect 168318 541245 168418 541255
rect 168318 539865 168338 541245
rect 168378 541215 168418 541245
rect 170338 541235 170448 541255
rect 170338 541215 170378 541235
rect 168378 541185 170378 541215
rect 168378 539915 168398 541185
rect 168512 541085 168528 541119
rect 168562 541085 168578 541119
rect 168815 541092 168831 541126
rect 168865 541092 168881 541126
rect 169007 541092 169023 541126
rect 169057 541092 169073 541126
rect 169199 541092 169215 541126
rect 169249 541092 169265 541126
rect 169391 541092 169407 541126
rect 169441 541092 169457 541126
rect 169583 541092 169599 541126
rect 169633 541092 169649 541126
rect 169775 541092 169791 541126
rect 169825 541092 169841 541126
rect 170192 541085 170208 541119
rect 170242 541085 170258 541119
rect 168484 541035 168518 541051
rect 168484 540043 168518 540059
rect 168572 541035 168606 541051
rect 168572 540043 168606 540059
rect 168687 541042 168721 541058
rect 168687 540050 168721 540066
rect 168783 541042 168817 541058
rect 168783 540050 168817 540066
rect 168879 541042 168913 541058
rect 168879 540050 168913 540066
rect 168975 541042 169009 541058
rect 168975 540050 169009 540066
rect 169071 541042 169105 541058
rect 169071 540050 169105 540066
rect 169167 541042 169201 541058
rect 169167 540050 169201 540066
rect 169263 541042 169297 541058
rect 169263 540050 169297 540066
rect 169359 541042 169393 541058
rect 169359 540050 169393 540066
rect 169455 541042 169489 541058
rect 169455 540050 169489 540066
rect 169551 541042 169585 541058
rect 169551 540050 169585 540066
rect 169647 541042 169681 541058
rect 169647 540050 169681 540066
rect 169743 541042 169777 541058
rect 169743 540050 169777 540066
rect 169839 541042 169873 541058
rect 170164 541035 170198 541051
rect 169992 540285 170008 540319
rect 170042 540285 170058 540319
rect 169839 540050 169873 540066
rect 169964 540235 169998 540251
rect 169964 540043 169998 540059
rect 170052 540235 170086 540251
rect 170052 540043 170086 540059
rect 170164 540043 170198 540059
rect 170252 541035 170286 541051
rect 170252 540043 170286 540059
rect 170358 540215 170378 541185
rect 170418 540215 170448 541235
rect 170358 540085 170368 540215
rect 170428 540085 170448 540215
rect 168512 539975 168528 540009
rect 168562 539975 168578 540009
rect 168719 539982 168735 540016
rect 168769 539982 168785 540016
rect 168911 539982 168927 540016
rect 168961 539982 168977 540016
rect 169103 539982 169119 540016
rect 169153 539982 169169 540016
rect 169295 539982 169311 540016
rect 169345 539982 169361 540016
rect 169487 539982 169503 540016
rect 169537 539982 169553 540016
rect 169679 539982 169695 540016
rect 169729 539982 169745 540016
rect 169992 539975 170008 540009
rect 170042 539975 170058 540009
rect 170192 539975 170208 540009
rect 170242 539975 170258 540009
rect 170358 539915 170378 540085
rect 168378 539895 170378 539915
rect 168378 539865 168418 539895
rect 168318 539855 168418 539865
rect 170338 539855 170378 539895
rect 170418 539855 170448 540085
rect 168318 539825 170448 539855
rect 172018 541255 174148 541275
rect 172018 541245 172118 541255
rect 172018 539865 172038 541245
rect 172078 541215 172118 541245
rect 174038 541235 174148 541255
rect 174038 541215 174078 541235
rect 172078 541185 174078 541215
rect 172078 539915 172098 541185
rect 172212 541085 172228 541119
rect 172262 541085 172278 541119
rect 172515 541092 172531 541126
rect 172565 541092 172581 541126
rect 172707 541092 172723 541126
rect 172757 541092 172773 541126
rect 172899 541092 172915 541126
rect 172949 541092 172965 541126
rect 173091 541092 173107 541126
rect 173141 541092 173157 541126
rect 173283 541092 173299 541126
rect 173333 541092 173349 541126
rect 173475 541092 173491 541126
rect 173525 541092 173541 541126
rect 173892 541085 173908 541119
rect 173942 541085 173958 541119
rect 172184 541035 172218 541051
rect 172184 540043 172218 540059
rect 172272 541035 172306 541051
rect 172272 540043 172306 540059
rect 172387 541042 172421 541058
rect 172387 540050 172421 540066
rect 172483 541042 172517 541058
rect 172483 540050 172517 540066
rect 172579 541042 172613 541058
rect 172579 540050 172613 540066
rect 172675 541042 172709 541058
rect 172675 540050 172709 540066
rect 172771 541042 172805 541058
rect 172771 540050 172805 540066
rect 172867 541042 172901 541058
rect 172867 540050 172901 540066
rect 172963 541042 172997 541058
rect 172963 540050 172997 540066
rect 173059 541042 173093 541058
rect 173059 540050 173093 540066
rect 173155 541042 173189 541058
rect 173155 540050 173189 540066
rect 173251 541042 173285 541058
rect 173251 540050 173285 540066
rect 173347 541042 173381 541058
rect 173347 540050 173381 540066
rect 173443 541042 173477 541058
rect 173443 540050 173477 540066
rect 173539 541042 173573 541058
rect 173864 541035 173898 541051
rect 173692 540285 173708 540319
rect 173742 540285 173758 540319
rect 173539 540050 173573 540066
rect 173664 540235 173698 540251
rect 173664 540043 173698 540059
rect 173752 540235 173786 540251
rect 173752 540043 173786 540059
rect 173864 540043 173898 540059
rect 173952 541035 173986 541051
rect 173952 540043 173986 540059
rect 174058 540215 174078 541185
rect 174118 540215 174148 541235
rect 174058 540085 174068 540215
rect 174128 540085 174148 540215
rect 172212 539975 172228 540009
rect 172262 539975 172278 540009
rect 172419 539982 172435 540016
rect 172469 539982 172485 540016
rect 172611 539982 172627 540016
rect 172661 539982 172677 540016
rect 172803 539982 172819 540016
rect 172853 539982 172869 540016
rect 172995 539982 173011 540016
rect 173045 539982 173061 540016
rect 173187 539982 173203 540016
rect 173237 539982 173253 540016
rect 173379 539982 173395 540016
rect 173429 539982 173445 540016
rect 173692 539975 173708 540009
rect 173742 539975 173758 540009
rect 173892 539975 173908 540009
rect 173942 539975 173958 540009
rect 174058 539915 174078 540085
rect 172078 539895 174078 539915
rect 172078 539865 172118 539895
rect 172018 539855 172118 539865
rect 174038 539855 174078 539895
rect 174118 539855 174148 540085
rect 172018 539825 174148 539855
rect 175518 541255 177648 541275
rect 175518 541245 175618 541255
rect 175518 539865 175538 541245
rect 175578 541215 175618 541245
rect 177538 541235 177648 541255
rect 177538 541215 177578 541235
rect 175578 541185 177578 541215
rect 175578 539915 175598 541185
rect 175712 541085 175728 541119
rect 175762 541085 175778 541119
rect 176015 541092 176031 541126
rect 176065 541092 176081 541126
rect 176207 541092 176223 541126
rect 176257 541092 176273 541126
rect 176399 541092 176415 541126
rect 176449 541092 176465 541126
rect 176591 541092 176607 541126
rect 176641 541092 176657 541126
rect 176783 541092 176799 541126
rect 176833 541092 176849 541126
rect 176975 541092 176991 541126
rect 177025 541092 177041 541126
rect 177392 541085 177408 541119
rect 177442 541085 177458 541119
rect 175684 541035 175718 541051
rect 175684 540043 175718 540059
rect 175772 541035 175806 541051
rect 175772 540043 175806 540059
rect 175887 541042 175921 541058
rect 175887 540050 175921 540066
rect 175983 541042 176017 541058
rect 175983 540050 176017 540066
rect 176079 541042 176113 541058
rect 176079 540050 176113 540066
rect 176175 541042 176209 541058
rect 176175 540050 176209 540066
rect 176271 541042 176305 541058
rect 176271 540050 176305 540066
rect 176367 541042 176401 541058
rect 176367 540050 176401 540066
rect 176463 541042 176497 541058
rect 176463 540050 176497 540066
rect 176559 541042 176593 541058
rect 176559 540050 176593 540066
rect 176655 541042 176689 541058
rect 176655 540050 176689 540066
rect 176751 541042 176785 541058
rect 176751 540050 176785 540066
rect 176847 541042 176881 541058
rect 176847 540050 176881 540066
rect 176943 541042 176977 541058
rect 176943 540050 176977 540066
rect 177039 541042 177073 541058
rect 177364 541035 177398 541051
rect 177192 540285 177208 540319
rect 177242 540285 177258 540319
rect 177039 540050 177073 540066
rect 177164 540235 177198 540251
rect 177164 540043 177198 540059
rect 177252 540235 177286 540251
rect 177252 540043 177286 540059
rect 177364 540043 177398 540059
rect 177452 541035 177486 541051
rect 177452 540043 177486 540059
rect 177558 540215 177578 541185
rect 177618 540215 177648 541235
rect 177558 540085 177568 540215
rect 177628 540085 177648 540215
rect 175712 539975 175728 540009
rect 175762 539975 175778 540009
rect 175919 539982 175935 540016
rect 175969 539982 175985 540016
rect 176111 539982 176127 540016
rect 176161 539982 176177 540016
rect 176303 539982 176319 540016
rect 176353 539982 176369 540016
rect 176495 539982 176511 540016
rect 176545 539982 176561 540016
rect 176687 539982 176703 540016
rect 176737 539982 176753 540016
rect 176879 539982 176895 540016
rect 176929 539982 176945 540016
rect 177192 539975 177208 540009
rect 177242 539975 177258 540009
rect 177392 539975 177408 540009
rect 177442 539975 177458 540009
rect 177558 539915 177578 540085
rect 175578 539895 177578 539915
rect 175578 539865 175618 539895
rect 175518 539855 175618 539865
rect 177538 539855 177578 539895
rect 177618 539855 177648 540085
rect 175518 539825 177648 539855
rect 179118 541255 181248 541275
rect 179118 541245 179218 541255
rect 179118 539865 179138 541245
rect 179178 541215 179218 541245
rect 181138 541235 181248 541255
rect 181138 541215 181178 541235
rect 179178 541185 181178 541215
rect 179178 539915 179198 541185
rect 179312 541085 179328 541119
rect 179362 541085 179378 541119
rect 179615 541092 179631 541126
rect 179665 541092 179681 541126
rect 179807 541092 179823 541126
rect 179857 541092 179873 541126
rect 179999 541092 180015 541126
rect 180049 541092 180065 541126
rect 180191 541092 180207 541126
rect 180241 541092 180257 541126
rect 180383 541092 180399 541126
rect 180433 541092 180449 541126
rect 180575 541092 180591 541126
rect 180625 541092 180641 541126
rect 180992 541085 181008 541119
rect 181042 541085 181058 541119
rect 179284 541035 179318 541051
rect 179284 540043 179318 540059
rect 179372 541035 179406 541051
rect 179372 540043 179406 540059
rect 179487 541042 179521 541058
rect 179487 540050 179521 540066
rect 179583 541042 179617 541058
rect 179583 540050 179617 540066
rect 179679 541042 179713 541058
rect 179679 540050 179713 540066
rect 179775 541042 179809 541058
rect 179775 540050 179809 540066
rect 179871 541042 179905 541058
rect 179871 540050 179905 540066
rect 179967 541042 180001 541058
rect 179967 540050 180001 540066
rect 180063 541042 180097 541058
rect 180063 540050 180097 540066
rect 180159 541042 180193 541058
rect 180159 540050 180193 540066
rect 180255 541042 180289 541058
rect 180255 540050 180289 540066
rect 180351 541042 180385 541058
rect 180351 540050 180385 540066
rect 180447 541042 180481 541058
rect 180447 540050 180481 540066
rect 180543 541042 180577 541058
rect 180543 540050 180577 540066
rect 180639 541042 180673 541058
rect 180964 541035 180998 541051
rect 180792 540285 180808 540319
rect 180842 540285 180858 540319
rect 180639 540050 180673 540066
rect 180764 540235 180798 540251
rect 180764 540043 180798 540059
rect 180852 540235 180886 540251
rect 180852 540043 180886 540059
rect 180964 540043 180998 540059
rect 181052 541035 181086 541051
rect 181052 540043 181086 540059
rect 181158 540215 181178 541185
rect 181218 540215 181248 541235
rect 181158 540085 181168 540215
rect 181228 540085 181248 540215
rect 179312 539975 179328 540009
rect 179362 539975 179378 540009
rect 179519 539982 179535 540016
rect 179569 539982 179585 540016
rect 179711 539982 179727 540016
rect 179761 539982 179777 540016
rect 179903 539982 179919 540016
rect 179953 539982 179969 540016
rect 180095 539982 180111 540016
rect 180145 539982 180161 540016
rect 180287 539982 180303 540016
rect 180337 539982 180353 540016
rect 180479 539982 180495 540016
rect 180529 539982 180545 540016
rect 180792 539975 180808 540009
rect 180842 539975 180858 540009
rect 180992 539975 181008 540009
rect 181042 539975 181058 540009
rect 181158 539915 181178 540085
rect 179178 539895 181178 539915
rect 179178 539865 179218 539895
rect 179118 539855 179218 539865
rect 181138 539855 181178 539895
rect 181218 539855 181248 540085
rect 179118 539825 181248 539855
rect 182418 541255 184548 541275
rect 182418 541245 182518 541255
rect 182418 539865 182438 541245
rect 182478 541215 182518 541245
rect 184438 541235 184548 541255
rect 184438 541215 184478 541235
rect 182478 541185 184478 541215
rect 182478 539915 182498 541185
rect 182612 541085 182628 541119
rect 182662 541085 182678 541119
rect 182915 541092 182931 541126
rect 182965 541092 182981 541126
rect 183107 541092 183123 541126
rect 183157 541092 183173 541126
rect 183299 541092 183315 541126
rect 183349 541092 183365 541126
rect 183491 541092 183507 541126
rect 183541 541092 183557 541126
rect 183683 541092 183699 541126
rect 183733 541092 183749 541126
rect 183875 541092 183891 541126
rect 183925 541092 183941 541126
rect 184292 541085 184308 541119
rect 184342 541085 184358 541119
rect 182584 541035 182618 541051
rect 182584 540043 182618 540059
rect 182672 541035 182706 541051
rect 182672 540043 182706 540059
rect 182787 541042 182821 541058
rect 182787 540050 182821 540066
rect 182883 541042 182917 541058
rect 182883 540050 182917 540066
rect 182979 541042 183013 541058
rect 182979 540050 183013 540066
rect 183075 541042 183109 541058
rect 183075 540050 183109 540066
rect 183171 541042 183205 541058
rect 183171 540050 183205 540066
rect 183267 541042 183301 541058
rect 183267 540050 183301 540066
rect 183363 541042 183397 541058
rect 183363 540050 183397 540066
rect 183459 541042 183493 541058
rect 183459 540050 183493 540066
rect 183555 541042 183589 541058
rect 183555 540050 183589 540066
rect 183651 541042 183685 541058
rect 183651 540050 183685 540066
rect 183747 541042 183781 541058
rect 183747 540050 183781 540066
rect 183843 541042 183877 541058
rect 183843 540050 183877 540066
rect 183939 541042 183973 541058
rect 184264 541035 184298 541051
rect 184092 540285 184108 540319
rect 184142 540285 184158 540319
rect 183939 540050 183973 540066
rect 184064 540235 184098 540251
rect 184064 540043 184098 540059
rect 184152 540235 184186 540251
rect 184152 540043 184186 540059
rect 184264 540043 184298 540059
rect 184352 541035 184386 541051
rect 184352 540043 184386 540059
rect 184458 540215 184478 541185
rect 184518 540215 184548 541235
rect 184458 540085 184468 540215
rect 184528 540085 184548 540215
rect 182612 539975 182628 540009
rect 182662 539975 182678 540009
rect 182819 539982 182835 540016
rect 182869 539982 182885 540016
rect 183011 539982 183027 540016
rect 183061 539982 183077 540016
rect 183203 539982 183219 540016
rect 183253 539982 183269 540016
rect 183395 539982 183411 540016
rect 183445 539982 183461 540016
rect 183587 539982 183603 540016
rect 183637 539982 183653 540016
rect 183779 539982 183795 540016
rect 183829 539982 183845 540016
rect 184092 539975 184108 540009
rect 184142 539975 184158 540009
rect 184292 539975 184308 540009
rect 184342 539975 184358 540009
rect 184458 539915 184478 540085
rect 182478 539895 184478 539915
rect 182478 539865 182518 539895
rect 182418 539855 182518 539865
rect 184438 539855 184478 539895
rect 184518 539855 184548 540085
rect 182418 539825 184548 539855
rect 185718 541255 187848 541275
rect 185718 541245 185818 541255
rect 185718 539865 185738 541245
rect 185778 541215 185818 541245
rect 187738 541235 187848 541255
rect 187738 541215 187778 541235
rect 185778 541185 187778 541215
rect 185778 539915 185798 541185
rect 185912 541085 185928 541119
rect 185962 541085 185978 541119
rect 186215 541092 186231 541126
rect 186265 541092 186281 541126
rect 186407 541092 186423 541126
rect 186457 541092 186473 541126
rect 186599 541092 186615 541126
rect 186649 541092 186665 541126
rect 186791 541092 186807 541126
rect 186841 541092 186857 541126
rect 186983 541092 186999 541126
rect 187033 541092 187049 541126
rect 187175 541092 187191 541126
rect 187225 541092 187241 541126
rect 187592 541085 187608 541119
rect 187642 541085 187658 541119
rect 185884 541035 185918 541051
rect 185884 540043 185918 540059
rect 185972 541035 186006 541051
rect 185972 540043 186006 540059
rect 186087 541042 186121 541058
rect 186087 540050 186121 540066
rect 186183 541042 186217 541058
rect 186183 540050 186217 540066
rect 186279 541042 186313 541058
rect 186279 540050 186313 540066
rect 186375 541042 186409 541058
rect 186375 540050 186409 540066
rect 186471 541042 186505 541058
rect 186471 540050 186505 540066
rect 186567 541042 186601 541058
rect 186567 540050 186601 540066
rect 186663 541042 186697 541058
rect 186663 540050 186697 540066
rect 186759 541042 186793 541058
rect 186759 540050 186793 540066
rect 186855 541042 186889 541058
rect 186855 540050 186889 540066
rect 186951 541042 186985 541058
rect 186951 540050 186985 540066
rect 187047 541042 187081 541058
rect 187047 540050 187081 540066
rect 187143 541042 187177 541058
rect 187143 540050 187177 540066
rect 187239 541042 187273 541058
rect 187564 541035 187598 541051
rect 187392 540285 187408 540319
rect 187442 540285 187458 540319
rect 187239 540050 187273 540066
rect 187364 540235 187398 540251
rect 187364 540043 187398 540059
rect 187452 540235 187486 540251
rect 187452 540043 187486 540059
rect 187564 540043 187598 540059
rect 187652 541035 187686 541051
rect 187652 540043 187686 540059
rect 187758 540215 187778 541185
rect 187818 540215 187848 541235
rect 187758 540085 187768 540215
rect 187828 540085 187848 540215
rect 185912 539975 185928 540009
rect 185962 539975 185978 540009
rect 186119 539982 186135 540016
rect 186169 539982 186185 540016
rect 186311 539982 186327 540016
rect 186361 539982 186377 540016
rect 186503 539982 186519 540016
rect 186553 539982 186569 540016
rect 186695 539982 186711 540016
rect 186745 539982 186761 540016
rect 186887 539982 186903 540016
rect 186937 539982 186953 540016
rect 187079 539982 187095 540016
rect 187129 539982 187145 540016
rect 187392 539975 187408 540009
rect 187442 539975 187458 540009
rect 187592 539975 187608 540009
rect 187642 539975 187658 540009
rect 187758 539915 187778 540085
rect 185778 539895 187778 539915
rect 185778 539865 185818 539895
rect 185718 539855 185818 539865
rect 187738 539855 187778 539895
rect 187818 539855 187848 540085
rect 185718 539825 187848 539855
rect 189018 541255 191148 541275
rect 189018 541245 189118 541255
rect 189018 539865 189038 541245
rect 189078 541215 189118 541245
rect 191038 541235 191148 541255
rect 191038 541215 191078 541235
rect 189078 541185 191078 541215
rect 189078 539915 189098 541185
rect 189212 541085 189228 541119
rect 189262 541085 189278 541119
rect 189515 541092 189531 541126
rect 189565 541092 189581 541126
rect 189707 541092 189723 541126
rect 189757 541092 189773 541126
rect 189899 541092 189915 541126
rect 189949 541092 189965 541126
rect 190091 541092 190107 541126
rect 190141 541092 190157 541126
rect 190283 541092 190299 541126
rect 190333 541092 190349 541126
rect 190475 541092 190491 541126
rect 190525 541092 190541 541126
rect 190892 541085 190908 541119
rect 190942 541085 190958 541119
rect 189184 541035 189218 541051
rect 189184 540043 189218 540059
rect 189272 541035 189306 541051
rect 189272 540043 189306 540059
rect 189387 541042 189421 541058
rect 189387 540050 189421 540066
rect 189483 541042 189517 541058
rect 189483 540050 189517 540066
rect 189579 541042 189613 541058
rect 189579 540050 189613 540066
rect 189675 541042 189709 541058
rect 189675 540050 189709 540066
rect 189771 541042 189805 541058
rect 189771 540050 189805 540066
rect 189867 541042 189901 541058
rect 189867 540050 189901 540066
rect 189963 541042 189997 541058
rect 189963 540050 189997 540066
rect 190059 541042 190093 541058
rect 190059 540050 190093 540066
rect 190155 541042 190189 541058
rect 190155 540050 190189 540066
rect 190251 541042 190285 541058
rect 190251 540050 190285 540066
rect 190347 541042 190381 541058
rect 190347 540050 190381 540066
rect 190443 541042 190477 541058
rect 190443 540050 190477 540066
rect 190539 541042 190573 541058
rect 190864 541035 190898 541051
rect 190692 540285 190708 540319
rect 190742 540285 190758 540319
rect 190539 540050 190573 540066
rect 190664 540235 190698 540251
rect 190664 540043 190698 540059
rect 190752 540235 190786 540251
rect 190752 540043 190786 540059
rect 190864 540043 190898 540059
rect 190952 541035 190986 541051
rect 190952 540043 190986 540059
rect 191058 540215 191078 541185
rect 191118 540215 191148 541235
rect 191058 540085 191068 540215
rect 191128 540085 191148 540215
rect 189212 539975 189228 540009
rect 189262 539975 189278 540009
rect 189419 539982 189435 540016
rect 189469 539982 189485 540016
rect 189611 539982 189627 540016
rect 189661 539982 189677 540016
rect 189803 539982 189819 540016
rect 189853 539982 189869 540016
rect 189995 539982 190011 540016
rect 190045 539982 190061 540016
rect 190187 539982 190203 540016
rect 190237 539982 190253 540016
rect 190379 539982 190395 540016
rect 190429 539982 190445 540016
rect 190692 539975 190708 540009
rect 190742 539975 190758 540009
rect 190892 539975 190908 540009
rect 190942 539975 190958 540009
rect 191058 539915 191078 540085
rect 189078 539895 191078 539915
rect 189078 539865 189118 539895
rect 189018 539855 189118 539865
rect 191038 539855 191078 539895
rect 191118 539855 191148 540085
rect 191808 540245 191988 540261
rect 191808 540049 191988 540065
rect 189018 539825 191148 539855
rect 164518 539735 166638 539755
rect 164518 539715 164618 539735
rect 157628 538705 162868 538725
rect 157628 538665 157708 538705
rect 162768 538665 162868 538705
rect 157628 538645 162868 538665
rect 157628 538625 157708 538645
rect 157628 537965 157648 538625
rect 157688 538005 157708 538625
rect 158710 538435 158726 538469
rect 158894 538435 158910 538469
rect 159086 538435 159102 538469
rect 159270 538435 159286 538469
rect 159344 538435 159360 538469
rect 159528 538435 159544 538469
rect 159602 538435 159618 538469
rect 159786 538435 159802 538469
rect 159860 538435 159876 538469
rect 160044 538435 160060 538469
rect 160118 538435 160134 538469
rect 160302 538435 160318 538469
rect 160376 538435 160392 538469
rect 160560 538435 160576 538469
rect 160634 538435 160650 538469
rect 160818 538435 160834 538469
rect 160892 538435 160908 538469
rect 161076 538435 161092 538469
rect 161150 538435 161166 538469
rect 161334 538435 161350 538469
rect 161530 538435 161546 538469
rect 161714 538435 161730 538469
rect 161930 538435 161946 538469
rect 162114 538435 162130 538469
rect 162310 538435 162326 538469
rect 162494 538435 162510 538469
rect 158664 538385 158698 538401
rect 158664 538193 158698 538209
rect 158922 538385 158956 538401
rect 158922 538193 158956 538209
rect 159040 538385 159074 538401
rect 159040 538193 159074 538209
rect 159298 538385 159332 538401
rect 159298 538193 159332 538209
rect 159556 538385 159590 538401
rect 159556 538193 159590 538209
rect 159814 538385 159848 538401
rect 159814 538193 159848 538209
rect 160072 538385 160106 538401
rect 160072 538193 160106 538209
rect 160330 538385 160364 538401
rect 160330 538193 160364 538209
rect 160588 538385 160622 538401
rect 160588 538193 160622 538209
rect 160846 538385 160880 538401
rect 160846 538193 160880 538209
rect 161104 538385 161138 538401
rect 161104 538193 161138 538209
rect 161362 538385 161396 538401
rect 161362 538193 161396 538209
rect 161484 538385 161518 538401
rect 161484 538193 161518 538209
rect 161742 538385 161776 538401
rect 161742 538193 161776 538209
rect 161884 538385 161918 538401
rect 161884 538193 161918 538209
rect 162142 538385 162176 538401
rect 162142 538193 162176 538209
rect 162264 538385 162298 538401
rect 162264 538193 162298 538209
rect 162522 538385 162556 538401
rect 162522 538193 162556 538209
rect 158710 538125 158726 538159
rect 158894 538125 158910 538159
rect 159086 538125 159102 538159
rect 159270 538125 159286 538159
rect 159344 538125 159360 538159
rect 159528 538125 159544 538159
rect 159602 538125 159618 538159
rect 159786 538125 159802 538159
rect 159860 538125 159876 538159
rect 160044 538125 160060 538159
rect 160118 538125 160134 538159
rect 160302 538125 160318 538159
rect 160376 538125 160392 538159
rect 160560 538125 160576 538159
rect 160634 538125 160650 538159
rect 160818 538125 160834 538159
rect 160892 538125 160908 538159
rect 161076 538125 161092 538159
rect 161150 538125 161166 538159
rect 161334 538125 161350 538159
rect 161530 538125 161546 538159
rect 161714 538125 161730 538159
rect 161930 538125 161946 538159
rect 162114 538125 162130 538159
rect 162310 538125 162326 538159
rect 162494 538125 162510 538159
rect 162788 538005 162808 538645
rect 162848 538005 162868 538645
rect 164518 538315 164538 539715
rect 164578 539695 164618 539715
rect 166538 539715 166638 539735
rect 166538 539695 166578 539715
rect 164578 539675 166578 539695
rect 164578 538355 164598 539675
rect 166538 539655 166578 539675
rect 164696 539572 164712 539606
rect 164746 539572 164762 539606
rect 165019 539579 165035 539613
rect 165069 539579 165085 539613
rect 165211 539579 165227 539613
rect 165261 539579 165277 539613
rect 165403 539579 165419 539613
rect 165453 539579 165469 539613
rect 165595 539579 165611 539613
rect 165645 539579 165661 539613
rect 165787 539579 165803 539613
rect 165837 539579 165853 539613
rect 165979 539579 165995 539613
rect 166029 539579 166045 539613
rect 166196 539572 166212 539606
rect 166246 539572 166262 539606
rect 166396 539572 166412 539606
rect 166446 539572 166462 539606
rect 164668 539513 164702 539529
rect 164668 538521 164702 538537
rect 164756 539513 164790 539529
rect 164756 538521 164790 538537
rect 164891 539520 164925 539536
rect 164891 538528 164925 538544
rect 164987 539520 165021 539536
rect 164987 538528 165021 538544
rect 165083 539520 165117 539536
rect 165083 538528 165117 538544
rect 165179 539520 165213 539536
rect 165179 538528 165213 538544
rect 165275 539520 165309 539536
rect 165275 538528 165309 538544
rect 165371 539520 165405 539536
rect 165371 538528 165405 538544
rect 165467 539520 165501 539536
rect 165467 538528 165501 538544
rect 165563 539520 165597 539536
rect 165563 538528 165597 538544
rect 165659 539520 165693 539536
rect 165659 538528 165693 538544
rect 165755 539520 165789 539536
rect 165755 538528 165789 538544
rect 165851 539520 165885 539536
rect 165851 538528 165885 538544
rect 165947 539520 165981 539536
rect 165947 538528 165981 538544
rect 166043 539520 166077 539536
rect 166168 539513 166202 539529
rect 166168 538921 166202 538937
rect 166256 539513 166290 539529
rect 166256 538921 166290 538937
rect 166368 539513 166402 539529
rect 166196 538844 166212 538878
rect 166246 538844 166262 538878
rect 166043 538528 166077 538544
rect 166368 538521 166402 538537
rect 166456 539513 166490 539529
rect 166456 538521 166490 538537
rect 166558 539265 166578 539655
rect 166558 539175 166568 539265
rect 164696 538444 164712 538478
rect 164746 538444 164762 538478
rect 164923 538451 164939 538485
rect 164973 538451 164989 538485
rect 165115 538451 165131 538485
rect 165165 538451 165181 538485
rect 165307 538451 165323 538485
rect 165357 538451 165373 538485
rect 165499 538451 165515 538485
rect 165549 538451 165565 538485
rect 165691 538451 165707 538485
rect 165741 538451 165757 538485
rect 165883 538451 165899 538485
rect 165933 538451 165949 538485
rect 166396 538444 166412 538478
rect 166446 538444 166462 538478
rect 166558 538355 166578 539175
rect 164578 538335 166578 538355
rect 164578 538315 164618 538335
rect 164518 538295 164618 538315
rect 166538 538315 166578 538335
rect 166618 538315 166638 539715
rect 166538 538295 166638 538315
rect 164518 538275 166638 538295
rect 168318 539735 170438 539755
rect 168318 539715 168418 539735
rect 168318 538315 168338 539715
rect 168378 539695 168418 539715
rect 170338 539715 170438 539735
rect 170338 539695 170378 539715
rect 168378 539675 170378 539695
rect 168378 538355 168398 539675
rect 170338 539655 170378 539675
rect 168496 539572 168512 539606
rect 168546 539572 168562 539606
rect 168819 539579 168835 539613
rect 168869 539579 168885 539613
rect 169011 539579 169027 539613
rect 169061 539579 169077 539613
rect 169203 539579 169219 539613
rect 169253 539579 169269 539613
rect 169395 539579 169411 539613
rect 169445 539579 169461 539613
rect 169587 539579 169603 539613
rect 169637 539579 169653 539613
rect 169779 539579 169795 539613
rect 169829 539579 169845 539613
rect 169996 539572 170012 539606
rect 170046 539572 170062 539606
rect 170196 539572 170212 539606
rect 170246 539572 170262 539606
rect 168468 539513 168502 539529
rect 168468 538521 168502 538537
rect 168556 539513 168590 539529
rect 168556 538521 168590 538537
rect 168691 539520 168725 539536
rect 168691 538528 168725 538544
rect 168787 539520 168821 539536
rect 168787 538528 168821 538544
rect 168883 539520 168917 539536
rect 168883 538528 168917 538544
rect 168979 539520 169013 539536
rect 168979 538528 169013 538544
rect 169075 539520 169109 539536
rect 169075 538528 169109 538544
rect 169171 539520 169205 539536
rect 169171 538528 169205 538544
rect 169267 539520 169301 539536
rect 169267 538528 169301 538544
rect 169363 539520 169397 539536
rect 169363 538528 169397 538544
rect 169459 539520 169493 539536
rect 169459 538528 169493 538544
rect 169555 539520 169589 539536
rect 169555 538528 169589 538544
rect 169651 539520 169685 539536
rect 169651 538528 169685 538544
rect 169747 539520 169781 539536
rect 169747 538528 169781 538544
rect 169843 539520 169877 539536
rect 169968 539513 170002 539529
rect 169968 538921 170002 538937
rect 170056 539513 170090 539529
rect 170056 538921 170090 538937
rect 170168 539513 170202 539529
rect 169996 538844 170012 538878
rect 170046 538844 170062 538878
rect 169843 538528 169877 538544
rect 170168 538521 170202 538537
rect 170256 539513 170290 539529
rect 170256 538521 170290 538537
rect 170358 539265 170378 539655
rect 170358 539175 170368 539265
rect 168496 538444 168512 538478
rect 168546 538444 168562 538478
rect 168723 538451 168739 538485
rect 168773 538451 168789 538485
rect 168915 538451 168931 538485
rect 168965 538451 168981 538485
rect 169107 538451 169123 538485
rect 169157 538451 169173 538485
rect 169299 538451 169315 538485
rect 169349 538451 169365 538485
rect 169491 538451 169507 538485
rect 169541 538451 169557 538485
rect 169683 538451 169699 538485
rect 169733 538451 169749 538485
rect 170196 538444 170212 538478
rect 170246 538444 170262 538478
rect 170358 538355 170378 539175
rect 168378 538335 170378 538355
rect 168378 538315 168418 538335
rect 168318 538295 168418 538315
rect 170338 538315 170378 538335
rect 170418 538315 170438 539715
rect 170338 538295 170438 538315
rect 168318 538275 170438 538295
rect 172018 539735 174138 539755
rect 172018 539715 172118 539735
rect 172018 538315 172038 539715
rect 172078 539695 172118 539715
rect 174038 539715 174138 539735
rect 174038 539695 174078 539715
rect 172078 539675 174078 539695
rect 172078 538355 172098 539675
rect 174038 539655 174078 539675
rect 172196 539572 172212 539606
rect 172246 539572 172262 539606
rect 172519 539579 172535 539613
rect 172569 539579 172585 539613
rect 172711 539579 172727 539613
rect 172761 539579 172777 539613
rect 172903 539579 172919 539613
rect 172953 539579 172969 539613
rect 173095 539579 173111 539613
rect 173145 539579 173161 539613
rect 173287 539579 173303 539613
rect 173337 539579 173353 539613
rect 173479 539579 173495 539613
rect 173529 539579 173545 539613
rect 173696 539572 173712 539606
rect 173746 539572 173762 539606
rect 173896 539572 173912 539606
rect 173946 539572 173962 539606
rect 172168 539513 172202 539529
rect 172168 538521 172202 538537
rect 172256 539513 172290 539529
rect 172256 538521 172290 538537
rect 172391 539520 172425 539536
rect 172391 538528 172425 538544
rect 172487 539520 172521 539536
rect 172487 538528 172521 538544
rect 172583 539520 172617 539536
rect 172583 538528 172617 538544
rect 172679 539520 172713 539536
rect 172679 538528 172713 538544
rect 172775 539520 172809 539536
rect 172775 538528 172809 538544
rect 172871 539520 172905 539536
rect 172871 538528 172905 538544
rect 172967 539520 173001 539536
rect 172967 538528 173001 538544
rect 173063 539520 173097 539536
rect 173063 538528 173097 538544
rect 173159 539520 173193 539536
rect 173159 538528 173193 538544
rect 173255 539520 173289 539536
rect 173255 538528 173289 538544
rect 173351 539520 173385 539536
rect 173351 538528 173385 538544
rect 173447 539520 173481 539536
rect 173447 538528 173481 538544
rect 173543 539520 173577 539536
rect 173668 539513 173702 539529
rect 173668 538921 173702 538937
rect 173756 539513 173790 539529
rect 173756 538921 173790 538937
rect 173868 539513 173902 539529
rect 173696 538844 173712 538878
rect 173746 538844 173762 538878
rect 173543 538528 173577 538544
rect 173868 538521 173902 538537
rect 173956 539513 173990 539529
rect 173956 538521 173990 538537
rect 174058 539265 174078 539655
rect 174058 539175 174068 539265
rect 172196 538444 172212 538478
rect 172246 538444 172262 538478
rect 172423 538451 172439 538485
rect 172473 538451 172489 538485
rect 172615 538451 172631 538485
rect 172665 538451 172681 538485
rect 172807 538451 172823 538485
rect 172857 538451 172873 538485
rect 172999 538451 173015 538485
rect 173049 538451 173065 538485
rect 173191 538451 173207 538485
rect 173241 538451 173257 538485
rect 173383 538451 173399 538485
rect 173433 538451 173449 538485
rect 173896 538444 173912 538478
rect 173946 538444 173962 538478
rect 174058 538355 174078 539175
rect 172078 538335 174078 538355
rect 172078 538315 172118 538335
rect 172018 538295 172118 538315
rect 174038 538315 174078 538335
rect 174118 538315 174138 539715
rect 174038 538295 174138 538315
rect 172018 538275 174138 538295
rect 175518 539735 177638 539755
rect 175518 539715 175618 539735
rect 175518 538315 175538 539715
rect 175578 539695 175618 539715
rect 177538 539715 177638 539735
rect 177538 539695 177578 539715
rect 175578 539675 177578 539695
rect 175578 538355 175598 539675
rect 177538 539655 177578 539675
rect 175696 539572 175712 539606
rect 175746 539572 175762 539606
rect 176019 539579 176035 539613
rect 176069 539579 176085 539613
rect 176211 539579 176227 539613
rect 176261 539579 176277 539613
rect 176403 539579 176419 539613
rect 176453 539579 176469 539613
rect 176595 539579 176611 539613
rect 176645 539579 176661 539613
rect 176787 539579 176803 539613
rect 176837 539579 176853 539613
rect 176979 539579 176995 539613
rect 177029 539579 177045 539613
rect 177196 539572 177212 539606
rect 177246 539572 177262 539606
rect 177396 539572 177412 539606
rect 177446 539572 177462 539606
rect 175668 539513 175702 539529
rect 175668 538521 175702 538537
rect 175756 539513 175790 539529
rect 175756 538521 175790 538537
rect 175891 539520 175925 539536
rect 175891 538528 175925 538544
rect 175987 539520 176021 539536
rect 175987 538528 176021 538544
rect 176083 539520 176117 539536
rect 176083 538528 176117 538544
rect 176179 539520 176213 539536
rect 176179 538528 176213 538544
rect 176275 539520 176309 539536
rect 176275 538528 176309 538544
rect 176371 539520 176405 539536
rect 176371 538528 176405 538544
rect 176467 539520 176501 539536
rect 176467 538528 176501 538544
rect 176563 539520 176597 539536
rect 176563 538528 176597 538544
rect 176659 539520 176693 539536
rect 176659 538528 176693 538544
rect 176755 539520 176789 539536
rect 176755 538528 176789 538544
rect 176851 539520 176885 539536
rect 176851 538528 176885 538544
rect 176947 539520 176981 539536
rect 176947 538528 176981 538544
rect 177043 539520 177077 539536
rect 177168 539513 177202 539529
rect 177168 538921 177202 538937
rect 177256 539513 177290 539529
rect 177256 538921 177290 538937
rect 177368 539513 177402 539529
rect 177196 538844 177212 538878
rect 177246 538844 177262 538878
rect 177043 538528 177077 538544
rect 177368 538521 177402 538537
rect 177456 539513 177490 539529
rect 177456 538521 177490 538537
rect 177558 539265 177578 539655
rect 177558 539175 177568 539265
rect 175696 538444 175712 538478
rect 175746 538444 175762 538478
rect 175923 538451 175939 538485
rect 175973 538451 175989 538485
rect 176115 538451 176131 538485
rect 176165 538451 176181 538485
rect 176307 538451 176323 538485
rect 176357 538451 176373 538485
rect 176499 538451 176515 538485
rect 176549 538451 176565 538485
rect 176691 538451 176707 538485
rect 176741 538451 176757 538485
rect 176883 538451 176899 538485
rect 176933 538451 176949 538485
rect 177396 538444 177412 538478
rect 177446 538444 177462 538478
rect 177558 538355 177578 539175
rect 175578 538335 177578 538355
rect 175578 538315 175618 538335
rect 175518 538295 175618 538315
rect 177538 538315 177578 538335
rect 177618 538315 177638 539715
rect 177538 538295 177638 538315
rect 175518 538275 177638 538295
rect 179118 539735 181238 539755
rect 179118 539715 179218 539735
rect 179118 538315 179138 539715
rect 179178 539695 179218 539715
rect 181138 539715 181238 539735
rect 181138 539695 181178 539715
rect 179178 539675 181178 539695
rect 179178 538355 179198 539675
rect 181138 539655 181178 539675
rect 179296 539572 179312 539606
rect 179346 539572 179362 539606
rect 179619 539579 179635 539613
rect 179669 539579 179685 539613
rect 179811 539579 179827 539613
rect 179861 539579 179877 539613
rect 180003 539579 180019 539613
rect 180053 539579 180069 539613
rect 180195 539579 180211 539613
rect 180245 539579 180261 539613
rect 180387 539579 180403 539613
rect 180437 539579 180453 539613
rect 180579 539579 180595 539613
rect 180629 539579 180645 539613
rect 180796 539572 180812 539606
rect 180846 539572 180862 539606
rect 180996 539572 181012 539606
rect 181046 539572 181062 539606
rect 179268 539513 179302 539529
rect 179268 538521 179302 538537
rect 179356 539513 179390 539529
rect 179356 538521 179390 538537
rect 179491 539520 179525 539536
rect 179491 538528 179525 538544
rect 179587 539520 179621 539536
rect 179587 538528 179621 538544
rect 179683 539520 179717 539536
rect 179683 538528 179717 538544
rect 179779 539520 179813 539536
rect 179779 538528 179813 538544
rect 179875 539520 179909 539536
rect 179875 538528 179909 538544
rect 179971 539520 180005 539536
rect 179971 538528 180005 538544
rect 180067 539520 180101 539536
rect 180067 538528 180101 538544
rect 180163 539520 180197 539536
rect 180163 538528 180197 538544
rect 180259 539520 180293 539536
rect 180259 538528 180293 538544
rect 180355 539520 180389 539536
rect 180355 538528 180389 538544
rect 180451 539520 180485 539536
rect 180451 538528 180485 538544
rect 180547 539520 180581 539536
rect 180547 538528 180581 538544
rect 180643 539520 180677 539536
rect 180768 539513 180802 539529
rect 180768 538921 180802 538937
rect 180856 539513 180890 539529
rect 180856 538921 180890 538937
rect 180968 539513 181002 539529
rect 180796 538844 180812 538878
rect 180846 538844 180862 538878
rect 180643 538528 180677 538544
rect 180968 538521 181002 538537
rect 181056 539513 181090 539529
rect 181056 538521 181090 538537
rect 181158 539265 181178 539655
rect 181158 539175 181168 539265
rect 179296 538444 179312 538478
rect 179346 538444 179362 538478
rect 179523 538451 179539 538485
rect 179573 538451 179589 538485
rect 179715 538451 179731 538485
rect 179765 538451 179781 538485
rect 179907 538451 179923 538485
rect 179957 538451 179973 538485
rect 180099 538451 180115 538485
rect 180149 538451 180165 538485
rect 180291 538451 180307 538485
rect 180341 538451 180357 538485
rect 180483 538451 180499 538485
rect 180533 538451 180549 538485
rect 180996 538444 181012 538478
rect 181046 538444 181062 538478
rect 181158 538355 181178 539175
rect 179178 538335 181178 538355
rect 179178 538315 179218 538335
rect 179118 538295 179218 538315
rect 181138 538315 181178 538335
rect 181218 538315 181238 539715
rect 181138 538295 181238 538315
rect 179118 538275 181238 538295
rect 182418 539735 184538 539755
rect 182418 539715 182518 539735
rect 182418 538315 182438 539715
rect 182478 539695 182518 539715
rect 184438 539715 184538 539735
rect 184438 539695 184478 539715
rect 182478 539675 184478 539695
rect 182478 538355 182498 539675
rect 184438 539655 184478 539675
rect 182596 539572 182612 539606
rect 182646 539572 182662 539606
rect 182919 539579 182935 539613
rect 182969 539579 182985 539613
rect 183111 539579 183127 539613
rect 183161 539579 183177 539613
rect 183303 539579 183319 539613
rect 183353 539579 183369 539613
rect 183495 539579 183511 539613
rect 183545 539579 183561 539613
rect 183687 539579 183703 539613
rect 183737 539579 183753 539613
rect 183879 539579 183895 539613
rect 183929 539579 183945 539613
rect 184096 539572 184112 539606
rect 184146 539572 184162 539606
rect 184296 539572 184312 539606
rect 184346 539572 184362 539606
rect 182568 539513 182602 539529
rect 182568 538521 182602 538537
rect 182656 539513 182690 539529
rect 182656 538521 182690 538537
rect 182791 539520 182825 539536
rect 182791 538528 182825 538544
rect 182887 539520 182921 539536
rect 182887 538528 182921 538544
rect 182983 539520 183017 539536
rect 182983 538528 183017 538544
rect 183079 539520 183113 539536
rect 183079 538528 183113 538544
rect 183175 539520 183209 539536
rect 183175 538528 183209 538544
rect 183271 539520 183305 539536
rect 183271 538528 183305 538544
rect 183367 539520 183401 539536
rect 183367 538528 183401 538544
rect 183463 539520 183497 539536
rect 183463 538528 183497 538544
rect 183559 539520 183593 539536
rect 183559 538528 183593 538544
rect 183655 539520 183689 539536
rect 183655 538528 183689 538544
rect 183751 539520 183785 539536
rect 183751 538528 183785 538544
rect 183847 539520 183881 539536
rect 183847 538528 183881 538544
rect 183943 539520 183977 539536
rect 184068 539513 184102 539529
rect 184068 538921 184102 538937
rect 184156 539513 184190 539529
rect 184156 538921 184190 538937
rect 184268 539513 184302 539529
rect 184096 538844 184112 538878
rect 184146 538844 184162 538878
rect 183943 538528 183977 538544
rect 184268 538521 184302 538537
rect 184356 539513 184390 539529
rect 184356 538521 184390 538537
rect 184458 539265 184478 539655
rect 184458 539175 184468 539265
rect 182596 538444 182612 538478
rect 182646 538444 182662 538478
rect 182823 538451 182839 538485
rect 182873 538451 182889 538485
rect 183015 538451 183031 538485
rect 183065 538451 183081 538485
rect 183207 538451 183223 538485
rect 183257 538451 183273 538485
rect 183399 538451 183415 538485
rect 183449 538451 183465 538485
rect 183591 538451 183607 538485
rect 183641 538451 183657 538485
rect 183783 538451 183799 538485
rect 183833 538451 183849 538485
rect 184296 538444 184312 538478
rect 184346 538444 184362 538478
rect 184458 538355 184478 539175
rect 182478 538335 184478 538355
rect 182478 538315 182518 538335
rect 182418 538295 182518 538315
rect 184438 538315 184478 538335
rect 184518 538315 184538 539715
rect 184438 538295 184538 538315
rect 182418 538275 184538 538295
rect 185718 539735 187838 539755
rect 185718 539715 185818 539735
rect 185718 538315 185738 539715
rect 185778 539695 185818 539715
rect 187738 539715 187838 539735
rect 187738 539695 187778 539715
rect 185778 539675 187778 539695
rect 185778 538355 185798 539675
rect 187738 539655 187778 539675
rect 185896 539572 185912 539606
rect 185946 539572 185962 539606
rect 186219 539579 186235 539613
rect 186269 539579 186285 539613
rect 186411 539579 186427 539613
rect 186461 539579 186477 539613
rect 186603 539579 186619 539613
rect 186653 539579 186669 539613
rect 186795 539579 186811 539613
rect 186845 539579 186861 539613
rect 186987 539579 187003 539613
rect 187037 539579 187053 539613
rect 187179 539579 187195 539613
rect 187229 539579 187245 539613
rect 187396 539572 187412 539606
rect 187446 539572 187462 539606
rect 187596 539572 187612 539606
rect 187646 539572 187662 539606
rect 185868 539513 185902 539529
rect 185868 538521 185902 538537
rect 185956 539513 185990 539529
rect 185956 538521 185990 538537
rect 186091 539520 186125 539536
rect 186091 538528 186125 538544
rect 186187 539520 186221 539536
rect 186187 538528 186221 538544
rect 186283 539520 186317 539536
rect 186283 538528 186317 538544
rect 186379 539520 186413 539536
rect 186379 538528 186413 538544
rect 186475 539520 186509 539536
rect 186475 538528 186509 538544
rect 186571 539520 186605 539536
rect 186571 538528 186605 538544
rect 186667 539520 186701 539536
rect 186667 538528 186701 538544
rect 186763 539520 186797 539536
rect 186763 538528 186797 538544
rect 186859 539520 186893 539536
rect 186859 538528 186893 538544
rect 186955 539520 186989 539536
rect 186955 538528 186989 538544
rect 187051 539520 187085 539536
rect 187051 538528 187085 538544
rect 187147 539520 187181 539536
rect 187147 538528 187181 538544
rect 187243 539520 187277 539536
rect 187368 539513 187402 539529
rect 187368 538921 187402 538937
rect 187456 539513 187490 539529
rect 187456 538921 187490 538937
rect 187568 539513 187602 539529
rect 187396 538844 187412 538878
rect 187446 538844 187462 538878
rect 187243 538528 187277 538544
rect 187568 538521 187602 538537
rect 187656 539513 187690 539529
rect 187656 538521 187690 538537
rect 187758 539265 187778 539655
rect 187758 539175 187768 539265
rect 185896 538444 185912 538478
rect 185946 538444 185962 538478
rect 186123 538451 186139 538485
rect 186173 538451 186189 538485
rect 186315 538451 186331 538485
rect 186365 538451 186381 538485
rect 186507 538451 186523 538485
rect 186557 538451 186573 538485
rect 186699 538451 186715 538485
rect 186749 538451 186765 538485
rect 186891 538451 186907 538485
rect 186941 538451 186957 538485
rect 187083 538451 187099 538485
rect 187133 538451 187149 538485
rect 187596 538444 187612 538478
rect 187646 538444 187662 538478
rect 187758 538355 187778 539175
rect 185778 538335 187778 538355
rect 185778 538315 185818 538335
rect 185718 538295 185818 538315
rect 187738 538315 187778 538335
rect 187818 538315 187838 539715
rect 187738 538295 187838 538315
rect 185718 538275 187838 538295
rect 189018 539735 191138 539755
rect 189018 539715 189118 539735
rect 189018 538315 189038 539715
rect 189078 539695 189118 539715
rect 191038 539715 191138 539735
rect 191038 539695 191078 539715
rect 189078 539675 191078 539695
rect 189078 538355 189098 539675
rect 191038 539655 191078 539675
rect 189196 539572 189212 539606
rect 189246 539572 189262 539606
rect 189519 539579 189535 539613
rect 189569 539579 189585 539613
rect 189711 539579 189727 539613
rect 189761 539579 189777 539613
rect 189903 539579 189919 539613
rect 189953 539579 189969 539613
rect 190095 539579 190111 539613
rect 190145 539579 190161 539613
rect 190287 539579 190303 539613
rect 190337 539579 190353 539613
rect 190479 539579 190495 539613
rect 190529 539579 190545 539613
rect 190696 539572 190712 539606
rect 190746 539572 190762 539606
rect 190896 539572 190912 539606
rect 190946 539572 190962 539606
rect 189168 539513 189202 539529
rect 189168 538521 189202 538537
rect 189256 539513 189290 539529
rect 189256 538521 189290 538537
rect 189391 539520 189425 539536
rect 189391 538528 189425 538544
rect 189487 539520 189521 539536
rect 189487 538528 189521 538544
rect 189583 539520 189617 539536
rect 189583 538528 189617 538544
rect 189679 539520 189713 539536
rect 189679 538528 189713 538544
rect 189775 539520 189809 539536
rect 189775 538528 189809 538544
rect 189871 539520 189905 539536
rect 189871 538528 189905 538544
rect 189967 539520 190001 539536
rect 189967 538528 190001 538544
rect 190063 539520 190097 539536
rect 190063 538528 190097 538544
rect 190159 539520 190193 539536
rect 190159 538528 190193 538544
rect 190255 539520 190289 539536
rect 190255 538528 190289 538544
rect 190351 539520 190385 539536
rect 190351 538528 190385 538544
rect 190447 539520 190481 539536
rect 190447 538528 190481 538544
rect 190543 539520 190577 539536
rect 190668 539513 190702 539529
rect 190668 538921 190702 538937
rect 190756 539513 190790 539529
rect 190756 538921 190790 538937
rect 190868 539513 190902 539529
rect 190696 538844 190712 538878
rect 190746 538844 190762 538878
rect 190543 538528 190577 538544
rect 190868 538521 190902 538537
rect 190956 539513 190990 539529
rect 190956 538521 190990 538537
rect 191058 539265 191078 539655
rect 191058 539175 191068 539265
rect 189196 538444 189212 538478
rect 189246 538444 189262 538478
rect 189423 538451 189439 538485
rect 189473 538451 189489 538485
rect 189615 538451 189631 538485
rect 189665 538451 189681 538485
rect 189807 538451 189823 538485
rect 189857 538451 189873 538485
rect 189999 538451 190015 538485
rect 190049 538451 190065 538485
rect 190191 538451 190207 538485
rect 190241 538451 190257 538485
rect 190383 538451 190399 538485
rect 190433 538451 190449 538485
rect 190896 538444 190912 538478
rect 190946 538444 190962 538478
rect 191058 538355 191078 539175
rect 189078 538335 191078 538355
rect 189078 538315 189118 538335
rect 189018 538295 189118 538315
rect 191038 538315 191078 538335
rect 191118 538315 191138 539715
rect 191038 538295 191138 538315
rect 189018 538275 191138 538295
rect 157688 537985 162868 538005
rect 157688 537965 157728 537985
rect 157628 537945 157728 537965
rect 162768 537945 162868 537985
rect 157628 537925 162868 537945
rect 164186 538045 164282 538079
rect 166646 538045 166742 538079
rect 164186 537983 164220 538045
rect 157588 537825 162848 537845
rect 157588 537785 157648 537825
rect 162748 537785 162848 537825
rect 157588 537765 162788 537785
rect 157588 537725 157668 537765
rect 157588 535785 157608 537725
rect 157648 535785 157668 537725
rect 161286 537672 161302 537706
rect 161336 537672 161352 537706
rect 161490 537672 161506 537706
rect 161540 537672 161556 537706
rect 161682 537672 161698 537706
rect 161732 537672 161748 537706
rect 161890 537672 161906 537706
rect 161940 537672 161956 537706
rect 162082 537672 162098 537706
rect 162132 537672 162148 537706
rect 162306 537672 162322 537706
rect 162356 537672 162372 537706
rect 161258 537613 161292 537629
rect 161258 537021 161292 537037
rect 161346 537613 161380 537629
rect 161346 537021 161380 537037
rect 161458 537613 161492 537629
rect 161458 537021 161492 537037
rect 161554 537613 161588 537629
rect 161554 537021 161588 537037
rect 161650 537613 161684 537629
rect 161650 537021 161684 537037
rect 161746 537613 161780 537629
rect 161746 537021 161780 537037
rect 161858 537613 161892 537629
rect 161858 537021 161892 537037
rect 161954 537613 161988 537629
rect 161954 537021 161988 537037
rect 162050 537613 162084 537629
rect 162050 537021 162084 537037
rect 162146 537613 162180 537629
rect 162146 537021 162180 537037
rect 162278 537613 162312 537629
rect 162278 537021 162312 537037
rect 162366 537613 162400 537629
rect 162366 537021 162400 537037
rect 161286 536944 161302 536978
rect 161336 536944 161352 536978
rect 161586 536944 161602 536978
rect 161636 536944 161652 536978
rect 161986 536944 162002 536978
rect 162036 536944 162052 536978
rect 162306 536944 162322 536978
rect 162356 536944 162372 536978
rect 157794 536652 157810 536686
rect 157978 536652 157994 536686
rect 158172 536652 158188 536686
rect 158356 536652 158372 536686
rect 158430 536652 158446 536686
rect 158614 536652 158630 536686
rect 158688 536652 158704 536686
rect 158872 536652 158888 536686
rect 158946 536652 158962 536686
rect 159130 536652 159146 536686
rect 159204 536652 159220 536686
rect 159388 536652 159404 536686
rect 159462 536652 159478 536686
rect 159646 536652 159662 536686
rect 159720 536652 159736 536686
rect 159904 536652 159920 536686
rect 159978 536652 159994 536686
rect 160162 536652 160178 536686
rect 160236 536652 160252 536686
rect 160420 536652 160436 536686
rect 160494 536652 160510 536686
rect 160678 536652 160694 536686
rect 160878 536652 160894 536686
rect 161062 536652 161078 536686
rect 161136 536652 161152 536686
rect 161320 536652 161336 536686
rect 161394 536652 161410 536686
rect 161578 536652 161594 536686
rect 161776 536652 161792 536686
rect 161960 536652 161976 536686
rect 162034 536652 162050 536686
rect 162218 536652 162234 536686
rect 162414 536652 162430 536686
rect 162598 536652 162614 536686
rect 157748 536593 157782 536609
rect 157748 536001 157782 536017
rect 158006 536593 158040 536609
rect 158006 536001 158040 536017
rect 158126 536593 158160 536609
rect 158126 536001 158160 536017
rect 158384 536593 158418 536609
rect 158384 536001 158418 536017
rect 158642 536593 158676 536609
rect 158642 536001 158676 536017
rect 158900 536593 158934 536609
rect 158900 536001 158934 536017
rect 159158 536593 159192 536609
rect 159158 536001 159192 536017
rect 159416 536593 159450 536609
rect 159416 536001 159450 536017
rect 159674 536593 159708 536609
rect 159674 536001 159708 536017
rect 159932 536593 159966 536609
rect 159932 536001 159966 536017
rect 160190 536593 160224 536609
rect 160190 536001 160224 536017
rect 160448 536593 160482 536609
rect 160448 536001 160482 536017
rect 160706 536593 160740 536609
rect 160706 536001 160740 536017
rect 160832 536593 160866 536609
rect 160832 536001 160866 536017
rect 161090 536593 161124 536609
rect 161090 536001 161124 536017
rect 161348 536593 161382 536609
rect 161348 536001 161382 536017
rect 161606 536593 161640 536609
rect 161606 536001 161640 536017
rect 161730 536593 161764 536609
rect 161730 536001 161764 536017
rect 161988 536593 162022 536609
rect 161988 536001 162022 536017
rect 162246 536593 162280 536609
rect 162246 536001 162280 536017
rect 162368 536593 162402 536609
rect 162368 536001 162402 536017
rect 162626 536593 162660 536609
rect 162626 536001 162660 536017
rect 157794 535924 157810 535958
rect 157978 535924 157994 535958
rect 158172 535924 158188 535958
rect 158356 535924 158372 535958
rect 158430 535924 158446 535958
rect 158614 535924 158630 535958
rect 158688 535924 158704 535958
rect 158872 535924 158888 535958
rect 158946 535924 158962 535958
rect 159130 535924 159146 535958
rect 159204 535924 159220 535958
rect 159388 535924 159404 535958
rect 159462 535924 159478 535958
rect 159646 535924 159662 535958
rect 159720 535924 159736 535958
rect 159904 535924 159920 535958
rect 159978 535924 159994 535958
rect 160162 535924 160178 535958
rect 160236 535924 160252 535958
rect 160420 535924 160436 535958
rect 160494 535924 160510 535958
rect 160678 535924 160694 535958
rect 160878 535924 160894 535958
rect 161062 535924 161078 535958
rect 161136 535924 161152 535958
rect 161320 535924 161336 535958
rect 161394 535924 161410 535958
rect 161578 535924 161594 535958
rect 161776 535924 161792 535958
rect 161960 535924 161976 535958
rect 162034 535924 162050 535958
rect 162218 535924 162234 535958
rect 162414 535924 162430 535958
rect 162598 535924 162614 535958
rect 157588 535765 157668 535785
rect 162768 535765 162788 537765
rect 162828 535765 162848 537785
rect 166708 537983 166742 538045
rect 164186 535905 164220 535967
rect 166708 535905 166742 535967
rect 164186 535871 164282 535905
rect 166646 535871 166742 535905
rect 167958 538045 168054 538079
rect 169146 538045 169242 538079
rect 167958 537983 167992 538045
rect 169208 537983 169242 538045
rect 167958 535905 167992 535967
rect 169208 535905 169242 535967
rect 167958 535871 168054 535905
rect 169146 535871 169242 535905
rect 171694 538045 171790 538079
rect 172246 538045 172342 538079
rect 171694 537983 171728 538045
rect 172308 537983 172342 538045
rect 171694 535905 171728 535967
rect 172308 535905 172342 535967
rect 171694 535871 171790 535905
rect 172246 535871 172342 535905
rect 175212 538045 175308 538079
rect 175446 538045 175542 538079
rect 175212 537983 175246 538045
rect 175508 537983 175542 538045
rect 175212 535905 175246 535967
rect 178812 538045 178908 538079
rect 179046 538045 179142 538079
rect 178812 537983 178846 538045
rect 179108 537983 179142 538045
rect 178812 536465 178846 536527
rect 182112 538045 182208 538079
rect 182346 538045 182442 538079
rect 182112 537983 182146 538045
rect 182408 537983 182442 538045
rect 182112 536745 182146 536807
rect 185412 538045 185508 538079
rect 185646 538045 185742 538079
rect 185412 537983 185446 538045
rect 185708 537983 185742 538045
rect 185412 536885 185446 536947
rect 185708 536885 185742 536947
rect 185412 536851 185508 536885
rect 185646 536851 185742 536885
rect 188712 538045 188808 538079
rect 188946 538045 189042 538079
rect 188712 537983 188746 538045
rect 189008 537983 189042 538045
rect 182408 536745 182442 536807
rect 188712 536789 188746 536851
rect 189008 536789 189042 536851
rect 188712 536755 188808 536789
rect 188946 536755 189042 536789
rect 182112 536711 182208 536745
rect 182346 536711 182442 536745
rect 179108 536465 179142 536527
rect 178812 536431 178908 536465
rect 179046 536431 179142 536465
rect 175508 535905 175542 535967
rect 175212 535871 175308 535905
rect 175446 535871 175542 535905
rect 157588 535745 162848 535765
rect 157588 535705 157668 535745
rect 162748 535705 162848 535745
rect 157588 535685 162848 535705
rect 164156 535705 164252 535739
rect 166616 535705 166712 535739
rect 164156 535643 164190 535705
rect 166678 535643 166712 535705
rect 164156 533565 164190 533627
rect 166678 533565 166712 533627
rect 164156 533531 164252 533565
rect 166616 533531 166712 533565
rect 172208 530562 172237 530596
rect 172271 530562 172329 530596
rect 172363 530562 172421 530596
rect 172455 530562 172513 530596
rect 172547 530562 172605 530596
rect 172639 530562 172697 530596
rect 172731 530562 172789 530596
rect 172823 530562 172881 530596
rect 172915 530562 172973 530596
rect 173007 530562 173065 530596
rect 173099 530562 173157 530596
rect 173191 530562 173249 530596
rect 173283 530562 173341 530596
rect 173375 530562 173433 530596
rect 173467 530562 173525 530596
rect 173559 530562 173617 530596
rect 173651 530562 173709 530596
rect 173743 530562 173801 530596
rect 173835 530562 173893 530596
rect 173927 530562 173985 530596
rect 174019 530562 174077 530596
rect 174111 530562 174169 530596
rect 174203 530562 174261 530596
rect 174295 530562 174353 530596
rect 174387 530562 174445 530596
rect 174479 530562 174537 530596
rect 174571 530562 174629 530596
rect 174663 530562 174721 530596
rect 174755 530562 174813 530596
rect 174847 530562 174905 530596
rect 174939 530562 174997 530596
rect 175031 530562 175089 530596
rect 175123 530562 175181 530596
rect 175215 530562 175273 530596
rect 175307 530562 175365 530596
rect 175399 530562 175457 530596
rect 175491 530562 175549 530596
rect 175583 530562 175641 530596
rect 175675 530562 175733 530596
rect 175767 530562 175825 530596
rect 175859 530562 175917 530596
rect 175951 530562 176009 530596
rect 176043 530562 176101 530596
rect 176135 530562 176193 530596
rect 176227 530562 176285 530596
rect 176319 530562 176377 530596
rect 176411 530562 176469 530596
rect 176503 530562 176561 530596
rect 176595 530562 176653 530596
rect 176687 530562 176745 530596
rect 176779 530562 176837 530596
rect 176871 530562 176929 530596
rect 176963 530562 177021 530596
rect 177055 530562 177113 530596
rect 177147 530562 177205 530596
rect 177239 530562 177297 530596
rect 177331 530562 177389 530596
rect 177423 530562 177481 530596
rect 177515 530562 177573 530596
rect 177607 530562 177665 530596
rect 177699 530562 177757 530596
rect 177791 530562 177849 530596
rect 177883 530562 177941 530596
rect 177975 530562 178033 530596
rect 178067 530562 178125 530596
rect 178159 530562 178217 530596
rect 178251 530562 178309 530596
rect 178343 530562 178401 530596
rect 178435 530562 178493 530596
rect 178527 530562 178585 530596
rect 178619 530562 178677 530596
rect 178711 530562 178769 530596
rect 178803 530562 178861 530596
rect 178895 530562 178953 530596
rect 178987 530562 179045 530596
rect 179079 530562 179137 530596
rect 179171 530562 179229 530596
rect 179263 530562 179321 530596
rect 179355 530562 179413 530596
rect 179447 530562 179505 530596
rect 179539 530562 179597 530596
rect 179631 530562 179689 530596
rect 179723 530562 179781 530596
rect 179815 530562 179873 530596
rect 179907 530562 179965 530596
rect 179999 530562 180057 530596
rect 180091 530562 180149 530596
rect 180183 530562 180241 530596
rect 180275 530562 180333 530596
rect 180367 530562 180425 530596
rect 180459 530562 180517 530596
rect 180551 530562 180609 530596
rect 180643 530562 180701 530596
rect 180735 530562 180793 530596
rect 180827 530562 180885 530596
rect 180919 530562 180977 530596
rect 181011 530562 181069 530596
rect 181103 530562 181161 530596
rect 181195 530562 181253 530596
rect 181287 530562 181345 530596
rect 181379 530562 181437 530596
rect 181471 530562 181529 530596
rect 181563 530562 181621 530596
rect 181655 530562 181713 530596
rect 181747 530562 181805 530596
rect 181839 530562 181897 530596
rect 181931 530562 181989 530596
rect 182023 530562 182081 530596
rect 182115 530562 182173 530596
rect 182207 530562 182265 530596
rect 182299 530562 182357 530596
rect 182391 530562 182449 530596
rect 182483 530562 182541 530596
rect 182575 530562 182633 530596
rect 182667 530562 182725 530596
rect 182759 530562 182817 530596
rect 182851 530562 182909 530596
rect 182943 530562 183001 530596
rect 183035 530562 183093 530596
rect 183127 530562 183185 530596
rect 183219 530562 183277 530596
rect 183311 530562 183369 530596
rect 183403 530562 183461 530596
rect 183495 530562 183553 530596
rect 183587 530562 183645 530596
rect 183679 530562 183737 530596
rect 183771 530562 183829 530596
rect 183863 530562 183921 530596
rect 183955 530562 184013 530596
rect 184047 530562 184105 530596
rect 184139 530562 184197 530596
rect 184231 530562 184289 530596
rect 184323 530562 184381 530596
rect 184415 530562 184473 530596
rect 184507 530562 184565 530596
rect 184599 530562 184657 530596
rect 184691 530562 184749 530596
rect 184783 530562 184841 530596
rect 184875 530562 184933 530596
rect 184967 530562 185025 530596
rect 185059 530562 185117 530596
rect 185151 530562 185209 530596
rect 185243 530562 185301 530596
rect 185335 530562 185393 530596
rect 185427 530562 185485 530596
rect 185519 530562 185577 530596
rect 185611 530562 185669 530596
rect 185703 530562 185761 530596
rect 185795 530562 185853 530596
rect 185887 530562 185945 530596
rect 185979 530562 186037 530596
rect 186071 530562 186129 530596
rect 186163 530562 186221 530596
rect 186255 530562 186313 530596
rect 186347 530562 186405 530596
rect 186439 530562 186497 530596
rect 186531 530562 186589 530596
rect 186623 530562 186681 530596
rect 186715 530562 186773 530596
rect 186807 530562 186865 530596
rect 186899 530562 186957 530596
rect 186991 530562 187049 530596
rect 187083 530562 187141 530596
rect 187175 530562 187233 530596
rect 187267 530562 187325 530596
rect 187359 530562 187417 530596
rect 187451 530562 187480 530596
rect 172225 530499 172467 530562
rect 172225 530465 172243 530499
rect 172277 530465 172415 530499
rect 172449 530465 172467 530499
rect 172513 530516 172569 530562
rect 172513 530482 172526 530516
rect 172560 530482 172569 530516
rect 172690 530516 172741 530562
rect 172513 530466 172569 530482
rect 172603 530494 172655 530510
rect 172225 530412 172467 530465
rect 172603 530460 172612 530494
rect 172646 530460 172655 530494
rect 172690 530482 172698 530516
rect 172732 530482 172741 530516
rect 172870 530516 172925 530562
rect 172690 530466 172741 530482
rect 172775 530494 172834 530510
rect 172603 530432 172655 530460
rect 172775 530460 172784 530494
rect 172818 530460 172834 530494
rect 172870 530482 172881 530516
rect 172915 530482 172925 530516
rect 172870 530466 172925 530482
rect 172959 530512 173019 530528
rect 172959 530478 172967 530512
rect 173001 530478 173019 530512
rect 172959 530462 173019 530478
rect 172775 530432 172834 530460
rect 172504 530426 172834 530432
rect 172225 530338 172329 530412
rect 172504 530392 172513 530426
rect 172547 530398 172834 530426
rect 172547 530392 172585 530398
rect 172225 530304 172275 530338
rect 172309 530304 172329 530338
rect 172363 530344 172383 530378
rect 172417 530344 172467 530378
rect 172363 530270 172467 530344
rect 172225 530223 172467 530270
rect 172504 530296 172585 530392
rect 172881 530364 172951 530428
rect 172619 530330 172635 530364
rect 172669 530330 172703 530364
rect 172737 530330 172771 530364
rect 172805 530330 172847 530364
rect 172504 530272 172655 530296
rect 172504 530262 172613 530272
rect 172603 530238 172613 530262
rect 172647 530238 172655 530272
rect 172813 530280 172847 530330
rect 172881 530358 172917 530364
rect 172915 530330 172917 530358
rect 172915 530324 172951 530330
rect 172881 530314 172951 530324
rect 172985 530280 173019 530462
rect 173053 530501 174122 530562
rect 173053 530467 173071 530501
rect 173105 530467 174071 530501
rect 174105 530467 174122 530501
rect 173053 530453 174122 530467
rect 174157 530501 174675 530562
rect 174157 530467 174175 530501
rect 174209 530467 174623 530501
rect 174657 530467 174675 530501
rect 173370 530338 173438 530453
rect 174157 530408 174675 530467
rect 174801 530468 174859 530562
rect 174801 530434 174813 530468
rect 174847 530434 174859 530468
rect 174905 530516 174961 530562
rect 174905 530482 174918 530516
rect 174952 530482 174961 530516
rect 175082 530516 175133 530562
rect 174905 530466 174961 530482
rect 174995 530494 175047 530510
rect 174801 530417 174859 530434
rect 174995 530460 175004 530494
rect 175038 530460 175047 530494
rect 175082 530482 175090 530516
rect 175124 530482 175133 530516
rect 175262 530516 175317 530562
rect 175082 530466 175133 530482
rect 175167 530494 175226 530510
rect 174995 530432 175047 530460
rect 175167 530460 175176 530494
rect 175210 530460 175226 530494
rect 175262 530482 175273 530516
rect 175307 530482 175317 530516
rect 175262 530466 175317 530482
rect 175351 530512 175411 530528
rect 175351 530478 175359 530512
rect 175393 530478 175411 530512
rect 175351 530462 175411 530478
rect 175167 530432 175226 530460
rect 174896 530426 175226 530432
rect 173370 530304 173387 530338
rect 173421 530304 173438 530338
rect 173370 530287 173438 530304
rect 173734 530374 173804 530389
rect 173734 530340 173751 530374
rect 173785 530340 173804 530374
rect 172813 530258 173019 530280
rect 172813 530246 172967 530258
rect 172225 530189 172243 530223
rect 172277 530189 172415 530223
rect 172449 530189 172467 530223
rect 172225 530128 172467 530189
rect 172225 530094 172243 530128
rect 172277 530094 172415 530128
rect 172449 530094 172467 530128
rect 172225 530052 172467 530094
rect 172512 530210 172569 530226
rect 172512 530176 172527 530210
rect 172561 530176 172569 530210
rect 172512 530142 172569 530176
rect 172512 530108 172527 530142
rect 172561 530108 172569 530142
rect 172512 530052 172569 530108
rect 172603 530212 172655 530238
rect 172957 530224 172967 530246
rect 173001 530224 173019 530258
rect 172603 530204 172827 530212
rect 172603 530170 172613 530204
rect 172647 530178 172827 530204
rect 172647 530170 172655 530178
rect 172603 530136 172655 530170
rect 172775 530163 172827 530178
rect 172603 530102 172613 530136
rect 172647 530102 172655 530136
rect 172603 530086 172655 530102
rect 172690 530128 172741 530144
rect 172690 530094 172699 530128
rect 172733 530094 172741 530128
rect 172690 530052 172741 530094
rect 172775 530129 172785 530163
rect 172819 530129 172827 530163
rect 172775 530086 172827 530129
rect 172861 530196 172923 530212
rect 172861 530162 172881 530196
rect 172915 530162 172923 530196
rect 172861 530128 172923 530162
rect 172861 530094 172881 530128
rect 172915 530094 172923 530128
rect 172861 530052 172923 530094
rect 172957 530136 173019 530224
rect 173734 530139 173804 530340
rect 174157 530338 174399 530408
rect 174896 530392 174905 530426
rect 174939 530398 175226 530426
rect 174939 530392 174977 530398
rect 174157 530304 174235 530338
rect 174269 530304 174345 530338
rect 174379 530304 174399 530338
rect 174433 530340 174453 530374
rect 174487 530340 174563 530374
rect 174597 530340 174675 530374
rect 174433 530270 174675 530340
rect 174896 530296 174977 530392
rect 175273 530364 175343 530428
rect 175011 530330 175027 530364
rect 175061 530330 175095 530364
rect 175129 530330 175163 530364
rect 175197 530330 175239 530364
rect 174157 530230 174675 530270
rect 174157 530196 174175 530230
rect 174209 530196 174623 530230
rect 174657 530196 174675 530230
rect 172957 530102 172967 530136
rect 173001 530102 173019 530136
rect 172957 530086 173019 530102
rect 173053 530128 174122 530139
rect 173053 530094 173071 530128
rect 173105 530094 174071 530128
rect 174105 530094 174122 530128
rect 173053 530052 174122 530094
rect 174157 530128 174675 530196
rect 174157 530094 174175 530128
rect 174209 530094 174623 530128
rect 174657 530094 174675 530128
rect 174157 530052 174675 530094
rect 174801 530250 174859 530285
rect 174896 530272 175047 530296
rect 174896 530262 175005 530272
rect 174801 530216 174813 530250
rect 174847 530216 174859 530250
rect 174995 530238 175005 530262
rect 175039 530238 175047 530272
rect 175205 530280 175239 530330
rect 175273 530358 175309 530364
rect 175307 530330 175309 530358
rect 175307 530324 175343 530330
rect 175273 530314 175343 530324
rect 175377 530280 175411 530462
rect 175205 530258 175411 530280
rect 175205 530246 175359 530258
rect 174801 530157 174859 530216
rect 174801 530123 174813 530157
rect 174847 530123 174859 530157
rect 174801 530052 174859 530123
rect 174904 530210 174961 530226
rect 174904 530176 174919 530210
rect 174953 530176 174961 530210
rect 174904 530142 174961 530176
rect 174904 530108 174919 530142
rect 174953 530108 174961 530142
rect 174904 530052 174961 530108
rect 174995 530212 175047 530238
rect 175349 530224 175359 530246
rect 175393 530224 175411 530258
rect 174995 530204 175219 530212
rect 174995 530170 175005 530204
rect 175039 530178 175219 530204
rect 175039 530170 175047 530178
rect 174995 530136 175047 530170
rect 175167 530163 175219 530178
rect 174995 530102 175005 530136
rect 175039 530102 175047 530136
rect 174995 530086 175047 530102
rect 175082 530128 175133 530144
rect 175082 530094 175091 530128
rect 175125 530094 175133 530128
rect 175082 530052 175133 530094
rect 175167 530129 175177 530163
rect 175211 530129 175219 530163
rect 175167 530086 175219 530129
rect 175253 530196 175315 530212
rect 175253 530162 175273 530196
rect 175307 530162 175315 530196
rect 175253 530128 175315 530162
rect 175253 530094 175273 530128
rect 175307 530094 175315 530128
rect 175253 530052 175315 530094
rect 175349 530136 175411 530224
rect 175349 530102 175359 530136
rect 175393 530102 175411 530136
rect 175538 530470 175589 530526
rect 175623 530520 175684 530562
rect 175981 530524 176019 530562
rect 175623 530486 175639 530520
rect 175673 530486 175684 530520
rect 175623 530470 175684 530486
rect 175733 530504 175947 530520
rect 175733 530470 175763 530504
rect 175797 530486 175947 530504
rect 175538 530436 175555 530470
rect 175538 530420 175589 530436
rect 175538 530290 175580 530420
rect 175733 530415 175797 530470
rect 175732 530380 175797 530415
rect 175614 530364 175797 530380
rect 175648 530330 175797 530364
rect 175614 530320 175797 530330
rect 175831 530426 175879 530452
rect 175831 530392 175845 530426
rect 175913 530440 175947 530486
rect 176015 530490 176019 530524
rect 175981 530474 176019 530490
rect 176053 530520 176243 530528
rect 176053 530486 176193 530520
rect 176227 530486 176243 530520
rect 176287 530490 176303 530524
rect 176337 530490 176357 530524
rect 176053 530472 176243 530486
rect 175913 530406 176019 530440
rect 175831 530372 175879 530392
rect 175975 530400 176019 530406
rect 175831 530338 175889 530372
rect 175923 530363 175939 530372
rect 175975 530366 175985 530400
rect 175975 530350 176019 530366
rect 175831 530329 175905 530338
rect 175614 530314 175762 530320
rect 175538 530256 175549 530290
rect 175583 530256 175589 530290
rect 175538 530232 175589 530256
rect 175538 530198 175555 530232
rect 175538 530164 175589 530198
rect 175538 530130 175555 530164
rect 175538 530114 175589 530130
rect 175623 530196 175684 530280
rect 175623 530162 175639 530196
rect 175673 530162 175684 530196
rect 175728 530196 175762 530314
rect 175831 530298 175939 530329
rect 176053 530316 176087 530472
rect 176006 530282 176087 530316
rect 176121 530374 176191 530438
rect 176121 530358 176129 530374
rect 176163 530340 176191 530374
rect 176155 530324 176191 530340
rect 176121 530314 176191 530324
rect 176225 530422 176267 530438
rect 176259 530388 176267 530422
rect 176006 530264 176040 530282
rect 176225 530280 176267 530388
rect 175796 530230 175812 530264
rect 175846 530230 176040 530264
rect 176132 530248 176267 530280
rect 175728 530162 175888 530196
rect 175623 530128 175684 530162
rect 175854 530154 175888 530162
rect 175349 530086 175411 530102
rect 175623 530094 175639 530128
rect 175673 530094 175684 530128
rect 175623 530052 175684 530094
rect 175752 530094 175768 530128
rect 175802 530094 175818 530128
rect 176006 530154 176040 530230
rect 176074 530214 176090 530248
rect 176124 530246 176267 530248
rect 176305 530412 176357 530490
rect 176399 530520 176465 530562
rect 176399 530486 176415 530520
rect 176449 530486 176465 530520
rect 176985 530524 177051 530562
rect 176399 530470 176465 530486
rect 176640 530484 176761 530518
rect 176795 530484 176811 530518
rect 176852 530484 176868 530518
rect 176902 530484 176951 530518
rect 176985 530490 177001 530524
rect 177035 530490 177051 530524
rect 177191 530520 177257 530562
rect 177123 530494 177157 530510
rect 176305 530274 176339 530412
rect 176441 530410 176493 530426
rect 176373 530362 176407 530378
rect 176441 530376 176469 530410
rect 176527 530392 176565 530426
rect 176503 530376 176599 530392
rect 176640 530342 176674 530484
rect 176708 530416 176779 530426
rect 176708 530382 176724 530416
rect 176758 530382 176779 530416
rect 176407 530328 176711 530342
rect 176373 530308 176711 530328
rect 176124 530222 176166 530246
rect 176074 530188 176121 530214
rect 176155 530188 176166 530222
rect 176305 530240 176555 530274
rect 176589 530240 176605 530274
rect 176305 530212 176339 530240
rect 176227 530178 176339 530212
rect 175854 530104 175888 530120
rect 175922 530128 175972 530144
rect 175752 530052 175818 530094
rect 175922 530094 175938 530128
rect 175922 530052 175972 530094
rect 176006 530129 176180 530154
rect 176006 530095 176130 530129
rect 176164 530095 176180 530129
rect 176006 530086 176180 530095
rect 176227 530136 176261 530178
rect 176428 530172 176643 530206
rect 176428 530154 176462 530172
rect 176227 530086 176261 530102
rect 176295 530128 176369 530144
rect 176295 530094 176315 530128
rect 176349 530094 176369 530128
rect 176609 530154 176643 530172
rect 176428 530104 176462 530120
rect 176496 530104 176512 530138
rect 176546 530104 176562 530138
rect 176609 530104 176643 530120
rect 176677 530152 176711 530308
rect 176745 530264 176779 530382
rect 176813 530410 176883 530426
rect 176813 530376 176826 530410
rect 176860 530376 176883 530410
rect 176813 530358 176883 530376
rect 176813 530324 176837 530358
rect 176871 530324 176883 530358
rect 176813 530302 176883 530324
rect 176745 530248 176838 530264
rect 176745 530222 176804 530248
rect 176779 530214 176804 530222
rect 176779 530188 176838 530214
rect 176917 530212 176951 530484
rect 177191 530486 177207 530520
rect 177241 530486 177257 530520
rect 177291 530494 177342 530510
rect 176985 530303 177077 530456
rect 177019 530290 177077 530303
rect 177019 530269 177021 530290
rect 176985 530256 177021 530269
rect 177055 530256 177077 530290
rect 176985 530246 177077 530256
rect 176745 530186 176838 530188
rect 176872 530178 176951 530212
rect 176872 530152 176906 530178
rect 176677 530130 176813 530152
rect 176295 530052 176369 530094
rect 176496 530052 176562 530104
rect 176677 530096 176763 530130
rect 176797 530096 176813 530130
rect 176677 530086 176813 530096
rect 176856 530136 176906 530152
rect 176890 530102 176906 530136
rect 176856 530086 176906 530102
rect 176940 530128 176990 530144
rect 176974 530094 176990 530128
rect 176940 530052 176990 530094
rect 177024 530089 177089 530246
rect 177123 530222 177157 530460
rect 177325 530460 177342 530494
rect 177291 530452 177342 530460
rect 177192 530418 177342 530452
rect 177377 530468 177435 530562
rect 177377 530434 177389 530468
rect 177423 530434 177435 530468
rect 177192 530358 177238 530418
rect 177377 530417 177435 530434
rect 177653 530494 177730 530528
rect 177653 530460 177690 530494
rect 177724 530460 177730 530494
rect 177764 530520 177829 530562
rect 177764 530486 177780 530520
rect 177814 530486 177829 530520
rect 177764 530470 177829 530486
rect 177933 530494 177989 530528
rect 177653 530414 177730 530460
rect 177933 530460 177939 530494
rect 177973 530460 177989 530494
rect 177933 530436 177989 530460
rect 177192 530349 177204 530358
rect 177226 530315 177238 530324
rect 177192 530220 177238 530315
rect 177272 530364 177342 530384
rect 177272 530330 177294 530364
rect 177328 530330 177342 530364
rect 177272 530290 177342 530330
rect 177272 530256 177297 530290
rect 177331 530256 177342 530290
rect 177272 530254 177342 530256
rect 177377 530250 177435 530285
rect 177192 530204 177342 530220
rect 177192 530186 177291 530204
rect 177123 530136 177157 530170
rect 177325 530170 177342 530204
rect 177123 530086 177157 530102
rect 177191 530118 177207 530152
rect 177241 530118 177257 530152
rect 177191 530052 177257 530118
rect 177291 530136 177342 530170
rect 177325 530102 177342 530136
rect 177291 530086 177342 530102
rect 177377 530216 177389 530250
rect 177423 530216 177435 530250
rect 177377 530157 177435 530216
rect 177377 530123 177389 530157
rect 177423 530123 177435 530157
rect 177377 530052 177435 530123
rect 177653 530280 177709 530414
rect 177764 530402 177989 530436
rect 178027 530494 178107 530528
rect 178027 530460 178043 530494
rect 178077 530460 178107 530494
rect 178187 530520 178241 530562
rect 178187 530486 178197 530520
rect 178231 530486 178241 530520
rect 178187 530470 178241 530486
rect 178275 530494 178332 530528
rect 177764 530380 177854 530402
rect 177743 530364 177854 530380
rect 178027 530368 178107 530460
rect 178275 530460 178281 530494
rect 178315 530460 178332 530494
rect 178275 530436 178332 530460
rect 177777 530330 177854 530364
rect 177743 530314 177854 530330
rect 177653 530154 177730 530280
rect 177764 530222 177854 530314
rect 177888 530364 178107 530368
rect 177888 530330 177939 530364
rect 177973 530330 178107 530364
rect 177888 530256 178107 530330
rect 177764 530178 177989 530222
rect 177653 530120 177665 530154
rect 177724 530120 177730 530154
rect 177933 530154 177989 530178
rect 177653 530086 177730 530120
rect 177764 530128 177829 530144
rect 177764 530094 177780 530128
rect 177814 530094 177829 530128
rect 177764 530052 177829 530094
rect 177933 530120 177939 530154
rect 177973 530120 177989 530154
rect 177933 530086 177989 530120
rect 178027 530154 178107 530256
rect 178141 530402 178332 530436
rect 178389 530490 178441 530528
rect 178389 530456 178407 530490
rect 178477 530520 178543 530562
rect 178477 530486 178493 530520
rect 178527 530486 178543 530520
rect 178579 530507 178613 530528
rect 178389 530427 178441 530456
rect 178579 530452 178613 530473
rect 178677 530516 178733 530562
rect 178677 530482 178690 530516
rect 178724 530482 178733 530516
rect 178854 530516 178905 530562
rect 178677 530466 178733 530482
rect 178767 530494 178819 530510
rect 178141 530364 178183 530402
rect 178141 530330 178143 530364
rect 178177 530330 178183 530364
rect 178141 530222 178183 530330
rect 178217 530364 178355 530368
rect 178217 530330 178257 530364
rect 178291 530330 178355 530364
rect 178217 530290 178355 530330
rect 178251 530256 178355 530290
rect 178389 530267 178423 530427
rect 178480 530418 178613 530452
rect 178767 530460 178769 530494
rect 178810 530460 178819 530494
rect 178854 530482 178862 530516
rect 178896 530482 178905 530516
rect 179034 530516 179089 530562
rect 178854 530466 178905 530482
rect 178939 530494 178998 530510
rect 178767 530432 178819 530460
rect 178939 530460 178948 530494
rect 178982 530460 178998 530494
rect 179034 530482 179045 530516
rect 179079 530482 179089 530516
rect 179034 530466 179089 530482
rect 179123 530512 179183 530528
rect 179123 530478 179131 530512
rect 179165 530478 179183 530512
rect 179123 530462 179183 530478
rect 178939 530432 178998 530460
rect 178480 530367 178514 530418
rect 178668 530398 178998 530432
rect 178457 530351 178514 530367
rect 178491 530317 178514 530351
rect 178457 530301 178514 530317
rect 178561 530364 178627 530382
rect 178561 530330 178577 530364
rect 178611 530358 178627 530364
rect 178561 530324 178585 530330
rect 178619 530324 178627 530358
rect 178561 530308 178627 530324
rect 178480 530272 178514 530301
rect 178668 530296 178749 530398
rect 179045 530364 179115 530428
rect 178783 530330 178799 530364
rect 178833 530330 178867 530364
rect 178901 530330 178935 530364
rect 178969 530330 179011 530364
rect 178668 530272 178819 530296
rect 178141 530178 178332 530222
rect 178027 530120 178043 530154
rect 178077 530120 178107 530154
rect 178275 530154 178332 530178
rect 178027 530086 178107 530120
rect 178187 530128 178241 530144
rect 178187 530094 178197 530128
rect 178231 530094 178241 530128
rect 178187 530052 178241 530094
rect 178275 530120 178281 530154
rect 178315 530120 178332 530154
rect 178275 530086 178332 530120
rect 178389 530217 178443 530267
rect 178480 530238 178613 530272
rect 178668 530262 178777 530272
rect 178389 530183 178407 530217
rect 178441 530183 178443 530217
rect 178579 530204 178613 530238
rect 178767 530238 178777 530262
rect 178811 530238 178819 530272
rect 178977 530280 179011 530330
rect 179045 530358 179081 530364
rect 179079 530330 179081 530358
rect 179079 530324 179115 530330
rect 179045 530314 179115 530324
rect 179149 530280 179183 530462
rect 178977 530258 179183 530280
rect 178977 530246 179131 530258
rect 178389 530154 178443 530183
rect 178389 530120 178401 530154
rect 178435 530136 178443 530154
rect 178389 530102 178407 530120
rect 178441 530102 178443 530136
rect 178389 530086 178443 530102
rect 178477 530170 178493 530204
rect 178527 530170 178543 530204
rect 178477 530136 178543 530170
rect 178477 530102 178493 530136
rect 178527 530102 178543 530136
rect 178477 530052 178543 530102
rect 178579 530136 178613 530170
rect 178579 530086 178613 530102
rect 178676 530210 178733 530226
rect 178676 530176 178691 530210
rect 178725 530176 178733 530210
rect 178676 530142 178733 530176
rect 178676 530108 178691 530142
rect 178725 530108 178733 530142
rect 178676 530052 178733 530108
rect 178767 530212 178819 530238
rect 179121 530224 179131 530246
rect 179165 530224 179183 530258
rect 178767 530204 178991 530212
rect 178767 530170 178777 530204
rect 178811 530178 178991 530204
rect 178811 530170 178819 530178
rect 178767 530136 178819 530170
rect 178939 530163 178991 530178
rect 178767 530102 178777 530136
rect 178811 530102 178819 530136
rect 178767 530086 178819 530102
rect 178854 530128 178905 530144
rect 178854 530094 178863 530128
rect 178897 530094 178905 530128
rect 178854 530052 178905 530094
rect 178939 530129 178949 530163
rect 178983 530129 178991 530163
rect 178939 530086 178991 530129
rect 179025 530196 179087 530212
rect 179025 530162 179045 530196
rect 179079 530162 179087 530196
rect 179025 530128 179087 530162
rect 179025 530094 179045 530128
rect 179079 530094 179087 530128
rect 179025 530052 179087 530094
rect 179121 530136 179183 530224
rect 179121 530102 179131 530136
rect 179165 530102 179183 530136
rect 179121 530086 179183 530102
rect 179217 530512 179277 530528
rect 179217 530478 179235 530512
rect 179269 530478 179277 530512
rect 179217 530462 179277 530478
rect 179311 530516 179366 530562
rect 179311 530482 179321 530516
rect 179355 530482 179366 530516
rect 179495 530516 179546 530562
rect 179311 530466 179366 530482
rect 179402 530494 179461 530510
rect 179217 530280 179251 530462
rect 179402 530460 179413 530494
rect 179452 530460 179461 530494
rect 179495 530482 179504 530516
rect 179538 530482 179546 530516
rect 179667 530516 179723 530562
rect 179495 530466 179546 530482
rect 179581 530494 179633 530510
rect 179402 530432 179461 530460
rect 179581 530460 179590 530494
rect 179624 530460 179633 530494
rect 179667 530482 179676 530516
rect 179710 530482 179723 530516
rect 179667 530466 179723 530482
rect 179953 530468 180011 530562
rect 179581 530432 179633 530460
rect 179953 530434 179965 530468
rect 179999 530434 180011 530468
rect 179285 530364 179355 530428
rect 179402 530398 179732 530432
rect 179953 530417 180011 530434
rect 180230 530501 180281 530528
rect 180230 530467 180247 530501
rect 180315 530520 180381 530562
rect 180315 530486 180331 530520
rect 180365 530486 180381 530520
rect 180315 530482 180381 530486
rect 180466 530505 180572 530528
rect 179319 530358 179355 530364
rect 179319 530330 179321 530358
rect 179285 530324 179321 530330
rect 179285 530314 179355 530324
rect 179389 530330 179431 530364
rect 179465 530330 179499 530364
rect 179533 530330 179567 530364
rect 179601 530330 179617 530364
rect 179389 530280 179423 530330
rect 179651 530296 179732 530398
rect 179217 530258 179423 530280
rect 179217 530224 179235 530258
rect 179269 530246 179423 530258
rect 179581 530272 179732 530296
rect 180230 530414 180281 530467
rect 180466 530471 180538 530505
rect 180466 530455 180572 530471
rect 180466 530448 180501 530455
rect 180315 530414 180501 530448
rect 179269 530224 179279 530246
rect 179217 530136 179279 530224
rect 179581 530238 179589 530272
rect 179623 530262 179732 530272
rect 179623 530238 179633 530262
rect 179581 530212 179633 530238
rect 179953 530250 180011 530285
rect 179217 530102 179235 530136
rect 179269 530102 179279 530136
rect 179217 530086 179279 530102
rect 179313 530196 179375 530212
rect 179313 530162 179321 530196
rect 179355 530162 179375 530196
rect 179313 530128 179375 530162
rect 179313 530094 179321 530128
rect 179355 530094 179375 530128
rect 179313 530052 179375 530094
rect 179409 530204 179633 530212
rect 179409 530178 179589 530204
rect 179409 530163 179461 530178
rect 179409 530129 179417 530163
rect 179451 530129 179461 530163
rect 179581 530170 179589 530178
rect 179623 530170 179633 530204
rect 179409 530086 179461 530129
rect 179495 530128 179546 530144
rect 179495 530094 179503 530128
rect 179537 530094 179546 530128
rect 179495 530052 179546 530094
rect 179581 530136 179633 530170
rect 179581 530102 179589 530136
rect 179623 530102 179633 530136
rect 179581 530086 179633 530102
rect 179667 530210 179724 530226
rect 179667 530176 179675 530210
rect 179709 530176 179724 530210
rect 179667 530142 179724 530176
rect 179667 530108 179675 530142
rect 179709 530108 179724 530142
rect 179667 530052 179724 530108
rect 179953 530216 179965 530250
rect 179999 530216 180011 530250
rect 179953 530157 180011 530216
rect 179953 530123 179965 530157
rect 179999 530123 180011 530157
rect 179953 530052 180011 530123
rect 180230 530280 180264 530414
rect 180315 530380 180349 530414
rect 180298 530364 180349 530380
rect 180332 530330 180349 530364
rect 180298 530314 180349 530330
rect 180394 530364 180433 530380
rect 180428 530330 180433 530364
rect 180394 530314 180433 530330
rect 180230 530264 180297 530280
rect 180230 530230 180247 530264
rect 180281 530230 180297 530264
rect 180230 530196 180297 530230
rect 180230 530162 180247 530196
rect 180281 530162 180297 530196
rect 180230 530154 180297 530162
rect 180230 530120 180241 530154
rect 180275 530128 180297 530154
rect 180230 530094 180247 530120
rect 180281 530094 180297 530128
rect 180230 530086 180297 530094
rect 180331 530264 180365 530280
rect 180331 530196 180365 530230
rect 180331 530128 180365 530162
rect 180331 530052 180365 530094
rect 180399 530120 180433 530314
rect 180467 530188 180501 530414
rect 180535 530400 180569 530416
rect 180535 530256 180569 530366
rect 180610 530400 180665 530528
rect 180610 530366 180631 530400
rect 180610 530358 180665 530366
rect 180643 530324 180665 530358
rect 180610 530296 180665 530324
rect 180699 530494 180737 530528
rect 180699 530460 180701 530494
rect 180735 530460 180737 530494
rect 180699 530287 180737 530460
rect 180773 530505 180875 530562
rect 180807 530471 180841 530505
rect 180773 530455 180875 530471
rect 180919 530505 180968 530521
rect 180919 530471 180925 530505
rect 180959 530471 180968 530505
rect 180919 530400 180968 530471
rect 181204 530505 181253 530521
rect 181204 530471 181213 530505
rect 181247 530471 181253 530505
rect 181204 530400 181253 530471
rect 181297 530505 181399 530562
rect 181331 530471 181365 530505
rect 181297 530455 181399 530471
rect 180777 530366 180793 530400
rect 180827 530366 181023 530400
rect 180699 530256 180703 530287
rect 180535 530253 180703 530256
rect 180535 530222 180737 530253
rect 180771 530290 180921 530291
rect 180771 530256 180793 530290
rect 180827 530287 180921 530290
rect 180827 530256 180871 530287
rect 180771 530253 180871 530256
rect 180905 530253 180921 530287
rect 180467 530154 180567 530188
rect 180601 530154 180642 530188
rect 180676 530154 180692 530188
rect 180771 530120 180805 530253
rect 180955 530204 181023 530366
rect 180399 530086 180805 530120
rect 180839 530188 180873 530204
rect 180839 530052 180873 530154
rect 180920 530188 181023 530204
rect 180920 530154 180925 530188
rect 180959 530154 181023 530188
rect 180920 530122 181023 530154
rect 181149 530366 181345 530400
rect 181379 530366 181395 530400
rect 181149 530204 181217 530366
rect 181251 530290 181401 530291
rect 181251 530256 181253 530290
rect 181287 530287 181401 530290
rect 181251 530253 181267 530256
rect 181301 530253 181401 530287
rect 181149 530188 181252 530204
rect 181149 530154 181213 530188
rect 181247 530154 181252 530188
rect 181149 530122 181252 530154
rect 181299 530188 181333 530204
rect 181299 530052 181333 530154
rect 181367 530120 181401 530253
rect 181435 530290 181473 530528
rect 181507 530400 181562 530528
rect 181600 530505 181706 530528
rect 181634 530471 181706 530505
rect 181791 530520 181857 530562
rect 181791 530486 181807 530520
rect 181841 530486 181857 530520
rect 181791 530482 181857 530486
rect 181891 530501 181942 530528
rect 181600 530455 181706 530471
rect 181671 530448 181706 530455
rect 181925 530467 181942 530501
rect 181541 530366 181562 530400
rect 181507 530358 181562 530366
rect 181603 530400 181637 530416
rect 181507 530324 181529 530358
rect 181507 530296 181562 530324
rect 181435 530287 181437 530290
rect 181471 530256 181473 530290
rect 181603 530256 181637 530366
rect 181469 530253 181637 530256
rect 181435 530222 181637 530253
rect 181671 530414 181857 530448
rect 181891 530414 181942 530467
rect 181671 530188 181705 530414
rect 181823 530380 181857 530414
rect 181480 530154 181496 530188
rect 181530 530154 181571 530188
rect 181605 530154 181705 530188
rect 181739 530364 181778 530380
rect 181739 530330 181744 530364
rect 181739 530314 181778 530330
rect 181823 530364 181874 530380
rect 181823 530330 181840 530364
rect 181823 530314 181874 530330
rect 181739 530120 181773 530314
rect 181908 530280 181942 530414
rect 181367 530086 181773 530120
rect 181807 530264 181841 530280
rect 181807 530196 181841 530230
rect 181807 530128 181841 530162
rect 181807 530052 181841 530094
rect 181875 530264 181942 530280
rect 181875 530230 181891 530264
rect 181925 530230 181942 530264
rect 181875 530222 181942 530230
rect 181875 530196 181897 530222
rect 181875 530162 181891 530196
rect 181931 530188 181942 530222
rect 181925 530162 181942 530188
rect 181875 530128 181942 530162
rect 181875 530094 181891 530128
rect 181925 530094 181942 530128
rect 181875 530086 181942 530094
rect 181977 530512 182037 530528
rect 181977 530478 181995 530512
rect 182029 530478 182037 530512
rect 181977 530462 182037 530478
rect 182071 530516 182126 530562
rect 182071 530482 182081 530516
rect 182115 530482 182126 530516
rect 182255 530516 182306 530562
rect 182071 530466 182126 530482
rect 182162 530494 182221 530510
rect 181977 530280 182011 530462
rect 182162 530460 182178 530494
rect 182212 530460 182221 530494
rect 182255 530482 182264 530516
rect 182298 530482 182306 530516
rect 182427 530516 182483 530562
rect 182255 530466 182306 530482
rect 182341 530494 182393 530510
rect 182162 530432 182221 530460
rect 182341 530460 182350 530494
rect 182384 530460 182393 530494
rect 182427 530482 182436 530516
rect 182470 530482 182483 530516
rect 182427 530466 182483 530482
rect 182529 530468 182587 530562
rect 182341 530432 182393 530460
rect 182529 530434 182541 530468
rect 182575 530434 182587 530468
rect 182045 530426 182115 530428
rect 182045 530392 182081 530426
rect 182162 530398 182492 530432
rect 182529 530417 182587 530434
rect 182621 530494 182955 530562
rect 182621 530460 182639 530494
rect 182673 530460 182903 530494
rect 182937 530460 182955 530494
rect 182045 530364 182115 530392
rect 182079 530330 182115 530364
rect 182045 530314 182115 530330
rect 182149 530330 182191 530364
rect 182225 530330 182259 530364
rect 182293 530330 182327 530364
rect 182361 530330 182377 530364
rect 182149 530280 182183 530330
rect 182411 530296 182492 530398
rect 182621 530408 182955 530460
rect 183081 530512 183141 530528
rect 183081 530478 183099 530512
rect 183133 530478 183141 530512
rect 183081 530462 183141 530478
rect 183175 530516 183230 530562
rect 183175 530482 183185 530516
rect 183219 530482 183230 530516
rect 183359 530516 183410 530562
rect 183175 530466 183230 530482
rect 183266 530494 183325 530510
rect 182621 530338 182771 530408
rect 182621 530304 182641 530338
rect 182675 530304 182771 530338
rect 182805 530340 182901 530374
rect 182935 530340 182955 530374
rect 181977 530258 182183 530280
rect 181977 530224 181995 530258
rect 182029 530246 182183 530258
rect 182341 530272 182492 530296
rect 182029 530224 182039 530246
rect 181977 530136 182039 530224
rect 182341 530238 182349 530272
rect 182383 530262 182492 530272
rect 182383 530238 182393 530262
rect 182341 530212 182393 530238
rect 182529 530250 182587 530285
rect 182805 530270 182955 530340
rect 181977 530102 181995 530136
rect 182029 530102 182039 530136
rect 181977 530086 182039 530102
rect 182073 530196 182135 530212
rect 182073 530162 182081 530196
rect 182115 530162 182135 530196
rect 182073 530128 182135 530162
rect 182073 530094 182081 530128
rect 182115 530094 182135 530128
rect 182073 530052 182135 530094
rect 182169 530204 182393 530212
rect 182169 530178 182349 530204
rect 182169 530163 182221 530178
rect 182169 530154 182177 530163
rect 182169 530120 182173 530154
rect 182211 530129 182221 530163
rect 182341 530170 182349 530178
rect 182383 530170 182393 530204
rect 182207 530120 182221 530129
rect 182169 530086 182221 530120
rect 182255 530128 182306 530144
rect 182255 530094 182263 530128
rect 182297 530094 182306 530128
rect 182255 530052 182306 530094
rect 182341 530136 182393 530170
rect 182341 530102 182349 530136
rect 182383 530102 182393 530136
rect 182341 530086 182393 530102
rect 182427 530210 182484 530226
rect 182427 530176 182435 530210
rect 182469 530176 182484 530210
rect 182427 530142 182484 530176
rect 182427 530108 182435 530142
rect 182469 530108 182484 530142
rect 182427 530052 182484 530108
rect 182529 530216 182541 530250
rect 182575 530216 182587 530250
rect 182529 530157 182587 530216
rect 182529 530123 182541 530157
rect 182575 530123 182587 530157
rect 182529 530052 182587 530123
rect 182621 530230 182955 530270
rect 182621 530196 182639 530230
rect 182673 530196 182903 530230
rect 182937 530196 182955 530230
rect 182621 530128 182955 530196
rect 182621 530094 182639 530128
rect 182673 530094 182903 530128
rect 182937 530094 182955 530128
rect 182621 530052 182955 530094
rect 183081 530280 183115 530462
rect 183266 530460 183277 530494
rect 183316 530460 183325 530494
rect 183359 530482 183368 530516
rect 183402 530482 183410 530516
rect 183531 530516 183587 530562
rect 183359 530466 183410 530482
rect 183445 530494 183497 530510
rect 183266 530432 183325 530460
rect 183445 530460 183454 530494
rect 183488 530460 183497 530494
rect 183531 530482 183540 530516
rect 183574 530482 183587 530516
rect 183531 530466 183587 530482
rect 183633 530501 184702 530562
rect 183633 530467 183651 530501
rect 183685 530467 184651 530501
rect 184685 530467 184702 530501
rect 183445 530432 183497 530460
rect 183633 530453 184702 530467
rect 184737 530494 185071 530562
rect 184737 530460 184755 530494
rect 184789 530460 185019 530494
rect 185053 530460 185071 530494
rect 183149 530364 183219 530428
rect 183266 530398 183596 530432
rect 183183 530358 183219 530364
rect 183183 530330 183185 530358
rect 183149 530324 183185 530330
rect 183149 530314 183219 530324
rect 183253 530330 183295 530364
rect 183329 530330 183363 530364
rect 183397 530330 183431 530364
rect 183465 530330 183481 530364
rect 183253 530280 183287 530330
rect 183515 530296 183596 530398
rect 183081 530258 183287 530280
rect 183081 530224 183099 530258
rect 183133 530246 183287 530258
rect 183445 530272 183596 530296
rect 183950 530338 184018 530453
rect 184737 530408 185071 530460
rect 185105 530468 185163 530562
rect 185105 530434 185117 530468
rect 185151 530434 185163 530468
rect 185105 530417 185163 530434
rect 185197 530512 185257 530528
rect 185197 530478 185215 530512
rect 185249 530478 185257 530512
rect 185197 530462 185257 530478
rect 185291 530516 185346 530562
rect 185291 530482 185301 530516
rect 185335 530482 185346 530516
rect 185475 530516 185526 530562
rect 185291 530466 185346 530482
rect 185382 530494 185441 530510
rect 183950 530304 183967 530338
rect 184001 530304 184018 530338
rect 183950 530287 184018 530304
rect 184314 530374 184384 530389
rect 184314 530340 184331 530374
rect 184365 530340 184384 530374
rect 183133 530224 183143 530246
rect 183081 530136 183143 530224
rect 183445 530238 183453 530272
rect 183487 530262 183596 530272
rect 183487 530238 183497 530262
rect 183445 530212 183497 530238
rect 183081 530102 183099 530136
rect 183133 530102 183143 530136
rect 183081 530086 183143 530102
rect 183177 530196 183239 530212
rect 183177 530162 183185 530196
rect 183219 530162 183239 530196
rect 183177 530128 183239 530162
rect 183177 530094 183185 530128
rect 183219 530094 183239 530128
rect 183177 530052 183239 530094
rect 183273 530204 183497 530212
rect 183273 530178 183453 530204
rect 183273 530163 183325 530178
rect 183273 530129 183281 530163
rect 183315 530129 183325 530163
rect 183445 530170 183453 530178
rect 183487 530170 183497 530204
rect 183273 530086 183325 530129
rect 183359 530128 183410 530144
rect 183359 530094 183367 530128
rect 183401 530094 183410 530128
rect 183359 530052 183410 530094
rect 183445 530136 183497 530170
rect 183445 530102 183453 530136
rect 183487 530102 183497 530136
rect 183445 530086 183497 530102
rect 183531 530210 183588 530226
rect 183531 530176 183539 530210
rect 183573 530176 183588 530210
rect 183531 530142 183588 530176
rect 183531 530108 183539 530142
rect 183573 530108 183588 530142
rect 184314 530139 184384 530340
rect 184737 530338 184887 530408
rect 184737 530304 184757 530338
rect 184791 530304 184887 530338
rect 184921 530340 185017 530374
rect 185051 530340 185071 530374
rect 184921 530270 185071 530340
rect 184737 530230 185071 530270
rect 184737 530196 184755 530230
rect 184789 530196 185019 530230
rect 185053 530196 185071 530230
rect 183531 530052 183588 530108
rect 183633 530128 184702 530139
rect 183633 530094 183651 530128
rect 183685 530094 184651 530128
rect 184685 530094 184702 530128
rect 183633 530052 184702 530094
rect 184737 530128 185071 530196
rect 184737 530094 184755 530128
rect 184789 530094 185019 530128
rect 185053 530094 185071 530128
rect 184737 530052 185071 530094
rect 185105 530250 185163 530285
rect 185105 530216 185117 530250
rect 185151 530216 185163 530250
rect 185105 530157 185163 530216
rect 185105 530123 185117 530157
rect 185151 530123 185163 530157
rect 185105 530052 185163 530123
rect 185197 530280 185231 530462
rect 185382 530460 185393 530494
rect 185432 530460 185441 530494
rect 185475 530482 185484 530516
rect 185518 530482 185526 530516
rect 185647 530516 185703 530562
rect 185475 530466 185526 530482
rect 185561 530494 185613 530510
rect 185382 530432 185441 530460
rect 185561 530460 185570 530494
rect 185604 530460 185613 530494
rect 185647 530482 185656 530516
rect 185690 530482 185703 530516
rect 185647 530466 185703 530482
rect 185749 530501 186818 530562
rect 187083 530532 187151 530562
rect 185749 530467 185767 530501
rect 185801 530467 186767 530501
rect 186801 530467 186818 530501
rect 185561 530432 185613 530460
rect 185749 530453 186818 530467
rect 186945 530494 186999 530528
rect 187033 530494 187049 530528
rect 186945 530460 187049 530494
rect 185265 530426 185335 530428
rect 185265 530392 185301 530426
rect 185382 530398 185712 530432
rect 185265 530364 185335 530392
rect 185299 530330 185335 530364
rect 185265 530314 185335 530330
rect 185369 530330 185411 530364
rect 185445 530330 185479 530364
rect 185513 530330 185547 530364
rect 185581 530330 185597 530364
rect 185369 530280 185403 530330
rect 185631 530296 185712 530398
rect 185197 530258 185403 530280
rect 185197 530224 185215 530258
rect 185249 530246 185403 530258
rect 185561 530272 185712 530296
rect 186066 530338 186134 530453
rect 186945 530426 186999 530460
rect 187033 530426 187049 530460
rect 187083 530498 187099 530532
rect 187133 530498 187151 530532
rect 187083 530464 187151 530498
rect 187083 530430 187099 530464
rect 187133 530430 187151 530464
rect 187221 530499 187463 530562
rect 187221 530465 187239 530499
rect 187273 530465 187411 530499
rect 187445 530465 187463 530499
rect 186066 530304 186083 530338
rect 186117 530304 186134 530338
rect 186066 530287 186134 530304
rect 186430 530374 186500 530389
rect 186430 530340 186447 530374
rect 186481 530340 186500 530374
rect 185249 530224 185259 530246
rect 185197 530136 185259 530224
rect 185561 530238 185569 530272
rect 185603 530262 185712 530272
rect 185603 530238 185613 530262
rect 185561 530212 185613 530238
rect 185197 530102 185215 530136
rect 185249 530102 185259 530136
rect 185197 530086 185259 530102
rect 185293 530196 185355 530212
rect 185293 530162 185301 530196
rect 185335 530162 185355 530196
rect 185293 530128 185355 530162
rect 185293 530094 185301 530128
rect 185335 530094 185355 530128
rect 185293 530052 185355 530094
rect 185389 530204 185613 530212
rect 185389 530178 185569 530204
rect 185389 530163 185441 530178
rect 185389 530129 185397 530163
rect 185431 530129 185441 530163
rect 185561 530170 185569 530178
rect 185603 530170 185613 530204
rect 185389 530086 185441 530129
rect 185475 530128 185526 530144
rect 185475 530094 185483 530128
rect 185517 530094 185526 530128
rect 185475 530052 185526 530094
rect 185561 530136 185613 530170
rect 185561 530102 185569 530136
rect 185603 530102 185613 530136
rect 185561 530086 185613 530102
rect 185647 530210 185704 530226
rect 185647 530176 185655 530210
rect 185689 530176 185704 530210
rect 185647 530142 185704 530176
rect 185647 530108 185655 530142
rect 185689 530108 185704 530142
rect 186430 530139 186500 530340
rect 186945 530231 187049 530426
rect 187221 530412 187463 530465
rect 187083 530358 187187 530396
rect 187083 530324 187141 530358
rect 187175 530324 187187 530358
rect 187083 530197 187187 530324
rect 186983 530163 186999 530197
rect 187033 530163 187049 530197
rect 185647 530052 185704 530108
rect 185749 530128 186818 530139
rect 185749 530094 185767 530128
rect 185801 530094 186767 530128
rect 186801 530094 186818 530128
rect 185749 530052 186818 530094
rect 186983 530129 187049 530163
rect 186983 530095 186999 530129
rect 187033 530095 187049 530129
rect 186983 530052 187049 530095
rect 187083 530163 187099 530197
rect 187133 530163 187187 530197
rect 187083 530129 187187 530163
rect 187083 530095 187099 530129
rect 187133 530095 187187 530129
rect 187083 530086 187187 530095
rect 187221 530344 187271 530378
rect 187305 530344 187325 530378
rect 187221 530270 187325 530344
rect 187359 530338 187463 530412
rect 187359 530304 187379 530338
rect 187413 530304 187463 530338
rect 187221 530223 187463 530270
rect 187221 530189 187239 530223
rect 187273 530189 187411 530223
rect 187445 530189 187463 530223
rect 187221 530128 187463 530189
rect 187221 530094 187239 530128
rect 187273 530094 187411 530128
rect 187445 530094 187463 530128
rect 187221 530052 187463 530094
rect 172208 530018 172237 530052
rect 172271 530018 172329 530052
rect 172363 530018 172421 530052
rect 172455 530018 172513 530052
rect 172547 530018 172605 530052
rect 172639 530018 172697 530052
rect 172731 530018 172789 530052
rect 172823 530018 172881 530052
rect 172915 530018 172973 530052
rect 173007 530018 173065 530052
rect 173099 530018 173157 530052
rect 173191 530018 173249 530052
rect 173283 530018 173341 530052
rect 173375 530018 173433 530052
rect 173467 530018 173525 530052
rect 173559 530018 173617 530052
rect 173651 530018 173709 530052
rect 173743 530018 173801 530052
rect 173835 530018 173893 530052
rect 173927 530018 173985 530052
rect 174019 530018 174077 530052
rect 174111 530018 174169 530052
rect 174203 530018 174261 530052
rect 174295 530018 174353 530052
rect 174387 530018 174445 530052
rect 174479 530018 174537 530052
rect 174571 530018 174629 530052
rect 174663 530018 174721 530052
rect 174755 530018 174813 530052
rect 174847 530018 174905 530052
rect 174939 530018 174997 530052
rect 175031 530018 175089 530052
rect 175123 530018 175181 530052
rect 175215 530018 175273 530052
rect 175307 530018 175365 530052
rect 175399 530018 175457 530052
rect 175491 530018 175549 530052
rect 175583 530018 175641 530052
rect 175675 530018 175733 530052
rect 175767 530018 175825 530052
rect 175859 530018 175917 530052
rect 175951 530018 176009 530052
rect 176043 530018 176101 530052
rect 176135 530018 176193 530052
rect 176227 530018 176285 530052
rect 176319 530018 176377 530052
rect 176411 530018 176469 530052
rect 176503 530018 176561 530052
rect 176595 530018 176653 530052
rect 176687 530018 176745 530052
rect 176779 530018 176837 530052
rect 176871 530018 176929 530052
rect 176963 530018 177021 530052
rect 177055 530018 177113 530052
rect 177147 530018 177205 530052
rect 177239 530018 177297 530052
rect 177331 530018 177389 530052
rect 177423 530018 177481 530052
rect 177515 530018 177573 530052
rect 177607 530018 177665 530052
rect 177699 530018 177757 530052
rect 177791 530018 177849 530052
rect 177883 530018 177941 530052
rect 177975 530018 178033 530052
rect 178067 530018 178125 530052
rect 178159 530018 178217 530052
rect 178251 530018 178309 530052
rect 178343 530018 178401 530052
rect 178435 530018 178493 530052
rect 178527 530018 178585 530052
rect 178619 530018 178677 530052
rect 178711 530018 178769 530052
rect 178803 530018 178861 530052
rect 178895 530018 178953 530052
rect 178987 530018 179045 530052
rect 179079 530018 179137 530052
rect 179171 530018 179229 530052
rect 179263 530018 179321 530052
rect 179355 530018 179413 530052
rect 179447 530018 179505 530052
rect 179539 530018 179597 530052
rect 179631 530018 179689 530052
rect 179723 530018 179781 530052
rect 179815 530018 179873 530052
rect 179907 530018 179965 530052
rect 179999 530018 180057 530052
rect 180091 530018 180149 530052
rect 180183 530018 180241 530052
rect 180275 530018 180333 530052
rect 180367 530018 180425 530052
rect 180459 530018 180517 530052
rect 180551 530018 180609 530052
rect 180643 530018 180701 530052
rect 180735 530018 180793 530052
rect 180827 530018 180885 530052
rect 180919 530018 180977 530052
rect 181011 530018 181069 530052
rect 181103 530018 181161 530052
rect 181195 530018 181253 530052
rect 181287 530018 181345 530052
rect 181379 530018 181437 530052
rect 181471 530018 181529 530052
rect 181563 530018 181621 530052
rect 181655 530018 181713 530052
rect 181747 530018 181805 530052
rect 181839 530018 181897 530052
rect 181931 530018 181989 530052
rect 182023 530018 182081 530052
rect 182115 530018 182173 530052
rect 182207 530018 182265 530052
rect 182299 530018 182357 530052
rect 182391 530018 182449 530052
rect 182483 530018 182541 530052
rect 182575 530018 182633 530052
rect 182667 530018 182725 530052
rect 182759 530018 182817 530052
rect 182851 530018 182909 530052
rect 182943 530018 183001 530052
rect 183035 530018 183093 530052
rect 183127 530018 183185 530052
rect 183219 530018 183277 530052
rect 183311 530018 183369 530052
rect 183403 530018 183461 530052
rect 183495 530018 183553 530052
rect 183587 530018 183645 530052
rect 183679 530018 183737 530052
rect 183771 530018 183829 530052
rect 183863 530018 183921 530052
rect 183955 530018 184013 530052
rect 184047 530018 184105 530052
rect 184139 530018 184197 530052
rect 184231 530018 184289 530052
rect 184323 530018 184381 530052
rect 184415 530018 184473 530052
rect 184507 530018 184565 530052
rect 184599 530018 184657 530052
rect 184691 530018 184749 530052
rect 184783 530018 184841 530052
rect 184875 530018 184933 530052
rect 184967 530018 185025 530052
rect 185059 530018 185117 530052
rect 185151 530018 185209 530052
rect 185243 530018 185301 530052
rect 185335 530018 185393 530052
rect 185427 530018 185485 530052
rect 185519 530018 185577 530052
rect 185611 530018 185669 530052
rect 185703 530018 185761 530052
rect 185795 530018 185853 530052
rect 185887 530018 185945 530052
rect 185979 530018 186037 530052
rect 186071 530018 186129 530052
rect 186163 530018 186221 530052
rect 186255 530018 186313 530052
rect 186347 530018 186405 530052
rect 186439 530018 186497 530052
rect 186531 530018 186589 530052
rect 186623 530018 186681 530052
rect 186715 530018 186773 530052
rect 186807 530018 186865 530052
rect 186899 530018 186957 530052
rect 186991 530018 187049 530052
rect 187083 530018 187141 530052
rect 187175 530018 187233 530052
rect 187267 530018 187325 530052
rect 187359 530018 187417 530052
rect 187451 530018 187480 530052
rect 172225 529976 172467 530018
rect 172225 529942 172243 529976
rect 172277 529942 172415 529976
rect 172449 529942 172467 529976
rect 172225 529881 172467 529942
rect 172501 529976 173570 530018
rect 172501 529942 172519 529976
rect 172553 529942 173519 529976
rect 173553 529942 173570 529976
rect 172501 529931 173570 529942
rect 173605 529976 174674 530018
rect 173605 529942 173623 529976
rect 173657 529942 174623 529976
rect 174657 529942 174674 529976
rect 173605 529931 174674 529942
rect 174824 529950 174881 529984
rect 172225 529847 172243 529881
rect 172277 529847 172415 529881
rect 172449 529847 172467 529881
rect 172225 529800 172467 529847
rect 172225 529732 172275 529766
rect 172309 529732 172329 529766
rect 172225 529658 172329 529732
rect 172363 529726 172467 529800
rect 172363 529692 172383 529726
rect 172417 529692 172467 529726
rect 172818 529766 172886 529783
rect 172818 529732 172835 529766
rect 172869 529732 172886 529766
rect 172225 529605 172467 529658
rect 172818 529617 172886 529732
rect 173182 529730 173252 529931
rect 173182 529696 173199 529730
rect 173233 529696 173252 529730
rect 173182 529681 173252 529696
rect 173922 529766 173990 529783
rect 173922 529732 173939 529766
rect 173973 529732 173990 529766
rect 173922 529617 173990 529732
rect 174286 529730 174356 529931
rect 174824 529916 174841 529950
rect 174875 529916 174881 529950
rect 174915 529976 174969 530018
rect 174915 529942 174925 529976
rect 174959 529942 174969 529976
rect 174915 529926 174969 529942
rect 175049 529950 175129 529984
rect 174824 529892 174881 529916
rect 175049 529916 175079 529950
rect 175113 529916 175129 529950
rect 174824 529848 175015 529892
rect 174286 529696 174303 529730
rect 174337 529696 174356 529730
rect 174801 529780 174813 529814
rect 174847 529780 174939 529814
rect 174801 529740 174939 529780
rect 174801 529706 174865 529740
rect 174899 529706 174939 529740
rect 174801 529702 174939 529706
rect 174973 529740 175015 529848
rect 174973 529706 174979 529740
rect 175013 529706 175015 529740
rect 174286 529681 174356 529696
rect 174973 529668 175015 529706
rect 174824 529634 175015 529668
rect 175049 529814 175129 529916
rect 175167 529950 175223 529984
rect 175167 529916 175183 529950
rect 175217 529916 175223 529950
rect 175327 529976 175392 530018
rect 175327 529942 175342 529976
rect 175376 529942 175392 529976
rect 175327 529926 175392 529942
rect 175426 529950 175503 529984
rect 175167 529892 175223 529916
rect 175426 529916 175432 529950
rect 175466 529916 175503 529950
rect 175167 529848 175392 529892
rect 175049 529740 175268 529814
rect 175049 529706 175183 529740
rect 175217 529706 175268 529740
rect 175049 529702 175268 529706
rect 175302 529756 175392 529848
rect 175426 529790 175503 529916
rect 175538 529968 175589 529984
rect 175538 529934 175555 529968
rect 175538 529900 175589 529934
rect 175623 529952 175689 530018
rect 175623 529918 175639 529952
rect 175673 529918 175689 529952
rect 175723 529968 175757 529984
rect 175538 529866 175555 529900
rect 175723 529900 175757 529934
rect 175589 529866 175688 529884
rect 175538 529850 175688 529866
rect 175302 529740 175413 529756
rect 175302 529706 175379 529740
rect 172225 529571 172243 529605
rect 172277 529571 172415 529605
rect 172449 529571 172467 529605
rect 172225 529508 172467 529571
rect 172501 529603 173570 529617
rect 172501 529569 172519 529603
rect 172553 529569 173519 529603
rect 173553 529569 173570 529603
rect 172501 529508 173570 529569
rect 173605 529603 174674 529617
rect 173605 529569 173623 529603
rect 173657 529569 174623 529603
rect 174657 529569 174674 529603
rect 173605 529508 174674 529569
rect 174824 529610 174881 529634
rect 174824 529576 174841 529610
rect 174875 529576 174881 529610
rect 175049 529610 175129 529702
rect 175302 529690 175413 529706
rect 175302 529668 175392 529690
rect 174824 529542 174881 529576
rect 174915 529584 174969 529600
rect 174915 529550 174925 529584
rect 174959 529550 174969 529584
rect 174915 529508 174969 529550
rect 175049 529576 175079 529610
rect 175113 529576 175129 529610
rect 175049 529542 175129 529576
rect 175167 529634 175392 529668
rect 175447 529656 175503 529790
rect 175538 529746 175608 529816
rect 175538 529712 175549 529746
rect 175583 529740 175608 529746
rect 175538 529706 175552 529712
rect 175586 529706 175608 529740
rect 175538 529686 175608 529706
rect 175642 529755 175688 529850
rect 175642 529746 175654 529755
rect 175676 529712 175688 529721
rect 175167 529610 175223 529634
rect 175167 529576 175183 529610
rect 175217 529576 175223 529610
rect 175426 529610 175503 529656
rect 175642 529652 175688 529712
rect 175167 529542 175223 529576
rect 175327 529584 175392 529600
rect 175327 529550 175342 529584
rect 175376 529550 175392 529584
rect 175327 529508 175392 529550
rect 175426 529576 175432 529610
rect 175491 529576 175503 529610
rect 175426 529542 175503 529576
rect 175538 529618 175688 529652
rect 175538 529610 175589 529618
rect 175538 529576 175555 529610
rect 175723 529610 175757 529848
rect 175791 529824 175856 529981
rect 175890 529976 175940 530018
rect 175890 529942 175906 529976
rect 175890 529926 175940 529942
rect 175974 529968 176024 529984
rect 175974 529934 175990 529968
rect 175974 529918 176024 529934
rect 176067 529974 176203 529984
rect 176067 529940 176083 529974
rect 176117 529940 176203 529974
rect 176318 529966 176384 530018
rect 176511 529976 176585 530018
rect 176067 529918 176203 529940
rect 175974 529892 176008 529918
rect 175929 529858 176008 529892
rect 176042 529882 176135 529884
rect 175803 529814 175895 529824
rect 175803 529780 175825 529814
rect 175859 529801 175895 529814
rect 175859 529780 175861 529801
rect 175803 529767 175861 529780
rect 175803 529614 175895 529767
rect 175538 529560 175589 529576
rect 175623 529550 175639 529584
rect 175673 529550 175689 529584
rect 175929 529586 175963 529858
rect 176042 529856 176101 529882
rect 176076 529848 176101 529856
rect 176076 529822 176135 529848
rect 176042 529806 176135 529822
rect 175997 529746 176067 529768
rect 175997 529712 176009 529746
rect 176043 529712 176067 529746
rect 175997 529694 176067 529712
rect 175997 529660 176020 529694
rect 176054 529660 176067 529694
rect 175997 529644 176067 529660
rect 176101 529688 176135 529806
rect 176169 529762 176203 529918
rect 176237 529950 176271 529966
rect 176318 529932 176334 529966
rect 176368 529932 176384 529966
rect 176418 529950 176452 529966
rect 176237 529898 176271 529916
rect 176511 529942 176531 529976
rect 176565 529942 176585 529976
rect 176511 529926 176585 529942
rect 176619 529968 176653 529984
rect 176418 529898 176452 529916
rect 176237 529864 176452 529898
rect 176619 529892 176653 529934
rect 176700 529975 176874 529984
rect 176700 529941 176716 529975
rect 176750 529941 176874 529975
rect 176700 529916 176874 529941
rect 176908 529976 176958 530018
rect 176942 529942 176958 529976
rect 177062 529976 177128 530018
rect 176908 529926 176958 529942
rect 176992 529950 177026 529966
rect 176541 529858 176653 529892
rect 176541 529830 176575 529858
rect 176275 529796 176291 529830
rect 176325 529796 176575 529830
rect 176714 529848 176725 529882
rect 176759 529856 176806 529882
rect 176714 529824 176756 529848
rect 176169 529742 176507 529762
rect 176169 529728 176473 529742
rect 176101 529654 176122 529688
rect 176156 529654 176172 529688
rect 176101 529644 176172 529654
rect 176206 529586 176240 529728
rect 176281 529678 176377 529694
rect 176315 529644 176353 529678
rect 176411 529660 176439 529694
rect 176473 529692 176507 529708
rect 176387 529644 176439 529660
rect 176541 529658 176575 529796
rect 175723 529560 175757 529576
rect 175623 529508 175689 529550
rect 175829 529546 175845 529580
rect 175879 529546 175895 529580
rect 175929 529552 175978 529586
rect 176012 529552 176028 529586
rect 176069 529552 176085 529586
rect 176119 529552 176240 529586
rect 176415 529584 176481 529600
rect 175829 529508 175895 529546
rect 176415 529550 176431 529584
rect 176465 529550 176481 529584
rect 176415 529508 176481 529550
rect 176523 529580 176575 529658
rect 176613 529822 176756 529824
rect 176790 529822 176806 529856
rect 176840 529840 176874 529916
rect 177062 529942 177078 529976
rect 177112 529942 177128 529976
rect 177196 529976 177257 530018
rect 177196 529942 177207 529976
rect 177241 529942 177257 529976
rect 176992 529908 177026 529916
rect 177196 529908 177257 529942
rect 176992 529874 177152 529908
rect 176613 529790 176748 529822
rect 176840 529806 177034 529840
rect 177068 529806 177084 529840
rect 176613 529682 176655 529790
rect 176840 529788 176874 529806
rect 176613 529648 176621 529682
rect 176613 529632 176655 529648
rect 176689 529746 176759 529756
rect 176689 529730 176725 529746
rect 176689 529696 176717 529730
rect 176751 529696 176759 529712
rect 176689 529632 176759 529696
rect 176793 529754 176874 529788
rect 176793 529598 176827 529754
rect 176941 529741 177049 529772
rect 177118 529756 177152 529874
rect 177196 529874 177207 529908
rect 177241 529874 177257 529908
rect 177196 529790 177257 529874
rect 177291 529950 177342 529956
rect 177291 529940 177297 529950
rect 177331 529916 177342 529950
rect 177325 529906 177342 529916
rect 177291 529872 177342 529906
rect 177325 529838 177342 529872
rect 177291 529780 177342 529838
rect 177377 529947 177435 530018
rect 177377 529913 177389 529947
rect 177423 529913 177435 529947
rect 177377 529854 177435 529913
rect 177377 529820 177389 529854
rect 177423 529820 177435 529854
rect 177377 529785 177435 529820
rect 177561 529916 177664 529948
rect 177561 529882 177625 529916
rect 177659 529882 177664 529916
rect 177561 529866 177664 529882
rect 177711 529916 177745 530018
rect 177711 529866 177745 529882
rect 177779 529950 178185 529984
rect 177118 529750 177266 529756
rect 176975 529732 177049 529741
rect 176861 529704 176905 529720
rect 176895 529670 176905 529704
rect 176941 529698 176957 529707
rect 176991 529698 177049 529732
rect 176861 529664 176905 529670
rect 177001 529678 177049 529698
rect 176861 529630 176967 529664
rect 176637 529584 176827 529598
rect 176523 529546 176543 529580
rect 176577 529546 176593 529580
rect 176637 529550 176653 529584
rect 176687 529550 176827 529584
rect 176637 529542 176827 529550
rect 176861 529580 176899 529596
rect 176861 529546 176865 529580
rect 176933 529584 176967 529630
rect 177035 529644 177049 529678
rect 177001 529618 177049 529644
rect 177083 529740 177266 529750
rect 177083 529706 177232 529740
rect 177083 529690 177266 529706
rect 177083 529655 177148 529690
rect 177083 529600 177147 529655
rect 177300 529650 177342 529780
rect 177561 529704 177629 529866
rect 177779 529817 177813 529950
rect 177892 529882 177908 529916
rect 177942 529882 177983 529916
rect 178017 529882 178117 529916
rect 177663 529814 177679 529817
rect 177663 529780 177665 529814
rect 177713 529783 177813 529817
rect 177699 529780 177813 529783
rect 177663 529779 177813 529780
rect 177847 529817 178049 529848
rect 177881 529814 178049 529817
rect 177881 529783 177885 529814
rect 177561 529670 177757 529704
rect 177791 529670 177807 529704
rect 177847 529678 177885 529783
rect 177291 529634 177342 529650
rect 177325 529600 177342 529634
rect 176933 529566 177083 529584
rect 177117 529566 177147 529600
rect 176933 529550 177147 529566
rect 177196 529584 177257 529600
rect 177196 529550 177207 529584
rect 177241 529550 177257 529584
rect 176861 529508 176899 529546
rect 177196 529508 177257 529550
rect 177291 529544 177342 529600
rect 177377 529636 177435 529653
rect 177377 529602 177389 529636
rect 177423 529602 177435 529636
rect 177377 529508 177435 529602
rect 177616 529599 177665 529670
rect 177847 529644 177849 529678
rect 177883 529644 177885 529678
rect 177616 529565 177625 529599
rect 177659 529565 177665 529599
rect 177616 529549 177665 529565
rect 177709 529599 177811 529615
rect 177743 529565 177777 529599
rect 177709 529508 177811 529565
rect 177847 529542 177885 529644
rect 177919 529746 177974 529774
rect 177919 529712 177941 529746
rect 177919 529704 177974 529712
rect 177953 529670 177974 529704
rect 177919 529542 177974 529670
rect 178015 529704 178049 529814
rect 178015 529654 178049 529670
rect 178083 529656 178117 529882
rect 178151 529756 178185 529950
rect 178219 529976 178253 530018
rect 178219 529908 178253 529942
rect 178219 529840 178253 529874
rect 178219 529790 178253 529806
rect 178287 529976 178354 529984
rect 178287 529942 178303 529976
rect 178337 529942 178354 529976
rect 178475 529976 178536 530018
rect 178287 529908 178354 529942
rect 178287 529874 178303 529908
rect 178337 529882 178354 529908
rect 178287 529848 178309 529874
rect 178343 529848 178354 529882
rect 178287 529840 178354 529848
rect 178287 529806 178303 529840
rect 178337 529806 178354 529840
rect 178287 529790 178354 529806
rect 178151 529740 178190 529756
rect 178151 529706 178156 529740
rect 178151 529690 178190 529706
rect 178235 529740 178286 529756
rect 178235 529706 178252 529740
rect 178235 529690 178286 529706
rect 178235 529656 178269 529690
rect 178320 529656 178354 529790
rect 178083 529622 178269 529656
rect 178083 529615 178118 529622
rect 178012 529599 178118 529615
rect 178046 529565 178118 529599
rect 178303 529603 178354 529656
rect 178012 529542 178118 529565
rect 178203 529584 178269 529588
rect 178203 529550 178219 529584
rect 178253 529550 178269 529584
rect 178203 529508 178269 529550
rect 178337 529569 178354 529603
rect 178303 529542 178354 529569
rect 178390 529950 178441 529956
rect 178390 529916 178401 529950
rect 178435 529940 178441 529950
rect 178390 529906 178407 529916
rect 178390 529872 178441 529906
rect 178390 529838 178407 529872
rect 178390 529780 178441 529838
rect 178475 529942 178491 529976
rect 178525 529942 178536 529976
rect 178604 529976 178670 530018
rect 178604 529942 178620 529976
rect 178654 529942 178670 529976
rect 178774 529976 178824 530018
rect 178706 529950 178740 529966
rect 178475 529908 178536 529942
rect 178774 529942 178790 529976
rect 178774 529926 178824 529942
rect 178858 529975 179032 529984
rect 178858 529941 178982 529975
rect 179016 529941 179032 529975
rect 178706 529908 178740 529916
rect 178475 529874 178491 529908
rect 178525 529874 178536 529908
rect 178475 529790 178536 529874
rect 178580 529874 178740 529908
rect 178858 529916 179032 529941
rect 179079 529968 179113 529984
rect 178390 529650 178432 529780
rect 178580 529756 178614 529874
rect 178858 529840 178892 529916
rect 179079 529892 179113 529934
rect 179147 529976 179221 530018
rect 179147 529942 179167 529976
rect 179201 529942 179221 529976
rect 179348 529966 179414 530018
rect 179529 529974 179665 529984
rect 179147 529926 179221 529942
rect 179280 529950 179314 529966
rect 179348 529932 179364 529966
rect 179398 529932 179414 529966
rect 179461 529950 179495 529966
rect 179280 529898 179314 529916
rect 179461 529898 179495 529916
rect 178648 529806 178664 529840
rect 178698 529806 178892 529840
rect 178926 529856 178973 529882
rect 178926 529822 178942 529856
rect 179007 529848 179018 529882
rect 179079 529858 179191 529892
rect 179280 529864 179495 529898
rect 179529 529940 179615 529974
rect 179649 529940 179665 529974
rect 179529 529918 179665 529940
rect 179708 529968 179758 529984
rect 179742 529934 179758 529968
rect 179708 529918 179758 529934
rect 179792 529976 179842 530018
rect 179826 529942 179842 529976
rect 179792 529926 179842 529942
rect 178976 529824 179018 529848
rect 179157 529830 179191 529858
rect 178976 529822 179119 529824
rect 178858 529788 178892 529806
rect 178984 529790 179119 529822
rect 178466 529750 178614 529756
rect 178466 529740 178649 529750
rect 178500 529706 178649 529740
rect 178466 529690 178649 529706
rect 178584 529655 178649 529690
rect 178390 529634 178441 529650
rect 178390 529600 178407 529634
rect 178585 529600 178649 529655
rect 178683 529741 178791 529772
rect 178858 529754 178939 529788
rect 178683 529732 178757 529741
rect 178683 529698 178741 529732
rect 178775 529698 178791 529707
rect 178827 529704 178871 529720
rect 178683 529678 178731 529698
rect 178683 529644 178697 529678
rect 178827 529670 178837 529704
rect 178827 529664 178871 529670
rect 178683 529618 178731 529644
rect 178765 529630 178871 529664
rect 178390 529544 178441 529600
rect 178475 529584 178536 529600
rect 178475 529550 178491 529584
rect 178525 529550 178536 529584
rect 178585 529566 178615 529600
rect 178765 529584 178799 529630
rect 178905 529598 178939 529754
rect 178973 529746 179043 529756
rect 179007 529730 179043 529746
rect 178973 529696 178981 529712
rect 179015 529696 179043 529730
rect 178973 529632 179043 529696
rect 179077 529682 179119 529790
rect 179111 529648 179119 529682
rect 179077 529632 179119 529648
rect 179157 529796 179407 529830
rect 179441 529796 179457 529830
rect 179157 529658 179191 529796
rect 179529 529762 179563 529918
rect 179724 529892 179758 529918
rect 179225 529742 179563 529762
rect 179259 529728 179563 529742
rect 179597 529882 179690 529884
rect 179631 529856 179690 529882
rect 179724 529858 179803 529892
rect 179631 529848 179656 529856
rect 179597 529822 179656 529848
rect 179597 529806 179690 529822
rect 179225 529692 179259 529708
rect 179293 529660 179321 529694
rect 179355 529678 179451 529694
rect 178649 529566 178799 529584
rect 178585 529550 178799 529566
rect 178833 529580 178871 529596
rect 178475 529508 178536 529550
rect 178867 529546 178871 529580
rect 178833 529508 178871 529546
rect 178905 529584 179095 529598
rect 178905 529550 179045 529584
rect 179079 529550 179095 529584
rect 179157 529580 179209 529658
rect 179293 529644 179345 529660
rect 179379 529644 179417 529678
rect 178905 529542 179095 529550
rect 179139 529546 179155 529580
rect 179189 529546 179209 529580
rect 179251 529584 179317 529600
rect 179251 529550 179267 529584
rect 179301 529550 179317 529584
rect 179492 529586 179526 529728
rect 179597 529688 179631 529806
rect 179560 529654 179576 529688
rect 179610 529654 179631 529688
rect 179560 529644 179631 529654
rect 179665 529746 179735 529768
rect 179665 529712 179689 529746
rect 179723 529712 179735 529746
rect 179665 529694 179735 529712
rect 179665 529660 179678 529694
rect 179712 529660 179735 529694
rect 179665 529644 179735 529660
rect 179769 529586 179803 529858
rect 179876 529824 179941 529981
rect 179975 529968 180009 529984
rect 179975 529900 180009 529934
rect 180043 529952 180109 530018
rect 180043 529918 180059 529952
rect 180093 529918 180109 529952
rect 180143 529968 180194 529984
rect 180177 529934 180194 529968
rect 180143 529900 180194 529934
rect 179837 529814 179929 529824
rect 179837 529801 179873 529814
rect 179871 529780 179873 529801
rect 179907 529780 179929 529814
rect 179871 529767 179929 529780
rect 179837 529614 179929 529767
rect 179492 529552 179613 529586
rect 179647 529552 179663 529586
rect 179704 529552 179720 529586
rect 179754 529552 179803 529586
rect 179975 529610 180009 529848
rect 180044 529866 180143 529884
rect 180177 529866 180194 529900
rect 180044 529850 180194 529866
rect 180230 529968 180281 529984
rect 180230 529934 180247 529968
rect 180230 529900 180281 529934
rect 180315 529952 180381 530018
rect 180315 529918 180331 529952
rect 180365 529918 180381 529952
rect 180415 529968 180449 529984
rect 180230 529866 180247 529900
rect 180415 529900 180449 529934
rect 180281 529866 180380 529884
rect 180230 529850 180380 529866
rect 180044 529755 180090 529850
rect 180078 529746 180090 529755
rect 180044 529712 180056 529721
rect 180044 529652 180090 529712
rect 180124 529746 180194 529816
rect 180124 529740 180149 529746
rect 180124 529706 180146 529740
rect 180183 529712 180194 529746
rect 180180 529706 180194 529712
rect 180124 529686 180194 529706
rect 180230 529746 180300 529816
rect 180230 529712 180241 529746
rect 180275 529740 180300 529746
rect 180230 529706 180244 529712
rect 180278 529706 180300 529740
rect 180230 529686 180300 529706
rect 180334 529755 180380 529850
rect 180334 529746 180346 529755
rect 180368 529712 180380 529721
rect 180334 529652 180380 529712
rect 180044 529618 180194 529652
rect 179251 529508 179317 529550
rect 179837 529546 179853 529580
rect 179887 529546 179903 529580
rect 180143 529610 180194 529618
rect 179975 529560 180009 529576
rect 179837 529508 179903 529546
rect 180043 529550 180059 529584
rect 180093 529550 180109 529584
rect 180177 529576 180194 529610
rect 180143 529560 180194 529576
rect 180230 529618 180380 529652
rect 180230 529610 180281 529618
rect 180230 529576 180247 529610
rect 180415 529610 180449 529848
rect 180483 529824 180548 529981
rect 180582 529976 180632 530018
rect 180582 529942 180598 529976
rect 180582 529926 180632 529942
rect 180666 529968 180716 529984
rect 180666 529934 180682 529968
rect 180666 529918 180716 529934
rect 180759 529974 180895 529984
rect 180759 529940 180775 529974
rect 180809 529940 180895 529974
rect 181010 529966 181076 530018
rect 181203 529976 181277 530018
rect 180759 529918 180895 529940
rect 180666 529892 180700 529918
rect 180621 529858 180700 529892
rect 180734 529882 180827 529884
rect 180495 529814 180587 529824
rect 180495 529780 180517 529814
rect 180551 529801 180587 529814
rect 180551 529780 180553 529801
rect 180495 529767 180553 529780
rect 180495 529614 180587 529767
rect 180230 529560 180281 529576
rect 180043 529508 180109 529550
rect 180315 529550 180331 529584
rect 180365 529550 180381 529584
rect 180621 529586 180655 529858
rect 180734 529856 180793 529882
rect 180768 529848 180793 529856
rect 180768 529822 180827 529848
rect 180734 529806 180827 529822
rect 180689 529746 180759 529768
rect 180689 529712 180701 529746
rect 180735 529712 180759 529746
rect 180689 529694 180759 529712
rect 180689 529660 180712 529694
rect 180746 529660 180759 529694
rect 180689 529644 180759 529660
rect 180793 529688 180827 529806
rect 180861 529762 180895 529918
rect 180929 529950 180963 529966
rect 181010 529932 181026 529966
rect 181060 529932 181076 529966
rect 181110 529950 181144 529966
rect 180929 529898 180963 529916
rect 181203 529942 181223 529976
rect 181257 529942 181277 529976
rect 181203 529926 181277 529942
rect 181311 529968 181345 529984
rect 181110 529898 181144 529916
rect 180929 529864 181144 529898
rect 181311 529892 181345 529934
rect 181392 529975 181566 529984
rect 181392 529941 181408 529975
rect 181442 529941 181566 529975
rect 181392 529916 181566 529941
rect 181600 529976 181650 530018
rect 181634 529942 181650 529976
rect 181754 529976 181820 530018
rect 181600 529926 181650 529942
rect 181684 529950 181718 529966
rect 181233 529858 181345 529892
rect 181233 529830 181267 529858
rect 180967 529796 180983 529830
rect 181017 529796 181267 529830
rect 181406 529848 181417 529882
rect 181451 529856 181498 529882
rect 181406 529824 181448 529848
rect 180861 529742 181199 529762
rect 180861 529728 181165 529742
rect 180793 529654 180814 529688
rect 180848 529654 180864 529688
rect 180793 529644 180864 529654
rect 180898 529586 180932 529728
rect 180973 529678 181069 529694
rect 181007 529644 181045 529678
rect 181103 529660 181131 529694
rect 181165 529692 181199 529708
rect 181079 529644 181131 529660
rect 181233 529658 181267 529796
rect 180415 529560 180449 529576
rect 180315 529508 180381 529550
rect 180521 529546 180537 529580
rect 180571 529546 180587 529580
rect 180621 529552 180670 529586
rect 180704 529552 180720 529586
rect 180761 529552 180777 529586
rect 180811 529552 180932 529586
rect 181107 529584 181173 529600
rect 180521 529508 180587 529546
rect 181107 529550 181123 529584
rect 181157 529550 181173 529584
rect 181107 529508 181173 529550
rect 181215 529580 181267 529658
rect 181305 529822 181448 529824
rect 181482 529822 181498 529856
rect 181532 529840 181566 529916
rect 181754 529942 181770 529976
rect 181804 529942 181820 529976
rect 181888 529976 181949 530018
rect 181888 529942 181899 529976
rect 181933 529942 181949 529976
rect 182069 529976 182403 530018
rect 181684 529908 181718 529916
rect 181888 529908 181949 529942
rect 181684 529874 181844 529908
rect 181305 529790 181440 529822
rect 181532 529806 181726 529840
rect 181760 529806 181776 529840
rect 181305 529682 181347 529790
rect 181532 529788 181566 529806
rect 181305 529648 181313 529682
rect 181305 529632 181347 529648
rect 181381 529746 181451 529756
rect 181381 529730 181417 529746
rect 181381 529696 181409 529730
rect 181443 529696 181451 529712
rect 181381 529632 181451 529696
rect 181485 529754 181566 529788
rect 181485 529598 181519 529754
rect 181633 529741 181741 529772
rect 181810 529756 181844 529874
rect 181888 529874 181899 529908
rect 181933 529874 181949 529908
rect 181888 529790 181949 529874
rect 181983 529940 182034 529956
rect 182017 529906 182034 529940
rect 181983 529872 182034 529906
rect 182017 529838 182034 529872
rect 181983 529814 182034 529838
rect 181983 529780 181989 529814
rect 182023 529780 182034 529814
rect 182069 529942 182087 529976
rect 182121 529942 182351 529976
rect 182385 529942 182403 529976
rect 182069 529874 182403 529942
rect 182069 529840 182087 529874
rect 182121 529840 182351 529874
rect 182385 529840 182403 529874
rect 182069 529800 182403 529840
rect 181810 529750 181958 529756
rect 181667 529732 181741 529741
rect 181553 529704 181597 529720
rect 181587 529670 181597 529704
rect 181633 529698 181649 529707
rect 181683 529698 181741 529732
rect 181553 529664 181597 529670
rect 181693 529678 181741 529698
rect 181553 529630 181659 529664
rect 181329 529584 181519 529598
rect 181215 529546 181235 529580
rect 181269 529546 181285 529580
rect 181329 529550 181345 529584
rect 181379 529550 181519 529584
rect 181329 529542 181519 529550
rect 181553 529580 181591 529596
rect 181553 529546 181557 529580
rect 181625 529584 181659 529630
rect 181727 529644 181741 529678
rect 181693 529618 181741 529644
rect 181775 529740 181958 529750
rect 181775 529706 181924 529740
rect 181775 529690 181958 529706
rect 181775 529655 181840 529690
rect 181775 529600 181839 529655
rect 181992 529650 182034 529780
rect 181983 529634 182034 529650
rect 182017 529600 182034 529634
rect 181625 529566 181775 529584
rect 181809 529566 181839 529600
rect 181625 529550 181839 529566
rect 181888 529584 181949 529600
rect 181888 529550 181899 529584
rect 181933 529550 181949 529584
rect 181553 529508 181591 529546
rect 181888 529508 181949 529550
rect 181983 529544 182034 529600
rect 182069 529732 182089 529766
rect 182123 529732 182219 529766
rect 182069 529662 182219 529732
rect 182253 529730 182403 529800
rect 182529 529947 182587 530018
rect 182529 529913 182541 529947
rect 182575 529913 182587 529947
rect 182529 529854 182587 529913
rect 182529 529820 182541 529854
rect 182575 529820 182587 529854
rect 182529 529785 182587 529820
rect 182621 529950 182698 529984
rect 182621 529916 182633 529950
rect 182692 529916 182698 529950
rect 182732 529976 182797 530018
rect 182732 529942 182748 529976
rect 182782 529942 182797 529976
rect 182732 529926 182797 529942
rect 182901 529950 182957 529984
rect 182621 529790 182698 529916
rect 182901 529916 182907 529950
rect 182941 529916 182957 529950
rect 182901 529892 182957 529916
rect 182732 529848 182957 529892
rect 182995 529950 183075 529984
rect 182995 529916 183011 529950
rect 183045 529916 183075 529950
rect 183155 529976 183209 530018
rect 183155 529942 183165 529976
rect 183199 529942 183209 529976
rect 183155 529926 183209 529942
rect 183243 529950 183300 529984
rect 182253 529696 182349 529730
rect 182383 529696 182403 529730
rect 182069 529610 182403 529662
rect 182621 529656 182677 529790
rect 182732 529756 182822 529848
rect 182995 529814 183075 529916
rect 183243 529916 183249 529950
rect 183283 529916 183300 529950
rect 183357 529976 184426 530018
rect 183357 529942 183375 529976
rect 183409 529942 184375 529976
rect 184409 529942 184426 529976
rect 183357 529931 184426 529942
rect 184461 529976 185530 530018
rect 184461 529942 184479 529976
rect 184513 529942 185479 529976
rect 185513 529942 185530 529976
rect 184461 529931 185530 529942
rect 185565 529976 186634 530018
rect 185565 529942 185583 529976
rect 185617 529942 186583 529976
rect 186617 529942 186634 529976
rect 185565 529931 186634 529942
rect 186669 529976 187187 530018
rect 186669 529942 186687 529976
rect 186721 529942 187135 529976
rect 187169 529942 187187 529976
rect 183243 529892 183300 529916
rect 182711 529740 182822 529756
rect 182745 529706 182822 529740
rect 182711 529690 182822 529706
rect 182856 529740 183075 529814
rect 182856 529706 182907 529740
rect 182941 529706 183075 529740
rect 182856 529702 183075 529706
rect 182732 529668 182822 529690
rect 182069 529576 182087 529610
rect 182121 529576 182351 529610
rect 182385 529576 182403 529610
rect 182069 529508 182403 529576
rect 182529 529636 182587 529653
rect 182529 529602 182541 529636
rect 182575 529602 182587 529636
rect 182529 529508 182587 529602
rect 182621 529610 182698 529656
rect 182732 529634 182957 529668
rect 182621 529576 182658 529610
rect 182692 529576 182698 529610
rect 182901 529610 182957 529634
rect 182621 529542 182698 529576
rect 182732 529584 182797 529600
rect 182732 529550 182748 529584
rect 182782 529550 182797 529584
rect 182732 529508 182797 529550
rect 182901 529576 182907 529610
rect 182941 529576 182957 529610
rect 182901 529542 182957 529576
rect 182995 529610 183075 529702
rect 183109 529848 183300 529892
rect 183109 529740 183151 529848
rect 183109 529706 183111 529740
rect 183145 529706 183151 529740
rect 183109 529668 183151 529706
rect 183219 529780 183323 529814
rect 183185 529740 183323 529780
rect 183185 529706 183225 529740
rect 183259 529706 183323 529740
rect 183185 529702 183323 529706
rect 183674 529766 183742 529783
rect 183674 529732 183691 529766
rect 183725 529732 183742 529766
rect 183109 529634 183300 529668
rect 182995 529576 183011 529610
rect 183045 529576 183075 529610
rect 183243 529610 183300 529634
rect 183674 529617 183742 529732
rect 184038 529730 184108 529931
rect 184038 529696 184055 529730
rect 184089 529696 184108 529730
rect 184038 529681 184108 529696
rect 184778 529766 184846 529783
rect 184778 529732 184795 529766
rect 184829 529732 184846 529766
rect 184778 529617 184846 529732
rect 185142 529730 185212 529931
rect 185142 529696 185159 529730
rect 185193 529696 185212 529730
rect 185142 529681 185212 529696
rect 185882 529766 185950 529783
rect 185882 529732 185899 529766
rect 185933 529732 185950 529766
rect 185882 529617 185950 529732
rect 186246 529730 186316 529931
rect 186669 529874 187187 529942
rect 186669 529840 186687 529874
rect 186721 529840 187135 529874
rect 187169 529840 187187 529874
rect 186669 529800 187187 529840
rect 186246 529696 186263 529730
rect 186297 529696 186316 529730
rect 186246 529681 186316 529696
rect 186669 529732 186747 529766
rect 186781 529732 186857 529766
rect 186891 529732 186911 529766
rect 186669 529662 186911 529732
rect 186945 529730 187187 529800
rect 186945 529696 186965 529730
rect 186999 529696 187075 529730
rect 187109 529696 187187 529730
rect 187221 529976 187463 530018
rect 187221 529942 187239 529976
rect 187273 529942 187411 529976
rect 187445 529942 187463 529976
rect 187221 529881 187463 529942
rect 187221 529847 187239 529881
rect 187273 529847 187411 529881
rect 187445 529847 187463 529881
rect 187221 529800 187463 529847
rect 187221 529726 187325 529800
rect 187221 529692 187271 529726
rect 187305 529692 187325 529726
rect 187359 529732 187379 529766
rect 187413 529732 187463 529766
rect 182995 529542 183075 529576
rect 183155 529584 183209 529600
rect 183155 529550 183165 529584
rect 183199 529550 183209 529584
rect 183155 529508 183209 529550
rect 183243 529576 183249 529610
rect 183283 529576 183300 529610
rect 183243 529542 183300 529576
rect 183357 529603 184426 529617
rect 183357 529569 183375 529603
rect 183409 529569 184375 529603
rect 184409 529569 184426 529603
rect 183357 529508 184426 529569
rect 184461 529603 185530 529617
rect 184461 529569 184479 529603
rect 184513 529569 185479 529603
rect 185513 529569 185530 529603
rect 184461 529508 185530 529569
rect 185565 529603 186634 529617
rect 185565 529569 185583 529603
rect 185617 529569 186583 529603
rect 186617 529569 186634 529603
rect 185565 529508 186634 529569
rect 186669 529603 187187 529662
rect 187359 529658 187463 529732
rect 186669 529569 186687 529603
rect 186721 529569 187135 529603
rect 187169 529569 187187 529603
rect 186669 529508 187187 529569
rect 187221 529605 187463 529658
rect 187221 529571 187239 529605
rect 187273 529571 187411 529605
rect 187445 529571 187463 529605
rect 187221 529508 187463 529571
rect 172208 529474 172237 529508
rect 172271 529474 172329 529508
rect 172363 529474 172421 529508
rect 172455 529474 172513 529508
rect 172547 529474 172605 529508
rect 172639 529474 172697 529508
rect 172731 529474 172789 529508
rect 172823 529474 172881 529508
rect 172915 529474 172973 529508
rect 173007 529474 173065 529508
rect 173099 529474 173157 529508
rect 173191 529474 173249 529508
rect 173283 529474 173341 529508
rect 173375 529474 173433 529508
rect 173467 529474 173525 529508
rect 173559 529474 173617 529508
rect 173651 529474 173709 529508
rect 173743 529474 173801 529508
rect 173835 529474 173893 529508
rect 173927 529474 173985 529508
rect 174019 529474 174077 529508
rect 174111 529474 174169 529508
rect 174203 529474 174261 529508
rect 174295 529474 174353 529508
rect 174387 529474 174445 529508
rect 174479 529474 174537 529508
rect 174571 529474 174629 529508
rect 174663 529474 174721 529508
rect 174755 529474 174813 529508
rect 174847 529474 174905 529508
rect 174939 529474 174997 529508
rect 175031 529474 175089 529508
rect 175123 529474 175181 529508
rect 175215 529474 175273 529508
rect 175307 529474 175365 529508
rect 175399 529474 175457 529508
rect 175491 529474 175549 529508
rect 175583 529474 175641 529508
rect 175675 529474 175733 529508
rect 175767 529474 175825 529508
rect 175859 529474 175917 529508
rect 175951 529474 176009 529508
rect 176043 529474 176101 529508
rect 176135 529474 176193 529508
rect 176227 529474 176285 529508
rect 176319 529474 176377 529508
rect 176411 529474 176469 529508
rect 176503 529474 176561 529508
rect 176595 529474 176653 529508
rect 176687 529474 176745 529508
rect 176779 529474 176837 529508
rect 176871 529474 176929 529508
rect 176963 529474 177021 529508
rect 177055 529474 177113 529508
rect 177147 529474 177205 529508
rect 177239 529474 177297 529508
rect 177331 529474 177389 529508
rect 177423 529474 177481 529508
rect 177515 529474 177573 529508
rect 177607 529474 177665 529508
rect 177699 529474 177757 529508
rect 177791 529474 177849 529508
rect 177883 529474 177941 529508
rect 177975 529474 178033 529508
rect 178067 529474 178125 529508
rect 178159 529474 178217 529508
rect 178251 529474 178309 529508
rect 178343 529474 178401 529508
rect 178435 529474 178493 529508
rect 178527 529474 178585 529508
rect 178619 529474 178677 529508
rect 178711 529474 178769 529508
rect 178803 529474 178861 529508
rect 178895 529474 178953 529508
rect 178987 529474 179045 529508
rect 179079 529474 179137 529508
rect 179171 529474 179229 529508
rect 179263 529474 179321 529508
rect 179355 529474 179413 529508
rect 179447 529474 179505 529508
rect 179539 529474 179597 529508
rect 179631 529474 179689 529508
rect 179723 529474 179781 529508
rect 179815 529474 179873 529508
rect 179907 529474 179965 529508
rect 179999 529474 180057 529508
rect 180091 529474 180149 529508
rect 180183 529474 180241 529508
rect 180275 529474 180333 529508
rect 180367 529474 180425 529508
rect 180459 529474 180517 529508
rect 180551 529474 180609 529508
rect 180643 529474 180701 529508
rect 180735 529474 180793 529508
rect 180827 529474 180885 529508
rect 180919 529474 180977 529508
rect 181011 529474 181069 529508
rect 181103 529474 181161 529508
rect 181195 529474 181253 529508
rect 181287 529474 181345 529508
rect 181379 529474 181437 529508
rect 181471 529474 181529 529508
rect 181563 529474 181621 529508
rect 181655 529474 181713 529508
rect 181747 529474 181805 529508
rect 181839 529474 181897 529508
rect 181931 529474 181989 529508
rect 182023 529474 182081 529508
rect 182115 529474 182173 529508
rect 182207 529474 182265 529508
rect 182299 529474 182357 529508
rect 182391 529474 182449 529508
rect 182483 529474 182541 529508
rect 182575 529474 182633 529508
rect 182667 529474 182725 529508
rect 182759 529474 182817 529508
rect 182851 529474 182909 529508
rect 182943 529474 183001 529508
rect 183035 529474 183093 529508
rect 183127 529474 183185 529508
rect 183219 529474 183277 529508
rect 183311 529474 183369 529508
rect 183403 529474 183461 529508
rect 183495 529474 183553 529508
rect 183587 529474 183645 529508
rect 183679 529474 183737 529508
rect 183771 529474 183829 529508
rect 183863 529474 183921 529508
rect 183955 529474 184013 529508
rect 184047 529474 184105 529508
rect 184139 529474 184197 529508
rect 184231 529474 184289 529508
rect 184323 529474 184381 529508
rect 184415 529474 184473 529508
rect 184507 529474 184565 529508
rect 184599 529474 184657 529508
rect 184691 529474 184749 529508
rect 184783 529474 184841 529508
rect 184875 529474 184933 529508
rect 184967 529474 185025 529508
rect 185059 529474 185117 529508
rect 185151 529474 185209 529508
rect 185243 529474 185301 529508
rect 185335 529474 185393 529508
rect 185427 529474 185485 529508
rect 185519 529474 185577 529508
rect 185611 529474 185669 529508
rect 185703 529474 185761 529508
rect 185795 529474 185853 529508
rect 185887 529474 185945 529508
rect 185979 529474 186037 529508
rect 186071 529474 186129 529508
rect 186163 529474 186221 529508
rect 186255 529474 186313 529508
rect 186347 529474 186405 529508
rect 186439 529474 186497 529508
rect 186531 529474 186589 529508
rect 186623 529474 186681 529508
rect 186715 529474 186773 529508
rect 186807 529474 186865 529508
rect 186899 529474 186957 529508
rect 186991 529474 187049 529508
rect 187083 529474 187141 529508
rect 187175 529474 187233 529508
rect 187267 529474 187325 529508
rect 187359 529474 187417 529508
rect 187451 529474 187480 529508
rect 172225 529411 172467 529474
rect 172225 529377 172243 529411
rect 172277 529377 172415 529411
rect 172449 529377 172467 529411
rect 172225 529324 172467 529377
rect 172501 529413 173570 529474
rect 172501 529379 172519 529413
rect 172553 529379 173519 529413
rect 173553 529379 173570 529413
rect 172501 529365 173570 529379
rect 173605 529413 174674 529474
rect 173605 529379 173623 529413
rect 173657 529379 174623 529413
rect 174657 529379 174674 529413
rect 173605 529365 174674 529379
rect 174801 529380 174859 529474
rect 172225 529250 172329 529324
rect 172225 529216 172275 529250
rect 172309 529216 172329 529250
rect 172363 529256 172383 529290
rect 172417 529256 172467 529290
rect 172363 529182 172467 529256
rect 172818 529250 172886 529365
rect 172818 529216 172835 529250
rect 172869 529216 172886 529250
rect 172818 529199 172886 529216
rect 173182 529286 173252 529301
rect 173182 529252 173199 529286
rect 173233 529252 173252 529286
rect 172225 529135 172467 529182
rect 172225 529101 172243 529135
rect 172277 529101 172415 529135
rect 172449 529101 172467 529135
rect 172225 529040 172467 529101
rect 173182 529051 173252 529252
rect 173922 529250 173990 529365
rect 174801 529346 174813 529380
rect 174847 529346 174859 529380
rect 174801 529329 174859 529346
rect 175132 529417 175181 529433
rect 175132 529383 175141 529417
rect 175175 529383 175181 529417
rect 175132 529312 175181 529383
rect 175225 529417 175327 529474
rect 175259 529383 175293 529417
rect 175225 529367 175327 529383
rect 175363 529406 175401 529440
rect 175363 529372 175365 529406
rect 175399 529372 175401 529406
rect 173922 529216 173939 529250
rect 173973 529216 173990 529250
rect 173922 529199 173990 529216
rect 174286 529286 174356 529301
rect 174286 529252 174303 529286
rect 174337 529252 174356 529286
rect 174286 529051 174356 529252
rect 175077 529278 175273 529312
rect 175307 529278 175323 529312
rect 174801 529162 174859 529197
rect 174801 529128 174813 529162
rect 174847 529128 174859 529162
rect 174801 529069 174859 529128
rect 172225 529006 172243 529040
rect 172277 529006 172415 529040
rect 172449 529006 172467 529040
rect 172225 528964 172467 529006
rect 172501 529040 173570 529051
rect 172501 529006 172519 529040
rect 172553 529006 173519 529040
rect 173553 529006 173570 529040
rect 172501 528964 173570 529006
rect 173605 529040 174674 529051
rect 173605 529006 173623 529040
rect 173657 529006 174623 529040
rect 174657 529006 174674 529040
rect 173605 528964 174674 529006
rect 174801 529035 174813 529069
rect 174847 529035 174859 529069
rect 174801 528964 174859 529035
rect 175077 529116 175145 529278
rect 175179 529202 175329 529203
rect 175179 529199 175273 529202
rect 175179 529165 175195 529199
rect 175229 529168 175273 529199
rect 175307 529168 175329 529202
rect 175229 529165 175329 529168
rect 175077 529100 175180 529116
rect 175077 529066 175141 529100
rect 175175 529066 175180 529100
rect 175077 529034 175180 529066
rect 175227 529100 175261 529116
rect 175227 528964 175261 529066
rect 175295 529032 175329 529165
rect 175363 529199 175401 529372
rect 175435 529312 175490 529440
rect 175528 529417 175634 529440
rect 175562 529383 175634 529417
rect 175719 529432 175785 529474
rect 175719 529398 175735 529432
rect 175769 529398 175785 529432
rect 175719 529394 175785 529398
rect 175819 529413 175870 529440
rect 175528 529367 175634 529383
rect 175599 529360 175634 529367
rect 175853 529379 175870 529413
rect 175469 529278 175490 529312
rect 175435 529270 175490 529278
rect 175531 529312 175565 529328
rect 175435 529236 175457 529270
rect 175435 529208 175490 529236
rect 175397 529168 175401 529199
rect 175531 529168 175565 529278
rect 175397 529165 175565 529168
rect 175363 529134 175565 529165
rect 175599 529326 175785 529360
rect 175819 529326 175870 529379
rect 175923 529428 175983 529474
rect 175923 529394 175940 529428
rect 175974 529394 175983 529428
rect 175923 529378 175983 529394
rect 176017 529419 176069 529435
rect 176017 529385 176026 529419
rect 176060 529385 176069 529419
rect 176017 529344 176069 529385
rect 176103 529428 176155 529474
rect 176103 529394 176112 529428
rect 176146 529394 176155 529428
rect 176103 529378 176155 529394
rect 176191 529419 176243 529435
rect 176191 529385 176198 529419
rect 176232 529385 176243 529419
rect 176191 529344 176243 529385
rect 176277 529428 176327 529474
rect 176277 529394 176284 529428
rect 176318 529394 176327 529428
rect 176277 529378 176327 529394
rect 176363 529419 176415 529435
rect 176363 529385 176370 529419
rect 176404 529385 176415 529419
rect 176363 529344 176415 529385
rect 176449 529428 176499 529474
rect 176449 529394 176456 529428
rect 176490 529394 176499 529428
rect 176449 529378 176499 529394
rect 176535 529419 176587 529435
rect 176535 529385 176542 529419
rect 176576 529385 176587 529419
rect 176535 529344 176587 529385
rect 176621 529428 176670 529474
rect 176621 529394 176627 529428
rect 176661 529394 176670 529428
rect 176621 529378 176670 529394
rect 176704 529419 176759 529435
rect 176704 529385 176713 529419
rect 176747 529385 176759 529419
rect 176704 529344 176759 529385
rect 176793 529428 176842 529474
rect 176793 529394 176799 529428
rect 176833 529394 176842 529428
rect 176793 529378 176842 529394
rect 176876 529419 176928 529435
rect 176876 529385 176885 529419
rect 176919 529385 176928 529419
rect 176876 529344 176928 529385
rect 176962 529428 177014 529474
rect 176962 529394 176971 529428
rect 177005 529394 177014 529428
rect 176962 529378 177014 529394
rect 177048 529419 177100 529435
rect 177048 529385 177057 529419
rect 177091 529385 177100 529419
rect 177048 529344 177100 529385
rect 177134 529428 177186 529474
rect 177134 529394 177143 529428
rect 177177 529394 177186 529428
rect 177134 529378 177186 529394
rect 177220 529419 177272 529435
rect 177220 529385 177229 529419
rect 177263 529385 177272 529419
rect 177220 529344 177272 529385
rect 177306 529419 177358 529474
rect 177306 529385 177315 529419
rect 177349 529385 177358 529419
rect 177306 529362 177358 529385
rect 177392 529419 177442 529438
rect 177392 529385 177401 529419
rect 177435 529385 177442 529419
rect 175599 529100 175633 529326
rect 175751 529292 175785 529326
rect 175408 529066 175424 529100
rect 175458 529066 175499 529100
rect 175533 529066 175633 529100
rect 175667 529276 175706 529292
rect 175667 529242 175672 529276
rect 175667 529226 175706 529242
rect 175751 529276 175802 529292
rect 175751 529242 175768 529276
rect 175751 529226 175802 529242
rect 175667 529032 175701 529226
rect 175836 529192 175870 529326
rect 175295 528998 175701 529032
rect 175735 529176 175769 529192
rect 175735 529108 175769 529142
rect 175735 529040 175769 529074
rect 175735 528964 175769 529006
rect 175803 529176 175870 529192
rect 175803 529142 175819 529176
rect 175853 529142 175870 529176
rect 175923 529310 177272 529344
rect 175923 529192 176156 529310
rect 177392 529276 177442 529385
rect 177478 529419 177530 529474
rect 177478 529385 177487 529419
rect 177521 529385 177530 529419
rect 177478 529369 177530 529385
rect 177564 529419 177614 529438
rect 177564 529385 177573 529419
rect 177607 529385 177614 529419
rect 177564 529276 177614 529385
rect 177650 529432 177711 529474
rect 177650 529398 177659 529432
rect 177693 529398 177711 529432
rect 177831 529432 177897 529474
rect 177650 529372 177711 529398
rect 177746 529406 177797 529422
rect 177746 529372 177763 529406
rect 177831 529398 177847 529432
rect 177881 529398 177897 529432
rect 178037 529436 178103 529474
rect 177931 529406 177965 529422
rect 177746 529364 177797 529372
rect 178037 529402 178053 529436
rect 178087 529402 178103 529436
rect 178623 529432 178689 529474
rect 176190 529242 176210 529276
rect 176244 529242 176278 529276
rect 176312 529242 176346 529276
rect 176380 529242 176414 529276
rect 176448 529242 176482 529276
rect 176516 529242 176550 529276
rect 176584 529242 176618 529276
rect 176652 529242 176686 529276
rect 176720 529242 176754 529276
rect 176788 529242 176822 529276
rect 176856 529242 176890 529276
rect 176924 529242 176958 529276
rect 176992 529242 177026 529276
rect 177060 529242 177094 529276
rect 177128 529242 177162 529276
rect 177196 529242 177230 529276
rect 177264 529242 177614 529276
rect 176190 529226 177614 529242
rect 177648 529276 177711 529338
rect 177746 529330 177896 529364
rect 177648 529242 177657 529276
rect 177691 529270 177711 529276
rect 177648 529236 177665 529242
rect 177699 529236 177711 529270
rect 177648 529226 177711 529236
rect 177746 529276 177816 529296
rect 177746 529242 177760 529276
rect 177794 529242 177816 529276
rect 175923 529170 177272 529192
rect 175923 529147 176026 529170
rect 175803 529108 175870 529142
rect 176011 529136 176026 529147
rect 176060 529147 176198 529170
rect 176060 529136 176069 529147
rect 175803 529074 175819 529108
rect 175853 529074 175870 529108
rect 175803 529066 175870 529074
rect 175803 529040 175825 529066
rect 175803 529006 175819 529040
rect 175859 529032 175870 529066
rect 175853 529006 175870 529032
rect 175803 528998 175870 529006
rect 175923 529064 175977 529113
rect 175923 529030 175940 529064
rect 175974 529030 175977 529064
rect 175923 528964 175977 529030
rect 176011 529084 176069 529136
rect 176191 529136 176198 529147
rect 176232 529144 176370 529170
rect 176232 529136 176243 529144
rect 176011 529050 176026 529084
rect 176060 529050 176069 529084
rect 176011 528999 176069 529050
rect 176103 529064 176154 529110
rect 176103 529030 176112 529064
rect 176146 529030 176154 529064
rect 176103 528965 176154 529030
rect 176191 529084 176243 529136
rect 176363 529136 176370 529144
rect 176404 529144 176542 529170
rect 176404 529136 176415 529144
rect 176191 529066 176198 529084
rect 176191 529032 176193 529066
rect 176232 529050 176243 529084
rect 176227 529032 176243 529050
rect 176191 528999 176243 529032
rect 176277 529064 176326 529110
rect 176277 529030 176284 529064
rect 176318 529030 176326 529064
rect 176277 528965 176326 529030
rect 176363 529084 176415 529136
rect 176535 529136 176542 529144
rect 176576 529144 176713 529170
rect 176576 529136 176587 529144
rect 176363 529050 176370 529084
rect 176404 529050 176415 529084
rect 176363 528999 176415 529050
rect 176449 529064 176498 529110
rect 176449 529030 176456 529064
rect 176490 529030 176498 529064
rect 176449 528965 176498 529030
rect 176535 529084 176587 529136
rect 176704 529136 176713 529144
rect 176747 529144 176885 529170
rect 176747 529136 176756 529144
rect 176535 529050 176542 529084
rect 176576 529050 176587 529084
rect 176535 528999 176587 529050
rect 176621 529064 176670 529110
rect 176621 529030 176627 529064
rect 176661 529030 176670 529064
rect 176621 528965 176670 529030
rect 176704 529084 176756 529136
rect 176876 529136 176885 529144
rect 176919 529144 177057 529170
rect 176919 529136 176928 529144
rect 176704 529050 176713 529084
rect 176747 529050 176756 529084
rect 176704 528999 176756 529050
rect 176790 529064 176842 529110
rect 176790 529030 176799 529064
rect 176833 529030 176842 529064
rect 176790 528965 176842 529030
rect 176876 529084 176928 529136
rect 177048 529136 177057 529144
rect 177091 529144 177229 529170
rect 177091 529136 177100 529144
rect 176876 529050 176885 529084
rect 176919 529050 176928 529084
rect 176876 528999 176928 529050
rect 176962 529064 177014 529110
rect 176962 529030 176971 529064
rect 177005 529030 177014 529064
rect 176962 528965 177014 529030
rect 177048 529084 177100 529136
rect 177220 529136 177229 529144
rect 177263 529136 177272 529170
rect 177048 529050 177057 529084
rect 177091 529050 177100 529084
rect 177048 528999 177100 529050
rect 177134 529064 177186 529110
rect 177134 529030 177143 529064
rect 177177 529030 177186 529064
rect 177134 528965 177186 529030
rect 177220 529084 177272 529136
rect 177392 529124 177442 529226
rect 177220 529050 177229 529084
rect 177263 529050 177272 529084
rect 177220 528999 177272 529050
rect 177306 529108 177358 529124
rect 177306 529074 177315 529108
rect 177349 529074 177358 529108
rect 177306 529040 177358 529074
rect 177306 529006 177315 529040
rect 177349 529006 177358 529040
rect 177306 528965 177358 529006
rect 177392 529090 177401 529124
rect 177435 529090 177442 529124
rect 177392 529056 177442 529090
rect 177392 529022 177401 529056
rect 177435 529022 177442 529056
rect 177392 528999 177442 529022
rect 177478 529108 177530 529126
rect 177478 529074 177487 529108
rect 177521 529074 177530 529108
rect 177478 529040 177530 529074
rect 177478 529006 177487 529040
rect 177521 529006 177530 529040
rect 176103 528964 177358 528965
rect 177478 528964 177530 529006
rect 177565 529116 177614 529226
rect 177746 529202 177816 529242
rect 177746 529168 177757 529202
rect 177791 529168 177816 529202
rect 177746 529166 177816 529168
rect 177850 529270 177896 529330
rect 177884 529261 177896 529270
rect 177850 529227 177862 529236
rect 177850 529132 177896 529227
rect 177565 529082 177573 529116
rect 177607 529082 177614 529116
rect 177565 529048 177614 529082
rect 177565 529014 177573 529048
rect 177607 529014 177614 529048
rect 177565 528998 177614 529014
rect 177650 529108 177709 529126
rect 177650 529074 177659 529108
rect 177693 529074 177709 529108
rect 177650 529040 177709 529074
rect 177650 529006 177659 529040
rect 177693 529006 177709 529040
rect 177650 528964 177709 529006
rect 177746 529116 177896 529132
rect 177746 529082 177763 529116
rect 177797 529098 177896 529116
rect 177931 529134 177965 529372
rect 178137 529396 178186 529430
rect 178220 529396 178236 529430
rect 178277 529396 178293 529430
rect 178327 529396 178448 529430
rect 178011 529338 178103 529368
rect 178011 529304 178033 529338
rect 178067 529304 178103 529338
rect 178011 529215 178103 529304
rect 178011 529181 178069 529215
rect 178011 529158 178103 529181
rect 177746 529048 177797 529082
rect 177746 529014 177763 529048
rect 177746 528998 177797 529014
rect 177831 529030 177847 529064
rect 177881 529030 177897 529064
rect 177831 528964 177897 529030
rect 177931 529048 177965 529082
rect 177931 528998 177965 529014
rect 177999 529001 178064 529158
rect 178137 529124 178171 529396
rect 178205 529322 178275 529338
rect 178205 529288 178228 529322
rect 178262 529288 178275 529322
rect 178205 529270 178275 529288
rect 178205 529236 178217 529270
rect 178251 529236 178275 529270
rect 178205 529214 178275 529236
rect 178309 529328 178380 529338
rect 178309 529294 178330 529328
rect 178364 529294 178380 529328
rect 178309 529176 178343 529294
rect 178414 529254 178448 529396
rect 178623 529398 178639 529432
rect 178673 529398 178689 529432
rect 178623 529382 178689 529398
rect 178731 529402 178751 529436
rect 178785 529402 178801 529436
rect 178845 529432 179035 529440
rect 178523 529304 178561 529338
rect 178595 529322 178647 529338
rect 178731 529324 178783 529402
rect 178845 529398 178861 529432
rect 178895 529398 179035 529432
rect 178845 529384 179035 529398
rect 179069 529436 179107 529474
rect 179069 529402 179073 529436
rect 179404 529432 179465 529474
rect 179069 529386 179107 529402
rect 179141 529416 179355 529432
rect 179141 529398 179291 529416
rect 178489 529288 178585 529304
rect 178619 529288 178647 529322
rect 178681 529274 178715 529290
rect 178250 529160 178343 529176
rect 178284 529134 178343 529160
rect 178284 529126 178309 529134
rect 178137 529090 178216 529124
rect 178250 529100 178309 529126
rect 178250 529098 178343 529100
rect 178377 529240 178681 529254
rect 178377 529220 178715 529240
rect 178182 529064 178216 529090
rect 178377 529064 178411 529220
rect 178749 529186 178783 529324
rect 178483 529152 178499 529186
rect 178533 529152 178783 529186
rect 178821 529334 178863 529350
rect 178821 529300 178829 529334
rect 178821 529192 178863 529300
rect 178897 529286 178967 529350
rect 178897 529252 178925 529286
rect 178959 529270 178967 529286
rect 178897 529236 178933 529252
rect 178897 529226 178967 529236
rect 179001 529228 179035 529384
rect 179141 529352 179175 529398
rect 179325 529382 179355 529416
rect 179404 529398 179415 529432
rect 179449 529398 179465 529432
rect 179404 529382 179465 529398
rect 179499 529382 179550 529438
rect 179069 529318 179175 529352
rect 179209 529338 179257 529364
rect 179069 529312 179113 529318
rect 179103 529278 179113 529312
rect 179243 529304 179257 529338
rect 179209 529284 179257 529304
rect 179069 529262 179113 529278
rect 179149 529275 179165 529284
rect 179199 529250 179257 529284
rect 179183 529241 179257 529250
rect 179001 529194 179082 529228
rect 179149 529210 179257 529241
rect 179291 529327 179355 529382
rect 179533 529348 179550 529382
rect 179499 529332 179550 529348
rect 179291 529292 179356 529327
rect 179291 529276 179474 529292
rect 179291 529242 179440 529276
rect 179291 529232 179474 529242
rect 179326 529226 179474 529232
rect 178821 529160 178956 529192
rect 179048 529176 179082 529194
rect 178821 529158 178964 529160
rect 178749 529124 178783 529152
rect 178922 529134 178964 529158
rect 178098 529040 178148 529056
rect 178098 529006 178114 529040
rect 178098 528964 178148 529006
rect 178182 529048 178232 529064
rect 178182 529014 178198 529048
rect 178182 528998 178232 529014
rect 178275 529042 178411 529064
rect 178275 529008 178291 529042
rect 178325 529008 178411 529042
rect 178445 529084 178660 529118
rect 178749 529090 178861 529124
rect 178922 529100 178933 529134
rect 178998 529126 179014 529160
rect 178967 529100 179014 529126
rect 179048 529142 179242 529176
rect 179276 529142 179292 529176
rect 178445 529066 178479 529084
rect 178626 529066 178660 529084
rect 178445 529016 178479 529032
rect 178526 529016 178542 529050
rect 178576 529016 178592 529050
rect 178626 529016 178660 529032
rect 178719 529040 178793 529056
rect 178275 528998 178411 529008
rect 178526 528964 178592 529016
rect 178719 529006 178739 529040
rect 178773 529006 178793 529040
rect 178719 528964 178793 529006
rect 178827 529048 178861 529090
rect 179048 529066 179082 529142
rect 179326 529108 179360 529226
rect 179508 529202 179550 529332
rect 179695 529419 179729 529440
rect 179765 529432 179831 529474
rect 179765 529398 179781 529432
rect 179815 529398 179831 529432
rect 179867 529406 179919 529440
rect 179867 529402 179873 529406
rect 179695 529364 179729 529385
rect 179907 529372 179919 529406
rect 179901 529368 179919 529372
rect 179695 529330 179828 529364
rect 179867 529339 179919 529368
rect 179681 529276 179747 529294
rect 179681 529270 179697 529276
rect 179681 529236 179689 529270
rect 179731 529242 179747 529276
rect 179723 529236 179747 529242
rect 179681 529220 179747 529236
rect 179794 529279 179828 529330
rect 179794 529263 179851 529279
rect 179794 529229 179817 529263
rect 178827 528998 178861 529014
rect 178908 529041 179082 529066
rect 179200 529074 179360 529108
rect 179404 529108 179465 529192
rect 179404 529074 179415 529108
rect 179449 529074 179465 529108
rect 179200 529066 179234 529074
rect 178908 529007 178924 529041
rect 178958 529007 179082 529041
rect 178908 528998 179082 529007
rect 179116 529040 179166 529056
rect 179150 529006 179166 529040
rect 179404 529040 179465 529074
rect 179200 529016 179234 529032
rect 179116 528964 179166 529006
rect 179270 529006 179286 529040
rect 179320 529006 179336 529040
rect 179270 528964 179336 529006
rect 179404 529006 179415 529040
rect 179449 529006 179465 529040
rect 179499 529144 179550 529202
rect 179794 529213 179851 529229
rect 179794 529184 179828 529213
rect 179533 529110 179550 529144
rect 179499 529076 179550 529110
rect 179533 529066 179550 529076
rect 179499 529032 179505 529042
rect 179539 529032 179550 529066
rect 179499 529026 179550 529032
rect 179695 529150 179828 529184
rect 179885 529179 179919 529339
rect 179953 529380 180011 529474
rect 179953 529346 179965 529380
rect 179999 529346 180011 529380
rect 179953 529329 180011 529346
rect 180045 529413 180563 529474
rect 180045 529379 180063 529413
rect 180097 529379 180511 529413
rect 180545 529379 180563 529413
rect 180045 529320 180563 529379
rect 180689 529432 180750 529474
rect 180689 529398 180707 529432
rect 180741 529398 180750 529432
rect 180689 529372 180750 529398
rect 180786 529419 180836 529438
rect 180786 529385 180793 529419
rect 180827 529385 180836 529419
rect 180045 529250 180287 529320
rect 180045 529216 180123 529250
rect 180157 529216 180233 529250
rect 180267 529216 180287 529250
rect 180321 529252 180341 529286
rect 180375 529252 180451 529286
rect 180485 529252 180563 529286
rect 179695 529116 179729 529150
rect 179865 529129 179919 529179
rect 179695 529048 179729 529082
rect 179404 528964 179465 529006
rect 179695 528998 179729 529014
rect 179765 529082 179781 529116
rect 179815 529082 179831 529116
rect 179765 529048 179831 529082
rect 179765 529014 179781 529048
rect 179815 529014 179831 529048
rect 179765 528964 179831 529014
rect 179865 529095 179867 529129
rect 179901 529095 179919 529129
rect 179865 529048 179919 529095
rect 179865 529014 179867 529048
rect 179901 529014 179919 529048
rect 179865 528998 179919 529014
rect 179953 529162 180011 529197
rect 180321 529182 180563 529252
rect 180689 529276 180752 529338
rect 180689 529270 180709 529276
rect 180689 529236 180701 529270
rect 180743 529242 180752 529276
rect 180735 529236 180752 529242
rect 180689 529226 180752 529236
rect 180786 529276 180836 529385
rect 180870 529419 180922 529474
rect 180870 529385 180879 529419
rect 180913 529385 180922 529419
rect 180870 529369 180922 529385
rect 180958 529419 181008 529438
rect 180958 529385 180965 529419
rect 180999 529385 181008 529419
rect 180958 529276 181008 529385
rect 181042 529419 181094 529474
rect 181042 529385 181051 529419
rect 181085 529385 181094 529419
rect 181042 529362 181094 529385
rect 181128 529419 181180 529435
rect 181128 529385 181137 529419
rect 181171 529385 181180 529419
rect 181128 529344 181180 529385
rect 181214 529428 181266 529474
rect 181214 529394 181223 529428
rect 181257 529394 181266 529428
rect 181214 529378 181266 529394
rect 181300 529419 181352 529435
rect 181300 529385 181309 529419
rect 181343 529385 181352 529419
rect 181300 529344 181352 529385
rect 181386 529428 181438 529474
rect 181386 529394 181395 529428
rect 181429 529394 181438 529428
rect 181386 529378 181438 529394
rect 181472 529419 181524 529435
rect 181472 529385 181481 529419
rect 181515 529385 181524 529419
rect 181472 529344 181524 529385
rect 181558 529428 181607 529474
rect 181558 529394 181567 529428
rect 181601 529394 181607 529428
rect 181558 529378 181607 529394
rect 181641 529419 181696 529435
rect 181641 529385 181653 529419
rect 181687 529385 181696 529419
rect 181641 529344 181696 529385
rect 181730 529428 181779 529474
rect 181730 529394 181739 529428
rect 181773 529394 181779 529428
rect 181730 529378 181779 529394
rect 181813 529419 181865 529435
rect 181813 529385 181824 529419
rect 181858 529385 181865 529419
rect 181813 529344 181865 529385
rect 181901 529428 181951 529474
rect 181901 529394 181910 529428
rect 181944 529394 181951 529428
rect 181901 529378 181951 529394
rect 181985 529419 182037 529435
rect 181985 529385 181996 529419
rect 182030 529385 182037 529419
rect 181985 529344 182037 529385
rect 182073 529428 182123 529474
rect 182073 529394 182082 529428
rect 182116 529394 182123 529428
rect 182073 529378 182123 529394
rect 182157 529419 182209 529435
rect 182157 529385 182168 529419
rect 182202 529385 182209 529419
rect 182157 529344 182209 529385
rect 182245 529428 182297 529474
rect 182245 529394 182254 529428
rect 182288 529394 182297 529428
rect 182245 529378 182297 529394
rect 182331 529419 182383 529435
rect 182331 529385 182340 529419
rect 182374 529385 182383 529419
rect 182331 529344 182383 529385
rect 182417 529428 182477 529474
rect 182417 529394 182426 529428
rect 182460 529394 182477 529428
rect 182417 529378 182477 529394
rect 182529 529406 182581 529440
rect 182529 529372 182541 529406
rect 182575 529402 182581 529406
rect 182617 529432 182683 529474
rect 182617 529398 182633 529432
rect 182667 529398 182683 529432
rect 182719 529419 182753 529440
rect 182529 529368 182547 529372
rect 181128 529310 182477 529344
rect 180786 529242 181136 529276
rect 181170 529242 181204 529276
rect 181238 529242 181272 529276
rect 181306 529242 181340 529276
rect 181374 529242 181408 529276
rect 181442 529242 181476 529276
rect 181510 529242 181544 529276
rect 181578 529242 181612 529276
rect 181646 529242 181680 529276
rect 181714 529242 181748 529276
rect 181782 529242 181816 529276
rect 181850 529242 181884 529276
rect 181918 529242 181952 529276
rect 181986 529242 182020 529276
rect 182054 529242 182088 529276
rect 182122 529242 182156 529276
rect 182190 529242 182210 529276
rect 180786 529226 182210 529242
rect 179953 529128 179965 529162
rect 179999 529128 180011 529162
rect 179953 529069 180011 529128
rect 179953 529035 179965 529069
rect 179999 529035 180011 529069
rect 179953 528964 180011 529035
rect 180045 529142 180563 529182
rect 180045 529108 180063 529142
rect 180097 529108 180511 529142
rect 180545 529108 180563 529142
rect 180045 529040 180563 529108
rect 180045 529006 180063 529040
rect 180097 529006 180511 529040
rect 180545 529006 180563 529040
rect 180045 528964 180563 529006
rect 180691 529108 180750 529126
rect 180691 529074 180707 529108
rect 180741 529074 180750 529108
rect 180691 529040 180750 529074
rect 180691 529006 180707 529040
rect 180741 529006 180750 529040
rect 180691 528964 180750 529006
rect 180786 529116 180835 529226
rect 180786 529082 180793 529116
rect 180827 529082 180835 529116
rect 180786 529048 180835 529082
rect 180786 529014 180793 529048
rect 180827 529014 180835 529048
rect 180786 528998 180835 529014
rect 180870 529108 180922 529126
rect 180870 529074 180879 529108
rect 180913 529074 180922 529108
rect 180870 529040 180922 529074
rect 180870 529006 180879 529040
rect 180913 529006 180922 529040
rect 180870 528964 180922 529006
rect 180958 529124 181008 529226
rect 182244 529192 182477 529310
rect 181128 529170 182477 529192
rect 181128 529136 181137 529170
rect 181171 529144 181309 529170
rect 181171 529136 181180 529144
rect 180958 529090 180965 529124
rect 180999 529090 181008 529124
rect 180958 529056 181008 529090
rect 180958 529022 180965 529056
rect 180999 529022 181008 529056
rect 180958 528999 181008 529022
rect 181042 529108 181094 529124
rect 181042 529074 181051 529108
rect 181085 529074 181094 529108
rect 181042 529040 181094 529074
rect 181042 529006 181051 529040
rect 181085 529006 181094 529040
rect 181042 528965 181094 529006
rect 181128 529084 181180 529136
rect 181300 529136 181309 529144
rect 181343 529144 181481 529170
rect 181343 529136 181352 529144
rect 181128 529050 181137 529084
rect 181171 529050 181180 529084
rect 181128 528999 181180 529050
rect 181214 529064 181266 529110
rect 181214 529030 181223 529064
rect 181257 529030 181266 529064
rect 181214 528965 181266 529030
rect 181300 529084 181352 529136
rect 181472 529136 181481 529144
rect 181515 529144 181653 529170
rect 181515 529136 181524 529144
rect 181300 529050 181309 529084
rect 181343 529050 181352 529084
rect 181300 528999 181352 529050
rect 181386 529064 181438 529110
rect 181386 529030 181395 529064
rect 181429 529030 181438 529064
rect 181386 528965 181438 529030
rect 181472 529084 181524 529136
rect 181644 529136 181653 529144
rect 181687 529144 181824 529170
rect 181687 529136 181696 529144
rect 181472 529050 181481 529084
rect 181515 529050 181524 529084
rect 181472 528999 181524 529050
rect 181558 529064 181610 529110
rect 181558 529030 181567 529064
rect 181601 529030 181610 529064
rect 181558 528965 181610 529030
rect 181644 529084 181696 529136
rect 181813 529136 181824 529144
rect 181858 529144 181996 529170
rect 181858 529136 181865 529144
rect 181644 529050 181653 529084
rect 181687 529050 181696 529084
rect 181644 528999 181696 529050
rect 181730 529064 181779 529110
rect 181730 529030 181739 529064
rect 181773 529030 181779 529064
rect 181730 528965 181779 529030
rect 181813 529084 181865 529136
rect 181985 529136 181996 529144
rect 182030 529144 182168 529170
rect 182030 529136 182037 529144
rect 181813 529050 181824 529084
rect 181858 529050 181865 529084
rect 181813 528999 181865 529050
rect 181902 529064 181951 529110
rect 181902 529030 181910 529064
rect 181944 529030 181951 529064
rect 181902 528965 181951 529030
rect 181985 529084 182037 529136
rect 182157 529136 182168 529144
rect 182202 529147 182340 529170
rect 182202 529136 182209 529147
rect 181985 529066 181996 529084
rect 181985 529032 181989 529066
rect 182030 529050 182037 529084
rect 182023 529032 182037 529050
rect 181985 528999 182037 529032
rect 182074 529064 182123 529110
rect 182074 529030 182082 529064
rect 182116 529030 182123 529064
rect 182074 528965 182123 529030
rect 182157 529084 182209 529136
rect 182331 529136 182340 529147
rect 182374 529147 182477 529170
rect 182529 529339 182581 529368
rect 182719 529364 182753 529385
rect 182805 529413 183874 529474
rect 182805 529379 182823 529413
rect 182857 529379 183823 529413
rect 183857 529379 183874 529413
rect 182805 529365 183874 529379
rect 183909 529413 184978 529474
rect 183909 529379 183927 529413
rect 183961 529379 184927 529413
rect 184961 529379 184978 529413
rect 183909 529365 184978 529379
rect 185105 529380 185163 529474
rect 182529 529179 182563 529339
rect 182620 529330 182753 529364
rect 182620 529279 182654 529330
rect 182597 529263 182654 529279
rect 182631 529229 182654 529263
rect 182597 529213 182654 529229
rect 182701 529276 182767 529294
rect 182701 529242 182717 529276
rect 182751 529270 182767 529276
rect 182701 529236 182725 529242
rect 182759 529236 182767 529270
rect 182701 529220 182767 529236
rect 183122 529250 183190 529365
rect 182620 529184 182654 529213
rect 183122 529216 183139 529250
rect 183173 529216 183190 529250
rect 183122 529199 183190 529216
rect 183486 529286 183556 529301
rect 183486 529252 183503 529286
rect 183537 529252 183556 529286
rect 182374 529136 182389 529147
rect 182157 529050 182168 529084
rect 182202 529050 182209 529084
rect 182157 528999 182209 529050
rect 182246 529064 182297 529110
rect 182246 529030 182254 529064
rect 182288 529030 182297 529064
rect 182246 528965 182297 529030
rect 182331 529084 182389 529136
rect 182529 529129 182583 529179
rect 182620 529150 182753 529184
rect 182331 529050 182340 529084
rect 182374 529050 182389 529084
rect 182331 528999 182389 529050
rect 182423 529064 182477 529113
rect 182423 529030 182426 529064
rect 182460 529030 182477 529064
rect 181042 528964 182297 528965
rect 182423 528964 182477 529030
rect 182529 529095 182547 529129
rect 182581 529095 182583 529129
rect 182719 529116 182753 529150
rect 182529 529048 182583 529095
rect 182529 529014 182547 529048
rect 182581 529014 182583 529048
rect 182529 528998 182583 529014
rect 182617 529082 182633 529116
rect 182667 529082 182683 529116
rect 182617 529048 182683 529082
rect 182617 529014 182633 529048
rect 182667 529014 182683 529048
rect 182617 528964 182683 529014
rect 182719 529048 182753 529082
rect 183486 529051 183556 529252
rect 184226 529250 184294 529365
rect 185105 529346 185117 529380
rect 185151 529346 185163 529380
rect 185197 529413 186266 529474
rect 185197 529379 185215 529413
rect 185249 529379 186215 529413
rect 186249 529379 186266 529413
rect 185197 529365 186266 529379
rect 186301 529413 187003 529474
rect 186301 529379 186319 529413
rect 186353 529379 186951 529413
rect 186985 529379 187003 529413
rect 185105 529329 185163 529346
rect 184226 529216 184243 529250
rect 184277 529216 184294 529250
rect 184226 529199 184294 529216
rect 184590 529286 184660 529301
rect 184590 529252 184607 529286
rect 184641 529252 184660 529286
rect 184590 529051 184660 529252
rect 185514 529250 185582 529365
rect 186301 529320 187003 529379
rect 187221 529411 187463 529474
rect 187221 529377 187239 529411
rect 187273 529377 187411 529411
rect 187445 529377 187463 529411
rect 187221 529324 187463 529377
rect 185514 529216 185531 529250
rect 185565 529216 185582 529250
rect 185514 529199 185582 529216
rect 185878 529286 185948 529301
rect 185878 529252 185895 529286
rect 185929 529252 185948 529286
rect 185105 529162 185163 529197
rect 185105 529128 185117 529162
rect 185151 529128 185163 529162
rect 185105 529069 185163 529128
rect 182719 528998 182753 529014
rect 182805 529040 183874 529051
rect 182805 529006 182823 529040
rect 182857 529006 183823 529040
rect 183857 529006 183874 529040
rect 182805 528964 183874 529006
rect 183909 529040 184978 529051
rect 183909 529006 183927 529040
rect 183961 529006 184927 529040
rect 184961 529006 184978 529040
rect 183909 528964 184978 529006
rect 185105 529035 185117 529069
rect 185151 529035 185163 529069
rect 185878 529051 185948 529252
rect 186301 529250 186631 529320
rect 186301 529216 186379 529250
rect 186413 529216 186478 529250
rect 186512 529216 186577 529250
rect 186611 529216 186631 529250
rect 186665 529252 186685 529286
rect 186719 529252 186788 529286
rect 186822 529252 186891 529286
rect 186925 529252 187003 529286
rect 186665 529182 187003 529252
rect 186301 529142 187003 529182
rect 186301 529108 186319 529142
rect 186353 529108 186951 529142
rect 186985 529108 187003 529142
rect 185105 528964 185163 529035
rect 185197 529040 186266 529051
rect 185197 529006 185215 529040
rect 185249 529006 186215 529040
rect 186249 529006 186266 529040
rect 185197 528964 186266 529006
rect 186301 529040 187003 529108
rect 186301 529006 186319 529040
rect 186353 529006 186951 529040
rect 186985 529006 187003 529040
rect 186301 528964 187003 529006
rect 187221 529256 187271 529290
rect 187305 529256 187325 529290
rect 187221 529182 187325 529256
rect 187359 529250 187463 529324
rect 187359 529216 187379 529250
rect 187413 529216 187463 529250
rect 187221 529135 187463 529182
rect 187221 529101 187239 529135
rect 187273 529101 187411 529135
rect 187445 529101 187463 529135
rect 187221 529040 187463 529101
rect 187221 529006 187239 529040
rect 187273 529006 187411 529040
rect 187445 529006 187463 529040
rect 187221 528964 187463 529006
rect 172208 528930 172237 528964
rect 172271 528930 172329 528964
rect 172363 528930 172421 528964
rect 172455 528930 172513 528964
rect 172547 528930 172605 528964
rect 172639 528930 172697 528964
rect 172731 528930 172789 528964
rect 172823 528930 172881 528964
rect 172915 528930 172973 528964
rect 173007 528930 173065 528964
rect 173099 528930 173157 528964
rect 173191 528930 173249 528964
rect 173283 528930 173341 528964
rect 173375 528930 173433 528964
rect 173467 528930 173525 528964
rect 173559 528930 173617 528964
rect 173651 528930 173709 528964
rect 173743 528930 173801 528964
rect 173835 528930 173893 528964
rect 173927 528930 173985 528964
rect 174019 528930 174077 528964
rect 174111 528930 174169 528964
rect 174203 528930 174261 528964
rect 174295 528930 174353 528964
rect 174387 528930 174445 528964
rect 174479 528930 174537 528964
rect 174571 528930 174629 528964
rect 174663 528930 174721 528964
rect 174755 528930 174813 528964
rect 174847 528930 174905 528964
rect 174939 528930 174997 528964
rect 175031 528930 175089 528964
rect 175123 528930 175181 528964
rect 175215 528930 175273 528964
rect 175307 528930 175365 528964
rect 175399 528930 175457 528964
rect 175491 528930 175549 528964
rect 175583 528930 175641 528964
rect 175675 528930 175733 528964
rect 175767 528930 175825 528964
rect 175859 528930 175917 528964
rect 175951 528930 176009 528964
rect 176043 528930 176101 528964
rect 176135 528930 176193 528964
rect 176227 528930 176285 528964
rect 176319 528930 176377 528964
rect 176411 528930 176469 528964
rect 176503 528930 176561 528964
rect 176595 528930 176653 528964
rect 176687 528930 176745 528964
rect 176779 528930 176837 528964
rect 176871 528930 176929 528964
rect 176963 528930 177021 528964
rect 177055 528930 177113 528964
rect 177147 528930 177205 528964
rect 177239 528930 177297 528964
rect 177331 528930 177389 528964
rect 177423 528930 177481 528964
rect 177515 528930 177573 528964
rect 177607 528930 177665 528964
rect 177699 528930 177757 528964
rect 177791 528930 177849 528964
rect 177883 528930 177941 528964
rect 177975 528930 178033 528964
rect 178067 528930 178125 528964
rect 178159 528930 178217 528964
rect 178251 528930 178309 528964
rect 178343 528930 178401 528964
rect 178435 528930 178493 528964
rect 178527 528930 178585 528964
rect 178619 528930 178677 528964
rect 178711 528930 178769 528964
rect 178803 528930 178861 528964
rect 178895 528930 178953 528964
rect 178987 528930 179045 528964
rect 179079 528930 179137 528964
rect 179171 528930 179229 528964
rect 179263 528930 179321 528964
rect 179355 528930 179413 528964
rect 179447 528930 179505 528964
rect 179539 528930 179597 528964
rect 179631 528930 179689 528964
rect 179723 528930 179781 528964
rect 179815 528930 179873 528964
rect 179907 528930 179965 528964
rect 179999 528930 180057 528964
rect 180091 528930 180149 528964
rect 180183 528930 180241 528964
rect 180275 528930 180333 528964
rect 180367 528930 180425 528964
rect 180459 528930 180517 528964
rect 180551 528930 180609 528964
rect 180643 528930 180701 528964
rect 180735 528930 180793 528964
rect 180827 528930 180885 528964
rect 180919 528930 180977 528964
rect 181011 528930 181069 528964
rect 181103 528930 181161 528964
rect 181195 528930 181253 528964
rect 181287 528930 181345 528964
rect 181379 528930 181437 528964
rect 181471 528930 181529 528964
rect 181563 528930 181621 528964
rect 181655 528930 181713 528964
rect 181747 528930 181805 528964
rect 181839 528930 181897 528964
rect 181931 528930 181989 528964
rect 182023 528930 182081 528964
rect 182115 528930 182173 528964
rect 182207 528930 182265 528964
rect 182299 528930 182357 528964
rect 182391 528930 182449 528964
rect 182483 528930 182541 528964
rect 182575 528930 182633 528964
rect 182667 528930 182725 528964
rect 182759 528930 182817 528964
rect 182851 528930 182909 528964
rect 182943 528930 183001 528964
rect 183035 528930 183093 528964
rect 183127 528930 183185 528964
rect 183219 528930 183277 528964
rect 183311 528930 183369 528964
rect 183403 528930 183461 528964
rect 183495 528930 183553 528964
rect 183587 528930 183645 528964
rect 183679 528930 183737 528964
rect 183771 528930 183829 528964
rect 183863 528930 183921 528964
rect 183955 528930 184013 528964
rect 184047 528930 184105 528964
rect 184139 528930 184197 528964
rect 184231 528930 184289 528964
rect 184323 528930 184381 528964
rect 184415 528930 184473 528964
rect 184507 528930 184565 528964
rect 184599 528930 184657 528964
rect 184691 528930 184749 528964
rect 184783 528930 184841 528964
rect 184875 528930 184933 528964
rect 184967 528930 185025 528964
rect 185059 528930 185117 528964
rect 185151 528930 185209 528964
rect 185243 528930 185301 528964
rect 185335 528930 185393 528964
rect 185427 528930 185485 528964
rect 185519 528930 185577 528964
rect 185611 528930 185669 528964
rect 185703 528930 185761 528964
rect 185795 528930 185853 528964
rect 185887 528930 185945 528964
rect 185979 528930 186037 528964
rect 186071 528930 186129 528964
rect 186163 528930 186221 528964
rect 186255 528930 186313 528964
rect 186347 528930 186405 528964
rect 186439 528930 186497 528964
rect 186531 528930 186589 528964
rect 186623 528930 186681 528964
rect 186715 528930 186773 528964
rect 186807 528930 186865 528964
rect 186899 528930 186957 528964
rect 186991 528930 187049 528964
rect 187083 528930 187141 528964
rect 187175 528930 187233 528964
rect 187267 528930 187325 528964
rect 187359 528930 187417 528964
rect 187451 528930 187480 528964
rect 172225 528888 172467 528930
rect 172225 528854 172243 528888
rect 172277 528854 172415 528888
rect 172449 528854 172467 528888
rect 172225 528793 172467 528854
rect 172501 528888 173570 528930
rect 172501 528854 172519 528888
rect 172553 528854 173519 528888
rect 173553 528854 173570 528888
rect 172501 528843 173570 528854
rect 173605 528888 174674 528930
rect 173605 528854 173623 528888
rect 173657 528854 174623 528888
rect 174657 528854 174674 528888
rect 173605 528843 174674 528854
rect 174709 528888 175778 528930
rect 174709 528854 174727 528888
rect 174761 528854 175727 528888
rect 175761 528854 175778 528888
rect 174709 528843 175778 528854
rect 175923 528880 175957 528896
rect 172225 528759 172243 528793
rect 172277 528759 172415 528793
rect 172449 528759 172467 528793
rect 172225 528712 172467 528759
rect 172225 528644 172275 528678
rect 172309 528644 172329 528678
rect 172225 528570 172329 528644
rect 172363 528638 172467 528712
rect 172363 528604 172383 528638
rect 172417 528604 172467 528638
rect 172818 528678 172886 528695
rect 172818 528644 172835 528678
rect 172869 528644 172886 528678
rect 172225 528517 172467 528570
rect 172818 528529 172886 528644
rect 173182 528642 173252 528843
rect 173182 528608 173199 528642
rect 173233 528608 173252 528642
rect 173182 528593 173252 528608
rect 173922 528678 173990 528695
rect 173922 528644 173939 528678
rect 173973 528644 173990 528678
rect 173922 528529 173990 528644
rect 174286 528642 174356 528843
rect 174286 528608 174303 528642
rect 174337 528608 174356 528642
rect 174286 528593 174356 528608
rect 175026 528678 175094 528695
rect 175026 528644 175043 528678
rect 175077 528644 175094 528678
rect 175026 528529 175094 528644
rect 175390 528642 175460 528843
rect 175923 528812 175957 528846
rect 175993 528880 176059 528930
rect 175993 528846 176009 528880
rect 176043 528846 176059 528880
rect 175993 528812 176059 528846
rect 175993 528778 176009 528812
rect 176043 528778 176059 528812
rect 176093 528880 176147 528896
rect 176093 528846 176095 528880
rect 176129 528862 176147 528880
rect 176093 528828 176101 528846
rect 176135 528828 176147 528862
rect 176093 528799 176147 528828
rect 175923 528744 175957 528778
rect 176093 528765 176095 528799
rect 176129 528765 176147 528799
rect 175923 528710 176056 528744
rect 176093 528715 176147 528765
rect 176022 528681 176056 528710
rect 175390 528608 175407 528642
rect 175441 528608 175460 528642
rect 175390 528593 175460 528608
rect 175909 528658 175975 528674
rect 175909 528624 175917 528658
rect 175951 528652 175975 528658
rect 175909 528618 175925 528624
rect 175959 528618 175975 528652
rect 175909 528600 175975 528618
rect 176022 528665 176079 528681
rect 176022 528631 176045 528665
rect 176022 528615 176079 528631
rect 176022 528564 176056 528615
rect 175923 528530 176056 528564
rect 176113 528555 176147 528715
rect 176199 528880 176233 528896
rect 176199 528812 176233 528846
rect 176269 528880 176335 528930
rect 176269 528846 176285 528880
rect 176319 528846 176335 528880
rect 176269 528812 176335 528846
rect 176269 528778 176285 528812
rect 176319 528778 176335 528812
rect 176369 528880 176423 528896
rect 176369 528846 176371 528880
rect 176405 528846 176423 528880
rect 176369 528799 176423 528846
rect 176199 528744 176233 528778
rect 176369 528765 176371 528799
rect 176405 528765 176423 528799
rect 176199 528710 176332 528744
rect 176369 528715 176423 528765
rect 176298 528681 176332 528710
rect 176185 528658 176251 528674
rect 176185 528624 176193 528658
rect 176227 528652 176251 528658
rect 176185 528618 176201 528624
rect 176235 528618 176251 528652
rect 176185 528600 176251 528618
rect 176298 528665 176355 528681
rect 176298 528631 176321 528665
rect 176298 528615 176355 528631
rect 176298 528564 176332 528615
rect 172225 528483 172243 528517
rect 172277 528483 172415 528517
rect 172449 528483 172467 528517
rect 172225 528420 172467 528483
rect 172501 528515 173570 528529
rect 172501 528481 172519 528515
rect 172553 528481 173519 528515
rect 173553 528481 173570 528515
rect 172501 528420 173570 528481
rect 173605 528515 174674 528529
rect 173605 528481 173623 528515
rect 173657 528481 174623 528515
rect 174657 528481 174674 528515
rect 173605 528420 174674 528481
rect 174709 528515 175778 528529
rect 174709 528481 174727 528515
rect 174761 528481 175727 528515
rect 175761 528481 175778 528515
rect 174709 528420 175778 528481
rect 175923 528509 175957 528530
rect 176095 528526 176147 528555
rect 175923 528454 175957 528475
rect 175993 528462 176009 528496
rect 176043 528462 176059 528496
rect 175993 528420 176059 528462
rect 176129 528492 176147 528526
rect 176095 528454 176147 528492
rect 176199 528530 176332 528564
rect 176389 528555 176423 528715
rect 176457 528828 176560 528860
rect 176457 528794 176521 528828
rect 176555 528794 176560 528828
rect 176457 528778 176560 528794
rect 176607 528828 176641 528930
rect 176607 528778 176641 528794
rect 176675 528862 177081 528896
rect 176457 528616 176525 528778
rect 176675 528729 176709 528862
rect 176788 528794 176804 528828
rect 176838 528794 176879 528828
rect 176913 528794 177013 528828
rect 176559 528726 176575 528729
rect 176559 528692 176561 528726
rect 176609 528695 176709 528729
rect 176595 528692 176709 528695
rect 176559 528691 176709 528692
rect 176743 528729 176945 528760
rect 176777 528726 176945 528729
rect 176777 528695 176781 528726
rect 176457 528582 176653 528616
rect 176687 528582 176703 528616
rect 176199 528509 176233 528530
rect 176371 528526 176423 528555
rect 176405 528522 176423 528526
rect 176199 528454 176233 528475
rect 176269 528462 176285 528496
rect 176319 528462 176335 528496
rect 176269 528420 176335 528462
rect 176371 528488 176377 528492
rect 176411 528488 176423 528522
rect 176371 528454 176423 528488
rect 176512 528511 176561 528582
rect 176512 528477 176521 528511
rect 176555 528477 176561 528511
rect 176512 528461 176561 528477
rect 176605 528511 176707 528527
rect 176639 528477 176673 528511
rect 176605 528420 176707 528477
rect 176743 528522 176781 528695
rect 176743 528488 176745 528522
rect 176779 528488 176781 528522
rect 176743 528454 176781 528488
rect 176815 528658 176870 528686
rect 176815 528624 176837 528658
rect 176815 528616 176870 528624
rect 176849 528582 176870 528616
rect 176815 528454 176870 528582
rect 176911 528616 176945 528726
rect 176911 528566 176945 528582
rect 176979 528568 177013 528794
rect 177047 528668 177081 528862
rect 177115 528888 177149 528930
rect 177115 528820 177149 528854
rect 177115 528752 177149 528786
rect 177115 528702 177149 528718
rect 177183 528888 177250 528896
rect 177183 528854 177199 528888
rect 177233 528854 177250 528888
rect 177183 528820 177250 528854
rect 177183 528786 177199 528820
rect 177233 528786 177250 528820
rect 177183 528752 177250 528786
rect 177183 528718 177199 528752
rect 177233 528718 177250 528752
rect 177183 528702 177250 528718
rect 177047 528652 177086 528668
rect 177047 528618 177052 528652
rect 177047 528602 177086 528618
rect 177131 528652 177182 528668
rect 177131 528618 177148 528652
rect 177131 528602 177182 528618
rect 177131 528568 177165 528602
rect 177216 528568 177250 528702
rect 177377 528859 177435 528930
rect 177377 528825 177389 528859
rect 177423 528825 177435 528859
rect 177377 528766 177435 528825
rect 177377 528732 177389 528766
rect 177423 528732 177435 528766
rect 177377 528697 177435 528732
rect 177469 528862 177546 528896
rect 177469 528828 177506 528862
rect 177540 528828 177546 528862
rect 177580 528888 177645 528930
rect 177580 528854 177596 528888
rect 177630 528854 177645 528888
rect 177580 528838 177645 528854
rect 177749 528862 177805 528896
rect 177469 528702 177546 528828
rect 177749 528828 177755 528862
rect 177789 528828 177805 528862
rect 177749 528804 177805 528828
rect 177580 528760 177805 528804
rect 177843 528862 177923 528896
rect 177843 528828 177859 528862
rect 177893 528828 177923 528862
rect 178003 528888 178057 528930
rect 178003 528854 178013 528888
rect 178047 528854 178057 528888
rect 178003 528838 178057 528854
rect 178091 528862 178148 528896
rect 176979 528534 177165 528568
rect 176979 528527 177014 528534
rect 176908 528511 177014 528527
rect 176942 528477 177014 528511
rect 177199 528522 177250 528568
rect 177469 528658 177525 528702
rect 177580 528668 177670 528760
rect 177843 528726 177923 528828
rect 178091 528828 178097 528862
rect 178131 528828 178148 528862
rect 178091 528804 178148 528828
rect 177469 528624 177481 528658
rect 177515 528624 177525 528658
rect 177469 528568 177525 528624
rect 177559 528652 177670 528668
rect 177593 528618 177670 528652
rect 177559 528602 177670 528618
rect 177704 528652 177923 528726
rect 177704 528618 177755 528652
rect 177789 528618 177923 528652
rect 177704 528614 177923 528618
rect 177580 528580 177670 528602
rect 177199 528515 177205 528522
rect 176908 528454 177014 528477
rect 177099 528496 177165 528500
rect 177099 528462 177115 528496
rect 177149 528462 177165 528496
rect 177099 528420 177165 528462
rect 177239 528488 177250 528522
rect 177233 528481 177250 528488
rect 177199 528454 177250 528481
rect 177377 528548 177435 528565
rect 177377 528514 177389 528548
rect 177423 528514 177435 528548
rect 177377 528420 177435 528514
rect 177469 528522 177546 528568
rect 177580 528546 177805 528580
rect 177469 528488 177506 528522
rect 177540 528488 177546 528522
rect 177749 528522 177805 528546
rect 177469 528454 177546 528488
rect 177580 528496 177645 528512
rect 177580 528462 177596 528496
rect 177630 528462 177645 528496
rect 177580 528420 177645 528462
rect 177749 528488 177755 528522
rect 177789 528488 177805 528522
rect 177749 528454 177805 528488
rect 177843 528522 177923 528614
rect 177957 528760 178148 528804
rect 178391 528888 178450 528930
rect 178391 528854 178407 528888
rect 178441 528854 178450 528888
rect 178391 528820 178450 528854
rect 178391 528786 178407 528820
rect 178441 528786 178450 528820
rect 178391 528768 178450 528786
rect 178486 528880 178535 528896
rect 178486 528846 178493 528880
rect 178527 528846 178535 528880
rect 178486 528812 178535 528846
rect 178486 528778 178493 528812
rect 178527 528778 178535 528812
rect 177957 528652 177999 528760
rect 177957 528618 177959 528652
rect 177993 528618 177999 528652
rect 177957 528580 177999 528618
rect 178033 528692 178125 528726
rect 178159 528692 178171 528726
rect 178033 528652 178171 528692
rect 178486 528668 178535 528778
rect 178570 528888 178622 528930
rect 178742 528929 179997 528930
rect 178570 528854 178579 528888
rect 178613 528854 178622 528888
rect 178570 528820 178622 528854
rect 178570 528786 178579 528820
rect 178613 528786 178622 528820
rect 178570 528768 178622 528786
rect 178658 528872 178708 528895
rect 178658 528838 178665 528872
rect 178699 528838 178708 528872
rect 178658 528804 178708 528838
rect 178658 528770 178665 528804
rect 178699 528770 178708 528804
rect 178742 528888 178794 528929
rect 178742 528854 178751 528888
rect 178785 528854 178794 528888
rect 178742 528820 178794 528854
rect 178742 528786 178751 528820
rect 178785 528786 178794 528820
rect 178742 528770 178794 528786
rect 178828 528844 178880 528895
rect 178828 528810 178837 528844
rect 178871 528810 178880 528844
rect 178658 528668 178708 528770
rect 178828 528758 178880 528810
rect 178914 528864 178966 528929
rect 178914 528830 178923 528864
rect 178957 528830 178966 528864
rect 178914 528784 178966 528830
rect 179000 528844 179052 528895
rect 179000 528810 179009 528844
rect 179043 528810 179052 528844
rect 178828 528724 178837 528758
rect 178871 528750 178880 528758
rect 179000 528758 179052 528810
rect 179086 528864 179138 528929
rect 179086 528830 179095 528864
rect 179129 528830 179138 528864
rect 179086 528784 179138 528830
rect 179172 528844 179224 528895
rect 179172 528810 179181 528844
rect 179215 528810 179224 528844
rect 179000 528750 179009 528758
rect 178871 528724 179009 528750
rect 179043 528750 179052 528758
rect 179172 528758 179224 528810
rect 179258 528864 179310 528929
rect 179258 528830 179267 528864
rect 179301 528830 179310 528864
rect 179258 528784 179310 528830
rect 179344 528844 179396 528895
rect 179344 528810 179353 528844
rect 179387 528810 179396 528844
rect 179172 528750 179181 528758
rect 179043 528724 179181 528750
rect 179215 528750 179224 528758
rect 179344 528758 179396 528810
rect 179430 528864 179479 528929
rect 179430 528830 179439 528864
rect 179473 528830 179479 528864
rect 179430 528784 179479 528830
rect 179513 528844 179565 528895
rect 179513 528810 179524 528844
rect 179558 528810 179565 528844
rect 179344 528750 179353 528758
rect 179215 528724 179353 528750
rect 179387 528750 179396 528758
rect 179513 528758 179565 528810
rect 179602 528864 179651 528929
rect 179602 528830 179610 528864
rect 179644 528830 179651 528864
rect 179602 528784 179651 528830
rect 179685 528862 179737 528895
rect 179685 528828 179689 528862
rect 179723 528844 179737 528862
rect 179685 528810 179696 528828
rect 179730 528810 179737 528844
rect 179513 528750 179524 528758
rect 179387 528724 179524 528750
rect 179558 528750 179565 528758
rect 179685 528758 179737 528810
rect 179774 528864 179823 528929
rect 179774 528830 179782 528864
rect 179816 528830 179823 528864
rect 179774 528784 179823 528830
rect 179857 528844 179909 528895
rect 179857 528810 179868 528844
rect 179902 528810 179909 528844
rect 179685 528750 179696 528758
rect 179558 528724 179696 528750
rect 179730 528750 179737 528758
rect 179857 528758 179909 528810
rect 179946 528864 179997 528929
rect 179946 528830 179954 528864
rect 179988 528830 179997 528864
rect 179946 528784 179997 528830
rect 180031 528844 180089 528895
rect 180031 528810 180040 528844
rect 180074 528810 180089 528844
rect 179857 528750 179868 528758
rect 179730 528724 179868 528750
rect 179902 528747 179909 528758
rect 180031 528758 180089 528810
rect 180123 528864 180177 528930
rect 180123 528830 180126 528864
rect 180160 528830 180177 528864
rect 180123 528781 180177 528830
rect 180247 528880 180281 528896
rect 180247 528812 180281 528846
rect 180031 528747 180040 528758
rect 179902 528724 180040 528747
rect 180074 528747 180089 528758
rect 180317 528880 180383 528930
rect 180317 528846 180333 528880
rect 180367 528846 180383 528880
rect 180317 528812 180383 528846
rect 180317 528778 180333 528812
rect 180367 528778 180383 528812
rect 180417 528880 180471 528896
rect 180417 528846 180419 528880
rect 180453 528846 180471 528880
rect 180417 528799 180471 528846
rect 180074 528724 180177 528747
rect 178828 528702 180177 528724
rect 180247 528744 180281 528778
rect 180417 528765 180419 528799
rect 180453 528794 180471 528799
rect 180417 528760 180425 528765
rect 180459 528760 180471 528794
rect 180506 528880 180557 528896
rect 180506 528846 180523 528880
rect 180506 528812 180557 528846
rect 180591 528864 180657 528930
rect 180591 528830 180607 528864
rect 180641 528830 180657 528864
rect 180691 528880 180725 528896
rect 180506 528778 180523 528812
rect 180691 528812 180725 528846
rect 180557 528778 180656 528796
rect 180506 528762 180656 528778
rect 180247 528710 180380 528744
rect 180417 528715 180471 528760
rect 178033 528618 178073 528652
rect 178107 528618 178171 528652
rect 178033 528614 178171 528618
rect 178389 528652 178452 528668
rect 178389 528618 178409 528652
rect 178443 528618 178452 528652
rect 178389 528590 178452 528618
rect 177957 528546 178148 528580
rect 178389 528556 178401 528590
rect 178435 528556 178452 528590
rect 178486 528652 179910 528668
rect 178486 528618 178836 528652
rect 178870 528618 178904 528652
rect 178938 528618 178972 528652
rect 179006 528618 179040 528652
rect 179074 528618 179108 528652
rect 179142 528618 179176 528652
rect 179210 528618 179244 528652
rect 179278 528618 179312 528652
rect 179346 528618 179380 528652
rect 179414 528618 179448 528652
rect 179482 528618 179516 528652
rect 179550 528618 179584 528652
rect 179618 528618 179652 528652
rect 179686 528618 179720 528652
rect 179754 528618 179788 528652
rect 179822 528618 179856 528652
rect 179890 528618 179910 528652
rect 177843 528488 177859 528522
rect 177893 528488 177923 528522
rect 178091 528522 178148 528546
rect 177843 528454 177923 528488
rect 178003 528496 178057 528512
rect 178003 528462 178013 528496
rect 178047 528462 178057 528496
rect 178003 528420 178057 528462
rect 178091 528488 178097 528522
rect 178131 528488 178148 528522
rect 178091 528454 178148 528488
rect 178389 528496 178450 528522
rect 178389 528462 178407 528496
rect 178441 528462 178450 528496
rect 178389 528420 178450 528462
rect 178486 528509 178536 528618
rect 178486 528475 178493 528509
rect 178527 528475 178536 528509
rect 178486 528456 178536 528475
rect 178570 528509 178622 528525
rect 178570 528475 178579 528509
rect 178613 528475 178622 528509
rect 178570 528420 178622 528475
rect 178658 528509 178708 528618
rect 179944 528584 180177 528702
rect 180346 528681 180380 528710
rect 180233 528658 180299 528674
rect 180233 528624 180241 528658
rect 180275 528652 180299 528658
rect 180233 528618 180249 528624
rect 180283 528618 180299 528652
rect 180233 528600 180299 528618
rect 180346 528665 180403 528681
rect 180346 528631 180369 528665
rect 180346 528615 180403 528631
rect 178828 528550 180177 528584
rect 180346 528564 180380 528615
rect 178658 528475 178665 528509
rect 178699 528475 178708 528509
rect 178658 528456 178708 528475
rect 178742 528509 178794 528532
rect 178742 528475 178751 528509
rect 178785 528475 178794 528509
rect 178742 528420 178794 528475
rect 178828 528509 178880 528550
rect 178828 528475 178837 528509
rect 178871 528475 178880 528509
rect 178828 528459 178880 528475
rect 178914 528500 178966 528516
rect 178914 528466 178923 528500
rect 178957 528466 178966 528500
rect 178914 528420 178966 528466
rect 179000 528509 179052 528550
rect 179000 528475 179009 528509
rect 179043 528475 179052 528509
rect 179000 528459 179052 528475
rect 179086 528500 179138 528516
rect 179086 528466 179095 528500
rect 179129 528466 179138 528500
rect 179086 528420 179138 528466
rect 179172 528509 179224 528550
rect 179172 528475 179181 528509
rect 179215 528475 179224 528509
rect 179172 528459 179224 528475
rect 179258 528500 179307 528516
rect 179258 528466 179267 528500
rect 179301 528466 179307 528500
rect 179258 528420 179307 528466
rect 179341 528509 179396 528550
rect 179341 528475 179353 528509
rect 179387 528475 179396 528509
rect 179341 528459 179396 528475
rect 179430 528500 179479 528516
rect 179430 528466 179439 528500
rect 179473 528466 179479 528500
rect 179430 528420 179479 528466
rect 179513 528509 179565 528550
rect 179513 528475 179524 528509
rect 179558 528475 179565 528509
rect 179513 528459 179565 528475
rect 179601 528500 179651 528516
rect 179601 528466 179610 528500
rect 179644 528466 179651 528500
rect 179601 528420 179651 528466
rect 179685 528509 179737 528550
rect 179685 528475 179696 528509
rect 179730 528475 179737 528509
rect 179685 528459 179737 528475
rect 179773 528500 179823 528516
rect 179773 528466 179782 528500
rect 179816 528466 179823 528500
rect 179773 528420 179823 528466
rect 179857 528509 179909 528550
rect 179857 528475 179868 528509
rect 179902 528475 179909 528509
rect 179857 528459 179909 528475
rect 179945 528500 179997 528516
rect 179945 528466 179954 528500
rect 179988 528466 179997 528500
rect 179945 528420 179997 528466
rect 180031 528509 180083 528550
rect 180247 528530 180380 528564
rect 180437 528555 180471 528715
rect 180506 528726 180576 528728
rect 180506 528692 180517 528726
rect 180551 528692 180576 528726
rect 180506 528652 180576 528692
rect 180506 528618 180520 528652
rect 180554 528618 180576 528652
rect 180506 528598 180576 528618
rect 180610 528667 180656 528762
rect 180610 528658 180622 528667
rect 180644 528624 180656 528633
rect 180610 528564 180656 528624
rect 180031 528475 180040 528509
rect 180074 528475 180083 528509
rect 180031 528459 180083 528475
rect 180117 528500 180177 528516
rect 180117 528466 180126 528500
rect 180160 528466 180177 528500
rect 180117 528420 180177 528466
rect 180247 528509 180281 528530
rect 180419 528526 180471 528555
rect 180247 528454 180281 528475
rect 180317 528462 180333 528496
rect 180367 528462 180383 528496
rect 180317 528420 180383 528462
rect 180453 528492 180471 528526
rect 180419 528454 180471 528492
rect 180506 528530 180656 528564
rect 180506 528522 180557 528530
rect 180506 528488 180523 528522
rect 180691 528522 180725 528760
rect 180759 528736 180824 528893
rect 180858 528888 180908 528930
rect 180858 528854 180874 528888
rect 180858 528838 180908 528854
rect 180942 528880 180992 528896
rect 180942 528846 180958 528880
rect 180942 528830 180992 528846
rect 181035 528886 181171 528896
rect 181035 528852 181051 528886
rect 181085 528852 181171 528886
rect 181286 528878 181352 528930
rect 181479 528888 181553 528930
rect 181035 528830 181171 528852
rect 180942 528804 180976 528830
rect 180897 528770 180976 528804
rect 181010 528794 181103 528796
rect 180771 528726 180863 528736
rect 180771 528692 180793 528726
rect 180827 528713 180863 528726
rect 180827 528692 180829 528713
rect 180771 528679 180829 528692
rect 180771 528526 180863 528679
rect 180506 528472 180557 528488
rect 180591 528462 180607 528496
rect 180641 528462 180657 528496
rect 180897 528498 180931 528770
rect 181010 528768 181069 528794
rect 181044 528760 181069 528768
rect 181044 528734 181103 528760
rect 181010 528718 181103 528734
rect 180965 528658 181035 528680
rect 180965 528624 180977 528658
rect 181011 528624 181035 528658
rect 180965 528606 181035 528624
rect 180965 528572 180988 528606
rect 181022 528572 181035 528606
rect 180965 528556 181035 528572
rect 181069 528600 181103 528718
rect 181137 528674 181171 528830
rect 181205 528862 181239 528878
rect 181286 528844 181302 528878
rect 181336 528844 181352 528878
rect 181386 528862 181420 528878
rect 181205 528810 181239 528828
rect 181479 528854 181499 528888
rect 181533 528854 181553 528888
rect 181479 528838 181553 528854
rect 181587 528880 181621 528896
rect 181386 528810 181420 528828
rect 181205 528776 181420 528810
rect 181587 528804 181621 528846
rect 181668 528887 181842 528896
rect 181668 528853 181684 528887
rect 181718 528853 181842 528887
rect 181668 528828 181842 528853
rect 181876 528888 181926 528930
rect 181910 528854 181926 528888
rect 182030 528888 182096 528930
rect 181876 528838 181926 528854
rect 181960 528862 181994 528878
rect 181509 528770 181621 528804
rect 181509 528742 181543 528770
rect 181243 528708 181259 528742
rect 181293 528708 181543 528742
rect 181682 528760 181693 528794
rect 181727 528768 181774 528794
rect 181682 528736 181724 528760
rect 181137 528654 181475 528674
rect 181137 528640 181441 528654
rect 181069 528566 181090 528600
rect 181124 528566 181140 528600
rect 181069 528556 181140 528566
rect 181174 528498 181208 528640
rect 181249 528590 181345 528606
rect 181283 528556 181321 528590
rect 181379 528572 181407 528606
rect 181441 528604 181475 528620
rect 181355 528556 181407 528572
rect 181509 528570 181543 528708
rect 180691 528472 180725 528488
rect 180591 528420 180657 528462
rect 180797 528458 180813 528492
rect 180847 528458 180863 528492
rect 180897 528464 180946 528498
rect 180980 528464 180996 528498
rect 181037 528464 181053 528498
rect 181087 528464 181208 528498
rect 181383 528496 181449 528512
rect 180797 528420 180863 528458
rect 181383 528462 181399 528496
rect 181433 528462 181449 528496
rect 181383 528420 181449 528462
rect 181491 528492 181543 528570
rect 181581 528734 181724 528736
rect 181758 528734 181774 528768
rect 181808 528752 181842 528828
rect 182030 528854 182046 528888
rect 182080 528854 182096 528888
rect 182164 528888 182225 528930
rect 182164 528854 182175 528888
rect 182209 528854 182225 528888
rect 181960 528820 181994 528828
rect 182164 528820 182225 528854
rect 181960 528786 182120 528820
rect 181581 528702 181716 528734
rect 181808 528718 182002 528752
rect 182036 528718 182052 528752
rect 181581 528594 181623 528702
rect 181808 528700 181842 528718
rect 181581 528560 181589 528594
rect 181581 528544 181623 528560
rect 181657 528658 181727 528668
rect 181657 528642 181693 528658
rect 181657 528608 181685 528642
rect 181719 528608 181727 528624
rect 181657 528544 181727 528608
rect 181761 528666 181842 528700
rect 181761 528510 181795 528666
rect 181909 528653 182017 528684
rect 182086 528668 182120 528786
rect 182164 528786 182175 528820
rect 182209 528786 182225 528820
rect 182164 528702 182225 528786
rect 182259 528862 182310 528868
rect 182259 528852 182265 528862
rect 182299 528828 182310 528862
rect 182293 528818 182310 528828
rect 182259 528784 182310 528818
rect 182293 528750 182310 528784
rect 182259 528692 182310 528750
rect 182529 528859 182587 528930
rect 182529 528825 182541 528859
rect 182575 528825 182587 528859
rect 182621 528888 183690 528930
rect 182621 528854 182639 528888
rect 182673 528854 183639 528888
rect 183673 528854 183690 528888
rect 182621 528843 183690 528854
rect 183725 528888 184794 528930
rect 183725 528854 183743 528888
rect 183777 528854 184743 528888
rect 184777 528854 184794 528888
rect 183725 528843 184794 528854
rect 184829 528888 185898 528930
rect 184829 528854 184847 528888
rect 184881 528854 185847 528888
rect 185881 528854 185898 528888
rect 184829 528843 185898 528854
rect 185933 528888 187002 528930
rect 185933 528854 185951 528888
rect 185985 528854 186951 528888
rect 186985 528854 187002 528888
rect 185933 528843 187002 528854
rect 187221 528888 187463 528930
rect 187221 528854 187239 528888
rect 187273 528854 187411 528888
rect 187445 528854 187463 528888
rect 182529 528766 182587 528825
rect 182529 528732 182541 528766
rect 182575 528732 182587 528766
rect 182529 528697 182587 528732
rect 182086 528662 182234 528668
rect 181943 528644 182017 528653
rect 181829 528616 181873 528632
rect 181863 528582 181873 528616
rect 181909 528610 181925 528619
rect 181959 528610 182017 528644
rect 181829 528576 181873 528582
rect 181969 528590 182017 528610
rect 181829 528542 181935 528576
rect 181605 528496 181795 528510
rect 181491 528458 181511 528492
rect 181545 528458 181561 528492
rect 181605 528462 181621 528496
rect 181655 528462 181795 528496
rect 181605 528454 181795 528462
rect 181829 528492 181867 528508
rect 181829 528458 181833 528492
rect 181901 528496 181935 528542
rect 182003 528556 182017 528590
rect 181969 528530 182017 528556
rect 182051 528652 182234 528662
rect 182051 528618 182200 528652
rect 182051 528602 182234 528618
rect 182051 528567 182116 528602
rect 182051 528512 182115 528567
rect 182268 528562 182310 528692
rect 182938 528678 183006 528695
rect 182938 528644 182955 528678
rect 182989 528644 183006 528678
rect 182259 528546 182310 528562
rect 182293 528512 182310 528546
rect 181901 528478 182051 528496
rect 182085 528478 182115 528512
rect 181901 528462 182115 528478
rect 182164 528496 182225 528512
rect 182164 528462 182175 528496
rect 182209 528462 182225 528496
rect 181829 528420 181867 528458
rect 182164 528420 182225 528462
rect 182259 528456 182310 528512
rect 182529 528548 182587 528565
rect 182529 528514 182541 528548
rect 182575 528514 182587 528548
rect 182938 528529 183006 528644
rect 183302 528642 183372 528843
rect 183302 528608 183319 528642
rect 183353 528608 183372 528642
rect 183302 528593 183372 528608
rect 184042 528678 184110 528695
rect 184042 528644 184059 528678
rect 184093 528644 184110 528678
rect 184042 528529 184110 528644
rect 184406 528642 184476 528843
rect 184406 528608 184423 528642
rect 184457 528608 184476 528642
rect 184406 528593 184476 528608
rect 185146 528678 185214 528695
rect 185146 528644 185163 528678
rect 185197 528644 185214 528678
rect 185146 528529 185214 528644
rect 185510 528642 185580 528843
rect 185510 528608 185527 528642
rect 185561 528608 185580 528642
rect 185510 528593 185580 528608
rect 186250 528678 186318 528695
rect 186250 528644 186267 528678
rect 186301 528644 186318 528678
rect 186250 528529 186318 528644
rect 186614 528642 186684 528843
rect 186614 528608 186631 528642
rect 186665 528608 186684 528642
rect 186614 528593 186684 528608
rect 187221 528793 187463 528854
rect 187221 528759 187239 528793
rect 187273 528759 187411 528793
rect 187445 528759 187463 528793
rect 187221 528712 187463 528759
rect 187221 528638 187325 528712
rect 187221 528604 187271 528638
rect 187305 528604 187325 528638
rect 187359 528644 187379 528678
rect 187413 528644 187463 528678
rect 187359 528570 187463 528644
rect 182529 528420 182587 528514
rect 182621 528515 183690 528529
rect 182621 528481 182639 528515
rect 182673 528481 183639 528515
rect 183673 528481 183690 528515
rect 182621 528420 183690 528481
rect 183725 528515 184794 528529
rect 183725 528481 183743 528515
rect 183777 528481 184743 528515
rect 184777 528481 184794 528515
rect 183725 528420 184794 528481
rect 184829 528515 185898 528529
rect 184829 528481 184847 528515
rect 184881 528481 185847 528515
rect 185881 528481 185898 528515
rect 184829 528420 185898 528481
rect 185933 528515 187002 528529
rect 185933 528481 185951 528515
rect 185985 528481 186951 528515
rect 186985 528481 187002 528515
rect 185933 528420 187002 528481
rect 187221 528517 187463 528570
rect 187221 528483 187239 528517
rect 187273 528483 187411 528517
rect 187445 528483 187463 528517
rect 187221 528420 187463 528483
rect 172208 528386 172237 528420
rect 172271 528386 172329 528420
rect 172363 528386 172421 528420
rect 172455 528386 172513 528420
rect 172547 528386 172605 528420
rect 172639 528386 172697 528420
rect 172731 528386 172789 528420
rect 172823 528386 172881 528420
rect 172915 528386 172973 528420
rect 173007 528386 173065 528420
rect 173099 528386 173157 528420
rect 173191 528386 173249 528420
rect 173283 528386 173341 528420
rect 173375 528386 173433 528420
rect 173467 528386 173525 528420
rect 173559 528386 173617 528420
rect 173651 528386 173709 528420
rect 173743 528386 173801 528420
rect 173835 528386 173893 528420
rect 173927 528386 173985 528420
rect 174019 528386 174077 528420
rect 174111 528386 174169 528420
rect 174203 528386 174261 528420
rect 174295 528386 174353 528420
rect 174387 528386 174445 528420
rect 174479 528386 174537 528420
rect 174571 528386 174629 528420
rect 174663 528386 174721 528420
rect 174755 528386 174813 528420
rect 174847 528386 174905 528420
rect 174939 528386 174997 528420
rect 175031 528386 175089 528420
rect 175123 528386 175181 528420
rect 175215 528386 175273 528420
rect 175307 528386 175365 528420
rect 175399 528386 175457 528420
rect 175491 528386 175549 528420
rect 175583 528386 175641 528420
rect 175675 528386 175733 528420
rect 175767 528386 175825 528420
rect 175859 528386 175917 528420
rect 175951 528386 176009 528420
rect 176043 528386 176101 528420
rect 176135 528386 176193 528420
rect 176227 528386 176285 528420
rect 176319 528386 176377 528420
rect 176411 528386 176469 528420
rect 176503 528386 176561 528420
rect 176595 528386 176653 528420
rect 176687 528386 176745 528420
rect 176779 528386 176837 528420
rect 176871 528386 176929 528420
rect 176963 528386 177021 528420
rect 177055 528386 177113 528420
rect 177147 528386 177205 528420
rect 177239 528386 177297 528420
rect 177331 528386 177389 528420
rect 177423 528386 177481 528420
rect 177515 528386 177573 528420
rect 177607 528386 177665 528420
rect 177699 528386 177757 528420
rect 177791 528386 177849 528420
rect 177883 528386 177941 528420
rect 177975 528386 178033 528420
rect 178067 528386 178125 528420
rect 178159 528386 178217 528420
rect 178251 528386 178309 528420
rect 178343 528386 178401 528420
rect 178435 528386 178493 528420
rect 178527 528386 178585 528420
rect 178619 528386 178677 528420
rect 178711 528386 178769 528420
rect 178803 528386 178861 528420
rect 178895 528386 178953 528420
rect 178987 528386 179045 528420
rect 179079 528386 179137 528420
rect 179171 528386 179229 528420
rect 179263 528386 179321 528420
rect 179355 528386 179413 528420
rect 179447 528386 179505 528420
rect 179539 528386 179597 528420
rect 179631 528386 179689 528420
rect 179723 528386 179781 528420
rect 179815 528386 179873 528420
rect 179907 528386 179965 528420
rect 179999 528386 180057 528420
rect 180091 528386 180149 528420
rect 180183 528386 180241 528420
rect 180275 528386 180333 528420
rect 180367 528386 180425 528420
rect 180459 528386 180517 528420
rect 180551 528386 180609 528420
rect 180643 528386 180701 528420
rect 180735 528386 180793 528420
rect 180827 528386 180885 528420
rect 180919 528386 180977 528420
rect 181011 528386 181069 528420
rect 181103 528386 181161 528420
rect 181195 528386 181253 528420
rect 181287 528386 181345 528420
rect 181379 528386 181437 528420
rect 181471 528386 181529 528420
rect 181563 528386 181621 528420
rect 181655 528386 181713 528420
rect 181747 528386 181805 528420
rect 181839 528386 181897 528420
rect 181931 528386 181989 528420
rect 182023 528386 182081 528420
rect 182115 528386 182173 528420
rect 182207 528386 182265 528420
rect 182299 528386 182357 528420
rect 182391 528386 182449 528420
rect 182483 528386 182541 528420
rect 182575 528386 182633 528420
rect 182667 528386 182725 528420
rect 182759 528386 182817 528420
rect 182851 528386 182909 528420
rect 182943 528386 183001 528420
rect 183035 528386 183093 528420
rect 183127 528386 183185 528420
rect 183219 528386 183277 528420
rect 183311 528386 183369 528420
rect 183403 528386 183461 528420
rect 183495 528386 183553 528420
rect 183587 528386 183645 528420
rect 183679 528386 183737 528420
rect 183771 528386 183829 528420
rect 183863 528386 183921 528420
rect 183955 528386 184013 528420
rect 184047 528386 184105 528420
rect 184139 528386 184197 528420
rect 184231 528386 184289 528420
rect 184323 528386 184381 528420
rect 184415 528386 184473 528420
rect 184507 528386 184565 528420
rect 184599 528386 184657 528420
rect 184691 528386 184749 528420
rect 184783 528386 184841 528420
rect 184875 528386 184933 528420
rect 184967 528386 185025 528420
rect 185059 528386 185117 528420
rect 185151 528386 185209 528420
rect 185243 528386 185301 528420
rect 185335 528386 185393 528420
rect 185427 528386 185485 528420
rect 185519 528386 185577 528420
rect 185611 528386 185669 528420
rect 185703 528386 185761 528420
rect 185795 528386 185853 528420
rect 185887 528386 185945 528420
rect 185979 528386 186037 528420
rect 186071 528386 186129 528420
rect 186163 528386 186221 528420
rect 186255 528386 186313 528420
rect 186347 528386 186405 528420
rect 186439 528386 186497 528420
rect 186531 528386 186589 528420
rect 186623 528386 186681 528420
rect 186715 528386 186773 528420
rect 186807 528386 186865 528420
rect 186899 528386 186957 528420
rect 186991 528386 187049 528420
rect 187083 528386 187141 528420
rect 187175 528386 187233 528420
rect 187267 528386 187325 528420
rect 187359 528386 187417 528420
rect 187451 528386 187480 528420
rect 172225 528323 172467 528386
rect 172225 528289 172243 528323
rect 172277 528289 172415 528323
rect 172449 528289 172467 528323
rect 172225 528236 172467 528289
rect 172501 528325 173570 528386
rect 172501 528291 172519 528325
rect 172553 528291 173519 528325
rect 173553 528291 173570 528325
rect 172501 528277 173570 528291
rect 173605 528325 174674 528386
rect 173605 528291 173623 528325
rect 173657 528291 174623 528325
rect 174657 528291 174674 528325
rect 173605 528277 174674 528291
rect 174801 528292 174859 528386
rect 172225 528162 172329 528236
rect 172225 528128 172275 528162
rect 172309 528128 172329 528162
rect 172363 528168 172383 528202
rect 172417 528168 172467 528202
rect 172363 528094 172467 528168
rect 172818 528162 172886 528277
rect 172818 528128 172835 528162
rect 172869 528128 172886 528162
rect 172818 528111 172886 528128
rect 173182 528198 173252 528213
rect 173182 528164 173199 528198
rect 173233 528164 173252 528198
rect 172225 528047 172467 528094
rect 172225 528013 172243 528047
rect 172277 528013 172415 528047
rect 172449 528013 172467 528047
rect 172225 527952 172467 528013
rect 173182 527963 173252 528164
rect 173922 528162 173990 528277
rect 174801 528258 174813 528292
rect 174847 528258 174859 528292
rect 174893 528325 175962 528386
rect 176175 528344 176241 528386
rect 174893 528291 174911 528325
rect 174945 528291 175911 528325
rect 175945 528291 175962 528325
rect 174893 528277 175962 528291
rect 176090 528318 176141 528334
rect 176090 528284 176107 528318
rect 176175 528310 176191 528344
rect 176225 528310 176241 528344
rect 176381 528348 176447 528386
rect 176275 528318 176309 528334
rect 174801 528241 174859 528258
rect 173922 528128 173939 528162
rect 173973 528128 173990 528162
rect 173922 528111 173990 528128
rect 174286 528198 174356 528213
rect 174286 528164 174303 528198
rect 174337 528164 174356 528198
rect 174286 527963 174356 528164
rect 175210 528162 175278 528277
rect 176090 528276 176141 528284
rect 176381 528314 176397 528348
rect 176431 528314 176447 528348
rect 176967 528344 177033 528386
rect 176090 528242 176240 528276
rect 175210 528128 175227 528162
rect 175261 528128 175278 528162
rect 175210 528111 175278 528128
rect 175574 528198 175644 528213
rect 175574 528164 175591 528198
rect 175625 528164 175644 528198
rect 174801 528074 174859 528109
rect 174801 528040 174813 528074
rect 174847 528040 174859 528074
rect 174801 527981 174859 528040
rect 172225 527918 172243 527952
rect 172277 527918 172415 527952
rect 172449 527918 172467 527952
rect 172225 527876 172467 527918
rect 172501 527952 173570 527963
rect 172501 527918 172519 527952
rect 172553 527918 173519 527952
rect 173553 527918 173570 527952
rect 172501 527876 173570 527918
rect 173605 527952 174674 527963
rect 173605 527918 173623 527952
rect 173657 527918 174623 527952
rect 174657 527918 174674 527952
rect 173605 527876 174674 527918
rect 174801 527947 174813 527981
rect 174847 527947 174859 527981
rect 175574 527963 175644 528164
rect 176090 528188 176160 528208
rect 176090 528182 176104 528188
rect 176090 528148 176101 528182
rect 176138 528154 176160 528188
rect 176135 528148 176160 528154
rect 176090 528078 176160 528148
rect 176194 528182 176240 528242
rect 176228 528173 176240 528182
rect 176194 528139 176206 528148
rect 176194 528044 176240 528139
rect 176090 528028 176240 528044
rect 176090 527994 176107 528028
rect 176141 528010 176240 528028
rect 176275 528046 176309 528284
rect 176481 528308 176530 528342
rect 176564 528308 176580 528342
rect 176621 528308 176637 528342
rect 176671 528308 176792 528342
rect 176355 528250 176447 528280
rect 176355 528216 176377 528250
rect 176411 528216 176447 528250
rect 176355 528127 176447 528216
rect 176355 528093 176413 528127
rect 176355 528070 176447 528093
rect 174801 527876 174859 527947
rect 174893 527952 175962 527963
rect 174893 527918 174911 527952
rect 174945 527918 175911 527952
rect 175945 527918 175962 527952
rect 174893 527876 175962 527918
rect 176090 527960 176141 527994
rect 176090 527926 176107 527960
rect 176090 527910 176141 527926
rect 176175 527942 176191 527976
rect 176225 527942 176241 527976
rect 176175 527876 176241 527942
rect 176275 527960 176309 527994
rect 176275 527910 176309 527926
rect 176343 527913 176408 528070
rect 176481 528036 176515 528308
rect 176549 528234 176619 528250
rect 176549 528200 176572 528234
rect 176606 528200 176619 528234
rect 176549 528182 176619 528200
rect 176549 528148 176561 528182
rect 176595 528148 176619 528182
rect 176549 528126 176619 528148
rect 176653 528240 176724 528250
rect 176653 528206 176674 528240
rect 176708 528206 176724 528240
rect 176653 528088 176687 528206
rect 176758 528166 176792 528308
rect 176967 528310 176983 528344
rect 177017 528310 177033 528344
rect 176967 528294 177033 528310
rect 177075 528314 177095 528348
rect 177129 528314 177145 528348
rect 177189 528344 177379 528352
rect 176867 528216 176905 528250
rect 176939 528234 176991 528250
rect 177075 528236 177127 528314
rect 177189 528310 177205 528344
rect 177239 528310 177379 528344
rect 177189 528296 177379 528310
rect 177413 528348 177451 528386
rect 177413 528314 177417 528348
rect 177748 528344 177809 528386
rect 177413 528298 177451 528314
rect 177485 528328 177699 528344
rect 177485 528310 177635 528328
rect 176833 528200 176929 528216
rect 176963 528200 176991 528234
rect 177025 528186 177059 528202
rect 176594 528072 176687 528088
rect 176628 528046 176687 528072
rect 176628 528038 176653 528046
rect 176481 528002 176560 528036
rect 176594 528012 176653 528038
rect 176594 528010 176687 528012
rect 176721 528152 177025 528166
rect 176721 528132 177059 528152
rect 176526 527976 176560 528002
rect 176721 527976 176755 528132
rect 177093 528098 177127 528236
rect 176827 528064 176843 528098
rect 176877 528064 177127 528098
rect 177165 528246 177207 528262
rect 177165 528212 177173 528246
rect 177165 528104 177207 528212
rect 177241 528198 177311 528262
rect 177241 528164 177269 528198
rect 177303 528182 177311 528198
rect 177241 528148 177277 528164
rect 177241 528138 177311 528148
rect 177345 528140 177379 528296
rect 177485 528264 177519 528310
rect 177669 528294 177699 528328
rect 177748 528310 177759 528344
rect 177793 528310 177809 528344
rect 177748 528294 177809 528310
rect 177843 528318 177894 528350
rect 177843 528294 177849 528318
rect 177413 528230 177519 528264
rect 177553 528250 177601 528276
rect 177413 528224 177457 528230
rect 177447 528190 177457 528224
rect 177587 528216 177601 528250
rect 177553 528196 177601 528216
rect 177413 528174 177457 528190
rect 177493 528187 177509 528196
rect 177543 528162 177601 528196
rect 177527 528153 177601 528162
rect 177345 528106 177426 528140
rect 177493 528122 177601 528153
rect 177635 528239 177699 528294
rect 177883 528284 177894 528318
rect 177877 528260 177894 528284
rect 177843 528244 177894 528260
rect 177635 528204 177700 528239
rect 177635 528188 177818 528204
rect 177635 528154 177784 528188
rect 177635 528144 177818 528154
rect 177670 528138 177818 528144
rect 177165 528072 177300 528104
rect 177392 528088 177426 528106
rect 177165 528070 177308 528072
rect 177093 528036 177127 528064
rect 177266 528046 177308 528070
rect 176442 527952 176492 527968
rect 176442 527918 176458 527952
rect 176442 527876 176492 527918
rect 176526 527960 176576 527976
rect 176526 527926 176542 527960
rect 176526 527910 176576 527926
rect 176619 527954 176755 527976
rect 176619 527920 176635 527954
rect 176669 527920 176755 527954
rect 176789 527996 177004 528030
rect 177093 528002 177205 528036
rect 177266 528012 177277 528046
rect 177342 528038 177358 528072
rect 177311 528012 177358 528038
rect 177392 528054 177586 528088
rect 177620 528054 177636 528088
rect 176789 527978 176823 527996
rect 176970 527978 177004 527996
rect 176789 527928 176823 527944
rect 176870 527928 176886 527962
rect 176920 527928 176936 527962
rect 176970 527928 177004 527944
rect 177063 527952 177137 527968
rect 176619 527910 176755 527920
rect 176870 527876 176936 527928
rect 177063 527918 177083 527952
rect 177117 527918 177137 527952
rect 177063 527876 177137 527918
rect 177171 527960 177205 528002
rect 177392 527978 177426 528054
rect 177670 528020 177704 528138
rect 177852 528114 177894 528244
rect 177171 527910 177205 527926
rect 177252 527953 177426 527978
rect 177544 527986 177704 528020
rect 177748 528020 177809 528104
rect 177748 527986 177759 528020
rect 177793 527986 177809 528020
rect 177544 527978 177578 527986
rect 177252 527919 177268 527953
rect 177302 527919 177426 527953
rect 177252 527910 177426 527919
rect 177460 527952 177510 527968
rect 177494 527918 177510 527952
rect 177748 527952 177809 527986
rect 177544 527928 177578 527944
rect 177460 527876 177510 527918
rect 177614 527918 177630 527952
rect 177664 527918 177680 527952
rect 177614 527876 177680 527918
rect 177748 527918 177759 527952
rect 177793 527918 177809 527952
rect 177843 528056 177894 528114
rect 177877 528022 177894 528056
rect 177843 527988 177894 528022
rect 177877 527954 177894 527988
rect 177843 527938 177894 527954
rect 177929 528314 177981 528352
rect 177929 528280 177947 528314
rect 178017 528344 178083 528386
rect 178017 528310 178033 528344
rect 178067 528310 178083 528344
rect 178119 528331 178153 528352
rect 177929 528251 177981 528280
rect 178119 528276 178153 528297
rect 177929 528091 177963 528251
rect 178020 528242 178153 528276
rect 178205 528325 178907 528386
rect 178205 528291 178223 528325
rect 178257 528291 178855 528325
rect 178889 528291 178907 528325
rect 178020 528191 178054 528242
rect 178205 528232 178907 528291
rect 178942 528325 178993 528352
rect 178942 528318 178959 528325
rect 178942 528284 178953 528318
rect 179027 528344 179093 528386
rect 179027 528310 179043 528344
rect 179077 528310 179093 528344
rect 179027 528306 179093 528310
rect 179178 528329 179284 528352
rect 178987 528284 178993 528291
rect 178942 528238 178993 528284
rect 179178 528295 179250 528329
rect 179178 528279 179284 528295
rect 179178 528272 179213 528279
rect 179027 528238 179213 528272
rect 177997 528175 178054 528191
rect 178031 528141 178054 528175
rect 177997 528125 178054 528141
rect 178101 528188 178167 528206
rect 178101 528154 178117 528188
rect 178151 528182 178167 528188
rect 178101 528148 178125 528154
rect 178159 528148 178167 528182
rect 178101 528132 178167 528148
rect 178205 528162 178535 528232
rect 178205 528128 178283 528162
rect 178317 528128 178382 528162
rect 178416 528128 178481 528162
rect 178515 528128 178535 528162
rect 178569 528164 178589 528198
rect 178623 528164 178692 528198
rect 178726 528164 178795 528198
rect 178829 528164 178907 528198
rect 178020 528096 178054 528125
rect 177929 528046 177983 528091
rect 178020 528062 178153 528096
rect 178569 528094 178907 528164
rect 177929 528012 177941 528046
rect 177975 528041 177983 528046
rect 177929 528007 177947 528012
rect 177981 528007 177983 528041
rect 178119 528028 178153 528062
rect 177929 527960 177983 528007
rect 177748 527876 177809 527918
rect 177929 527926 177947 527960
rect 177981 527926 177983 527960
rect 177929 527910 177983 527926
rect 178017 527994 178033 528028
rect 178067 527994 178083 528028
rect 178017 527960 178083 527994
rect 178017 527926 178033 527960
rect 178067 527926 178083 527960
rect 178017 527876 178083 527926
rect 178119 527960 178153 527994
rect 178119 527910 178153 527926
rect 178205 528054 178907 528094
rect 178205 528020 178223 528054
rect 178257 528020 178855 528054
rect 178889 528020 178907 528054
rect 178205 527952 178907 528020
rect 178205 527918 178223 527952
rect 178257 527918 178855 527952
rect 178889 527918 178907 527952
rect 178205 527876 178907 527918
rect 178942 528104 178976 528238
rect 179027 528204 179061 528238
rect 179010 528188 179061 528204
rect 179044 528154 179061 528188
rect 179010 528138 179061 528154
rect 179106 528188 179145 528204
rect 179140 528154 179145 528188
rect 179106 528138 179145 528154
rect 178942 528088 179009 528104
rect 178942 528054 178959 528088
rect 178993 528054 179009 528088
rect 178942 528020 179009 528054
rect 178942 527986 178959 528020
rect 178993 527986 179009 528020
rect 178942 527952 179009 527986
rect 178942 527918 178959 527952
rect 178993 527918 179009 527952
rect 178942 527910 179009 527918
rect 179043 528088 179077 528104
rect 179043 528020 179077 528054
rect 179043 527952 179077 527986
rect 179043 527876 179077 527918
rect 179111 527944 179145 528138
rect 179179 528012 179213 528238
rect 179247 528224 179281 528240
rect 179247 528080 179281 528190
rect 179322 528224 179377 528352
rect 179322 528190 179343 528224
rect 179322 528182 179377 528190
rect 179355 528148 179377 528182
rect 179322 528120 179377 528148
rect 179411 528318 179449 528352
rect 179411 528284 179413 528318
rect 179447 528284 179449 528318
rect 179411 528111 179449 528284
rect 179485 528329 179587 528386
rect 179519 528295 179553 528329
rect 179485 528279 179587 528295
rect 179631 528329 179680 528345
rect 179631 528295 179637 528329
rect 179671 528295 179680 528329
rect 179631 528224 179680 528295
rect 179953 528292 180011 528386
rect 179953 528258 179965 528292
rect 179999 528258 180011 528292
rect 179953 528241 180011 528258
rect 180045 528325 180747 528386
rect 180045 528291 180063 528325
rect 180097 528291 180695 528325
rect 180729 528291 180747 528325
rect 180045 528232 180747 528291
rect 180966 528325 181017 528352
rect 180966 528318 180983 528325
rect 180966 528284 180977 528318
rect 181051 528344 181117 528386
rect 181051 528310 181067 528344
rect 181101 528310 181117 528344
rect 181051 528306 181117 528310
rect 181202 528329 181308 528352
rect 181011 528284 181017 528291
rect 180966 528238 181017 528284
rect 181202 528295 181274 528329
rect 181202 528279 181308 528295
rect 181202 528272 181237 528279
rect 181051 528238 181237 528272
rect 179489 528190 179505 528224
rect 179539 528190 179735 528224
rect 179411 528080 179415 528111
rect 179247 528077 179415 528080
rect 179247 528046 179449 528077
rect 179483 528114 179633 528115
rect 179483 528080 179505 528114
rect 179539 528111 179633 528114
rect 179539 528080 179583 528111
rect 179483 528077 179583 528080
rect 179617 528077 179633 528111
rect 179179 527978 179279 528012
rect 179313 527978 179354 528012
rect 179388 527978 179404 528012
rect 179483 527944 179517 528077
rect 179667 528028 179735 528190
rect 180045 528162 180375 528232
rect 180045 528128 180123 528162
rect 180157 528128 180222 528162
rect 180256 528128 180321 528162
rect 180355 528128 180375 528162
rect 180409 528164 180429 528198
rect 180463 528164 180532 528198
rect 180566 528164 180635 528198
rect 180669 528164 180747 528198
rect 179111 527910 179517 527944
rect 179551 528012 179585 528028
rect 179551 527876 179585 527978
rect 179632 528012 179735 528028
rect 179632 527978 179637 528012
rect 179671 527978 179735 528012
rect 179632 527946 179735 527978
rect 179953 528074 180011 528109
rect 180409 528094 180747 528164
rect 179953 528040 179965 528074
rect 179999 528040 180011 528074
rect 179953 527981 180011 528040
rect 179953 527947 179965 527981
rect 179999 527947 180011 527981
rect 179953 527876 180011 527947
rect 180045 528054 180747 528094
rect 180045 528020 180063 528054
rect 180097 528020 180695 528054
rect 180729 528020 180747 528054
rect 180045 527952 180747 528020
rect 180045 527918 180063 527952
rect 180097 527918 180695 527952
rect 180729 527918 180747 527952
rect 180045 527876 180747 527918
rect 180966 528104 181000 528238
rect 181051 528204 181085 528238
rect 181034 528188 181085 528204
rect 181068 528154 181085 528188
rect 181034 528138 181085 528154
rect 181130 528188 181169 528204
rect 181164 528154 181169 528188
rect 181130 528138 181169 528154
rect 180966 528088 181033 528104
rect 180966 528054 180983 528088
rect 181017 528054 181033 528088
rect 180966 528020 181033 528054
rect 180966 527986 180983 528020
rect 181017 527986 181033 528020
rect 180966 527952 181033 527986
rect 180966 527918 180983 527952
rect 181017 527918 181033 527952
rect 180966 527910 181033 527918
rect 181067 528088 181101 528104
rect 181067 528020 181101 528054
rect 181067 527952 181101 527986
rect 181067 527876 181101 527918
rect 181135 527944 181169 528138
rect 181203 528012 181237 528238
rect 181271 528224 181305 528240
rect 181271 528080 181305 528190
rect 181346 528224 181401 528352
rect 181346 528190 181367 528224
rect 181346 528182 181401 528190
rect 181379 528148 181401 528182
rect 181346 528120 181401 528148
rect 181435 528318 181473 528352
rect 181435 528284 181437 528318
rect 181471 528284 181473 528318
rect 181435 528111 181473 528284
rect 181509 528329 181611 528386
rect 181543 528295 181577 528329
rect 181509 528279 181611 528295
rect 181655 528329 181704 528345
rect 181655 528295 181661 528329
rect 181695 528295 181704 528329
rect 181655 528224 181704 528295
rect 181793 528325 182862 528386
rect 181793 528291 181811 528325
rect 181845 528291 182811 528325
rect 182845 528291 182862 528325
rect 181793 528277 182862 528291
rect 182897 528325 183966 528386
rect 182897 528291 182915 528325
rect 182949 528291 183915 528325
rect 183949 528291 183966 528325
rect 182897 528277 183966 528291
rect 184001 528325 185070 528386
rect 184001 528291 184019 528325
rect 184053 528291 185019 528325
rect 185053 528291 185070 528325
rect 184001 528277 185070 528291
rect 185105 528292 185163 528386
rect 181513 528190 181529 528224
rect 181563 528190 181759 528224
rect 181435 528080 181439 528111
rect 181271 528077 181439 528080
rect 181271 528046 181473 528077
rect 181507 528114 181657 528115
rect 181507 528080 181529 528114
rect 181563 528111 181657 528114
rect 181563 528080 181607 528111
rect 181507 528077 181607 528080
rect 181641 528077 181657 528111
rect 181203 527978 181303 528012
rect 181337 527978 181378 528012
rect 181412 527978 181428 528012
rect 181507 527944 181541 528077
rect 181691 528028 181759 528190
rect 182110 528162 182178 528277
rect 182110 528128 182127 528162
rect 182161 528128 182178 528162
rect 182110 528111 182178 528128
rect 182474 528198 182544 528213
rect 182474 528164 182491 528198
rect 182525 528164 182544 528198
rect 181135 527910 181541 527944
rect 181575 528012 181609 528028
rect 181575 527876 181609 527978
rect 181656 528012 181759 528028
rect 181656 527978 181661 528012
rect 181695 527978 181759 528012
rect 181656 527946 181759 527978
rect 182474 527963 182544 528164
rect 183214 528162 183282 528277
rect 183214 528128 183231 528162
rect 183265 528128 183282 528162
rect 183214 528111 183282 528128
rect 183578 528198 183648 528213
rect 183578 528164 183595 528198
rect 183629 528164 183648 528198
rect 183578 527963 183648 528164
rect 184318 528162 184386 528277
rect 185105 528258 185117 528292
rect 185151 528258 185163 528292
rect 185197 528325 186266 528386
rect 185197 528291 185215 528325
rect 185249 528291 186215 528325
rect 186249 528291 186266 528325
rect 185197 528277 186266 528291
rect 186301 528325 187003 528386
rect 186301 528291 186319 528325
rect 186353 528291 186951 528325
rect 186985 528291 187003 528325
rect 185105 528241 185163 528258
rect 184318 528128 184335 528162
rect 184369 528128 184386 528162
rect 184318 528111 184386 528128
rect 184682 528198 184752 528213
rect 184682 528164 184699 528198
rect 184733 528164 184752 528198
rect 184682 527963 184752 528164
rect 185514 528162 185582 528277
rect 186301 528232 187003 528291
rect 187221 528323 187463 528386
rect 187221 528289 187239 528323
rect 187273 528289 187411 528323
rect 187445 528289 187463 528323
rect 187221 528236 187463 528289
rect 185514 528128 185531 528162
rect 185565 528128 185582 528162
rect 185514 528111 185582 528128
rect 185878 528198 185948 528213
rect 185878 528164 185895 528198
rect 185929 528164 185948 528198
rect 185105 528074 185163 528109
rect 185105 528040 185117 528074
rect 185151 528040 185163 528074
rect 185105 527981 185163 528040
rect 181793 527952 182862 527963
rect 181793 527918 181811 527952
rect 181845 527918 182811 527952
rect 182845 527918 182862 527952
rect 181793 527876 182862 527918
rect 182897 527952 183966 527963
rect 182897 527918 182915 527952
rect 182949 527918 183915 527952
rect 183949 527918 183966 527952
rect 182897 527876 183966 527918
rect 184001 527952 185070 527963
rect 184001 527918 184019 527952
rect 184053 527918 185019 527952
rect 185053 527918 185070 527952
rect 184001 527876 185070 527918
rect 185105 527947 185117 527981
rect 185151 527947 185163 527981
rect 185878 527963 185948 528164
rect 186301 528162 186631 528232
rect 186301 528128 186379 528162
rect 186413 528128 186478 528162
rect 186512 528128 186577 528162
rect 186611 528128 186631 528162
rect 186665 528164 186685 528198
rect 186719 528164 186788 528198
rect 186822 528164 186891 528198
rect 186925 528164 187003 528198
rect 186665 528094 187003 528164
rect 186301 528054 187003 528094
rect 186301 528020 186319 528054
rect 186353 528020 186951 528054
rect 186985 528020 187003 528054
rect 185105 527876 185163 527947
rect 185197 527952 186266 527963
rect 185197 527918 185215 527952
rect 185249 527918 186215 527952
rect 186249 527918 186266 527952
rect 185197 527876 186266 527918
rect 186301 527952 187003 528020
rect 186301 527918 186319 527952
rect 186353 527918 186951 527952
rect 186985 527918 187003 527952
rect 186301 527876 187003 527918
rect 187221 528168 187271 528202
rect 187305 528168 187325 528202
rect 187221 528094 187325 528168
rect 187359 528162 187463 528236
rect 187359 528128 187379 528162
rect 187413 528128 187463 528162
rect 187221 528047 187463 528094
rect 187221 528013 187239 528047
rect 187273 528013 187411 528047
rect 187445 528013 187463 528047
rect 187221 527952 187463 528013
rect 187221 527918 187239 527952
rect 187273 527918 187411 527952
rect 187445 527918 187463 527952
rect 187221 527876 187463 527918
rect 172208 527842 172237 527876
rect 172271 527842 172329 527876
rect 172363 527842 172421 527876
rect 172455 527842 172513 527876
rect 172547 527842 172605 527876
rect 172639 527842 172697 527876
rect 172731 527842 172789 527876
rect 172823 527842 172881 527876
rect 172915 527842 172973 527876
rect 173007 527842 173065 527876
rect 173099 527842 173157 527876
rect 173191 527842 173249 527876
rect 173283 527842 173341 527876
rect 173375 527842 173433 527876
rect 173467 527842 173525 527876
rect 173559 527842 173617 527876
rect 173651 527842 173709 527876
rect 173743 527842 173801 527876
rect 173835 527842 173893 527876
rect 173927 527842 173985 527876
rect 174019 527842 174077 527876
rect 174111 527842 174169 527876
rect 174203 527842 174261 527876
rect 174295 527842 174353 527876
rect 174387 527842 174445 527876
rect 174479 527842 174537 527876
rect 174571 527842 174629 527876
rect 174663 527842 174721 527876
rect 174755 527842 174813 527876
rect 174847 527842 174905 527876
rect 174939 527842 174997 527876
rect 175031 527842 175089 527876
rect 175123 527842 175181 527876
rect 175215 527842 175273 527876
rect 175307 527842 175365 527876
rect 175399 527842 175457 527876
rect 175491 527842 175549 527876
rect 175583 527842 175641 527876
rect 175675 527842 175733 527876
rect 175767 527842 175825 527876
rect 175859 527842 175917 527876
rect 175951 527842 176009 527876
rect 176043 527842 176101 527876
rect 176135 527842 176193 527876
rect 176227 527842 176285 527876
rect 176319 527842 176377 527876
rect 176411 527842 176469 527876
rect 176503 527842 176561 527876
rect 176595 527842 176653 527876
rect 176687 527842 176745 527876
rect 176779 527842 176837 527876
rect 176871 527842 176929 527876
rect 176963 527842 177021 527876
rect 177055 527842 177113 527876
rect 177147 527842 177205 527876
rect 177239 527842 177297 527876
rect 177331 527842 177389 527876
rect 177423 527842 177481 527876
rect 177515 527842 177573 527876
rect 177607 527842 177665 527876
rect 177699 527842 177757 527876
rect 177791 527842 177849 527876
rect 177883 527842 177941 527876
rect 177975 527842 178033 527876
rect 178067 527842 178125 527876
rect 178159 527842 178217 527876
rect 178251 527842 178309 527876
rect 178343 527842 178401 527876
rect 178435 527842 178493 527876
rect 178527 527842 178585 527876
rect 178619 527842 178677 527876
rect 178711 527842 178769 527876
rect 178803 527842 178861 527876
rect 178895 527842 178953 527876
rect 178987 527842 179045 527876
rect 179079 527842 179137 527876
rect 179171 527842 179229 527876
rect 179263 527842 179321 527876
rect 179355 527842 179413 527876
rect 179447 527842 179505 527876
rect 179539 527842 179597 527876
rect 179631 527842 179689 527876
rect 179723 527842 179781 527876
rect 179815 527842 179873 527876
rect 179907 527842 179965 527876
rect 179999 527842 180057 527876
rect 180091 527842 180149 527876
rect 180183 527842 180241 527876
rect 180275 527842 180333 527876
rect 180367 527842 180425 527876
rect 180459 527842 180517 527876
rect 180551 527842 180609 527876
rect 180643 527842 180701 527876
rect 180735 527842 180793 527876
rect 180827 527842 180885 527876
rect 180919 527842 180977 527876
rect 181011 527842 181069 527876
rect 181103 527842 181161 527876
rect 181195 527842 181253 527876
rect 181287 527842 181345 527876
rect 181379 527842 181437 527876
rect 181471 527842 181529 527876
rect 181563 527842 181621 527876
rect 181655 527842 181713 527876
rect 181747 527842 181805 527876
rect 181839 527842 181897 527876
rect 181931 527842 181989 527876
rect 182023 527842 182081 527876
rect 182115 527842 182173 527876
rect 182207 527842 182265 527876
rect 182299 527842 182357 527876
rect 182391 527842 182449 527876
rect 182483 527842 182541 527876
rect 182575 527842 182633 527876
rect 182667 527842 182725 527876
rect 182759 527842 182817 527876
rect 182851 527842 182909 527876
rect 182943 527842 183001 527876
rect 183035 527842 183093 527876
rect 183127 527842 183185 527876
rect 183219 527842 183277 527876
rect 183311 527842 183369 527876
rect 183403 527842 183461 527876
rect 183495 527842 183553 527876
rect 183587 527842 183645 527876
rect 183679 527842 183737 527876
rect 183771 527842 183829 527876
rect 183863 527842 183921 527876
rect 183955 527842 184013 527876
rect 184047 527842 184105 527876
rect 184139 527842 184197 527876
rect 184231 527842 184289 527876
rect 184323 527842 184381 527876
rect 184415 527842 184473 527876
rect 184507 527842 184565 527876
rect 184599 527842 184657 527876
rect 184691 527842 184749 527876
rect 184783 527842 184841 527876
rect 184875 527842 184933 527876
rect 184967 527842 185025 527876
rect 185059 527842 185117 527876
rect 185151 527842 185209 527876
rect 185243 527842 185301 527876
rect 185335 527842 185393 527876
rect 185427 527842 185485 527876
rect 185519 527842 185577 527876
rect 185611 527842 185669 527876
rect 185703 527842 185761 527876
rect 185795 527842 185853 527876
rect 185887 527842 185945 527876
rect 185979 527842 186037 527876
rect 186071 527842 186129 527876
rect 186163 527842 186221 527876
rect 186255 527842 186313 527876
rect 186347 527842 186405 527876
rect 186439 527842 186497 527876
rect 186531 527842 186589 527876
rect 186623 527842 186681 527876
rect 186715 527842 186773 527876
rect 186807 527842 186865 527876
rect 186899 527842 186957 527876
rect 186991 527842 187049 527876
rect 187083 527842 187141 527876
rect 187175 527842 187233 527876
rect 187267 527842 187325 527876
rect 187359 527842 187417 527876
rect 187451 527842 187480 527876
rect 172225 527800 172467 527842
rect 172225 527766 172243 527800
rect 172277 527766 172415 527800
rect 172449 527766 172467 527800
rect 172225 527705 172467 527766
rect 172501 527800 173570 527842
rect 172501 527766 172519 527800
rect 172553 527766 173519 527800
rect 173553 527766 173570 527800
rect 172501 527755 173570 527766
rect 173605 527800 174674 527842
rect 173605 527766 173623 527800
rect 173657 527766 174623 527800
rect 174657 527766 174674 527800
rect 173605 527755 174674 527766
rect 174709 527800 175778 527842
rect 174709 527766 174727 527800
rect 174761 527766 175727 527800
rect 175761 527766 175778 527800
rect 174709 527755 175778 527766
rect 175813 527800 176331 527842
rect 175813 527766 175831 527800
rect 175865 527766 176279 527800
rect 176313 527766 176331 527800
rect 172225 527671 172243 527705
rect 172277 527671 172415 527705
rect 172449 527671 172467 527705
rect 172225 527624 172467 527671
rect 172225 527556 172275 527590
rect 172309 527556 172329 527590
rect 172225 527482 172329 527556
rect 172363 527550 172467 527624
rect 172363 527516 172383 527550
rect 172417 527516 172467 527550
rect 172818 527590 172886 527607
rect 172818 527556 172835 527590
rect 172869 527556 172886 527590
rect 172225 527429 172467 527482
rect 172818 527441 172886 527556
rect 173182 527554 173252 527755
rect 173182 527520 173199 527554
rect 173233 527520 173252 527554
rect 173182 527505 173252 527520
rect 173922 527590 173990 527607
rect 173922 527556 173939 527590
rect 173973 527556 173990 527590
rect 173922 527441 173990 527556
rect 174286 527554 174356 527755
rect 174286 527520 174303 527554
rect 174337 527520 174356 527554
rect 174286 527505 174356 527520
rect 175026 527590 175094 527607
rect 175026 527556 175043 527590
rect 175077 527556 175094 527590
rect 175026 527441 175094 527556
rect 175390 527554 175460 527755
rect 175813 527698 176331 527766
rect 175813 527664 175831 527698
rect 175865 527664 176279 527698
rect 176313 527664 176331 527698
rect 175813 527624 176331 527664
rect 175390 527520 175407 527554
rect 175441 527520 175460 527554
rect 175390 527505 175460 527520
rect 175813 527556 175891 527590
rect 175925 527556 176001 527590
rect 176035 527556 176055 527590
rect 175813 527486 176055 527556
rect 176089 527554 176331 527624
rect 176089 527520 176109 527554
rect 176143 527520 176219 527554
rect 176253 527520 176331 527554
rect 176365 527774 176442 527808
rect 176365 527740 176377 527774
rect 176436 527740 176442 527774
rect 176476 527800 176541 527842
rect 176476 527766 176492 527800
rect 176526 527766 176541 527800
rect 176476 527750 176541 527766
rect 176645 527774 176701 527808
rect 176365 527614 176442 527740
rect 176645 527740 176651 527774
rect 176685 527740 176701 527774
rect 176645 527716 176701 527740
rect 176476 527672 176701 527716
rect 176739 527774 176819 527808
rect 176739 527740 176755 527774
rect 176789 527740 176819 527774
rect 176899 527800 176953 527842
rect 176899 527766 176909 527800
rect 176943 527766 176953 527800
rect 176899 527750 176953 527766
rect 176987 527774 177044 527808
rect 172225 527395 172243 527429
rect 172277 527395 172415 527429
rect 172449 527395 172467 527429
rect 172225 527332 172467 527395
rect 172501 527427 173570 527441
rect 172501 527393 172519 527427
rect 172553 527393 173519 527427
rect 173553 527393 173570 527427
rect 172501 527332 173570 527393
rect 173605 527427 174674 527441
rect 173605 527393 173623 527427
rect 173657 527393 174623 527427
rect 174657 527393 174674 527427
rect 173605 527332 174674 527393
rect 174709 527427 175778 527441
rect 174709 527393 174727 527427
rect 174761 527393 175727 527427
rect 175761 527393 175778 527427
rect 174709 527332 175778 527393
rect 175813 527427 176331 527486
rect 175813 527393 175831 527427
rect 175865 527393 176279 527427
rect 176313 527393 176331 527427
rect 175813 527332 176331 527393
rect 176365 527480 176421 527614
rect 176476 527580 176566 527672
rect 176739 527638 176819 527740
rect 176987 527740 176993 527774
rect 177027 527740 177044 527774
rect 176987 527716 177044 527740
rect 176455 527564 176566 527580
rect 176489 527530 176566 527564
rect 176455 527514 176566 527530
rect 176600 527564 176819 527638
rect 176600 527530 176651 527564
rect 176685 527530 176819 527564
rect 176600 527526 176819 527530
rect 176476 527492 176566 527514
rect 176365 527434 176442 527480
rect 176476 527458 176701 527492
rect 176365 527400 176402 527434
rect 176436 527400 176442 527434
rect 176645 527434 176701 527458
rect 176365 527366 176442 527400
rect 176476 527408 176541 527424
rect 176476 527374 176492 527408
rect 176526 527374 176541 527408
rect 176476 527332 176541 527374
rect 176645 527400 176651 527434
rect 176685 527400 176701 527434
rect 176645 527366 176701 527400
rect 176739 527434 176819 527526
rect 176853 527672 177044 527716
rect 177101 527800 177343 527842
rect 177101 527766 177119 527800
rect 177153 527766 177291 527800
rect 177325 527766 177343 527800
rect 177101 527705 177343 527766
rect 176853 527564 176895 527672
rect 177101 527671 177119 527705
rect 177153 527671 177291 527705
rect 177325 527671 177343 527705
rect 176853 527530 176855 527564
rect 176889 527530 176895 527564
rect 176853 527492 176895 527530
rect 176929 527604 177021 527638
rect 177055 527604 177067 527638
rect 177101 527624 177343 527671
rect 176929 527564 177067 527604
rect 176929 527530 176969 527564
rect 177003 527530 177067 527564
rect 176929 527526 177067 527530
rect 177101 527556 177151 527590
rect 177185 527556 177205 527590
rect 176853 527458 177044 527492
rect 176739 527400 176755 527434
rect 176789 527400 176819 527434
rect 176987 527434 177044 527458
rect 176739 527366 176819 527400
rect 176899 527408 176953 527424
rect 176899 527374 176909 527408
rect 176943 527374 176953 527408
rect 176899 527332 176953 527374
rect 176987 527400 176993 527434
rect 177027 527400 177044 527434
rect 176987 527366 177044 527400
rect 177101 527482 177205 527556
rect 177239 527550 177343 527624
rect 177377 527771 177435 527842
rect 177377 527737 177389 527771
rect 177423 527737 177435 527771
rect 177469 527800 178538 527842
rect 177469 527766 177487 527800
rect 177521 527766 178487 527800
rect 178521 527766 178538 527800
rect 177469 527755 178538 527766
rect 178573 527800 178907 527842
rect 178573 527766 178591 527800
rect 178625 527766 178855 527800
rect 178889 527766 178907 527800
rect 177377 527678 177435 527737
rect 177377 527644 177389 527678
rect 177423 527644 177435 527678
rect 177377 527609 177435 527644
rect 177239 527516 177259 527550
rect 177293 527516 177343 527550
rect 177786 527590 177854 527607
rect 177786 527556 177803 527590
rect 177837 527556 177854 527590
rect 177101 527429 177343 527482
rect 177101 527395 177119 527429
rect 177153 527395 177291 527429
rect 177325 527395 177343 527429
rect 177101 527332 177343 527395
rect 177377 527460 177435 527477
rect 177377 527426 177389 527460
rect 177423 527426 177435 527460
rect 177786 527441 177854 527556
rect 178150 527554 178220 527755
rect 178573 527698 178907 527766
rect 178573 527664 178591 527698
rect 178625 527664 178855 527698
rect 178889 527664 178907 527698
rect 178573 527624 178907 527664
rect 178150 527520 178167 527554
rect 178201 527520 178220 527554
rect 178150 527505 178220 527520
rect 178573 527556 178593 527590
rect 178627 527556 178723 527590
rect 178573 527486 178723 527556
rect 178757 527554 178907 527624
rect 178757 527520 178853 527554
rect 178887 527520 178907 527554
rect 178941 527774 179018 527808
rect 178941 527740 178953 527774
rect 179012 527740 179018 527774
rect 179052 527800 179117 527842
rect 179052 527766 179068 527800
rect 179102 527766 179117 527800
rect 179052 527750 179117 527766
rect 179221 527774 179277 527808
rect 178941 527614 179018 527740
rect 179221 527740 179227 527774
rect 179261 527740 179277 527774
rect 179221 527716 179277 527740
rect 179052 527672 179277 527716
rect 179315 527774 179395 527808
rect 179315 527740 179331 527774
rect 179365 527740 179395 527774
rect 179475 527800 179529 527842
rect 179475 527766 179485 527800
rect 179519 527766 179529 527800
rect 179475 527750 179529 527766
rect 179563 527774 179620 527808
rect 177377 527332 177435 527426
rect 177469 527427 178538 527441
rect 177469 527393 177487 527427
rect 177521 527393 178487 527427
rect 178521 527393 178538 527427
rect 177469 527332 178538 527393
rect 178573 527434 178907 527486
rect 178573 527400 178591 527434
rect 178625 527400 178855 527434
rect 178889 527400 178907 527434
rect 178573 527332 178907 527400
rect 178941 527480 178997 527614
rect 179052 527580 179142 527672
rect 179315 527638 179395 527740
rect 179563 527740 179569 527774
rect 179603 527740 179620 527774
rect 179677 527800 180746 527842
rect 179677 527766 179695 527800
rect 179729 527766 180695 527800
rect 180729 527766 180746 527800
rect 179677 527755 180746 527766
rect 180781 527800 181850 527842
rect 180781 527766 180799 527800
rect 180833 527766 181799 527800
rect 181833 527766 181850 527800
rect 180781 527755 181850 527766
rect 181885 527800 182403 527842
rect 181885 527766 181903 527800
rect 181937 527766 182351 527800
rect 182385 527766 182403 527800
rect 179563 527716 179620 527740
rect 179031 527564 179142 527580
rect 179065 527530 179142 527564
rect 179031 527514 179142 527530
rect 179176 527564 179395 527638
rect 179176 527530 179227 527564
rect 179261 527530 179395 527564
rect 179176 527526 179395 527530
rect 179052 527492 179142 527514
rect 178941 527434 179018 527480
rect 179052 527458 179277 527492
rect 178941 527400 178978 527434
rect 179012 527400 179018 527434
rect 179221 527434 179277 527458
rect 178941 527366 179018 527400
rect 179052 527408 179117 527424
rect 179052 527374 179068 527408
rect 179102 527374 179117 527408
rect 179052 527332 179117 527374
rect 179221 527400 179227 527434
rect 179261 527400 179277 527434
rect 179221 527366 179277 527400
rect 179315 527434 179395 527526
rect 179429 527672 179620 527716
rect 179429 527564 179471 527672
rect 179429 527530 179431 527564
rect 179465 527530 179471 527564
rect 179429 527492 179471 527530
rect 179539 527604 179643 527638
rect 179505 527564 179643 527604
rect 179505 527530 179545 527564
rect 179579 527530 179643 527564
rect 179505 527526 179643 527530
rect 179994 527590 180062 527607
rect 179994 527556 180011 527590
rect 180045 527556 180062 527590
rect 179429 527458 179620 527492
rect 179315 527400 179331 527434
rect 179365 527400 179395 527434
rect 179563 527434 179620 527458
rect 179994 527441 180062 527556
rect 180358 527554 180428 527755
rect 180358 527520 180375 527554
rect 180409 527520 180428 527554
rect 180358 527505 180428 527520
rect 181098 527590 181166 527607
rect 181098 527556 181115 527590
rect 181149 527556 181166 527590
rect 181098 527441 181166 527556
rect 181462 527554 181532 527755
rect 181885 527698 182403 527766
rect 181885 527664 181903 527698
rect 181937 527664 182351 527698
rect 182385 527664 182403 527698
rect 181885 527624 182403 527664
rect 181462 527520 181479 527554
rect 181513 527520 181532 527554
rect 181462 527505 181532 527520
rect 181885 527556 181963 527590
rect 181997 527556 182073 527590
rect 182107 527556 182127 527590
rect 181885 527486 182127 527556
rect 182161 527554 182403 527624
rect 182529 527771 182587 527842
rect 182529 527737 182541 527771
rect 182575 527737 182587 527771
rect 182621 527800 183690 527842
rect 182621 527766 182639 527800
rect 182673 527766 183639 527800
rect 183673 527766 183690 527800
rect 182621 527755 183690 527766
rect 183725 527800 184794 527842
rect 183725 527766 183743 527800
rect 183777 527766 184743 527800
rect 184777 527766 184794 527800
rect 183725 527755 184794 527766
rect 184829 527800 185898 527842
rect 184829 527766 184847 527800
rect 184881 527766 185847 527800
rect 185881 527766 185898 527800
rect 184829 527755 185898 527766
rect 185933 527800 187002 527842
rect 185933 527766 185951 527800
rect 185985 527766 186951 527800
rect 186985 527766 187002 527800
rect 185933 527755 187002 527766
rect 187221 527800 187463 527842
rect 187221 527766 187239 527800
rect 187273 527766 187411 527800
rect 187445 527766 187463 527800
rect 182529 527678 182587 527737
rect 182529 527644 182541 527678
rect 182575 527644 182587 527678
rect 182529 527609 182587 527644
rect 182161 527520 182181 527554
rect 182215 527520 182291 527554
rect 182325 527520 182403 527554
rect 182938 527590 183006 527607
rect 182938 527556 182955 527590
rect 182989 527556 183006 527590
rect 179315 527366 179395 527400
rect 179475 527408 179529 527424
rect 179475 527374 179485 527408
rect 179519 527374 179529 527408
rect 179475 527332 179529 527374
rect 179563 527400 179569 527434
rect 179603 527400 179620 527434
rect 179563 527366 179620 527400
rect 179677 527427 180746 527441
rect 179677 527393 179695 527427
rect 179729 527393 180695 527427
rect 180729 527393 180746 527427
rect 179677 527332 180746 527393
rect 180781 527427 181850 527441
rect 180781 527393 180799 527427
rect 180833 527393 181799 527427
rect 181833 527393 181850 527427
rect 180781 527332 181850 527393
rect 181885 527427 182403 527486
rect 181885 527393 181903 527427
rect 181937 527393 182351 527427
rect 182385 527393 182403 527427
rect 181885 527332 182403 527393
rect 182529 527460 182587 527477
rect 182529 527426 182541 527460
rect 182575 527426 182587 527460
rect 182938 527441 183006 527556
rect 183302 527554 183372 527755
rect 183302 527520 183319 527554
rect 183353 527520 183372 527554
rect 183302 527505 183372 527520
rect 184042 527590 184110 527607
rect 184042 527556 184059 527590
rect 184093 527556 184110 527590
rect 184042 527441 184110 527556
rect 184406 527554 184476 527755
rect 184406 527520 184423 527554
rect 184457 527520 184476 527554
rect 184406 527505 184476 527520
rect 185146 527590 185214 527607
rect 185146 527556 185163 527590
rect 185197 527556 185214 527590
rect 185146 527441 185214 527556
rect 185510 527554 185580 527755
rect 185510 527520 185527 527554
rect 185561 527520 185580 527554
rect 185510 527505 185580 527520
rect 186250 527590 186318 527607
rect 186250 527556 186267 527590
rect 186301 527556 186318 527590
rect 186250 527441 186318 527556
rect 186614 527554 186684 527755
rect 186614 527520 186631 527554
rect 186665 527520 186684 527554
rect 186614 527505 186684 527520
rect 187221 527705 187463 527766
rect 187221 527671 187239 527705
rect 187273 527671 187411 527705
rect 187445 527671 187463 527705
rect 187221 527624 187463 527671
rect 187221 527550 187325 527624
rect 187221 527516 187271 527550
rect 187305 527516 187325 527550
rect 187359 527556 187379 527590
rect 187413 527556 187463 527590
rect 187359 527482 187463 527556
rect 182529 527332 182587 527426
rect 182621 527427 183690 527441
rect 182621 527393 182639 527427
rect 182673 527393 183639 527427
rect 183673 527393 183690 527427
rect 182621 527332 183690 527393
rect 183725 527427 184794 527441
rect 183725 527393 183743 527427
rect 183777 527393 184743 527427
rect 184777 527393 184794 527427
rect 183725 527332 184794 527393
rect 184829 527427 185898 527441
rect 184829 527393 184847 527427
rect 184881 527393 185847 527427
rect 185881 527393 185898 527427
rect 184829 527332 185898 527393
rect 185933 527427 187002 527441
rect 185933 527393 185951 527427
rect 185985 527393 186951 527427
rect 186985 527393 187002 527427
rect 185933 527332 187002 527393
rect 187221 527429 187463 527482
rect 187221 527395 187239 527429
rect 187273 527395 187411 527429
rect 187445 527395 187463 527429
rect 187221 527332 187463 527395
rect 172208 527298 172237 527332
rect 172271 527298 172329 527332
rect 172363 527298 172421 527332
rect 172455 527298 172513 527332
rect 172547 527298 172605 527332
rect 172639 527298 172697 527332
rect 172731 527298 172789 527332
rect 172823 527298 172881 527332
rect 172915 527298 172973 527332
rect 173007 527298 173065 527332
rect 173099 527298 173157 527332
rect 173191 527298 173249 527332
rect 173283 527298 173341 527332
rect 173375 527298 173433 527332
rect 173467 527298 173525 527332
rect 173559 527298 173617 527332
rect 173651 527298 173709 527332
rect 173743 527298 173801 527332
rect 173835 527298 173893 527332
rect 173927 527298 173985 527332
rect 174019 527298 174077 527332
rect 174111 527298 174169 527332
rect 174203 527298 174261 527332
rect 174295 527298 174353 527332
rect 174387 527298 174445 527332
rect 174479 527298 174537 527332
rect 174571 527298 174629 527332
rect 174663 527298 174721 527332
rect 174755 527298 174813 527332
rect 174847 527298 174905 527332
rect 174939 527298 174997 527332
rect 175031 527298 175089 527332
rect 175123 527298 175181 527332
rect 175215 527298 175273 527332
rect 175307 527298 175365 527332
rect 175399 527298 175457 527332
rect 175491 527298 175549 527332
rect 175583 527298 175641 527332
rect 175675 527298 175733 527332
rect 175767 527298 175825 527332
rect 175859 527298 175917 527332
rect 175951 527298 176009 527332
rect 176043 527298 176101 527332
rect 176135 527298 176193 527332
rect 176227 527298 176285 527332
rect 176319 527298 176377 527332
rect 176411 527298 176469 527332
rect 176503 527298 176561 527332
rect 176595 527298 176653 527332
rect 176687 527298 176745 527332
rect 176779 527298 176837 527332
rect 176871 527298 176929 527332
rect 176963 527298 177021 527332
rect 177055 527298 177113 527332
rect 177147 527298 177205 527332
rect 177239 527298 177297 527332
rect 177331 527298 177389 527332
rect 177423 527298 177481 527332
rect 177515 527298 177573 527332
rect 177607 527298 177665 527332
rect 177699 527298 177757 527332
rect 177791 527298 177849 527332
rect 177883 527298 177941 527332
rect 177975 527298 178033 527332
rect 178067 527298 178125 527332
rect 178159 527298 178217 527332
rect 178251 527298 178309 527332
rect 178343 527298 178401 527332
rect 178435 527298 178493 527332
rect 178527 527298 178585 527332
rect 178619 527298 178677 527332
rect 178711 527298 178769 527332
rect 178803 527298 178861 527332
rect 178895 527298 178953 527332
rect 178987 527298 179045 527332
rect 179079 527298 179137 527332
rect 179171 527298 179229 527332
rect 179263 527298 179321 527332
rect 179355 527298 179413 527332
rect 179447 527298 179505 527332
rect 179539 527298 179597 527332
rect 179631 527298 179689 527332
rect 179723 527298 179781 527332
rect 179815 527298 179873 527332
rect 179907 527298 179965 527332
rect 179999 527298 180057 527332
rect 180091 527298 180149 527332
rect 180183 527298 180241 527332
rect 180275 527298 180333 527332
rect 180367 527298 180425 527332
rect 180459 527298 180517 527332
rect 180551 527298 180609 527332
rect 180643 527298 180701 527332
rect 180735 527298 180793 527332
rect 180827 527298 180885 527332
rect 180919 527298 180977 527332
rect 181011 527298 181069 527332
rect 181103 527298 181161 527332
rect 181195 527298 181253 527332
rect 181287 527298 181345 527332
rect 181379 527298 181437 527332
rect 181471 527298 181529 527332
rect 181563 527298 181621 527332
rect 181655 527298 181713 527332
rect 181747 527298 181805 527332
rect 181839 527298 181897 527332
rect 181931 527298 181989 527332
rect 182023 527298 182081 527332
rect 182115 527298 182173 527332
rect 182207 527298 182265 527332
rect 182299 527298 182357 527332
rect 182391 527298 182449 527332
rect 182483 527298 182541 527332
rect 182575 527298 182633 527332
rect 182667 527298 182725 527332
rect 182759 527298 182817 527332
rect 182851 527298 182909 527332
rect 182943 527298 183001 527332
rect 183035 527298 183093 527332
rect 183127 527298 183185 527332
rect 183219 527298 183277 527332
rect 183311 527298 183369 527332
rect 183403 527298 183461 527332
rect 183495 527298 183553 527332
rect 183587 527298 183645 527332
rect 183679 527298 183737 527332
rect 183771 527298 183829 527332
rect 183863 527298 183921 527332
rect 183955 527298 184013 527332
rect 184047 527298 184105 527332
rect 184139 527298 184197 527332
rect 184231 527298 184289 527332
rect 184323 527298 184381 527332
rect 184415 527298 184473 527332
rect 184507 527298 184565 527332
rect 184599 527298 184657 527332
rect 184691 527298 184749 527332
rect 184783 527298 184841 527332
rect 184875 527298 184933 527332
rect 184967 527298 185025 527332
rect 185059 527298 185117 527332
rect 185151 527298 185209 527332
rect 185243 527298 185301 527332
rect 185335 527298 185393 527332
rect 185427 527298 185485 527332
rect 185519 527298 185577 527332
rect 185611 527298 185669 527332
rect 185703 527298 185761 527332
rect 185795 527298 185853 527332
rect 185887 527298 185945 527332
rect 185979 527298 186037 527332
rect 186071 527298 186129 527332
rect 186163 527298 186221 527332
rect 186255 527298 186313 527332
rect 186347 527298 186405 527332
rect 186439 527298 186497 527332
rect 186531 527298 186589 527332
rect 186623 527298 186681 527332
rect 186715 527298 186773 527332
rect 186807 527298 186865 527332
rect 186899 527298 186957 527332
rect 186991 527298 187049 527332
rect 187083 527298 187141 527332
rect 187175 527298 187233 527332
rect 187267 527298 187325 527332
rect 187359 527298 187417 527332
rect 187451 527298 187480 527332
rect 172225 527235 172467 527298
rect 172225 527201 172243 527235
rect 172277 527201 172415 527235
rect 172449 527201 172467 527235
rect 172225 527148 172467 527201
rect 172501 527237 173570 527298
rect 172501 527203 172519 527237
rect 172553 527203 173519 527237
rect 173553 527203 173570 527237
rect 172501 527189 173570 527203
rect 173605 527237 174674 527298
rect 173605 527203 173623 527237
rect 173657 527203 174623 527237
rect 174657 527203 174674 527237
rect 173605 527189 174674 527203
rect 174801 527204 174859 527298
rect 172225 527074 172329 527148
rect 172225 527040 172275 527074
rect 172309 527040 172329 527074
rect 172363 527080 172383 527114
rect 172417 527080 172467 527114
rect 172363 527006 172467 527080
rect 172818 527074 172886 527189
rect 172818 527040 172835 527074
rect 172869 527040 172886 527074
rect 172818 527023 172886 527040
rect 173182 527110 173252 527125
rect 173182 527076 173199 527110
rect 173233 527076 173252 527110
rect 172225 526959 172467 527006
rect 172225 526925 172243 526959
rect 172277 526925 172415 526959
rect 172449 526925 172467 526959
rect 172225 526864 172467 526925
rect 173182 526875 173252 527076
rect 173922 527074 173990 527189
rect 174801 527170 174813 527204
rect 174847 527170 174859 527204
rect 174893 527237 175962 527298
rect 174893 527203 174911 527237
rect 174945 527203 175911 527237
rect 175945 527203 175962 527237
rect 174893 527189 175962 527203
rect 175997 527237 177066 527298
rect 175997 527203 176015 527237
rect 176049 527203 177015 527237
rect 177049 527203 177066 527237
rect 175997 527189 177066 527203
rect 177101 527237 178170 527298
rect 177101 527203 177119 527237
rect 177153 527203 178119 527237
rect 178153 527203 178170 527237
rect 177101 527189 178170 527203
rect 178205 527237 179274 527298
rect 178205 527203 178223 527237
rect 178257 527203 179223 527237
rect 179257 527203 179274 527237
rect 178205 527189 179274 527203
rect 179309 527237 179827 527298
rect 179309 527203 179327 527237
rect 179361 527203 179775 527237
rect 179809 527203 179827 527237
rect 174801 527153 174859 527170
rect 173922 527040 173939 527074
rect 173973 527040 173990 527074
rect 173922 527023 173990 527040
rect 174286 527110 174356 527125
rect 174286 527076 174303 527110
rect 174337 527076 174356 527110
rect 174286 526875 174356 527076
rect 175210 527074 175278 527189
rect 175210 527040 175227 527074
rect 175261 527040 175278 527074
rect 175210 527023 175278 527040
rect 175574 527110 175644 527125
rect 175574 527076 175591 527110
rect 175625 527076 175644 527110
rect 174801 526986 174859 527021
rect 174801 526952 174813 526986
rect 174847 526952 174859 526986
rect 174801 526893 174859 526952
rect 172225 526830 172243 526864
rect 172277 526830 172415 526864
rect 172449 526830 172467 526864
rect 172225 526788 172467 526830
rect 172501 526864 173570 526875
rect 172501 526830 172519 526864
rect 172553 526830 173519 526864
rect 173553 526830 173570 526864
rect 172501 526788 173570 526830
rect 173605 526864 174674 526875
rect 173605 526830 173623 526864
rect 173657 526830 174623 526864
rect 174657 526830 174674 526864
rect 173605 526788 174674 526830
rect 174801 526859 174813 526893
rect 174847 526859 174859 526893
rect 175574 526875 175644 527076
rect 176314 527074 176382 527189
rect 176314 527040 176331 527074
rect 176365 527040 176382 527074
rect 176314 527023 176382 527040
rect 176678 527110 176748 527125
rect 176678 527076 176695 527110
rect 176729 527076 176748 527110
rect 176678 526875 176748 527076
rect 177418 527074 177486 527189
rect 177418 527040 177435 527074
rect 177469 527040 177486 527074
rect 177418 527023 177486 527040
rect 177782 527110 177852 527125
rect 177782 527076 177799 527110
rect 177833 527076 177852 527110
rect 177782 526875 177852 527076
rect 178522 527074 178590 527189
rect 179309 527144 179827 527203
rect 179953 527204 180011 527298
rect 179953 527170 179965 527204
rect 179999 527170 180011 527204
rect 180045 527237 181114 527298
rect 180045 527203 180063 527237
rect 180097 527203 181063 527237
rect 181097 527203 181114 527237
rect 180045 527189 181114 527203
rect 181149 527237 182218 527298
rect 181149 527203 181167 527237
rect 181201 527203 182167 527237
rect 182201 527203 182218 527237
rect 181149 527189 182218 527203
rect 182253 527237 183322 527298
rect 182253 527203 182271 527237
rect 182305 527203 183271 527237
rect 183305 527203 183322 527237
rect 182253 527189 183322 527203
rect 183357 527237 184426 527298
rect 183357 527203 183375 527237
rect 183409 527203 184375 527237
rect 184409 527203 184426 527237
rect 183357 527189 184426 527203
rect 184461 527237 184979 527298
rect 184461 527203 184479 527237
rect 184513 527203 184927 527237
rect 184961 527203 184979 527237
rect 179953 527153 180011 527170
rect 178522 527040 178539 527074
rect 178573 527040 178590 527074
rect 178522 527023 178590 527040
rect 178886 527110 178956 527125
rect 178886 527076 178903 527110
rect 178937 527076 178956 527110
rect 178886 526875 178956 527076
rect 179309 527074 179551 527144
rect 179309 527040 179387 527074
rect 179421 527040 179497 527074
rect 179531 527040 179551 527074
rect 179585 527076 179605 527110
rect 179639 527076 179715 527110
rect 179749 527076 179827 527110
rect 179585 527006 179827 527076
rect 180362 527074 180430 527189
rect 180362 527040 180379 527074
rect 180413 527040 180430 527074
rect 180362 527023 180430 527040
rect 180726 527110 180796 527125
rect 180726 527076 180743 527110
rect 180777 527076 180796 527110
rect 179309 526966 179827 527006
rect 179309 526932 179327 526966
rect 179361 526932 179775 526966
rect 179809 526932 179827 526966
rect 174801 526788 174859 526859
rect 174893 526864 175962 526875
rect 174893 526830 174911 526864
rect 174945 526830 175911 526864
rect 175945 526830 175962 526864
rect 174893 526788 175962 526830
rect 175997 526864 177066 526875
rect 175997 526830 176015 526864
rect 176049 526830 177015 526864
rect 177049 526830 177066 526864
rect 175997 526788 177066 526830
rect 177101 526864 178170 526875
rect 177101 526830 177119 526864
rect 177153 526830 178119 526864
rect 178153 526830 178170 526864
rect 177101 526788 178170 526830
rect 178205 526864 179274 526875
rect 178205 526830 178223 526864
rect 178257 526830 179223 526864
rect 179257 526830 179274 526864
rect 178205 526788 179274 526830
rect 179309 526864 179827 526932
rect 179309 526830 179327 526864
rect 179361 526830 179775 526864
rect 179809 526830 179827 526864
rect 179309 526788 179827 526830
rect 179953 526986 180011 527021
rect 179953 526952 179965 526986
rect 179999 526952 180011 526986
rect 179953 526893 180011 526952
rect 179953 526859 179965 526893
rect 179999 526859 180011 526893
rect 180726 526875 180796 527076
rect 181466 527074 181534 527189
rect 181466 527040 181483 527074
rect 181517 527040 181534 527074
rect 181466 527023 181534 527040
rect 181830 527110 181900 527125
rect 181830 527076 181847 527110
rect 181881 527076 181900 527110
rect 181830 526875 181900 527076
rect 182570 527074 182638 527189
rect 182570 527040 182587 527074
rect 182621 527040 182638 527074
rect 182570 527023 182638 527040
rect 182934 527110 183004 527125
rect 182934 527076 182951 527110
rect 182985 527076 183004 527110
rect 182934 526875 183004 527076
rect 183674 527074 183742 527189
rect 184461 527144 184979 527203
rect 185105 527204 185163 527298
rect 185105 527170 185117 527204
rect 185151 527170 185163 527204
rect 185197 527237 186266 527298
rect 185197 527203 185215 527237
rect 185249 527203 186215 527237
rect 186249 527203 186266 527237
rect 185197 527189 186266 527203
rect 186301 527237 187003 527298
rect 186301 527203 186319 527237
rect 186353 527203 186951 527237
rect 186985 527203 187003 527237
rect 185105 527153 185163 527170
rect 183674 527040 183691 527074
rect 183725 527040 183742 527074
rect 183674 527023 183742 527040
rect 184038 527110 184108 527125
rect 184038 527076 184055 527110
rect 184089 527076 184108 527110
rect 184038 526875 184108 527076
rect 184461 527074 184703 527144
rect 184461 527040 184539 527074
rect 184573 527040 184649 527074
rect 184683 527040 184703 527074
rect 184737 527076 184757 527110
rect 184791 527076 184867 527110
rect 184901 527076 184979 527110
rect 184737 527006 184979 527076
rect 185514 527074 185582 527189
rect 186301 527144 187003 527203
rect 187221 527235 187463 527298
rect 187221 527201 187239 527235
rect 187273 527201 187411 527235
rect 187445 527201 187463 527235
rect 187221 527148 187463 527201
rect 185514 527040 185531 527074
rect 185565 527040 185582 527074
rect 185514 527023 185582 527040
rect 185878 527110 185948 527125
rect 185878 527076 185895 527110
rect 185929 527076 185948 527110
rect 184461 526966 184979 527006
rect 184461 526932 184479 526966
rect 184513 526932 184927 526966
rect 184961 526932 184979 526966
rect 179953 526788 180011 526859
rect 180045 526864 181114 526875
rect 180045 526830 180063 526864
rect 180097 526830 181063 526864
rect 181097 526830 181114 526864
rect 180045 526788 181114 526830
rect 181149 526864 182218 526875
rect 181149 526830 181167 526864
rect 181201 526830 182167 526864
rect 182201 526830 182218 526864
rect 181149 526788 182218 526830
rect 182253 526864 183322 526875
rect 182253 526830 182271 526864
rect 182305 526830 183271 526864
rect 183305 526830 183322 526864
rect 182253 526788 183322 526830
rect 183357 526864 184426 526875
rect 183357 526830 183375 526864
rect 183409 526830 184375 526864
rect 184409 526830 184426 526864
rect 183357 526788 184426 526830
rect 184461 526864 184979 526932
rect 184461 526830 184479 526864
rect 184513 526830 184927 526864
rect 184961 526830 184979 526864
rect 184461 526788 184979 526830
rect 185105 526986 185163 527021
rect 185105 526952 185117 526986
rect 185151 526952 185163 526986
rect 185105 526893 185163 526952
rect 185105 526859 185117 526893
rect 185151 526859 185163 526893
rect 185878 526875 185948 527076
rect 186301 527074 186631 527144
rect 186301 527040 186379 527074
rect 186413 527040 186478 527074
rect 186512 527040 186577 527074
rect 186611 527040 186631 527074
rect 186665 527076 186685 527110
rect 186719 527076 186788 527110
rect 186822 527076 186891 527110
rect 186925 527076 187003 527110
rect 186665 527006 187003 527076
rect 186301 526966 187003 527006
rect 186301 526932 186319 526966
rect 186353 526932 186951 526966
rect 186985 526932 187003 526966
rect 185105 526788 185163 526859
rect 185197 526864 186266 526875
rect 185197 526830 185215 526864
rect 185249 526830 186215 526864
rect 186249 526830 186266 526864
rect 185197 526788 186266 526830
rect 186301 526864 187003 526932
rect 186301 526830 186319 526864
rect 186353 526830 186951 526864
rect 186985 526830 187003 526864
rect 186301 526788 187003 526830
rect 187221 527080 187271 527114
rect 187305 527080 187325 527114
rect 187221 527006 187325 527080
rect 187359 527074 187463 527148
rect 187359 527040 187379 527074
rect 187413 527040 187463 527074
rect 187221 526959 187463 527006
rect 187221 526925 187239 526959
rect 187273 526925 187411 526959
rect 187445 526925 187463 526959
rect 187221 526864 187463 526925
rect 187221 526830 187239 526864
rect 187273 526830 187411 526864
rect 187445 526830 187463 526864
rect 187221 526788 187463 526830
rect 172208 526754 172237 526788
rect 172271 526754 172329 526788
rect 172363 526754 172421 526788
rect 172455 526754 172513 526788
rect 172547 526754 172605 526788
rect 172639 526754 172697 526788
rect 172731 526754 172789 526788
rect 172823 526754 172881 526788
rect 172915 526754 172973 526788
rect 173007 526754 173065 526788
rect 173099 526754 173157 526788
rect 173191 526754 173249 526788
rect 173283 526754 173341 526788
rect 173375 526754 173433 526788
rect 173467 526754 173525 526788
rect 173559 526754 173617 526788
rect 173651 526754 173709 526788
rect 173743 526754 173801 526788
rect 173835 526754 173893 526788
rect 173927 526754 173985 526788
rect 174019 526754 174077 526788
rect 174111 526754 174169 526788
rect 174203 526754 174261 526788
rect 174295 526754 174353 526788
rect 174387 526754 174445 526788
rect 174479 526754 174537 526788
rect 174571 526754 174629 526788
rect 174663 526754 174721 526788
rect 174755 526754 174813 526788
rect 174847 526754 174905 526788
rect 174939 526754 174997 526788
rect 175031 526754 175089 526788
rect 175123 526754 175181 526788
rect 175215 526754 175273 526788
rect 175307 526754 175365 526788
rect 175399 526754 175457 526788
rect 175491 526754 175549 526788
rect 175583 526754 175641 526788
rect 175675 526754 175733 526788
rect 175767 526754 175825 526788
rect 175859 526754 175917 526788
rect 175951 526754 176009 526788
rect 176043 526754 176101 526788
rect 176135 526754 176193 526788
rect 176227 526754 176285 526788
rect 176319 526754 176377 526788
rect 176411 526754 176469 526788
rect 176503 526754 176561 526788
rect 176595 526754 176653 526788
rect 176687 526754 176745 526788
rect 176779 526754 176837 526788
rect 176871 526754 176929 526788
rect 176963 526754 177021 526788
rect 177055 526754 177113 526788
rect 177147 526754 177205 526788
rect 177239 526754 177297 526788
rect 177331 526754 177389 526788
rect 177423 526754 177481 526788
rect 177515 526754 177573 526788
rect 177607 526754 177665 526788
rect 177699 526754 177757 526788
rect 177791 526754 177849 526788
rect 177883 526754 177941 526788
rect 177975 526754 178033 526788
rect 178067 526754 178125 526788
rect 178159 526754 178217 526788
rect 178251 526754 178309 526788
rect 178343 526754 178401 526788
rect 178435 526754 178493 526788
rect 178527 526754 178585 526788
rect 178619 526754 178677 526788
rect 178711 526754 178769 526788
rect 178803 526754 178861 526788
rect 178895 526754 178953 526788
rect 178987 526754 179045 526788
rect 179079 526754 179137 526788
rect 179171 526754 179229 526788
rect 179263 526754 179321 526788
rect 179355 526754 179413 526788
rect 179447 526754 179505 526788
rect 179539 526754 179597 526788
rect 179631 526754 179689 526788
rect 179723 526754 179781 526788
rect 179815 526754 179873 526788
rect 179907 526754 179965 526788
rect 179999 526754 180057 526788
rect 180091 526754 180149 526788
rect 180183 526754 180241 526788
rect 180275 526754 180333 526788
rect 180367 526754 180425 526788
rect 180459 526754 180517 526788
rect 180551 526754 180609 526788
rect 180643 526754 180701 526788
rect 180735 526754 180793 526788
rect 180827 526754 180885 526788
rect 180919 526754 180977 526788
rect 181011 526754 181069 526788
rect 181103 526754 181161 526788
rect 181195 526754 181253 526788
rect 181287 526754 181345 526788
rect 181379 526754 181437 526788
rect 181471 526754 181529 526788
rect 181563 526754 181621 526788
rect 181655 526754 181713 526788
rect 181747 526754 181805 526788
rect 181839 526754 181897 526788
rect 181931 526754 181989 526788
rect 182023 526754 182081 526788
rect 182115 526754 182173 526788
rect 182207 526754 182265 526788
rect 182299 526754 182357 526788
rect 182391 526754 182449 526788
rect 182483 526754 182541 526788
rect 182575 526754 182633 526788
rect 182667 526754 182725 526788
rect 182759 526754 182817 526788
rect 182851 526754 182909 526788
rect 182943 526754 183001 526788
rect 183035 526754 183093 526788
rect 183127 526754 183185 526788
rect 183219 526754 183277 526788
rect 183311 526754 183369 526788
rect 183403 526754 183461 526788
rect 183495 526754 183553 526788
rect 183587 526754 183645 526788
rect 183679 526754 183737 526788
rect 183771 526754 183829 526788
rect 183863 526754 183921 526788
rect 183955 526754 184013 526788
rect 184047 526754 184105 526788
rect 184139 526754 184197 526788
rect 184231 526754 184289 526788
rect 184323 526754 184381 526788
rect 184415 526754 184473 526788
rect 184507 526754 184565 526788
rect 184599 526754 184657 526788
rect 184691 526754 184749 526788
rect 184783 526754 184841 526788
rect 184875 526754 184933 526788
rect 184967 526754 185025 526788
rect 185059 526754 185117 526788
rect 185151 526754 185209 526788
rect 185243 526754 185301 526788
rect 185335 526754 185393 526788
rect 185427 526754 185485 526788
rect 185519 526754 185577 526788
rect 185611 526754 185669 526788
rect 185703 526754 185761 526788
rect 185795 526754 185853 526788
rect 185887 526754 185945 526788
rect 185979 526754 186037 526788
rect 186071 526754 186129 526788
rect 186163 526754 186221 526788
rect 186255 526754 186313 526788
rect 186347 526754 186405 526788
rect 186439 526754 186497 526788
rect 186531 526754 186589 526788
rect 186623 526754 186681 526788
rect 186715 526754 186773 526788
rect 186807 526754 186865 526788
rect 186899 526754 186957 526788
rect 186991 526754 187049 526788
rect 187083 526754 187141 526788
rect 187175 526754 187233 526788
rect 187267 526754 187325 526788
rect 187359 526754 187417 526788
rect 187451 526754 187480 526788
rect 172225 526712 172467 526754
rect 172225 526678 172243 526712
rect 172277 526678 172415 526712
rect 172449 526678 172467 526712
rect 172225 526617 172467 526678
rect 172501 526712 173570 526754
rect 172501 526678 172519 526712
rect 172553 526678 173519 526712
rect 173553 526678 173570 526712
rect 172501 526667 173570 526678
rect 173605 526712 174674 526754
rect 173605 526678 173623 526712
rect 173657 526678 174623 526712
rect 174657 526678 174674 526712
rect 173605 526667 174674 526678
rect 174709 526712 175778 526754
rect 174709 526678 174727 526712
rect 174761 526678 175727 526712
rect 175761 526678 175778 526712
rect 174709 526667 175778 526678
rect 175813 526712 176882 526754
rect 175813 526678 175831 526712
rect 175865 526678 176831 526712
rect 176865 526678 176882 526712
rect 175813 526667 176882 526678
rect 176917 526712 177251 526754
rect 176917 526678 176935 526712
rect 176969 526678 177199 526712
rect 177233 526678 177251 526712
rect 172225 526583 172243 526617
rect 172277 526583 172415 526617
rect 172449 526583 172467 526617
rect 172225 526536 172467 526583
rect 172225 526468 172275 526502
rect 172309 526468 172329 526502
rect 172225 526394 172329 526468
rect 172363 526462 172467 526536
rect 172363 526428 172383 526462
rect 172417 526428 172467 526462
rect 172818 526502 172886 526519
rect 172818 526468 172835 526502
rect 172869 526468 172886 526502
rect 172225 526341 172467 526394
rect 172818 526353 172886 526468
rect 173182 526466 173252 526667
rect 173182 526432 173199 526466
rect 173233 526432 173252 526466
rect 173182 526417 173252 526432
rect 173922 526502 173990 526519
rect 173922 526468 173939 526502
rect 173973 526468 173990 526502
rect 173922 526353 173990 526468
rect 174286 526466 174356 526667
rect 174286 526432 174303 526466
rect 174337 526432 174356 526466
rect 174286 526417 174356 526432
rect 175026 526502 175094 526519
rect 175026 526468 175043 526502
rect 175077 526468 175094 526502
rect 175026 526353 175094 526468
rect 175390 526466 175460 526667
rect 175390 526432 175407 526466
rect 175441 526432 175460 526466
rect 175390 526417 175460 526432
rect 176130 526502 176198 526519
rect 176130 526468 176147 526502
rect 176181 526468 176198 526502
rect 176130 526353 176198 526468
rect 176494 526466 176564 526667
rect 176917 526610 177251 526678
rect 176917 526576 176935 526610
rect 176969 526576 177199 526610
rect 177233 526576 177251 526610
rect 176917 526536 177251 526576
rect 176494 526432 176511 526466
rect 176545 526432 176564 526466
rect 176494 526417 176564 526432
rect 176917 526468 176937 526502
rect 176971 526468 177067 526502
rect 176917 526398 177067 526468
rect 177101 526466 177251 526536
rect 177377 526683 177435 526754
rect 177377 526649 177389 526683
rect 177423 526649 177435 526683
rect 177469 526712 178538 526754
rect 177469 526678 177487 526712
rect 177521 526678 178487 526712
rect 178521 526678 178538 526712
rect 177469 526667 178538 526678
rect 178573 526712 179642 526754
rect 178573 526678 178591 526712
rect 178625 526678 179591 526712
rect 179625 526678 179642 526712
rect 178573 526667 179642 526678
rect 179677 526712 180746 526754
rect 179677 526678 179695 526712
rect 179729 526678 180695 526712
rect 180729 526678 180746 526712
rect 179677 526667 180746 526678
rect 180781 526712 181850 526754
rect 180781 526678 180799 526712
rect 180833 526678 181799 526712
rect 181833 526678 181850 526712
rect 180781 526667 181850 526678
rect 181885 526712 182403 526754
rect 181885 526678 181903 526712
rect 181937 526678 182351 526712
rect 182385 526678 182403 526712
rect 177377 526590 177435 526649
rect 177377 526556 177389 526590
rect 177423 526556 177435 526590
rect 177377 526521 177435 526556
rect 177101 526432 177197 526466
rect 177231 526432 177251 526466
rect 177786 526502 177854 526519
rect 177786 526468 177803 526502
rect 177837 526468 177854 526502
rect 172225 526307 172243 526341
rect 172277 526307 172415 526341
rect 172449 526307 172467 526341
rect 172225 526244 172467 526307
rect 172501 526339 173570 526353
rect 172501 526305 172519 526339
rect 172553 526305 173519 526339
rect 173553 526305 173570 526339
rect 172501 526244 173570 526305
rect 173605 526339 174674 526353
rect 173605 526305 173623 526339
rect 173657 526305 174623 526339
rect 174657 526305 174674 526339
rect 173605 526244 174674 526305
rect 174709 526339 175778 526353
rect 174709 526305 174727 526339
rect 174761 526305 175727 526339
rect 175761 526305 175778 526339
rect 174709 526244 175778 526305
rect 175813 526339 176882 526353
rect 175813 526305 175831 526339
rect 175865 526305 176831 526339
rect 176865 526305 176882 526339
rect 175813 526244 176882 526305
rect 176917 526346 177251 526398
rect 176917 526312 176935 526346
rect 176969 526312 177199 526346
rect 177233 526312 177251 526346
rect 176917 526244 177251 526312
rect 177377 526372 177435 526389
rect 177377 526338 177389 526372
rect 177423 526338 177435 526372
rect 177786 526353 177854 526468
rect 178150 526466 178220 526667
rect 178150 526432 178167 526466
rect 178201 526432 178220 526466
rect 178150 526417 178220 526432
rect 178890 526502 178958 526519
rect 178890 526468 178907 526502
rect 178941 526468 178958 526502
rect 178890 526353 178958 526468
rect 179254 526466 179324 526667
rect 179254 526432 179271 526466
rect 179305 526432 179324 526466
rect 179254 526417 179324 526432
rect 179994 526502 180062 526519
rect 179994 526468 180011 526502
rect 180045 526468 180062 526502
rect 179994 526353 180062 526468
rect 180358 526466 180428 526667
rect 180358 526432 180375 526466
rect 180409 526432 180428 526466
rect 180358 526417 180428 526432
rect 181098 526502 181166 526519
rect 181098 526468 181115 526502
rect 181149 526468 181166 526502
rect 181098 526353 181166 526468
rect 181462 526466 181532 526667
rect 181885 526610 182403 526678
rect 181885 526576 181903 526610
rect 181937 526576 182351 526610
rect 182385 526576 182403 526610
rect 181885 526536 182403 526576
rect 181462 526432 181479 526466
rect 181513 526432 181532 526466
rect 181462 526417 181532 526432
rect 181885 526468 181963 526502
rect 181997 526468 182073 526502
rect 182107 526468 182127 526502
rect 181885 526398 182127 526468
rect 182161 526466 182403 526536
rect 182529 526683 182587 526754
rect 182529 526649 182541 526683
rect 182575 526649 182587 526683
rect 182621 526712 183690 526754
rect 182621 526678 182639 526712
rect 182673 526678 183639 526712
rect 183673 526678 183690 526712
rect 182621 526667 183690 526678
rect 183725 526712 184794 526754
rect 183725 526678 183743 526712
rect 183777 526678 184743 526712
rect 184777 526678 184794 526712
rect 183725 526667 184794 526678
rect 184829 526712 185898 526754
rect 184829 526678 184847 526712
rect 184881 526678 185847 526712
rect 185881 526678 185898 526712
rect 184829 526667 185898 526678
rect 185933 526712 187002 526754
rect 185933 526678 185951 526712
rect 185985 526678 186951 526712
rect 186985 526678 187002 526712
rect 185933 526667 187002 526678
rect 187221 526712 187463 526754
rect 187221 526678 187239 526712
rect 187273 526678 187411 526712
rect 187445 526678 187463 526712
rect 182529 526590 182587 526649
rect 182529 526556 182541 526590
rect 182575 526556 182587 526590
rect 182529 526521 182587 526556
rect 182161 526432 182181 526466
rect 182215 526432 182291 526466
rect 182325 526432 182403 526466
rect 182938 526502 183006 526519
rect 182938 526468 182955 526502
rect 182989 526468 183006 526502
rect 177377 526244 177435 526338
rect 177469 526339 178538 526353
rect 177469 526305 177487 526339
rect 177521 526305 178487 526339
rect 178521 526305 178538 526339
rect 177469 526244 178538 526305
rect 178573 526339 179642 526353
rect 178573 526305 178591 526339
rect 178625 526305 179591 526339
rect 179625 526305 179642 526339
rect 178573 526244 179642 526305
rect 179677 526339 180746 526353
rect 179677 526305 179695 526339
rect 179729 526305 180695 526339
rect 180729 526305 180746 526339
rect 179677 526244 180746 526305
rect 180781 526339 181850 526353
rect 180781 526305 180799 526339
rect 180833 526305 181799 526339
rect 181833 526305 181850 526339
rect 180781 526244 181850 526305
rect 181885 526339 182403 526398
rect 181885 526305 181903 526339
rect 181937 526305 182351 526339
rect 182385 526305 182403 526339
rect 181885 526244 182403 526305
rect 182529 526372 182587 526389
rect 182529 526338 182541 526372
rect 182575 526338 182587 526372
rect 182938 526353 183006 526468
rect 183302 526466 183372 526667
rect 183302 526432 183319 526466
rect 183353 526432 183372 526466
rect 183302 526417 183372 526432
rect 184042 526502 184110 526519
rect 184042 526468 184059 526502
rect 184093 526468 184110 526502
rect 184042 526353 184110 526468
rect 184406 526466 184476 526667
rect 184406 526432 184423 526466
rect 184457 526432 184476 526466
rect 184406 526417 184476 526432
rect 185146 526502 185214 526519
rect 185146 526468 185163 526502
rect 185197 526468 185214 526502
rect 185146 526353 185214 526468
rect 185510 526466 185580 526667
rect 185510 526432 185527 526466
rect 185561 526432 185580 526466
rect 185510 526417 185580 526432
rect 186250 526502 186318 526519
rect 186250 526468 186267 526502
rect 186301 526468 186318 526502
rect 186250 526353 186318 526468
rect 186614 526466 186684 526667
rect 186614 526432 186631 526466
rect 186665 526432 186684 526466
rect 186614 526417 186684 526432
rect 187221 526617 187463 526678
rect 187221 526583 187239 526617
rect 187273 526583 187411 526617
rect 187445 526583 187463 526617
rect 187221 526536 187463 526583
rect 187221 526462 187325 526536
rect 187221 526428 187271 526462
rect 187305 526428 187325 526462
rect 187359 526468 187379 526502
rect 187413 526468 187463 526502
rect 187359 526394 187463 526468
rect 182529 526244 182587 526338
rect 182621 526339 183690 526353
rect 182621 526305 182639 526339
rect 182673 526305 183639 526339
rect 183673 526305 183690 526339
rect 182621 526244 183690 526305
rect 183725 526339 184794 526353
rect 183725 526305 183743 526339
rect 183777 526305 184743 526339
rect 184777 526305 184794 526339
rect 183725 526244 184794 526305
rect 184829 526339 185898 526353
rect 184829 526305 184847 526339
rect 184881 526305 185847 526339
rect 185881 526305 185898 526339
rect 184829 526244 185898 526305
rect 185933 526339 187002 526353
rect 185933 526305 185951 526339
rect 185985 526305 186951 526339
rect 186985 526305 187002 526339
rect 185933 526244 187002 526305
rect 187221 526341 187463 526394
rect 187221 526307 187239 526341
rect 187273 526307 187411 526341
rect 187445 526307 187463 526341
rect 187221 526244 187463 526307
rect 172208 526210 172237 526244
rect 172271 526210 172329 526244
rect 172363 526210 172421 526244
rect 172455 526210 172513 526244
rect 172547 526210 172605 526244
rect 172639 526210 172697 526244
rect 172731 526210 172789 526244
rect 172823 526210 172881 526244
rect 172915 526210 172973 526244
rect 173007 526210 173065 526244
rect 173099 526210 173157 526244
rect 173191 526210 173249 526244
rect 173283 526210 173341 526244
rect 173375 526210 173433 526244
rect 173467 526210 173525 526244
rect 173559 526210 173617 526244
rect 173651 526210 173709 526244
rect 173743 526210 173801 526244
rect 173835 526210 173893 526244
rect 173927 526210 173985 526244
rect 174019 526210 174077 526244
rect 174111 526210 174169 526244
rect 174203 526210 174261 526244
rect 174295 526210 174353 526244
rect 174387 526210 174445 526244
rect 174479 526210 174537 526244
rect 174571 526210 174629 526244
rect 174663 526210 174721 526244
rect 174755 526210 174813 526244
rect 174847 526210 174905 526244
rect 174939 526210 174997 526244
rect 175031 526210 175089 526244
rect 175123 526210 175181 526244
rect 175215 526210 175273 526244
rect 175307 526210 175365 526244
rect 175399 526210 175457 526244
rect 175491 526210 175549 526244
rect 175583 526210 175641 526244
rect 175675 526210 175733 526244
rect 175767 526210 175825 526244
rect 175859 526210 175917 526244
rect 175951 526210 176009 526244
rect 176043 526210 176101 526244
rect 176135 526210 176193 526244
rect 176227 526210 176285 526244
rect 176319 526210 176377 526244
rect 176411 526210 176469 526244
rect 176503 526210 176561 526244
rect 176595 526210 176653 526244
rect 176687 526210 176745 526244
rect 176779 526210 176837 526244
rect 176871 526210 176929 526244
rect 176963 526210 177021 526244
rect 177055 526210 177113 526244
rect 177147 526210 177205 526244
rect 177239 526210 177297 526244
rect 177331 526210 177389 526244
rect 177423 526210 177481 526244
rect 177515 526210 177573 526244
rect 177607 526210 177665 526244
rect 177699 526210 177757 526244
rect 177791 526210 177849 526244
rect 177883 526210 177941 526244
rect 177975 526210 178033 526244
rect 178067 526210 178125 526244
rect 178159 526210 178217 526244
rect 178251 526210 178309 526244
rect 178343 526210 178401 526244
rect 178435 526210 178493 526244
rect 178527 526210 178585 526244
rect 178619 526210 178677 526244
rect 178711 526210 178769 526244
rect 178803 526210 178861 526244
rect 178895 526210 178953 526244
rect 178987 526210 179045 526244
rect 179079 526210 179137 526244
rect 179171 526210 179229 526244
rect 179263 526210 179321 526244
rect 179355 526210 179413 526244
rect 179447 526210 179505 526244
rect 179539 526210 179597 526244
rect 179631 526210 179689 526244
rect 179723 526210 179781 526244
rect 179815 526210 179873 526244
rect 179907 526210 179965 526244
rect 179999 526210 180057 526244
rect 180091 526210 180149 526244
rect 180183 526210 180241 526244
rect 180275 526210 180333 526244
rect 180367 526210 180425 526244
rect 180459 526210 180517 526244
rect 180551 526210 180609 526244
rect 180643 526210 180701 526244
rect 180735 526210 180793 526244
rect 180827 526210 180885 526244
rect 180919 526210 180977 526244
rect 181011 526210 181069 526244
rect 181103 526210 181161 526244
rect 181195 526210 181253 526244
rect 181287 526210 181345 526244
rect 181379 526210 181437 526244
rect 181471 526210 181529 526244
rect 181563 526210 181621 526244
rect 181655 526210 181713 526244
rect 181747 526210 181805 526244
rect 181839 526210 181897 526244
rect 181931 526210 181989 526244
rect 182023 526210 182081 526244
rect 182115 526210 182173 526244
rect 182207 526210 182265 526244
rect 182299 526210 182357 526244
rect 182391 526210 182449 526244
rect 182483 526210 182541 526244
rect 182575 526210 182633 526244
rect 182667 526210 182725 526244
rect 182759 526210 182817 526244
rect 182851 526210 182909 526244
rect 182943 526210 183001 526244
rect 183035 526210 183093 526244
rect 183127 526210 183185 526244
rect 183219 526210 183277 526244
rect 183311 526210 183369 526244
rect 183403 526210 183461 526244
rect 183495 526210 183553 526244
rect 183587 526210 183645 526244
rect 183679 526210 183737 526244
rect 183771 526210 183829 526244
rect 183863 526210 183921 526244
rect 183955 526210 184013 526244
rect 184047 526210 184105 526244
rect 184139 526210 184197 526244
rect 184231 526210 184289 526244
rect 184323 526210 184381 526244
rect 184415 526210 184473 526244
rect 184507 526210 184565 526244
rect 184599 526210 184657 526244
rect 184691 526210 184749 526244
rect 184783 526210 184841 526244
rect 184875 526210 184933 526244
rect 184967 526210 185025 526244
rect 185059 526210 185117 526244
rect 185151 526210 185209 526244
rect 185243 526210 185301 526244
rect 185335 526210 185393 526244
rect 185427 526210 185485 526244
rect 185519 526210 185577 526244
rect 185611 526210 185669 526244
rect 185703 526210 185761 526244
rect 185795 526210 185853 526244
rect 185887 526210 185945 526244
rect 185979 526210 186037 526244
rect 186071 526210 186129 526244
rect 186163 526210 186221 526244
rect 186255 526210 186313 526244
rect 186347 526210 186405 526244
rect 186439 526210 186497 526244
rect 186531 526210 186589 526244
rect 186623 526210 186681 526244
rect 186715 526210 186773 526244
rect 186807 526210 186865 526244
rect 186899 526210 186957 526244
rect 186991 526210 187049 526244
rect 187083 526210 187141 526244
rect 187175 526210 187233 526244
rect 187267 526210 187325 526244
rect 187359 526210 187417 526244
rect 187451 526210 187480 526244
rect 172225 526147 172467 526210
rect 172225 526113 172243 526147
rect 172277 526113 172415 526147
rect 172449 526113 172467 526147
rect 172225 526060 172467 526113
rect 172501 526149 173570 526210
rect 172501 526115 172519 526149
rect 172553 526115 173519 526149
rect 173553 526115 173570 526149
rect 172501 526101 173570 526115
rect 173605 526149 174674 526210
rect 173605 526115 173623 526149
rect 173657 526115 174623 526149
rect 174657 526115 174674 526149
rect 173605 526101 174674 526115
rect 174801 526116 174859 526210
rect 172225 525986 172329 526060
rect 172225 525952 172275 525986
rect 172309 525952 172329 525986
rect 172363 525992 172383 526026
rect 172417 525992 172467 526026
rect 172363 525918 172467 525992
rect 172818 525986 172886 526101
rect 172818 525952 172835 525986
rect 172869 525952 172886 525986
rect 172818 525935 172886 525952
rect 173182 526022 173252 526037
rect 173182 525988 173199 526022
rect 173233 525988 173252 526022
rect 172225 525871 172467 525918
rect 172225 525837 172243 525871
rect 172277 525837 172415 525871
rect 172449 525837 172467 525871
rect 172225 525776 172467 525837
rect 173182 525787 173252 525988
rect 173922 525986 173990 526101
rect 174801 526082 174813 526116
rect 174847 526082 174859 526116
rect 174893 526149 175962 526210
rect 174893 526115 174911 526149
rect 174945 526115 175911 526149
rect 175945 526115 175962 526149
rect 174893 526101 175962 526115
rect 175997 526149 177066 526210
rect 175997 526115 176015 526149
rect 176049 526115 177015 526149
rect 177049 526115 177066 526149
rect 175997 526101 177066 526115
rect 177101 526149 178170 526210
rect 177101 526115 177119 526149
rect 177153 526115 178119 526149
rect 178153 526115 178170 526149
rect 177101 526101 178170 526115
rect 178205 526149 179274 526210
rect 178205 526115 178223 526149
rect 178257 526115 179223 526149
rect 179257 526115 179274 526149
rect 178205 526101 179274 526115
rect 179309 526149 179827 526210
rect 179309 526115 179327 526149
rect 179361 526115 179775 526149
rect 179809 526115 179827 526149
rect 174801 526065 174859 526082
rect 173922 525952 173939 525986
rect 173973 525952 173990 525986
rect 173922 525935 173990 525952
rect 174286 526022 174356 526037
rect 174286 525988 174303 526022
rect 174337 525988 174356 526022
rect 174286 525787 174356 525988
rect 175210 525986 175278 526101
rect 175210 525952 175227 525986
rect 175261 525952 175278 525986
rect 175210 525935 175278 525952
rect 175574 526022 175644 526037
rect 175574 525988 175591 526022
rect 175625 525988 175644 526022
rect 174801 525898 174859 525933
rect 174801 525864 174813 525898
rect 174847 525864 174859 525898
rect 174801 525805 174859 525864
rect 172225 525742 172243 525776
rect 172277 525742 172415 525776
rect 172449 525742 172467 525776
rect 172225 525700 172467 525742
rect 172501 525776 173570 525787
rect 172501 525742 172519 525776
rect 172553 525742 173519 525776
rect 173553 525742 173570 525776
rect 172501 525700 173570 525742
rect 173605 525776 174674 525787
rect 173605 525742 173623 525776
rect 173657 525742 174623 525776
rect 174657 525742 174674 525776
rect 173605 525700 174674 525742
rect 174801 525771 174813 525805
rect 174847 525771 174859 525805
rect 175574 525787 175644 525988
rect 176314 525986 176382 526101
rect 176314 525952 176331 525986
rect 176365 525952 176382 525986
rect 176314 525935 176382 525952
rect 176678 526022 176748 526037
rect 176678 525988 176695 526022
rect 176729 525988 176748 526022
rect 176678 525787 176748 525988
rect 177418 525986 177486 526101
rect 177418 525952 177435 525986
rect 177469 525952 177486 525986
rect 177418 525935 177486 525952
rect 177782 526022 177852 526037
rect 177782 525988 177799 526022
rect 177833 525988 177852 526022
rect 177782 525787 177852 525988
rect 178522 525986 178590 526101
rect 179309 526056 179827 526115
rect 179953 526116 180011 526210
rect 179953 526082 179965 526116
rect 179999 526082 180011 526116
rect 180045 526149 181114 526210
rect 180045 526115 180063 526149
rect 180097 526115 181063 526149
rect 181097 526115 181114 526149
rect 180045 526101 181114 526115
rect 181149 526149 182218 526210
rect 181149 526115 181167 526149
rect 181201 526115 182167 526149
rect 182201 526115 182218 526149
rect 181149 526101 182218 526115
rect 182253 526149 183322 526210
rect 182253 526115 182271 526149
rect 182305 526115 183271 526149
rect 183305 526115 183322 526149
rect 182253 526101 183322 526115
rect 183357 526149 184426 526210
rect 183357 526115 183375 526149
rect 183409 526115 184375 526149
rect 184409 526115 184426 526149
rect 183357 526101 184426 526115
rect 184461 526149 184979 526210
rect 184461 526115 184479 526149
rect 184513 526115 184927 526149
rect 184961 526115 184979 526149
rect 179953 526065 180011 526082
rect 178522 525952 178539 525986
rect 178573 525952 178590 525986
rect 178522 525935 178590 525952
rect 178886 526022 178956 526037
rect 178886 525988 178903 526022
rect 178937 525988 178956 526022
rect 178886 525787 178956 525988
rect 179309 525986 179551 526056
rect 179309 525952 179387 525986
rect 179421 525952 179497 525986
rect 179531 525952 179551 525986
rect 179585 525988 179605 526022
rect 179639 525988 179715 526022
rect 179749 525988 179827 526022
rect 179585 525918 179827 525988
rect 180362 525986 180430 526101
rect 180362 525952 180379 525986
rect 180413 525952 180430 525986
rect 180362 525935 180430 525952
rect 180726 526022 180796 526037
rect 180726 525988 180743 526022
rect 180777 525988 180796 526022
rect 179309 525878 179827 525918
rect 179309 525844 179327 525878
rect 179361 525844 179775 525878
rect 179809 525844 179827 525878
rect 174801 525700 174859 525771
rect 174893 525776 175962 525787
rect 174893 525742 174911 525776
rect 174945 525742 175911 525776
rect 175945 525742 175962 525776
rect 174893 525700 175962 525742
rect 175997 525776 177066 525787
rect 175997 525742 176015 525776
rect 176049 525742 177015 525776
rect 177049 525742 177066 525776
rect 175997 525700 177066 525742
rect 177101 525776 178170 525787
rect 177101 525742 177119 525776
rect 177153 525742 178119 525776
rect 178153 525742 178170 525776
rect 177101 525700 178170 525742
rect 178205 525776 179274 525787
rect 178205 525742 178223 525776
rect 178257 525742 179223 525776
rect 179257 525742 179274 525776
rect 178205 525700 179274 525742
rect 179309 525776 179827 525844
rect 179309 525742 179327 525776
rect 179361 525742 179775 525776
rect 179809 525742 179827 525776
rect 179309 525700 179827 525742
rect 179953 525898 180011 525933
rect 179953 525864 179965 525898
rect 179999 525864 180011 525898
rect 179953 525805 180011 525864
rect 179953 525771 179965 525805
rect 179999 525771 180011 525805
rect 180726 525787 180796 525988
rect 181466 525986 181534 526101
rect 181466 525952 181483 525986
rect 181517 525952 181534 525986
rect 181466 525935 181534 525952
rect 181830 526022 181900 526037
rect 181830 525988 181847 526022
rect 181881 525988 181900 526022
rect 181830 525787 181900 525988
rect 182570 525986 182638 526101
rect 182570 525952 182587 525986
rect 182621 525952 182638 525986
rect 182570 525935 182638 525952
rect 182934 526022 183004 526037
rect 182934 525988 182951 526022
rect 182985 525988 183004 526022
rect 182934 525787 183004 525988
rect 183674 525986 183742 526101
rect 184461 526056 184979 526115
rect 185105 526116 185163 526210
rect 185105 526082 185117 526116
rect 185151 526082 185163 526116
rect 185197 526149 186266 526210
rect 185197 526115 185215 526149
rect 185249 526115 186215 526149
rect 186249 526115 186266 526149
rect 185197 526101 186266 526115
rect 186301 526149 187003 526210
rect 186301 526115 186319 526149
rect 186353 526115 186951 526149
rect 186985 526115 187003 526149
rect 185105 526065 185163 526082
rect 183674 525952 183691 525986
rect 183725 525952 183742 525986
rect 183674 525935 183742 525952
rect 184038 526022 184108 526037
rect 184038 525988 184055 526022
rect 184089 525988 184108 526022
rect 184038 525787 184108 525988
rect 184461 525986 184703 526056
rect 184461 525952 184539 525986
rect 184573 525952 184649 525986
rect 184683 525952 184703 525986
rect 184737 525988 184757 526022
rect 184791 525988 184867 526022
rect 184901 525988 184979 526022
rect 184737 525918 184979 525988
rect 185514 525986 185582 526101
rect 186301 526056 187003 526115
rect 187221 526147 187463 526210
rect 187221 526113 187239 526147
rect 187273 526113 187411 526147
rect 187445 526113 187463 526147
rect 187221 526060 187463 526113
rect 185514 525952 185531 525986
rect 185565 525952 185582 525986
rect 185514 525935 185582 525952
rect 185878 526022 185948 526037
rect 185878 525988 185895 526022
rect 185929 525988 185948 526022
rect 184461 525878 184979 525918
rect 184461 525844 184479 525878
rect 184513 525844 184927 525878
rect 184961 525844 184979 525878
rect 179953 525700 180011 525771
rect 180045 525776 181114 525787
rect 180045 525742 180063 525776
rect 180097 525742 181063 525776
rect 181097 525742 181114 525776
rect 180045 525700 181114 525742
rect 181149 525776 182218 525787
rect 181149 525742 181167 525776
rect 181201 525742 182167 525776
rect 182201 525742 182218 525776
rect 181149 525700 182218 525742
rect 182253 525776 183322 525787
rect 182253 525742 182271 525776
rect 182305 525742 183271 525776
rect 183305 525742 183322 525776
rect 182253 525700 183322 525742
rect 183357 525776 184426 525787
rect 183357 525742 183375 525776
rect 183409 525742 184375 525776
rect 184409 525742 184426 525776
rect 183357 525700 184426 525742
rect 184461 525776 184979 525844
rect 184461 525742 184479 525776
rect 184513 525742 184927 525776
rect 184961 525742 184979 525776
rect 184461 525700 184979 525742
rect 185105 525898 185163 525933
rect 185105 525864 185117 525898
rect 185151 525864 185163 525898
rect 185105 525805 185163 525864
rect 185105 525771 185117 525805
rect 185151 525771 185163 525805
rect 185878 525787 185948 525988
rect 186301 525986 186631 526056
rect 186301 525952 186379 525986
rect 186413 525952 186478 525986
rect 186512 525952 186577 525986
rect 186611 525952 186631 525986
rect 186665 525988 186685 526022
rect 186719 525988 186788 526022
rect 186822 525988 186891 526022
rect 186925 525988 187003 526022
rect 186665 525918 187003 525988
rect 186301 525878 187003 525918
rect 186301 525844 186319 525878
rect 186353 525844 186951 525878
rect 186985 525844 187003 525878
rect 185105 525700 185163 525771
rect 185197 525776 186266 525787
rect 185197 525742 185215 525776
rect 185249 525742 186215 525776
rect 186249 525742 186266 525776
rect 185197 525700 186266 525742
rect 186301 525776 187003 525844
rect 186301 525742 186319 525776
rect 186353 525742 186951 525776
rect 186985 525742 187003 525776
rect 186301 525700 187003 525742
rect 187221 525992 187271 526026
rect 187305 525992 187325 526026
rect 187221 525918 187325 525992
rect 187359 525986 187463 526060
rect 187359 525952 187379 525986
rect 187413 525952 187463 525986
rect 187221 525871 187463 525918
rect 187221 525837 187239 525871
rect 187273 525837 187411 525871
rect 187445 525837 187463 525871
rect 187221 525776 187463 525837
rect 187221 525742 187239 525776
rect 187273 525742 187411 525776
rect 187445 525742 187463 525776
rect 187221 525700 187463 525742
rect 172208 525666 172237 525700
rect 172271 525666 172329 525700
rect 172363 525666 172421 525700
rect 172455 525666 172513 525700
rect 172547 525666 172605 525700
rect 172639 525666 172697 525700
rect 172731 525666 172789 525700
rect 172823 525666 172881 525700
rect 172915 525666 172973 525700
rect 173007 525666 173065 525700
rect 173099 525666 173157 525700
rect 173191 525666 173249 525700
rect 173283 525666 173341 525700
rect 173375 525666 173433 525700
rect 173467 525666 173525 525700
rect 173559 525666 173617 525700
rect 173651 525666 173709 525700
rect 173743 525666 173801 525700
rect 173835 525666 173893 525700
rect 173927 525666 173985 525700
rect 174019 525666 174077 525700
rect 174111 525666 174169 525700
rect 174203 525666 174261 525700
rect 174295 525666 174353 525700
rect 174387 525666 174445 525700
rect 174479 525666 174537 525700
rect 174571 525666 174629 525700
rect 174663 525666 174721 525700
rect 174755 525666 174813 525700
rect 174847 525666 174905 525700
rect 174939 525666 174997 525700
rect 175031 525666 175089 525700
rect 175123 525666 175181 525700
rect 175215 525666 175273 525700
rect 175307 525666 175365 525700
rect 175399 525666 175457 525700
rect 175491 525666 175549 525700
rect 175583 525666 175641 525700
rect 175675 525666 175733 525700
rect 175767 525666 175825 525700
rect 175859 525666 175917 525700
rect 175951 525666 176009 525700
rect 176043 525666 176101 525700
rect 176135 525666 176193 525700
rect 176227 525666 176285 525700
rect 176319 525666 176377 525700
rect 176411 525666 176469 525700
rect 176503 525666 176561 525700
rect 176595 525666 176653 525700
rect 176687 525666 176745 525700
rect 176779 525666 176837 525700
rect 176871 525666 176929 525700
rect 176963 525666 177021 525700
rect 177055 525666 177113 525700
rect 177147 525666 177205 525700
rect 177239 525666 177297 525700
rect 177331 525666 177389 525700
rect 177423 525666 177481 525700
rect 177515 525666 177573 525700
rect 177607 525666 177665 525700
rect 177699 525666 177757 525700
rect 177791 525666 177849 525700
rect 177883 525666 177941 525700
rect 177975 525666 178033 525700
rect 178067 525666 178125 525700
rect 178159 525666 178217 525700
rect 178251 525666 178309 525700
rect 178343 525666 178401 525700
rect 178435 525666 178493 525700
rect 178527 525666 178585 525700
rect 178619 525666 178677 525700
rect 178711 525666 178769 525700
rect 178803 525666 178861 525700
rect 178895 525666 178953 525700
rect 178987 525666 179045 525700
rect 179079 525666 179137 525700
rect 179171 525666 179229 525700
rect 179263 525666 179321 525700
rect 179355 525666 179413 525700
rect 179447 525666 179505 525700
rect 179539 525666 179597 525700
rect 179631 525666 179689 525700
rect 179723 525666 179781 525700
rect 179815 525666 179873 525700
rect 179907 525666 179965 525700
rect 179999 525666 180057 525700
rect 180091 525666 180149 525700
rect 180183 525666 180241 525700
rect 180275 525666 180333 525700
rect 180367 525666 180425 525700
rect 180459 525666 180517 525700
rect 180551 525666 180609 525700
rect 180643 525666 180701 525700
rect 180735 525666 180793 525700
rect 180827 525666 180885 525700
rect 180919 525666 180977 525700
rect 181011 525666 181069 525700
rect 181103 525666 181161 525700
rect 181195 525666 181253 525700
rect 181287 525666 181345 525700
rect 181379 525666 181437 525700
rect 181471 525666 181529 525700
rect 181563 525666 181621 525700
rect 181655 525666 181713 525700
rect 181747 525666 181805 525700
rect 181839 525666 181897 525700
rect 181931 525666 181989 525700
rect 182023 525666 182081 525700
rect 182115 525666 182173 525700
rect 182207 525666 182265 525700
rect 182299 525666 182357 525700
rect 182391 525666 182449 525700
rect 182483 525666 182541 525700
rect 182575 525666 182633 525700
rect 182667 525666 182725 525700
rect 182759 525666 182817 525700
rect 182851 525666 182909 525700
rect 182943 525666 183001 525700
rect 183035 525666 183093 525700
rect 183127 525666 183185 525700
rect 183219 525666 183277 525700
rect 183311 525666 183369 525700
rect 183403 525666 183461 525700
rect 183495 525666 183553 525700
rect 183587 525666 183645 525700
rect 183679 525666 183737 525700
rect 183771 525666 183829 525700
rect 183863 525666 183921 525700
rect 183955 525666 184013 525700
rect 184047 525666 184105 525700
rect 184139 525666 184197 525700
rect 184231 525666 184289 525700
rect 184323 525666 184381 525700
rect 184415 525666 184473 525700
rect 184507 525666 184565 525700
rect 184599 525666 184657 525700
rect 184691 525666 184749 525700
rect 184783 525666 184841 525700
rect 184875 525666 184933 525700
rect 184967 525666 185025 525700
rect 185059 525666 185117 525700
rect 185151 525666 185209 525700
rect 185243 525666 185301 525700
rect 185335 525666 185393 525700
rect 185427 525666 185485 525700
rect 185519 525666 185577 525700
rect 185611 525666 185669 525700
rect 185703 525666 185761 525700
rect 185795 525666 185853 525700
rect 185887 525666 185945 525700
rect 185979 525666 186037 525700
rect 186071 525666 186129 525700
rect 186163 525666 186221 525700
rect 186255 525666 186313 525700
rect 186347 525666 186405 525700
rect 186439 525666 186497 525700
rect 186531 525666 186589 525700
rect 186623 525666 186681 525700
rect 186715 525666 186773 525700
rect 186807 525666 186865 525700
rect 186899 525666 186957 525700
rect 186991 525666 187049 525700
rect 187083 525666 187141 525700
rect 187175 525666 187233 525700
rect 187267 525666 187325 525700
rect 187359 525666 187417 525700
rect 187451 525666 187480 525700
rect 172225 525624 172467 525666
rect 172225 525590 172243 525624
rect 172277 525590 172415 525624
rect 172449 525590 172467 525624
rect 172225 525529 172467 525590
rect 172501 525624 173570 525666
rect 172501 525590 172519 525624
rect 172553 525590 173519 525624
rect 173553 525590 173570 525624
rect 172501 525579 173570 525590
rect 173605 525624 174674 525666
rect 173605 525590 173623 525624
rect 173657 525590 174623 525624
rect 174657 525590 174674 525624
rect 173605 525579 174674 525590
rect 174709 525624 175778 525666
rect 174709 525590 174727 525624
rect 174761 525590 175727 525624
rect 175761 525590 175778 525624
rect 174709 525579 175778 525590
rect 175813 525624 176882 525666
rect 175813 525590 175831 525624
rect 175865 525590 176831 525624
rect 176865 525590 176882 525624
rect 175813 525579 176882 525590
rect 176917 525624 177251 525666
rect 176917 525590 176935 525624
rect 176969 525590 177199 525624
rect 177233 525590 177251 525624
rect 172225 525495 172243 525529
rect 172277 525495 172415 525529
rect 172449 525495 172467 525529
rect 172225 525448 172467 525495
rect 172225 525380 172275 525414
rect 172309 525380 172329 525414
rect 172225 525306 172329 525380
rect 172363 525374 172467 525448
rect 172363 525340 172383 525374
rect 172417 525340 172467 525374
rect 172818 525414 172886 525431
rect 172818 525380 172835 525414
rect 172869 525380 172886 525414
rect 172225 525253 172467 525306
rect 172818 525265 172886 525380
rect 173182 525378 173252 525579
rect 173182 525344 173199 525378
rect 173233 525344 173252 525378
rect 173182 525329 173252 525344
rect 173922 525414 173990 525431
rect 173922 525380 173939 525414
rect 173973 525380 173990 525414
rect 173922 525265 173990 525380
rect 174286 525378 174356 525579
rect 174286 525344 174303 525378
rect 174337 525344 174356 525378
rect 174286 525329 174356 525344
rect 175026 525414 175094 525431
rect 175026 525380 175043 525414
rect 175077 525380 175094 525414
rect 175026 525265 175094 525380
rect 175390 525378 175460 525579
rect 175390 525344 175407 525378
rect 175441 525344 175460 525378
rect 175390 525329 175460 525344
rect 176130 525414 176198 525431
rect 176130 525380 176147 525414
rect 176181 525380 176198 525414
rect 176130 525265 176198 525380
rect 176494 525378 176564 525579
rect 176917 525522 177251 525590
rect 176917 525488 176935 525522
rect 176969 525488 177199 525522
rect 177233 525488 177251 525522
rect 176917 525448 177251 525488
rect 176494 525344 176511 525378
rect 176545 525344 176564 525378
rect 176494 525329 176564 525344
rect 176917 525380 176937 525414
rect 176971 525380 177067 525414
rect 176917 525310 177067 525380
rect 177101 525378 177251 525448
rect 177377 525595 177435 525666
rect 177377 525561 177389 525595
rect 177423 525561 177435 525595
rect 177469 525624 178538 525666
rect 177469 525590 177487 525624
rect 177521 525590 178487 525624
rect 178521 525590 178538 525624
rect 177469 525579 178538 525590
rect 178573 525624 179642 525666
rect 178573 525590 178591 525624
rect 178625 525590 179591 525624
rect 179625 525590 179642 525624
rect 178573 525579 179642 525590
rect 179677 525624 180746 525666
rect 179677 525590 179695 525624
rect 179729 525590 180695 525624
rect 180729 525590 180746 525624
rect 179677 525579 180746 525590
rect 180781 525624 181850 525666
rect 180781 525590 180799 525624
rect 180833 525590 181799 525624
rect 181833 525590 181850 525624
rect 180781 525579 181850 525590
rect 181885 525624 182403 525666
rect 181885 525590 181903 525624
rect 181937 525590 182351 525624
rect 182385 525590 182403 525624
rect 177377 525502 177435 525561
rect 177377 525468 177389 525502
rect 177423 525468 177435 525502
rect 177377 525433 177435 525468
rect 177101 525344 177197 525378
rect 177231 525344 177251 525378
rect 177786 525414 177854 525431
rect 177786 525380 177803 525414
rect 177837 525380 177854 525414
rect 172225 525219 172243 525253
rect 172277 525219 172415 525253
rect 172449 525219 172467 525253
rect 172225 525156 172467 525219
rect 172501 525251 173570 525265
rect 172501 525217 172519 525251
rect 172553 525217 173519 525251
rect 173553 525217 173570 525251
rect 172501 525156 173570 525217
rect 173605 525251 174674 525265
rect 173605 525217 173623 525251
rect 173657 525217 174623 525251
rect 174657 525217 174674 525251
rect 173605 525156 174674 525217
rect 174709 525251 175778 525265
rect 174709 525217 174727 525251
rect 174761 525217 175727 525251
rect 175761 525217 175778 525251
rect 174709 525156 175778 525217
rect 175813 525251 176882 525265
rect 175813 525217 175831 525251
rect 175865 525217 176831 525251
rect 176865 525217 176882 525251
rect 175813 525156 176882 525217
rect 176917 525258 177251 525310
rect 176917 525224 176935 525258
rect 176969 525224 177199 525258
rect 177233 525224 177251 525258
rect 176917 525156 177251 525224
rect 177377 525284 177435 525301
rect 177377 525250 177389 525284
rect 177423 525250 177435 525284
rect 177786 525265 177854 525380
rect 178150 525378 178220 525579
rect 178150 525344 178167 525378
rect 178201 525344 178220 525378
rect 178150 525329 178220 525344
rect 178890 525414 178958 525431
rect 178890 525380 178907 525414
rect 178941 525380 178958 525414
rect 178890 525265 178958 525380
rect 179254 525378 179324 525579
rect 179254 525344 179271 525378
rect 179305 525344 179324 525378
rect 179254 525329 179324 525344
rect 179994 525414 180062 525431
rect 179994 525380 180011 525414
rect 180045 525380 180062 525414
rect 179994 525265 180062 525380
rect 180358 525378 180428 525579
rect 180358 525344 180375 525378
rect 180409 525344 180428 525378
rect 180358 525329 180428 525344
rect 181098 525414 181166 525431
rect 181098 525380 181115 525414
rect 181149 525380 181166 525414
rect 181098 525265 181166 525380
rect 181462 525378 181532 525579
rect 181885 525522 182403 525590
rect 181885 525488 181903 525522
rect 181937 525488 182351 525522
rect 182385 525488 182403 525522
rect 181885 525448 182403 525488
rect 181462 525344 181479 525378
rect 181513 525344 181532 525378
rect 181462 525329 181532 525344
rect 181885 525380 181963 525414
rect 181997 525380 182073 525414
rect 182107 525380 182127 525414
rect 181885 525310 182127 525380
rect 182161 525378 182403 525448
rect 182529 525595 182587 525666
rect 182529 525561 182541 525595
rect 182575 525561 182587 525595
rect 182621 525624 183690 525666
rect 182621 525590 182639 525624
rect 182673 525590 183639 525624
rect 183673 525590 183690 525624
rect 182621 525579 183690 525590
rect 183725 525624 184794 525666
rect 183725 525590 183743 525624
rect 183777 525590 184743 525624
rect 184777 525590 184794 525624
rect 183725 525579 184794 525590
rect 184829 525624 185898 525666
rect 184829 525590 184847 525624
rect 184881 525590 185847 525624
rect 185881 525590 185898 525624
rect 184829 525579 185898 525590
rect 185933 525624 187002 525666
rect 185933 525590 185951 525624
rect 185985 525590 186951 525624
rect 186985 525590 187002 525624
rect 185933 525579 187002 525590
rect 187221 525624 187463 525666
rect 187221 525590 187239 525624
rect 187273 525590 187411 525624
rect 187445 525590 187463 525624
rect 182529 525502 182587 525561
rect 182529 525468 182541 525502
rect 182575 525468 182587 525502
rect 182529 525433 182587 525468
rect 182161 525344 182181 525378
rect 182215 525344 182291 525378
rect 182325 525344 182403 525378
rect 182938 525414 183006 525431
rect 182938 525380 182955 525414
rect 182989 525380 183006 525414
rect 177377 525156 177435 525250
rect 177469 525251 178538 525265
rect 177469 525217 177487 525251
rect 177521 525217 178487 525251
rect 178521 525217 178538 525251
rect 177469 525156 178538 525217
rect 178573 525251 179642 525265
rect 178573 525217 178591 525251
rect 178625 525217 179591 525251
rect 179625 525217 179642 525251
rect 178573 525156 179642 525217
rect 179677 525251 180746 525265
rect 179677 525217 179695 525251
rect 179729 525217 180695 525251
rect 180729 525217 180746 525251
rect 179677 525156 180746 525217
rect 180781 525251 181850 525265
rect 180781 525217 180799 525251
rect 180833 525217 181799 525251
rect 181833 525217 181850 525251
rect 180781 525156 181850 525217
rect 181885 525251 182403 525310
rect 181885 525217 181903 525251
rect 181937 525217 182351 525251
rect 182385 525217 182403 525251
rect 181885 525156 182403 525217
rect 182529 525284 182587 525301
rect 182529 525250 182541 525284
rect 182575 525250 182587 525284
rect 182938 525265 183006 525380
rect 183302 525378 183372 525579
rect 183302 525344 183319 525378
rect 183353 525344 183372 525378
rect 183302 525329 183372 525344
rect 184042 525414 184110 525431
rect 184042 525380 184059 525414
rect 184093 525380 184110 525414
rect 184042 525265 184110 525380
rect 184406 525378 184476 525579
rect 184406 525344 184423 525378
rect 184457 525344 184476 525378
rect 184406 525329 184476 525344
rect 185146 525414 185214 525431
rect 185146 525380 185163 525414
rect 185197 525380 185214 525414
rect 185146 525265 185214 525380
rect 185510 525378 185580 525579
rect 185510 525344 185527 525378
rect 185561 525344 185580 525378
rect 185510 525329 185580 525344
rect 186250 525414 186318 525431
rect 186250 525380 186267 525414
rect 186301 525380 186318 525414
rect 186250 525265 186318 525380
rect 186614 525378 186684 525579
rect 186614 525344 186631 525378
rect 186665 525344 186684 525378
rect 186614 525329 186684 525344
rect 187221 525529 187463 525590
rect 187221 525495 187239 525529
rect 187273 525495 187411 525529
rect 187445 525495 187463 525529
rect 187221 525448 187463 525495
rect 187221 525374 187325 525448
rect 187221 525340 187271 525374
rect 187305 525340 187325 525374
rect 187359 525380 187379 525414
rect 187413 525380 187463 525414
rect 187359 525306 187463 525380
rect 182529 525156 182587 525250
rect 182621 525251 183690 525265
rect 182621 525217 182639 525251
rect 182673 525217 183639 525251
rect 183673 525217 183690 525251
rect 182621 525156 183690 525217
rect 183725 525251 184794 525265
rect 183725 525217 183743 525251
rect 183777 525217 184743 525251
rect 184777 525217 184794 525251
rect 183725 525156 184794 525217
rect 184829 525251 185898 525265
rect 184829 525217 184847 525251
rect 184881 525217 185847 525251
rect 185881 525217 185898 525251
rect 184829 525156 185898 525217
rect 185933 525251 187002 525265
rect 185933 525217 185951 525251
rect 185985 525217 186951 525251
rect 186985 525217 187002 525251
rect 185933 525156 187002 525217
rect 187221 525253 187463 525306
rect 187221 525219 187239 525253
rect 187273 525219 187411 525253
rect 187445 525219 187463 525253
rect 187221 525156 187463 525219
rect 172208 525122 172237 525156
rect 172271 525122 172329 525156
rect 172363 525122 172421 525156
rect 172455 525122 172513 525156
rect 172547 525122 172605 525156
rect 172639 525122 172697 525156
rect 172731 525122 172789 525156
rect 172823 525122 172881 525156
rect 172915 525122 172973 525156
rect 173007 525122 173065 525156
rect 173099 525122 173157 525156
rect 173191 525122 173249 525156
rect 173283 525122 173341 525156
rect 173375 525122 173433 525156
rect 173467 525122 173525 525156
rect 173559 525122 173617 525156
rect 173651 525122 173709 525156
rect 173743 525122 173801 525156
rect 173835 525122 173893 525156
rect 173927 525122 173985 525156
rect 174019 525122 174077 525156
rect 174111 525122 174169 525156
rect 174203 525122 174261 525156
rect 174295 525122 174353 525156
rect 174387 525122 174445 525156
rect 174479 525122 174537 525156
rect 174571 525122 174629 525156
rect 174663 525122 174721 525156
rect 174755 525122 174813 525156
rect 174847 525122 174905 525156
rect 174939 525122 174997 525156
rect 175031 525122 175089 525156
rect 175123 525122 175181 525156
rect 175215 525122 175273 525156
rect 175307 525122 175365 525156
rect 175399 525122 175457 525156
rect 175491 525122 175549 525156
rect 175583 525122 175641 525156
rect 175675 525122 175733 525156
rect 175767 525122 175825 525156
rect 175859 525122 175917 525156
rect 175951 525122 176009 525156
rect 176043 525122 176101 525156
rect 176135 525122 176193 525156
rect 176227 525122 176285 525156
rect 176319 525122 176377 525156
rect 176411 525122 176469 525156
rect 176503 525122 176561 525156
rect 176595 525122 176653 525156
rect 176687 525122 176745 525156
rect 176779 525122 176837 525156
rect 176871 525122 176929 525156
rect 176963 525122 177021 525156
rect 177055 525122 177113 525156
rect 177147 525122 177205 525156
rect 177239 525122 177297 525156
rect 177331 525122 177389 525156
rect 177423 525122 177481 525156
rect 177515 525122 177573 525156
rect 177607 525122 177665 525156
rect 177699 525122 177757 525156
rect 177791 525122 177849 525156
rect 177883 525122 177941 525156
rect 177975 525122 178033 525156
rect 178067 525122 178125 525156
rect 178159 525122 178217 525156
rect 178251 525122 178309 525156
rect 178343 525122 178401 525156
rect 178435 525122 178493 525156
rect 178527 525122 178585 525156
rect 178619 525122 178677 525156
rect 178711 525122 178769 525156
rect 178803 525122 178861 525156
rect 178895 525122 178953 525156
rect 178987 525122 179045 525156
rect 179079 525122 179137 525156
rect 179171 525122 179229 525156
rect 179263 525122 179321 525156
rect 179355 525122 179413 525156
rect 179447 525122 179505 525156
rect 179539 525122 179597 525156
rect 179631 525122 179689 525156
rect 179723 525122 179781 525156
rect 179815 525122 179873 525156
rect 179907 525122 179965 525156
rect 179999 525122 180057 525156
rect 180091 525122 180149 525156
rect 180183 525122 180241 525156
rect 180275 525122 180333 525156
rect 180367 525122 180425 525156
rect 180459 525122 180517 525156
rect 180551 525122 180609 525156
rect 180643 525122 180701 525156
rect 180735 525122 180793 525156
rect 180827 525122 180885 525156
rect 180919 525122 180977 525156
rect 181011 525122 181069 525156
rect 181103 525122 181161 525156
rect 181195 525122 181253 525156
rect 181287 525122 181345 525156
rect 181379 525122 181437 525156
rect 181471 525122 181529 525156
rect 181563 525122 181621 525156
rect 181655 525122 181713 525156
rect 181747 525122 181805 525156
rect 181839 525122 181897 525156
rect 181931 525122 181989 525156
rect 182023 525122 182081 525156
rect 182115 525122 182173 525156
rect 182207 525122 182265 525156
rect 182299 525122 182357 525156
rect 182391 525122 182449 525156
rect 182483 525122 182541 525156
rect 182575 525122 182633 525156
rect 182667 525122 182725 525156
rect 182759 525122 182817 525156
rect 182851 525122 182909 525156
rect 182943 525122 183001 525156
rect 183035 525122 183093 525156
rect 183127 525122 183185 525156
rect 183219 525122 183277 525156
rect 183311 525122 183369 525156
rect 183403 525122 183461 525156
rect 183495 525122 183553 525156
rect 183587 525122 183645 525156
rect 183679 525122 183737 525156
rect 183771 525122 183829 525156
rect 183863 525122 183921 525156
rect 183955 525122 184013 525156
rect 184047 525122 184105 525156
rect 184139 525122 184197 525156
rect 184231 525122 184289 525156
rect 184323 525122 184381 525156
rect 184415 525122 184473 525156
rect 184507 525122 184565 525156
rect 184599 525122 184657 525156
rect 184691 525122 184749 525156
rect 184783 525122 184841 525156
rect 184875 525122 184933 525156
rect 184967 525122 185025 525156
rect 185059 525122 185117 525156
rect 185151 525122 185209 525156
rect 185243 525122 185301 525156
rect 185335 525122 185393 525156
rect 185427 525122 185485 525156
rect 185519 525122 185577 525156
rect 185611 525122 185669 525156
rect 185703 525122 185761 525156
rect 185795 525122 185853 525156
rect 185887 525122 185945 525156
rect 185979 525122 186037 525156
rect 186071 525122 186129 525156
rect 186163 525122 186221 525156
rect 186255 525122 186313 525156
rect 186347 525122 186405 525156
rect 186439 525122 186497 525156
rect 186531 525122 186589 525156
rect 186623 525122 186681 525156
rect 186715 525122 186773 525156
rect 186807 525122 186865 525156
rect 186899 525122 186957 525156
rect 186991 525122 187049 525156
rect 187083 525122 187141 525156
rect 187175 525122 187233 525156
rect 187267 525122 187325 525156
rect 187359 525122 187417 525156
rect 187451 525122 187480 525156
rect 172225 525059 172467 525122
rect 172225 525025 172243 525059
rect 172277 525025 172415 525059
rect 172449 525025 172467 525059
rect 172225 524972 172467 525025
rect 172501 525061 173570 525122
rect 172501 525027 172519 525061
rect 172553 525027 173519 525061
rect 173553 525027 173570 525061
rect 172501 525013 173570 525027
rect 173605 525061 174674 525122
rect 173605 525027 173623 525061
rect 173657 525027 174623 525061
rect 174657 525027 174674 525061
rect 173605 525013 174674 525027
rect 174801 525028 174859 525122
rect 172225 524898 172329 524972
rect 172225 524864 172275 524898
rect 172309 524864 172329 524898
rect 172363 524904 172383 524938
rect 172417 524904 172467 524938
rect 172363 524830 172467 524904
rect 172818 524898 172886 525013
rect 172818 524864 172835 524898
rect 172869 524864 172886 524898
rect 172818 524847 172886 524864
rect 173182 524934 173252 524949
rect 173182 524900 173199 524934
rect 173233 524900 173252 524934
rect 172225 524783 172467 524830
rect 172225 524749 172243 524783
rect 172277 524749 172415 524783
rect 172449 524749 172467 524783
rect 172225 524688 172467 524749
rect 173182 524699 173252 524900
rect 173922 524898 173990 525013
rect 174801 524994 174813 525028
rect 174847 524994 174859 525028
rect 174893 525061 175962 525122
rect 174893 525027 174911 525061
rect 174945 525027 175911 525061
rect 175945 525027 175962 525061
rect 174893 525013 175962 525027
rect 175997 525061 177066 525122
rect 175997 525027 176015 525061
rect 176049 525027 177015 525061
rect 177049 525027 177066 525061
rect 175997 525013 177066 525027
rect 177101 525061 178170 525122
rect 177101 525027 177119 525061
rect 177153 525027 178119 525061
rect 178153 525027 178170 525061
rect 177101 525013 178170 525027
rect 178205 525061 179274 525122
rect 178205 525027 178223 525061
rect 178257 525027 179223 525061
rect 179257 525027 179274 525061
rect 178205 525013 179274 525027
rect 179309 525061 179827 525122
rect 179309 525027 179327 525061
rect 179361 525027 179775 525061
rect 179809 525027 179827 525061
rect 174801 524977 174859 524994
rect 173922 524864 173939 524898
rect 173973 524864 173990 524898
rect 173922 524847 173990 524864
rect 174286 524934 174356 524949
rect 174286 524900 174303 524934
rect 174337 524900 174356 524934
rect 174286 524699 174356 524900
rect 175210 524898 175278 525013
rect 175210 524864 175227 524898
rect 175261 524864 175278 524898
rect 175210 524847 175278 524864
rect 175574 524934 175644 524949
rect 175574 524900 175591 524934
rect 175625 524900 175644 524934
rect 174801 524810 174859 524845
rect 174801 524776 174813 524810
rect 174847 524776 174859 524810
rect 174801 524717 174859 524776
rect 172225 524654 172243 524688
rect 172277 524654 172415 524688
rect 172449 524654 172467 524688
rect 172225 524612 172467 524654
rect 172501 524688 173570 524699
rect 172501 524654 172519 524688
rect 172553 524654 173519 524688
rect 173553 524654 173570 524688
rect 172501 524612 173570 524654
rect 173605 524688 174674 524699
rect 173605 524654 173623 524688
rect 173657 524654 174623 524688
rect 174657 524654 174674 524688
rect 173605 524612 174674 524654
rect 174801 524683 174813 524717
rect 174847 524683 174859 524717
rect 175574 524699 175644 524900
rect 176314 524898 176382 525013
rect 176314 524864 176331 524898
rect 176365 524864 176382 524898
rect 176314 524847 176382 524864
rect 176678 524934 176748 524949
rect 176678 524900 176695 524934
rect 176729 524900 176748 524934
rect 176678 524699 176748 524900
rect 177418 524898 177486 525013
rect 177418 524864 177435 524898
rect 177469 524864 177486 524898
rect 177418 524847 177486 524864
rect 177782 524934 177852 524949
rect 177782 524900 177799 524934
rect 177833 524900 177852 524934
rect 177782 524699 177852 524900
rect 178522 524898 178590 525013
rect 179309 524968 179827 525027
rect 179953 525028 180011 525122
rect 179953 524994 179965 525028
rect 179999 524994 180011 525028
rect 180045 525061 181114 525122
rect 180045 525027 180063 525061
rect 180097 525027 181063 525061
rect 181097 525027 181114 525061
rect 180045 525013 181114 525027
rect 181149 525061 182218 525122
rect 181149 525027 181167 525061
rect 181201 525027 182167 525061
rect 182201 525027 182218 525061
rect 181149 525013 182218 525027
rect 182253 525061 183322 525122
rect 182253 525027 182271 525061
rect 182305 525027 183271 525061
rect 183305 525027 183322 525061
rect 182253 525013 183322 525027
rect 183357 525061 184426 525122
rect 183357 525027 183375 525061
rect 183409 525027 184375 525061
rect 184409 525027 184426 525061
rect 183357 525013 184426 525027
rect 184461 525061 184979 525122
rect 184461 525027 184479 525061
rect 184513 525027 184927 525061
rect 184961 525027 184979 525061
rect 179953 524977 180011 524994
rect 178522 524864 178539 524898
rect 178573 524864 178590 524898
rect 178522 524847 178590 524864
rect 178886 524934 178956 524949
rect 178886 524900 178903 524934
rect 178937 524900 178956 524934
rect 178886 524699 178956 524900
rect 179309 524898 179551 524968
rect 179309 524864 179387 524898
rect 179421 524864 179497 524898
rect 179531 524864 179551 524898
rect 179585 524900 179605 524934
rect 179639 524900 179715 524934
rect 179749 524900 179827 524934
rect 179585 524830 179827 524900
rect 180362 524898 180430 525013
rect 180362 524864 180379 524898
rect 180413 524864 180430 524898
rect 180362 524847 180430 524864
rect 180726 524934 180796 524949
rect 180726 524900 180743 524934
rect 180777 524900 180796 524934
rect 179309 524790 179827 524830
rect 179309 524756 179327 524790
rect 179361 524756 179775 524790
rect 179809 524756 179827 524790
rect 174801 524612 174859 524683
rect 174893 524688 175962 524699
rect 174893 524654 174911 524688
rect 174945 524654 175911 524688
rect 175945 524654 175962 524688
rect 174893 524612 175962 524654
rect 175997 524688 177066 524699
rect 175997 524654 176015 524688
rect 176049 524654 177015 524688
rect 177049 524654 177066 524688
rect 175997 524612 177066 524654
rect 177101 524688 178170 524699
rect 177101 524654 177119 524688
rect 177153 524654 178119 524688
rect 178153 524654 178170 524688
rect 177101 524612 178170 524654
rect 178205 524688 179274 524699
rect 178205 524654 178223 524688
rect 178257 524654 179223 524688
rect 179257 524654 179274 524688
rect 178205 524612 179274 524654
rect 179309 524688 179827 524756
rect 179309 524654 179327 524688
rect 179361 524654 179775 524688
rect 179809 524654 179827 524688
rect 179309 524612 179827 524654
rect 179953 524810 180011 524845
rect 179953 524776 179965 524810
rect 179999 524776 180011 524810
rect 179953 524717 180011 524776
rect 179953 524683 179965 524717
rect 179999 524683 180011 524717
rect 180726 524699 180796 524900
rect 181466 524898 181534 525013
rect 181466 524864 181483 524898
rect 181517 524864 181534 524898
rect 181466 524847 181534 524864
rect 181830 524934 181900 524949
rect 181830 524900 181847 524934
rect 181881 524900 181900 524934
rect 181830 524699 181900 524900
rect 182570 524898 182638 525013
rect 182570 524864 182587 524898
rect 182621 524864 182638 524898
rect 182570 524847 182638 524864
rect 182934 524934 183004 524949
rect 182934 524900 182951 524934
rect 182985 524900 183004 524934
rect 182934 524699 183004 524900
rect 183674 524898 183742 525013
rect 184461 524968 184979 525027
rect 185105 525028 185163 525122
rect 185105 524994 185117 525028
rect 185151 524994 185163 525028
rect 185197 525061 186266 525122
rect 185197 525027 185215 525061
rect 185249 525027 186215 525061
rect 186249 525027 186266 525061
rect 185197 525013 186266 525027
rect 186301 525061 187003 525122
rect 186301 525027 186319 525061
rect 186353 525027 186951 525061
rect 186985 525027 187003 525061
rect 185105 524977 185163 524994
rect 183674 524864 183691 524898
rect 183725 524864 183742 524898
rect 183674 524847 183742 524864
rect 184038 524934 184108 524949
rect 184038 524900 184055 524934
rect 184089 524900 184108 524934
rect 184038 524699 184108 524900
rect 184461 524898 184703 524968
rect 184461 524864 184539 524898
rect 184573 524864 184649 524898
rect 184683 524864 184703 524898
rect 184737 524900 184757 524934
rect 184791 524900 184867 524934
rect 184901 524900 184979 524934
rect 184737 524830 184979 524900
rect 185514 524898 185582 525013
rect 186301 524968 187003 525027
rect 187221 525059 187463 525122
rect 187221 525025 187239 525059
rect 187273 525025 187411 525059
rect 187445 525025 187463 525059
rect 187221 524972 187463 525025
rect 185514 524864 185531 524898
rect 185565 524864 185582 524898
rect 185514 524847 185582 524864
rect 185878 524934 185948 524949
rect 185878 524900 185895 524934
rect 185929 524900 185948 524934
rect 184461 524790 184979 524830
rect 184461 524756 184479 524790
rect 184513 524756 184927 524790
rect 184961 524756 184979 524790
rect 179953 524612 180011 524683
rect 180045 524688 181114 524699
rect 180045 524654 180063 524688
rect 180097 524654 181063 524688
rect 181097 524654 181114 524688
rect 180045 524612 181114 524654
rect 181149 524688 182218 524699
rect 181149 524654 181167 524688
rect 181201 524654 182167 524688
rect 182201 524654 182218 524688
rect 181149 524612 182218 524654
rect 182253 524688 183322 524699
rect 182253 524654 182271 524688
rect 182305 524654 183271 524688
rect 183305 524654 183322 524688
rect 182253 524612 183322 524654
rect 183357 524688 184426 524699
rect 183357 524654 183375 524688
rect 183409 524654 184375 524688
rect 184409 524654 184426 524688
rect 183357 524612 184426 524654
rect 184461 524688 184979 524756
rect 184461 524654 184479 524688
rect 184513 524654 184927 524688
rect 184961 524654 184979 524688
rect 184461 524612 184979 524654
rect 185105 524810 185163 524845
rect 185105 524776 185117 524810
rect 185151 524776 185163 524810
rect 185105 524717 185163 524776
rect 185105 524683 185117 524717
rect 185151 524683 185163 524717
rect 185878 524699 185948 524900
rect 186301 524898 186631 524968
rect 186301 524864 186379 524898
rect 186413 524864 186478 524898
rect 186512 524864 186577 524898
rect 186611 524864 186631 524898
rect 186665 524900 186685 524934
rect 186719 524900 186788 524934
rect 186822 524900 186891 524934
rect 186925 524900 187003 524934
rect 186665 524830 187003 524900
rect 186301 524790 187003 524830
rect 186301 524756 186319 524790
rect 186353 524756 186951 524790
rect 186985 524756 187003 524790
rect 185105 524612 185163 524683
rect 185197 524688 186266 524699
rect 185197 524654 185215 524688
rect 185249 524654 186215 524688
rect 186249 524654 186266 524688
rect 185197 524612 186266 524654
rect 186301 524688 187003 524756
rect 186301 524654 186319 524688
rect 186353 524654 186951 524688
rect 186985 524654 187003 524688
rect 186301 524612 187003 524654
rect 187221 524904 187271 524938
rect 187305 524904 187325 524938
rect 187221 524830 187325 524904
rect 187359 524898 187463 524972
rect 187359 524864 187379 524898
rect 187413 524864 187463 524898
rect 187221 524783 187463 524830
rect 187221 524749 187239 524783
rect 187273 524749 187411 524783
rect 187445 524749 187463 524783
rect 187221 524688 187463 524749
rect 187221 524654 187239 524688
rect 187273 524654 187411 524688
rect 187445 524654 187463 524688
rect 187221 524612 187463 524654
rect 172208 524578 172237 524612
rect 172271 524578 172329 524612
rect 172363 524578 172421 524612
rect 172455 524578 172513 524612
rect 172547 524578 172605 524612
rect 172639 524578 172697 524612
rect 172731 524578 172789 524612
rect 172823 524578 172881 524612
rect 172915 524578 172973 524612
rect 173007 524578 173065 524612
rect 173099 524578 173157 524612
rect 173191 524578 173249 524612
rect 173283 524578 173341 524612
rect 173375 524578 173433 524612
rect 173467 524578 173525 524612
rect 173559 524578 173617 524612
rect 173651 524578 173709 524612
rect 173743 524578 173801 524612
rect 173835 524578 173893 524612
rect 173927 524578 173985 524612
rect 174019 524578 174077 524612
rect 174111 524578 174169 524612
rect 174203 524578 174261 524612
rect 174295 524578 174353 524612
rect 174387 524578 174445 524612
rect 174479 524578 174537 524612
rect 174571 524578 174629 524612
rect 174663 524578 174721 524612
rect 174755 524578 174813 524612
rect 174847 524578 174905 524612
rect 174939 524578 174997 524612
rect 175031 524578 175089 524612
rect 175123 524578 175181 524612
rect 175215 524578 175273 524612
rect 175307 524578 175365 524612
rect 175399 524578 175457 524612
rect 175491 524578 175549 524612
rect 175583 524578 175641 524612
rect 175675 524578 175733 524612
rect 175767 524578 175825 524612
rect 175859 524578 175917 524612
rect 175951 524578 176009 524612
rect 176043 524578 176101 524612
rect 176135 524578 176193 524612
rect 176227 524578 176285 524612
rect 176319 524578 176377 524612
rect 176411 524578 176469 524612
rect 176503 524578 176561 524612
rect 176595 524578 176653 524612
rect 176687 524578 176745 524612
rect 176779 524578 176837 524612
rect 176871 524578 176929 524612
rect 176963 524578 177021 524612
rect 177055 524578 177113 524612
rect 177147 524578 177205 524612
rect 177239 524578 177297 524612
rect 177331 524578 177389 524612
rect 177423 524578 177481 524612
rect 177515 524578 177573 524612
rect 177607 524578 177665 524612
rect 177699 524578 177757 524612
rect 177791 524578 177849 524612
rect 177883 524578 177941 524612
rect 177975 524578 178033 524612
rect 178067 524578 178125 524612
rect 178159 524578 178217 524612
rect 178251 524578 178309 524612
rect 178343 524578 178401 524612
rect 178435 524578 178493 524612
rect 178527 524578 178585 524612
rect 178619 524578 178677 524612
rect 178711 524578 178769 524612
rect 178803 524578 178861 524612
rect 178895 524578 178953 524612
rect 178987 524578 179045 524612
rect 179079 524578 179137 524612
rect 179171 524578 179229 524612
rect 179263 524578 179321 524612
rect 179355 524578 179413 524612
rect 179447 524578 179505 524612
rect 179539 524578 179597 524612
rect 179631 524578 179689 524612
rect 179723 524578 179781 524612
rect 179815 524578 179873 524612
rect 179907 524578 179965 524612
rect 179999 524578 180057 524612
rect 180091 524578 180149 524612
rect 180183 524578 180241 524612
rect 180275 524578 180333 524612
rect 180367 524578 180425 524612
rect 180459 524578 180517 524612
rect 180551 524578 180609 524612
rect 180643 524578 180701 524612
rect 180735 524578 180793 524612
rect 180827 524578 180885 524612
rect 180919 524578 180977 524612
rect 181011 524578 181069 524612
rect 181103 524578 181161 524612
rect 181195 524578 181253 524612
rect 181287 524578 181345 524612
rect 181379 524578 181437 524612
rect 181471 524578 181529 524612
rect 181563 524578 181621 524612
rect 181655 524578 181713 524612
rect 181747 524578 181805 524612
rect 181839 524578 181897 524612
rect 181931 524578 181989 524612
rect 182023 524578 182081 524612
rect 182115 524578 182173 524612
rect 182207 524578 182265 524612
rect 182299 524578 182357 524612
rect 182391 524578 182449 524612
rect 182483 524578 182541 524612
rect 182575 524578 182633 524612
rect 182667 524578 182725 524612
rect 182759 524578 182817 524612
rect 182851 524578 182909 524612
rect 182943 524578 183001 524612
rect 183035 524578 183093 524612
rect 183127 524578 183185 524612
rect 183219 524578 183277 524612
rect 183311 524578 183369 524612
rect 183403 524578 183461 524612
rect 183495 524578 183553 524612
rect 183587 524578 183645 524612
rect 183679 524578 183737 524612
rect 183771 524578 183829 524612
rect 183863 524578 183921 524612
rect 183955 524578 184013 524612
rect 184047 524578 184105 524612
rect 184139 524578 184197 524612
rect 184231 524578 184289 524612
rect 184323 524578 184381 524612
rect 184415 524578 184473 524612
rect 184507 524578 184565 524612
rect 184599 524578 184657 524612
rect 184691 524578 184749 524612
rect 184783 524578 184841 524612
rect 184875 524578 184933 524612
rect 184967 524578 185025 524612
rect 185059 524578 185117 524612
rect 185151 524578 185209 524612
rect 185243 524578 185301 524612
rect 185335 524578 185393 524612
rect 185427 524578 185485 524612
rect 185519 524578 185577 524612
rect 185611 524578 185669 524612
rect 185703 524578 185761 524612
rect 185795 524578 185853 524612
rect 185887 524578 185945 524612
rect 185979 524578 186037 524612
rect 186071 524578 186129 524612
rect 186163 524578 186221 524612
rect 186255 524578 186313 524612
rect 186347 524578 186405 524612
rect 186439 524578 186497 524612
rect 186531 524578 186589 524612
rect 186623 524578 186681 524612
rect 186715 524578 186773 524612
rect 186807 524578 186865 524612
rect 186899 524578 186957 524612
rect 186991 524578 187049 524612
rect 187083 524578 187141 524612
rect 187175 524578 187233 524612
rect 187267 524578 187325 524612
rect 187359 524578 187417 524612
rect 187451 524578 187480 524612
rect 172225 524536 172467 524578
rect 172225 524502 172243 524536
rect 172277 524502 172415 524536
rect 172449 524502 172467 524536
rect 172225 524441 172467 524502
rect 172501 524536 173570 524578
rect 172501 524502 172519 524536
rect 172553 524502 173519 524536
rect 173553 524502 173570 524536
rect 172501 524491 173570 524502
rect 173605 524536 174674 524578
rect 173605 524502 173623 524536
rect 173657 524502 174623 524536
rect 174657 524502 174674 524536
rect 173605 524491 174674 524502
rect 174709 524536 175778 524578
rect 174709 524502 174727 524536
rect 174761 524502 175727 524536
rect 175761 524502 175778 524536
rect 174709 524491 175778 524502
rect 175813 524536 176882 524578
rect 175813 524502 175831 524536
rect 175865 524502 176831 524536
rect 176865 524502 176882 524536
rect 175813 524491 176882 524502
rect 176917 524536 177251 524578
rect 176917 524502 176935 524536
rect 176969 524502 177199 524536
rect 177233 524502 177251 524536
rect 172225 524407 172243 524441
rect 172277 524407 172415 524441
rect 172449 524407 172467 524441
rect 172225 524360 172467 524407
rect 172225 524292 172275 524326
rect 172309 524292 172329 524326
rect 172225 524218 172329 524292
rect 172363 524286 172467 524360
rect 172363 524252 172383 524286
rect 172417 524252 172467 524286
rect 172818 524326 172886 524343
rect 172818 524292 172835 524326
rect 172869 524292 172886 524326
rect 172225 524165 172467 524218
rect 172818 524177 172886 524292
rect 173182 524290 173252 524491
rect 173182 524256 173199 524290
rect 173233 524256 173252 524290
rect 173182 524241 173252 524256
rect 173922 524326 173990 524343
rect 173922 524292 173939 524326
rect 173973 524292 173990 524326
rect 173922 524177 173990 524292
rect 174286 524290 174356 524491
rect 174286 524256 174303 524290
rect 174337 524256 174356 524290
rect 174286 524241 174356 524256
rect 175026 524326 175094 524343
rect 175026 524292 175043 524326
rect 175077 524292 175094 524326
rect 175026 524177 175094 524292
rect 175390 524290 175460 524491
rect 175390 524256 175407 524290
rect 175441 524256 175460 524290
rect 175390 524241 175460 524256
rect 176130 524326 176198 524343
rect 176130 524292 176147 524326
rect 176181 524292 176198 524326
rect 176130 524177 176198 524292
rect 176494 524290 176564 524491
rect 176917 524434 177251 524502
rect 176917 524400 176935 524434
rect 176969 524400 177199 524434
rect 177233 524400 177251 524434
rect 176917 524360 177251 524400
rect 176494 524256 176511 524290
rect 176545 524256 176564 524290
rect 176494 524241 176564 524256
rect 176917 524292 176937 524326
rect 176971 524292 177067 524326
rect 176917 524222 177067 524292
rect 177101 524290 177251 524360
rect 177377 524507 177435 524578
rect 177377 524473 177389 524507
rect 177423 524473 177435 524507
rect 177469 524536 178538 524578
rect 177469 524502 177487 524536
rect 177521 524502 178487 524536
rect 178521 524502 178538 524536
rect 177469 524491 178538 524502
rect 178573 524536 179642 524578
rect 178573 524502 178591 524536
rect 178625 524502 179591 524536
rect 179625 524502 179642 524536
rect 178573 524491 179642 524502
rect 179677 524536 180746 524578
rect 179677 524502 179695 524536
rect 179729 524502 180695 524536
rect 180729 524502 180746 524536
rect 179677 524491 180746 524502
rect 180781 524536 181850 524578
rect 180781 524502 180799 524536
rect 180833 524502 181799 524536
rect 181833 524502 181850 524536
rect 180781 524491 181850 524502
rect 181885 524536 182403 524578
rect 181885 524502 181903 524536
rect 181937 524502 182351 524536
rect 182385 524502 182403 524536
rect 177377 524414 177435 524473
rect 177377 524380 177389 524414
rect 177423 524380 177435 524414
rect 177377 524345 177435 524380
rect 177101 524256 177197 524290
rect 177231 524256 177251 524290
rect 177786 524326 177854 524343
rect 177786 524292 177803 524326
rect 177837 524292 177854 524326
rect 172225 524131 172243 524165
rect 172277 524131 172415 524165
rect 172449 524131 172467 524165
rect 172225 524068 172467 524131
rect 172501 524163 173570 524177
rect 172501 524129 172519 524163
rect 172553 524129 173519 524163
rect 173553 524129 173570 524163
rect 172501 524068 173570 524129
rect 173605 524163 174674 524177
rect 173605 524129 173623 524163
rect 173657 524129 174623 524163
rect 174657 524129 174674 524163
rect 173605 524068 174674 524129
rect 174709 524163 175778 524177
rect 174709 524129 174727 524163
rect 174761 524129 175727 524163
rect 175761 524129 175778 524163
rect 174709 524068 175778 524129
rect 175813 524163 176882 524177
rect 175813 524129 175831 524163
rect 175865 524129 176831 524163
rect 176865 524129 176882 524163
rect 175813 524068 176882 524129
rect 176917 524170 177251 524222
rect 176917 524136 176935 524170
rect 176969 524136 177199 524170
rect 177233 524136 177251 524170
rect 176917 524068 177251 524136
rect 177377 524196 177435 524213
rect 177377 524162 177389 524196
rect 177423 524162 177435 524196
rect 177786 524177 177854 524292
rect 178150 524290 178220 524491
rect 178150 524256 178167 524290
rect 178201 524256 178220 524290
rect 178150 524241 178220 524256
rect 178890 524326 178958 524343
rect 178890 524292 178907 524326
rect 178941 524292 178958 524326
rect 178890 524177 178958 524292
rect 179254 524290 179324 524491
rect 179254 524256 179271 524290
rect 179305 524256 179324 524290
rect 179254 524241 179324 524256
rect 179994 524326 180062 524343
rect 179994 524292 180011 524326
rect 180045 524292 180062 524326
rect 179994 524177 180062 524292
rect 180358 524290 180428 524491
rect 180358 524256 180375 524290
rect 180409 524256 180428 524290
rect 180358 524241 180428 524256
rect 181098 524326 181166 524343
rect 181098 524292 181115 524326
rect 181149 524292 181166 524326
rect 181098 524177 181166 524292
rect 181462 524290 181532 524491
rect 181885 524434 182403 524502
rect 181885 524400 181903 524434
rect 181937 524400 182351 524434
rect 182385 524400 182403 524434
rect 181885 524360 182403 524400
rect 181462 524256 181479 524290
rect 181513 524256 181532 524290
rect 181462 524241 181532 524256
rect 181885 524292 181963 524326
rect 181997 524292 182073 524326
rect 182107 524292 182127 524326
rect 181885 524222 182127 524292
rect 182161 524290 182403 524360
rect 182529 524507 182587 524578
rect 182529 524473 182541 524507
rect 182575 524473 182587 524507
rect 182621 524536 183690 524578
rect 182621 524502 182639 524536
rect 182673 524502 183639 524536
rect 183673 524502 183690 524536
rect 182621 524491 183690 524502
rect 183725 524536 184794 524578
rect 183725 524502 183743 524536
rect 183777 524502 184743 524536
rect 184777 524502 184794 524536
rect 183725 524491 184794 524502
rect 184829 524536 185898 524578
rect 184829 524502 184847 524536
rect 184881 524502 185847 524536
rect 185881 524502 185898 524536
rect 184829 524491 185898 524502
rect 185933 524536 187002 524578
rect 185933 524502 185951 524536
rect 185985 524502 186951 524536
rect 186985 524502 187002 524536
rect 185933 524491 187002 524502
rect 187221 524536 187463 524578
rect 187221 524502 187239 524536
rect 187273 524502 187411 524536
rect 187445 524502 187463 524536
rect 182529 524414 182587 524473
rect 182529 524380 182541 524414
rect 182575 524380 182587 524414
rect 182529 524345 182587 524380
rect 182161 524256 182181 524290
rect 182215 524256 182291 524290
rect 182325 524256 182403 524290
rect 182938 524326 183006 524343
rect 182938 524292 182955 524326
rect 182989 524292 183006 524326
rect 177377 524068 177435 524162
rect 177469 524163 178538 524177
rect 177469 524129 177487 524163
rect 177521 524129 178487 524163
rect 178521 524129 178538 524163
rect 177469 524068 178538 524129
rect 178573 524163 179642 524177
rect 178573 524129 178591 524163
rect 178625 524129 179591 524163
rect 179625 524129 179642 524163
rect 178573 524068 179642 524129
rect 179677 524163 180746 524177
rect 179677 524129 179695 524163
rect 179729 524129 180695 524163
rect 180729 524129 180746 524163
rect 179677 524068 180746 524129
rect 180781 524163 181850 524177
rect 180781 524129 180799 524163
rect 180833 524129 181799 524163
rect 181833 524129 181850 524163
rect 180781 524068 181850 524129
rect 181885 524163 182403 524222
rect 181885 524129 181903 524163
rect 181937 524129 182351 524163
rect 182385 524129 182403 524163
rect 181885 524068 182403 524129
rect 182529 524196 182587 524213
rect 182529 524162 182541 524196
rect 182575 524162 182587 524196
rect 182938 524177 183006 524292
rect 183302 524290 183372 524491
rect 183302 524256 183319 524290
rect 183353 524256 183372 524290
rect 183302 524241 183372 524256
rect 184042 524326 184110 524343
rect 184042 524292 184059 524326
rect 184093 524292 184110 524326
rect 184042 524177 184110 524292
rect 184406 524290 184476 524491
rect 184406 524256 184423 524290
rect 184457 524256 184476 524290
rect 184406 524241 184476 524256
rect 185146 524326 185214 524343
rect 185146 524292 185163 524326
rect 185197 524292 185214 524326
rect 185146 524177 185214 524292
rect 185510 524290 185580 524491
rect 185510 524256 185527 524290
rect 185561 524256 185580 524290
rect 185510 524241 185580 524256
rect 186250 524326 186318 524343
rect 186250 524292 186267 524326
rect 186301 524292 186318 524326
rect 186250 524177 186318 524292
rect 186614 524290 186684 524491
rect 186614 524256 186631 524290
rect 186665 524256 186684 524290
rect 186614 524241 186684 524256
rect 187221 524441 187463 524502
rect 187221 524407 187239 524441
rect 187273 524407 187411 524441
rect 187445 524407 187463 524441
rect 187221 524360 187463 524407
rect 187221 524286 187325 524360
rect 187221 524252 187271 524286
rect 187305 524252 187325 524286
rect 187359 524292 187379 524326
rect 187413 524292 187463 524326
rect 187359 524218 187463 524292
rect 182529 524068 182587 524162
rect 182621 524163 183690 524177
rect 182621 524129 182639 524163
rect 182673 524129 183639 524163
rect 183673 524129 183690 524163
rect 182621 524068 183690 524129
rect 183725 524163 184794 524177
rect 183725 524129 183743 524163
rect 183777 524129 184743 524163
rect 184777 524129 184794 524163
rect 183725 524068 184794 524129
rect 184829 524163 185898 524177
rect 184829 524129 184847 524163
rect 184881 524129 185847 524163
rect 185881 524129 185898 524163
rect 184829 524068 185898 524129
rect 185933 524163 187002 524177
rect 185933 524129 185951 524163
rect 185985 524129 186951 524163
rect 186985 524129 187002 524163
rect 185933 524068 187002 524129
rect 187221 524165 187463 524218
rect 187221 524131 187239 524165
rect 187273 524131 187411 524165
rect 187445 524131 187463 524165
rect 187221 524068 187463 524131
rect 172208 524034 172237 524068
rect 172271 524034 172329 524068
rect 172363 524034 172421 524068
rect 172455 524034 172513 524068
rect 172547 524034 172605 524068
rect 172639 524034 172697 524068
rect 172731 524034 172789 524068
rect 172823 524034 172881 524068
rect 172915 524034 172973 524068
rect 173007 524034 173065 524068
rect 173099 524034 173157 524068
rect 173191 524034 173249 524068
rect 173283 524034 173341 524068
rect 173375 524034 173433 524068
rect 173467 524034 173525 524068
rect 173559 524034 173617 524068
rect 173651 524034 173709 524068
rect 173743 524034 173801 524068
rect 173835 524034 173893 524068
rect 173927 524034 173985 524068
rect 174019 524034 174077 524068
rect 174111 524034 174169 524068
rect 174203 524034 174261 524068
rect 174295 524034 174353 524068
rect 174387 524034 174445 524068
rect 174479 524034 174537 524068
rect 174571 524034 174629 524068
rect 174663 524034 174721 524068
rect 174755 524034 174813 524068
rect 174847 524034 174905 524068
rect 174939 524034 174997 524068
rect 175031 524034 175089 524068
rect 175123 524034 175181 524068
rect 175215 524034 175273 524068
rect 175307 524034 175365 524068
rect 175399 524034 175457 524068
rect 175491 524034 175549 524068
rect 175583 524034 175641 524068
rect 175675 524034 175733 524068
rect 175767 524034 175825 524068
rect 175859 524034 175917 524068
rect 175951 524034 176009 524068
rect 176043 524034 176101 524068
rect 176135 524034 176193 524068
rect 176227 524034 176285 524068
rect 176319 524034 176377 524068
rect 176411 524034 176469 524068
rect 176503 524034 176561 524068
rect 176595 524034 176653 524068
rect 176687 524034 176745 524068
rect 176779 524034 176837 524068
rect 176871 524034 176929 524068
rect 176963 524034 177021 524068
rect 177055 524034 177113 524068
rect 177147 524034 177205 524068
rect 177239 524034 177297 524068
rect 177331 524034 177389 524068
rect 177423 524034 177481 524068
rect 177515 524034 177573 524068
rect 177607 524034 177665 524068
rect 177699 524034 177757 524068
rect 177791 524034 177849 524068
rect 177883 524034 177941 524068
rect 177975 524034 178033 524068
rect 178067 524034 178125 524068
rect 178159 524034 178217 524068
rect 178251 524034 178309 524068
rect 178343 524034 178401 524068
rect 178435 524034 178493 524068
rect 178527 524034 178585 524068
rect 178619 524034 178677 524068
rect 178711 524034 178769 524068
rect 178803 524034 178861 524068
rect 178895 524034 178953 524068
rect 178987 524034 179045 524068
rect 179079 524034 179137 524068
rect 179171 524034 179229 524068
rect 179263 524034 179321 524068
rect 179355 524034 179413 524068
rect 179447 524034 179505 524068
rect 179539 524034 179597 524068
rect 179631 524034 179689 524068
rect 179723 524034 179781 524068
rect 179815 524034 179873 524068
rect 179907 524034 179965 524068
rect 179999 524034 180057 524068
rect 180091 524034 180149 524068
rect 180183 524034 180241 524068
rect 180275 524034 180333 524068
rect 180367 524034 180425 524068
rect 180459 524034 180517 524068
rect 180551 524034 180609 524068
rect 180643 524034 180701 524068
rect 180735 524034 180793 524068
rect 180827 524034 180885 524068
rect 180919 524034 180977 524068
rect 181011 524034 181069 524068
rect 181103 524034 181161 524068
rect 181195 524034 181253 524068
rect 181287 524034 181345 524068
rect 181379 524034 181437 524068
rect 181471 524034 181529 524068
rect 181563 524034 181621 524068
rect 181655 524034 181713 524068
rect 181747 524034 181805 524068
rect 181839 524034 181897 524068
rect 181931 524034 181989 524068
rect 182023 524034 182081 524068
rect 182115 524034 182173 524068
rect 182207 524034 182265 524068
rect 182299 524034 182357 524068
rect 182391 524034 182449 524068
rect 182483 524034 182541 524068
rect 182575 524034 182633 524068
rect 182667 524034 182725 524068
rect 182759 524034 182817 524068
rect 182851 524034 182909 524068
rect 182943 524034 183001 524068
rect 183035 524034 183093 524068
rect 183127 524034 183185 524068
rect 183219 524034 183277 524068
rect 183311 524034 183369 524068
rect 183403 524034 183461 524068
rect 183495 524034 183553 524068
rect 183587 524034 183645 524068
rect 183679 524034 183737 524068
rect 183771 524034 183829 524068
rect 183863 524034 183921 524068
rect 183955 524034 184013 524068
rect 184047 524034 184105 524068
rect 184139 524034 184197 524068
rect 184231 524034 184289 524068
rect 184323 524034 184381 524068
rect 184415 524034 184473 524068
rect 184507 524034 184565 524068
rect 184599 524034 184657 524068
rect 184691 524034 184749 524068
rect 184783 524034 184841 524068
rect 184875 524034 184933 524068
rect 184967 524034 185025 524068
rect 185059 524034 185117 524068
rect 185151 524034 185209 524068
rect 185243 524034 185301 524068
rect 185335 524034 185393 524068
rect 185427 524034 185485 524068
rect 185519 524034 185577 524068
rect 185611 524034 185669 524068
rect 185703 524034 185761 524068
rect 185795 524034 185853 524068
rect 185887 524034 185945 524068
rect 185979 524034 186037 524068
rect 186071 524034 186129 524068
rect 186163 524034 186221 524068
rect 186255 524034 186313 524068
rect 186347 524034 186405 524068
rect 186439 524034 186497 524068
rect 186531 524034 186589 524068
rect 186623 524034 186681 524068
rect 186715 524034 186773 524068
rect 186807 524034 186865 524068
rect 186899 524034 186957 524068
rect 186991 524034 187049 524068
rect 187083 524034 187141 524068
rect 187175 524034 187233 524068
rect 187267 524034 187325 524068
rect 187359 524034 187417 524068
rect 187451 524034 187480 524068
rect 172225 523971 172467 524034
rect 172225 523937 172243 523971
rect 172277 523937 172415 523971
rect 172449 523937 172467 523971
rect 172225 523884 172467 523937
rect 172501 523973 173570 524034
rect 172501 523939 172519 523973
rect 172553 523939 173519 523973
rect 173553 523939 173570 523973
rect 172501 523925 173570 523939
rect 173605 523973 174674 524034
rect 173605 523939 173623 523973
rect 173657 523939 174623 523973
rect 174657 523939 174674 523973
rect 173605 523925 174674 523939
rect 174801 523940 174859 524034
rect 172225 523810 172329 523884
rect 172225 523776 172275 523810
rect 172309 523776 172329 523810
rect 172363 523816 172383 523850
rect 172417 523816 172467 523850
rect 172363 523742 172467 523816
rect 172818 523810 172886 523925
rect 172818 523776 172835 523810
rect 172869 523776 172886 523810
rect 172818 523759 172886 523776
rect 173182 523846 173252 523861
rect 173182 523812 173199 523846
rect 173233 523812 173252 523846
rect 172225 523695 172467 523742
rect 172225 523661 172243 523695
rect 172277 523661 172415 523695
rect 172449 523661 172467 523695
rect 172225 523600 172467 523661
rect 173182 523611 173252 523812
rect 173922 523810 173990 523925
rect 174801 523906 174813 523940
rect 174847 523906 174859 523940
rect 174893 523973 175962 524034
rect 174893 523939 174911 523973
rect 174945 523939 175911 523973
rect 175945 523939 175962 523973
rect 174893 523925 175962 523939
rect 175997 523973 177066 524034
rect 175997 523939 176015 523973
rect 176049 523939 177015 523973
rect 177049 523939 177066 523973
rect 175997 523925 177066 523939
rect 177101 523973 178170 524034
rect 177101 523939 177119 523973
rect 177153 523939 178119 523973
rect 178153 523939 178170 523973
rect 177101 523925 178170 523939
rect 178205 523973 179274 524034
rect 178205 523939 178223 523973
rect 178257 523939 179223 523973
rect 179257 523939 179274 523973
rect 178205 523925 179274 523939
rect 179309 523973 179827 524034
rect 179309 523939 179327 523973
rect 179361 523939 179775 523973
rect 179809 523939 179827 523973
rect 174801 523889 174859 523906
rect 173922 523776 173939 523810
rect 173973 523776 173990 523810
rect 173922 523759 173990 523776
rect 174286 523846 174356 523861
rect 174286 523812 174303 523846
rect 174337 523812 174356 523846
rect 174286 523611 174356 523812
rect 175210 523810 175278 523925
rect 175210 523776 175227 523810
rect 175261 523776 175278 523810
rect 175210 523759 175278 523776
rect 175574 523846 175644 523861
rect 175574 523812 175591 523846
rect 175625 523812 175644 523846
rect 174801 523722 174859 523757
rect 174801 523688 174813 523722
rect 174847 523688 174859 523722
rect 174801 523629 174859 523688
rect 172225 523566 172243 523600
rect 172277 523566 172415 523600
rect 172449 523566 172467 523600
rect 172225 523524 172467 523566
rect 172501 523600 173570 523611
rect 172501 523566 172519 523600
rect 172553 523566 173519 523600
rect 173553 523566 173570 523600
rect 172501 523524 173570 523566
rect 173605 523600 174674 523611
rect 173605 523566 173623 523600
rect 173657 523566 174623 523600
rect 174657 523566 174674 523600
rect 173605 523524 174674 523566
rect 174801 523595 174813 523629
rect 174847 523595 174859 523629
rect 175574 523611 175644 523812
rect 176314 523810 176382 523925
rect 176314 523776 176331 523810
rect 176365 523776 176382 523810
rect 176314 523759 176382 523776
rect 176678 523846 176748 523861
rect 176678 523812 176695 523846
rect 176729 523812 176748 523846
rect 176678 523611 176748 523812
rect 177418 523810 177486 523925
rect 177418 523776 177435 523810
rect 177469 523776 177486 523810
rect 177418 523759 177486 523776
rect 177782 523846 177852 523861
rect 177782 523812 177799 523846
rect 177833 523812 177852 523846
rect 177782 523611 177852 523812
rect 178522 523810 178590 523925
rect 179309 523880 179827 523939
rect 179953 523940 180011 524034
rect 179953 523906 179965 523940
rect 179999 523906 180011 523940
rect 180045 523973 181114 524034
rect 180045 523939 180063 523973
rect 180097 523939 181063 523973
rect 181097 523939 181114 523973
rect 180045 523925 181114 523939
rect 181149 523973 182218 524034
rect 181149 523939 181167 523973
rect 181201 523939 182167 523973
rect 182201 523939 182218 523973
rect 181149 523925 182218 523939
rect 182253 523973 183322 524034
rect 182253 523939 182271 523973
rect 182305 523939 183271 523973
rect 183305 523939 183322 523973
rect 182253 523925 183322 523939
rect 183357 523973 184426 524034
rect 183357 523939 183375 523973
rect 183409 523939 184375 523973
rect 184409 523939 184426 523973
rect 183357 523925 184426 523939
rect 184461 523973 184979 524034
rect 184461 523939 184479 523973
rect 184513 523939 184927 523973
rect 184961 523939 184979 523973
rect 179953 523889 180011 523906
rect 178522 523776 178539 523810
rect 178573 523776 178590 523810
rect 178522 523759 178590 523776
rect 178886 523846 178956 523861
rect 178886 523812 178903 523846
rect 178937 523812 178956 523846
rect 178886 523611 178956 523812
rect 179309 523810 179551 523880
rect 179309 523776 179387 523810
rect 179421 523776 179497 523810
rect 179531 523776 179551 523810
rect 179585 523812 179605 523846
rect 179639 523812 179715 523846
rect 179749 523812 179827 523846
rect 179585 523742 179827 523812
rect 180362 523810 180430 523925
rect 180362 523776 180379 523810
rect 180413 523776 180430 523810
rect 180362 523759 180430 523776
rect 180726 523846 180796 523861
rect 180726 523812 180743 523846
rect 180777 523812 180796 523846
rect 179309 523702 179827 523742
rect 179309 523668 179327 523702
rect 179361 523668 179775 523702
rect 179809 523668 179827 523702
rect 174801 523524 174859 523595
rect 174893 523600 175962 523611
rect 174893 523566 174911 523600
rect 174945 523566 175911 523600
rect 175945 523566 175962 523600
rect 174893 523524 175962 523566
rect 175997 523600 177066 523611
rect 175997 523566 176015 523600
rect 176049 523566 177015 523600
rect 177049 523566 177066 523600
rect 175997 523524 177066 523566
rect 177101 523600 178170 523611
rect 177101 523566 177119 523600
rect 177153 523566 178119 523600
rect 178153 523566 178170 523600
rect 177101 523524 178170 523566
rect 178205 523600 179274 523611
rect 178205 523566 178223 523600
rect 178257 523566 179223 523600
rect 179257 523566 179274 523600
rect 178205 523524 179274 523566
rect 179309 523600 179827 523668
rect 179309 523566 179327 523600
rect 179361 523566 179775 523600
rect 179809 523566 179827 523600
rect 179309 523524 179827 523566
rect 179953 523722 180011 523757
rect 179953 523688 179965 523722
rect 179999 523688 180011 523722
rect 179953 523629 180011 523688
rect 179953 523595 179965 523629
rect 179999 523595 180011 523629
rect 180726 523611 180796 523812
rect 181466 523810 181534 523925
rect 181466 523776 181483 523810
rect 181517 523776 181534 523810
rect 181466 523759 181534 523776
rect 181830 523846 181900 523861
rect 181830 523812 181847 523846
rect 181881 523812 181900 523846
rect 181830 523611 181900 523812
rect 182570 523810 182638 523925
rect 182570 523776 182587 523810
rect 182621 523776 182638 523810
rect 182570 523759 182638 523776
rect 182934 523846 183004 523861
rect 182934 523812 182951 523846
rect 182985 523812 183004 523846
rect 182934 523611 183004 523812
rect 183674 523810 183742 523925
rect 184461 523880 184979 523939
rect 185105 523940 185163 524034
rect 185105 523906 185117 523940
rect 185151 523906 185163 523940
rect 185197 523973 186266 524034
rect 185197 523939 185215 523973
rect 185249 523939 186215 523973
rect 186249 523939 186266 523973
rect 185197 523925 186266 523939
rect 186301 523973 187003 524034
rect 186301 523939 186319 523973
rect 186353 523939 186951 523973
rect 186985 523939 187003 523973
rect 185105 523889 185163 523906
rect 183674 523776 183691 523810
rect 183725 523776 183742 523810
rect 183674 523759 183742 523776
rect 184038 523846 184108 523861
rect 184038 523812 184055 523846
rect 184089 523812 184108 523846
rect 184038 523611 184108 523812
rect 184461 523810 184703 523880
rect 184461 523776 184539 523810
rect 184573 523776 184649 523810
rect 184683 523776 184703 523810
rect 184737 523812 184757 523846
rect 184791 523812 184867 523846
rect 184901 523812 184979 523846
rect 184737 523742 184979 523812
rect 185514 523810 185582 523925
rect 186301 523880 187003 523939
rect 187221 523971 187463 524034
rect 187221 523937 187239 523971
rect 187273 523937 187411 523971
rect 187445 523937 187463 523971
rect 187221 523884 187463 523937
rect 185514 523776 185531 523810
rect 185565 523776 185582 523810
rect 185514 523759 185582 523776
rect 185878 523846 185948 523861
rect 185878 523812 185895 523846
rect 185929 523812 185948 523846
rect 184461 523702 184979 523742
rect 184461 523668 184479 523702
rect 184513 523668 184927 523702
rect 184961 523668 184979 523702
rect 179953 523524 180011 523595
rect 180045 523600 181114 523611
rect 180045 523566 180063 523600
rect 180097 523566 181063 523600
rect 181097 523566 181114 523600
rect 180045 523524 181114 523566
rect 181149 523600 182218 523611
rect 181149 523566 181167 523600
rect 181201 523566 182167 523600
rect 182201 523566 182218 523600
rect 181149 523524 182218 523566
rect 182253 523600 183322 523611
rect 182253 523566 182271 523600
rect 182305 523566 183271 523600
rect 183305 523566 183322 523600
rect 182253 523524 183322 523566
rect 183357 523600 184426 523611
rect 183357 523566 183375 523600
rect 183409 523566 184375 523600
rect 184409 523566 184426 523600
rect 183357 523524 184426 523566
rect 184461 523600 184979 523668
rect 184461 523566 184479 523600
rect 184513 523566 184927 523600
rect 184961 523566 184979 523600
rect 184461 523524 184979 523566
rect 185105 523722 185163 523757
rect 185105 523688 185117 523722
rect 185151 523688 185163 523722
rect 185105 523629 185163 523688
rect 185105 523595 185117 523629
rect 185151 523595 185163 523629
rect 185878 523611 185948 523812
rect 186301 523810 186631 523880
rect 186301 523776 186379 523810
rect 186413 523776 186478 523810
rect 186512 523776 186577 523810
rect 186611 523776 186631 523810
rect 186665 523812 186685 523846
rect 186719 523812 186788 523846
rect 186822 523812 186891 523846
rect 186925 523812 187003 523846
rect 186665 523742 187003 523812
rect 186301 523702 187003 523742
rect 186301 523668 186319 523702
rect 186353 523668 186951 523702
rect 186985 523668 187003 523702
rect 185105 523524 185163 523595
rect 185197 523600 186266 523611
rect 185197 523566 185215 523600
rect 185249 523566 186215 523600
rect 186249 523566 186266 523600
rect 185197 523524 186266 523566
rect 186301 523600 187003 523668
rect 186301 523566 186319 523600
rect 186353 523566 186951 523600
rect 186985 523566 187003 523600
rect 186301 523524 187003 523566
rect 187221 523816 187271 523850
rect 187305 523816 187325 523850
rect 187221 523742 187325 523816
rect 187359 523810 187463 523884
rect 187359 523776 187379 523810
rect 187413 523776 187463 523810
rect 187221 523695 187463 523742
rect 187221 523661 187239 523695
rect 187273 523661 187411 523695
rect 187445 523661 187463 523695
rect 187221 523600 187463 523661
rect 187221 523566 187239 523600
rect 187273 523566 187411 523600
rect 187445 523566 187463 523600
rect 187221 523524 187463 523566
rect 172208 523490 172237 523524
rect 172271 523490 172329 523524
rect 172363 523490 172421 523524
rect 172455 523490 172513 523524
rect 172547 523490 172605 523524
rect 172639 523490 172697 523524
rect 172731 523490 172789 523524
rect 172823 523490 172881 523524
rect 172915 523490 172973 523524
rect 173007 523490 173065 523524
rect 173099 523490 173157 523524
rect 173191 523490 173249 523524
rect 173283 523490 173341 523524
rect 173375 523490 173433 523524
rect 173467 523490 173525 523524
rect 173559 523490 173617 523524
rect 173651 523490 173709 523524
rect 173743 523490 173801 523524
rect 173835 523490 173893 523524
rect 173927 523490 173985 523524
rect 174019 523490 174077 523524
rect 174111 523490 174169 523524
rect 174203 523490 174261 523524
rect 174295 523490 174353 523524
rect 174387 523490 174445 523524
rect 174479 523490 174537 523524
rect 174571 523490 174629 523524
rect 174663 523490 174721 523524
rect 174755 523490 174813 523524
rect 174847 523490 174905 523524
rect 174939 523490 174997 523524
rect 175031 523490 175089 523524
rect 175123 523490 175181 523524
rect 175215 523490 175273 523524
rect 175307 523490 175365 523524
rect 175399 523490 175457 523524
rect 175491 523490 175549 523524
rect 175583 523490 175641 523524
rect 175675 523490 175733 523524
rect 175767 523490 175825 523524
rect 175859 523490 175917 523524
rect 175951 523490 176009 523524
rect 176043 523490 176101 523524
rect 176135 523490 176193 523524
rect 176227 523490 176285 523524
rect 176319 523490 176377 523524
rect 176411 523490 176469 523524
rect 176503 523490 176561 523524
rect 176595 523490 176653 523524
rect 176687 523490 176745 523524
rect 176779 523490 176837 523524
rect 176871 523490 176929 523524
rect 176963 523490 177021 523524
rect 177055 523490 177113 523524
rect 177147 523490 177205 523524
rect 177239 523490 177297 523524
rect 177331 523490 177389 523524
rect 177423 523490 177481 523524
rect 177515 523490 177573 523524
rect 177607 523490 177665 523524
rect 177699 523490 177757 523524
rect 177791 523490 177849 523524
rect 177883 523490 177941 523524
rect 177975 523490 178033 523524
rect 178067 523490 178125 523524
rect 178159 523490 178217 523524
rect 178251 523490 178309 523524
rect 178343 523490 178401 523524
rect 178435 523490 178493 523524
rect 178527 523490 178585 523524
rect 178619 523490 178677 523524
rect 178711 523490 178769 523524
rect 178803 523490 178861 523524
rect 178895 523490 178953 523524
rect 178987 523490 179045 523524
rect 179079 523490 179137 523524
rect 179171 523490 179229 523524
rect 179263 523490 179321 523524
rect 179355 523490 179413 523524
rect 179447 523490 179505 523524
rect 179539 523490 179597 523524
rect 179631 523490 179689 523524
rect 179723 523490 179781 523524
rect 179815 523490 179873 523524
rect 179907 523490 179965 523524
rect 179999 523490 180057 523524
rect 180091 523490 180149 523524
rect 180183 523490 180241 523524
rect 180275 523490 180333 523524
rect 180367 523490 180425 523524
rect 180459 523490 180517 523524
rect 180551 523490 180609 523524
rect 180643 523490 180701 523524
rect 180735 523490 180793 523524
rect 180827 523490 180885 523524
rect 180919 523490 180977 523524
rect 181011 523490 181069 523524
rect 181103 523490 181161 523524
rect 181195 523490 181253 523524
rect 181287 523490 181345 523524
rect 181379 523490 181437 523524
rect 181471 523490 181529 523524
rect 181563 523490 181621 523524
rect 181655 523490 181713 523524
rect 181747 523490 181805 523524
rect 181839 523490 181897 523524
rect 181931 523490 181989 523524
rect 182023 523490 182081 523524
rect 182115 523490 182173 523524
rect 182207 523490 182265 523524
rect 182299 523490 182357 523524
rect 182391 523490 182449 523524
rect 182483 523490 182541 523524
rect 182575 523490 182633 523524
rect 182667 523490 182725 523524
rect 182759 523490 182817 523524
rect 182851 523490 182909 523524
rect 182943 523490 183001 523524
rect 183035 523490 183093 523524
rect 183127 523490 183185 523524
rect 183219 523490 183277 523524
rect 183311 523490 183369 523524
rect 183403 523490 183461 523524
rect 183495 523490 183553 523524
rect 183587 523490 183645 523524
rect 183679 523490 183737 523524
rect 183771 523490 183829 523524
rect 183863 523490 183921 523524
rect 183955 523490 184013 523524
rect 184047 523490 184105 523524
rect 184139 523490 184197 523524
rect 184231 523490 184289 523524
rect 184323 523490 184381 523524
rect 184415 523490 184473 523524
rect 184507 523490 184565 523524
rect 184599 523490 184657 523524
rect 184691 523490 184749 523524
rect 184783 523490 184841 523524
rect 184875 523490 184933 523524
rect 184967 523490 185025 523524
rect 185059 523490 185117 523524
rect 185151 523490 185209 523524
rect 185243 523490 185301 523524
rect 185335 523490 185393 523524
rect 185427 523490 185485 523524
rect 185519 523490 185577 523524
rect 185611 523490 185669 523524
rect 185703 523490 185761 523524
rect 185795 523490 185853 523524
rect 185887 523490 185945 523524
rect 185979 523490 186037 523524
rect 186071 523490 186129 523524
rect 186163 523490 186221 523524
rect 186255 523490 186313 523524
rect 186347 523490 186405 523524
rect 186439 523490 186497 523524
rect 186531 523490 186589 523524
rect 186623 523490 186681 523524
rect 186715 523490 186773 523524
rect 186807 523490 186865 523524
rect 186899 523490 186957 523524
rect 186991 523490 187049 523524
rect 187083 523490 187141 523524
rect 187175 523490 187233 523524
rect 187267 523490 187325 523524
rect 187359 523490 187417 523524
rect 187451 523490 187480 523524
rect 172225 523448 172467 523490
rect 172225 523414 172243 523448
rect 172277 523414 172415 523448
rect 172449 523414 172467 523448
rect 172225 523353 172467 523414
rect 172501 523448 173570 523490
rect 172501 523414 172519 523448
rect 172553 523414 173519 523448
rect 173553 523414 173570 523448
rect 172501 523403 173570 523414
rect 173605 523448 174674 523490
rect 173605 523414 173623 523448
rect 173657 523414 174623 523448
rect 174657 523414 174674 523448
rect 173605 523403 174674 523414
rect 174709 523448 175778 523490
rect 174709 523414 174727 523448
rect 174761 523414 175727 523448
rect 175761 523414 175778 523448
rect 174709 523403 175778 523414
rect 175813 523448 176882 523490
rect 175813 523414 175831 523448
rect 175865 523414 176831 523448
rect 176865 523414 176882 523448
rect 175813 523403 176882 523414
rect 176917 523448 177251 523490
rect 176917 523414 176935 523448
rect 176969 523414 177199 523448
rect 177233 523414 177251 523448
rect 172225 523319 172243 523353
rect 172277 523319 172415 523353
rect 172449 523319 172467 523353
rect 172225 523272 172467 523319
rect 172225 523204 172275 523238
rect 172309 523204 172329 523238
rect 172225 523130 172329 523204
rect 172363 523198 172467 523272
rect 172363 523164 172383 523198
rect 172417 523164 172467 523198
rect 172818 523238 172886 523255
rect 172818 523204 172835 523238
rect 172869 523204 172886 523238
rect 172225 523077 172467 523130
rect 172818 523089 172886 523204
rect 173182 523202 173252 523403
rect 173182 523168 173199 523202
rect 173233 523168 173252 523202
rect 173182 523153 173252 523168
rect 173922 523238 173990 523255
rect 173922 523204 173939 523238
rect 173973 523204 173990 523238
rect 173922 523089 173990 523204
rect 174286 523202 174356 523403
rect 174286 523168 174303 523202
rect 174337 523168 174356 523202
rect 174286 523153 174356 523168
rect 175026 523238 175094 523255
rect 175026 523204 175043 523238
rect 175077 523204 175094 523238
rect 175026 523089 175094 523204
rect 175390 523202 175460 523403
rect 175390 523168 175407 523202
rect 175441 523168 175460 523202
rect 175390 523153 175460 523168
rect 176130 523238 176198 523255
rect 176130 523204 176147 523238
rect 176181 523204 176198 523238
rect 176130 523089 176198 523204
rect 176494 523202 176564 523403
rect 176917 523346 177251 523414
rect 176917 523312 176935 523346
rect 176969 523312 177199 523346
rect 177233 523312 177251 523346
rect 176917 523272 177251 523312
rect 176494 523168 176511 523202
rect 176545 523168 176564 523202
rect 176494 523153 176564 523168
rect 176917 523204 176937 523238
rect 176971 523204 177067 523238
rect 176917 523134 177067 523204
rect 177101 523202 177251 523272
rect 177377 523419 177435 523490
rect 177377 523385 177389 523419
rect 177423 523385 177435 523419
rect 177469 523448 178538 523490
rect 177469 523414 177487 523448
rect 177521 523414 178487 523448
rect 178521 523414 178538 523448
rect 177469 523403 178538 523414
rect 178573 523448 179642 523490
rect 178573 523414 178591 523448
rect 178625 523414 179591 523448
rect 179625 523414 179642 523448
rect 178573 523403 179642 523414
rect 179677 523448 180746 523490
rect 179677 523414 179695 523448
rect 179729 523414 180695 523448
rect 180729 523414 180746 523448
rect 179677 523403 180746 523414
rect 180781 523448 181850 523490
rect 180781 523414 180799 523448
rect 180833 523414 181799 523448
rect 181833 523414 181850 523448
rect 180781 523403 181850 523414
rect 181885 523448 182403 523490
rect 181885 523414 181903 523448
rect 181937 523414 182351 523448
rect 182385 523414 182403 523448
rect 177377 523326 177435 523385
rect 177377 523292 177389 523326
rect 177423 523292 177435 523326
rect 177377 523257 177435 523292
rect 177101 523168 177197 523202
rect 177231 523168 177251 523202
rect 177786 523238 177854 523255
rect 177786 523204 177803 523238
rect 177837 523204 177854 523238
rect 172225 523043 172243 523077
rect 172277 523043 172415 523077
rect 172449 523043 172467 523077
rect 172225 522980 172467 523043
rect 172501 523075 173570 523089
rect 172501 523041 172519 523075
rect 172553 523041 173519 523075
rect 173553 523041 173570 523075
rect 172501 522980 173570 523041
rect 173605 523075 174674 523089
rect 173605 523041 173623 523075
rect 173657 523041 174623 523075
rect 174657 523041 174674 523075
rect 173605 522980 174674 523041
rect 174709 523075 175778 523089
rect 174709 523041 174727 523075
rect 174761 523041 175727 523075
rect 175761 523041 175778 523075
rect 174709 522980 175778 523041
rect 175813 523075 176882 523089
rect 175813 523041 175831 523075
rect 175865 523041 176831 523075
rect 176865 523041 176882 523075
rect 175813 522980 176882 523041
rect 176917 523082 177251 523134
rect 176917 523048 176935 523082
rect 176969 523048 177199 523082
rect 177233 523048 177251 523082
rect 176917 522980 177251 523048
rect 177377 523108 177435 523125
rect 177377 523074 177389 523108
rect 177423 523074 177435 523108
rect 177786 523089 177854 523204
rect 178150 523202 178220 523403
rect 178150 523168 178167 523202
rect 178201 523168 178220 523202
rect 178150 523153 178220 523168
rect 178890 523238 178958 523255
rect 178890 523204 178907 523238
rect 178941 523204 178958 523238
rect 178890 523089 178958 523204
rect 179254 523202 179324 523403
rect 179254 523168 179271 523202
rect 179305 523168 179324 523202
rect 179254 523153 179324 523168
rect 179994 523238 180062 523255
rect 179994 523204 180011 523238
rect 180045 523204 180062 523238
rect 179994 523089 180062 523204
rect 180358 523202 180428 523403
rect 180358 523168 180375 523202
rect 180409 523168 180428 523202
rect 180358 523153 180428 523168
rect 181098 523238 181166 523255
rect 181098 523204 181115 523238
rect 181149 523204 181166 523238
rect 181098 523089 181166 523204
rect 181462 523202 181532 523403
rect 181885 523346 182403 523414
rect 181885 523312 181903 523346
rect 181937 523312 182351 523346
rect 182385 523312 182403 523346
rect 181885 523272 182403 523312
rect 181462 523168 181479 523202
rect 181513 523168 181532 523202
rect 181462 523153 181532 523168
rect 181885 523204 181963 523238
rect 181997 523204 182073 523238
rect 182107 523204 182127 523238
rect 181885 523134 182127 523204
rect 182161 523202 182403 523272
rect 182529 523419 182587 523490
rect 182529 523385 182541 523419
rect 182575 523385 182587 523419
rect 182621 523448 183690 523490
rect 182621 523414 182639 523448
rect 182673 523414 183639 523448
rect 183673 523414 183690 523448
rect 182621 523403 183690 523414
rect 183725 523448 184794 523490
rect 183725 523414 183743 523448
rect 183777 523414 184743 523448
rect 184777 523414 184794 523448
rect 183725 523403 184794 523414
rect 184829 523448 185898 523490
rect 184829 523414 184847 523448
rect 184881 523414 185847 523448
rect 185881 523414 185898 523448
rect 184829 523403 185898 523414
rect 185933 523448 187002 523490
rect 185933 523414 185951 523448
rect 185985 523414 186951 523448
rect 186985 523414 187002 523448
rect 185933 523403 187002 523414
rect 187221 523448 187463 523490
rect 187221 523414 187239 523448
rect 187273 523414 187411 523448
rect 187445 523414 187463 523448
rect 182529 523326 182587 523385
rect 182529 523292 182541 523326
rect 182575 523292 182587 523326
rect 182529 523257 182587 523292
rect 182161 523168 182181 523202
rect 182215 523168 182291 523202
rect 182325 523168 182403 523202
rect 182938 523238 183006 523255
rect 182938 523204 182955 523238
rect 182989 523204 183006 523238
rect 177377 522980 177435 523074
rect 177469 523075 178538 523089
rect 177469 523041 177487 523075
rect 177521 523041 178487 523075
rect 178521 523041 178538 523075
rect 177469 522980 178538 523041
rect 178573 523075 179642 523089
rect 178573 523041 178591 523075
rect 178625 523041 179591 523075
rect 179625 523041 179642 523075
rect 178573 522980 179642 523041
rect 179677 523075 180746 523089
rect 179677 523041 179695 523075
rect 179729 523041 180695 523075
rect 180729 523041 180746 523075
rect 179677 522980 180746 523041
rect 180781 523075 181850 523089
rect 180781 523041 180799 523075
rect 180833 523041 181799 523075
rect 181833 523041 181850 523075
rect 180781 522980 181850 523041
rect 181885 523075 182403 523134
rect 181885 523041 181903 523075
rect 181937 523041 182351 523075
rect 182385 523041 182403 523075
rect 181885 522980 182403 523041
rect 182529 523108 182587 523125
rect 182529 523074 182541 523108
rect 182575 523074 182587 523108
rect 182938 523089 183006 523204
rect 183302 523202 183372 523403
rect 183302 523168 183319 523202
rect 183353 523168 183372 523202
rect 183302 523153 183372 523168
rect 184042 523238 184110 523255
rect 184042 523204 184059 523238
rect 184093 523204 184110 523238
rect 184042 523089 184110 523204
rect 184406 523202 184476 523403
rect 184406 523168 184423 523202
rect 184457 523168 184476 523202
rect 184406 523153 184476 523168
rect 185146 523238 185214 523255
rect 185146 523204 185163 523238
rect 185197 523204 185214 523238
rect 185146 523089 185214 523204
rect 185510 523202 185580 523403
rect 185510 523168 185527 523202
rect 185561 523168 185580 523202
rect 185510 523153 185580 523168
rect 186250 523238 186318 523255
rect 186250 523204 186267 523238
rect 186301 523204 186318 523238
rect 186250 523089 186318 523204
rect 186614 523202 186684 523403
rect 186614 523168 186631 523202
rect 186665 523168 186684 523202
rect 186614 523153 186684 523168
rect 187221 523353 187463 523414
rect 187221 523319 187239 523353
rect 187273 523319 187411 523353
rect 187445 523319 187463 523353
rect 187221 523272 187463 523319
rect 187221 523198 187325 523272
rect 187221 523164 187271 523198
rect 187305 523164 187325 523198
rect 187359 523204 187379 523238
rect 187413 523204 187463 523238
rect 187359 523130 187463 523204
rect 182529 522980 182587 523074
rect 182621 523075 183690 523089
rect 182621 523041 182639 523075
rect 182673 523041 183639 523075
rect 183673 523041 183690 523075
rect 182621 522980 183690 523041
rect 183725 523075 184794 523089
rect 183725 523041 183743 523075
rect 183777 523041 184743 523075
rect 184777 523041 184794 523075
rect 183725 522980 184794 523041
rect 184829 523075 185898 523089
rect 184829 523041 184847 523075
rect 184881 523041 185847 523075
rect 185881 523041 185898 523075
rect 184829 522980 185898 523041
rect 185933 523075 187002 523089
rect 185933 523041 185951 523075
rect 185985 523041 186951 523075
rect 186985 523041 187002 523075
rect 185933 522980 187002 523041
rect 187221 523077 187463 523130
rect 187221 523043 187239 523077
rect 187273 523043 187411 523077
rect 187445 523043 187463 523077
rect 187221 522980 187463 523043
rect 172208 522946 172237 522980
rect 172271 522946 172329 522980
rect 172363 522946 172421 522980
rect 172455 522946 172513 522980
rect 172547 522946 172605 522980
rect 172639 522946 172697 522980
rect 172731 522946 172789 522980
rect 172823 522946 172881 522980
rect 172915 522946 172973 522980
rect 173007 522946 173065 522980
rect 173099 522946 173157 522980
rect 173191 522946 173249 522980
rect 173283 522946 173341 522980
rect 173375 522946 173433 522980
rect 173467 522946 173525 522980
rect 173559 522946 173617 522980
rect 173651 522946 173709 522980
rect 173743 522946 173801 522980
rect 173835 522946 173893 522980
rect 173927 522946 173985 522980
rect 174019 522946 174077 522980
rect 174111 522946 174169 522980
rect 174203 522946 174261 522980
rect 174295 522946 174353 522980
rect 174387 522946 174445 522980
rect 174479 522946 174537 522980
rect 174571 522946 174629 522980
rect 174663 522946 174721 522980
rect 174755 522946 174813 522980
rect 174847 522946 174905 522980
rect 174939 522946 174997 522980
rect 175031 522946 175089 522980
rect 175123 522946 175181 522980
rect 175215 522946 175273 522980
rect 175307 522946 175365 522980
rect 175399 522946 175457 522980
rect 175491 522946 175549 522980
rect 175583 522946 175641 522980
rect 175675 522946 175733 522980
rect 175767 522946 175825 522980
rect 175859 522946 175917 522980
rect 175951 522946 176009 522980
rect 176043 522946 176101 522980
rect 176135 522946 176193 522980
rect 176227 522946 176285 522980
rect 176319 522946 176377 522980
rect 176411 522946 176469 522980
rect 176503 522946 176561 522980
rect 176595 522946 176653 522980
rect 176687 522946 176745 522980
rect 176779 522946 176837 522980
rect 176871 522946 176929 522980
rect 176963 522946 177021 522980
rect 177055 522946 177113 522980
rect 177147 522946 177205 522980
rect 177239 522946 177297 522980
rect 177331 522946 177389 522980
rect 177423 522946 177481 522980
rect 177515 522946 177573 522980
rect 177607 522946 177665 522980
rect 177699 522946 177757 522980
rect 177791 522946 177849 522980
rect 177883 522946 177941 522980
rect 177975 522946 178033 522980
rect 178067 522946 178125 522980
rect 178159 522946 178217 522980
rect 178251 522946 178309 522980
rect 178343 522946 178401 522980
rect 178435 522946 178493 522980
rect 178527 522946 178585 522980
rect 178619 522946 178677 522980
rect 178711 522946 178769 522980
rect 178803 522946 178861 522980
rect 178895 522946 178953 522980
rect 178987 522946 179045 522980
rect 179079 522946 179137 522980
rect 179171 522946 179229 522980
rect 179263 522946 179321 522980
rect 179355 522946 179413 522980
rect 179447 522946 179505 522980
rect 179539 522946 179597 522980
rect 179631 522946 179689 522980
rect 179723 522946 179781 522980
rect 179815 522946 179873 522980
rect 179907 522946 179965 522980
rect 179999 522946 180057 522980
rect 180091 522946 180149 522980
rect 180183 522946 180241 522980
rect 180275 522946 180333 522980
rect 180367 522946 180425 522980
rect 180459 522946 180517 522980
rect 180551 522946 180609 522980
rect 180643 522946 180701 522980
rect 180735 522946 180793 522980
rect 180827 522946 180885 522980
rect 180919 522946 180977 522980
rect 181011 522946 181069 522980
rect 181103 522946 181161 522980
rect 181195 522946 181253 522980
rect 181287 522946 181345 522980
rect 181379 522946 181437 522980
rect 181471 522946 181529 522980
rect 181563 522946 181621 522980
rect 181655 522946 181713 522980
rect 181747 522946 181805 522980
rect 181839 522946 181897 522980
rect 181931 522946 181989 522980
rect 182023 522946 182081 522980
rect 182115 522946 182173 522980
rect 182207 522946 182265 522980
rect 182299 522946 182357 522980
rect 182391 522946 182449 522980
rect 182483 522946 182541 522980
rect 182575 522946 182633 522980
rect 182667 522946 182725 522980
rect 182759 522946 182817 522980
rect 182851 522946 182909 522980
rect 182943 522946 183001 522980
rect 183035 522946 183093 522980
rect 183127 522946 183185 522980
rect 183219 522946 183277 522980
rect 183311 522946 183369 522980
rect 183403 522946 183461 522980
rect 183495 522946 183553 522980
rect 183587 522946 183645 522980
rect 183679 522946 183737 522980
rect 183771 522946 183829 522980
rect 183863 522946 183921 522980
rect 183955 522946 184013 522980
rect 184047 522946 184105 522980
rect 184139 522946 184197 522980
rect 184231 522946 184289 522980
rect 184323 522946 184381 522980
rect 184415 522946 184473 522980
rect 184507 522946 184565 522980
rect 184599 522946 184657 522980
rect 184691 522946 184749 522980
rect 184783 522946 184841 522980
rect 184875 522946 184933 522980
rect 184967 522946 185025 522980
rect 185059 522946 185117 522980
rect 185151 522946 185209 522980
rect 185243 522946 185301 522980
rect 185335 522946 185393 522980
rect 185427 522946 185485 522980
rect 185519 522946 185577 522980
rect 185611 522946 185669 522980
rect 185703 522946 185761 522980
rect 185795 522946 185853 522980
rect 185887 522946 185945 522980
rect 185979 522946 186037 522980
rect 186071 522946 186129 522980
rect 186163 522946 186221 522980
rect 186255 522946 186313 522980
rect 186347 522946 186405 522980
rect 186439 522946 186497 522980
rect 186531 522946 186589 522980
rect 186623 522946 186681 522980
rect 186715 522946 186773 522980
rect 186807 522946 186865 522980
rect 186899 522946 186957 522980
rect 186991 522946 187049 522980
rect 187083 522946 187141 522980
rect 187175 522946 187233 522980
rect 187267 522946 187325 522980
rect 187359 522946 187417 522980
rect 187451 522946 187480 522980
rect 172225 522883 172467 522946
rect 172225 522849 172243 522883
rect 172277 522849 172415 522883
rect 172449 522849 172467 522883
rect 172225 522796 172467 522849
rect 172501 522885 173570 522946
rect 172501 522851 172519 522885
rect 172553 522851 173519 522885
rect 173553 522851 173570 522885
rect 172501 522837 173570 522851
rect 173605 522885 174674 522946
rect 173605 522851 173623 522885
rect 173657 522851 174623 522885
rect 174657 522851 174674 522885
rect 173605 522837 174674 522851
rect 174801 522852 174859 522946
rect 172225 522722 172329 522796
rect 172225 522688 172275 522722
rect 172309 522688 172329 522722
rect 172363 522728 172383 522762
rect 172417 522728 172467 522762
rect 172363 522654 172467 522728
rect 172818 522722 172886 522837
rect 172818 522688 172835 522722
rect 172869 522688 172886 522722
rect 172818 522671 172886 522688
rect 173182 522758 173252 522773
rect 173182 522724 173199 522758
rect 173233 522724 173252 522758
rect 172225 522607 172467 522654
rect 172225 522573 172243 522607
rect 172277 522573 172415 522607
rect 172449 522573 172467 522607
rect 172225 522512 172467 522573
rect 173182 522523 173252 522724
rect 173922 522722 173990 522837
rect 174801 522818 174813 522852
rect 174847 522818 174859 522852
rect 174893 522885 175962 522946
rect 174893 522851 174911 522885
rect 174945 522851 175911 522885
rect 175945 522851 175962 522885
rect 174893 522837 175962 522851
rect 175997 522885 177066 522946
rect 175997 522851 176015 522885
rect 176049 522851 177015 522885
rect 177049 522851 177066 522885
rect 175997 522837 177066 522851
rect 177101 522885 178170 522946
rect 177101 522851 177119 522885
rect 177153 522851 178119 522885
rect 178153 522851 178170 522885
rect 177101 522837 178170 522851
rect 178205 522885 179274 522946
rect 178205 522851 178223 522885
rect 178257 522851 179223 522885
rect 179257 522851 179274 522885
rect 178205 522837 179274 522851
rect 179309 522885 179827 522946
rect 179309 522851 179327 522885
rect 179361 522851 179775 522885
rect 179809 522851 179827 522885
rect 174801 522801 174859 522818
rect 173922 522688 173939 522722
rect 173973 522688 173990 522722
rect 173922 522671 173990 522688
rect 174286 522758 174356 522773
rect 174286 522724 174303 522758
rect 174337 522724 174356 522758
rect 174286 522523 174356 522724
rect 175210 522722 175278 522837
rect 175210 522688 175227 522722
rect 175261 522688 175278 522722
rect 175210 522671 175278 522688
rect 175574 522758 175644 522773
rect 175574 522724 175591 522758
rect 175625 522724 175644 522758
rect 174801 522634 174859 522669
rect 174801 522600 174813 522634
rect 174847 522600 174859 522634
rect 174801 522541 174859 522600
rect 172225 522478 172243 522512
rect 172277 522478 172415 522512
rect 172449 522478 172467 522512
rect 172225 522436 172467 522478
rect 172501 522512 173570 522523
rect 172501 522478 172519 522512
rect 172553 522478 173519 522512
rect 173553 522478 173570 522512
rect 172501 522436 173570 522478
rect 173605 522512 174674 522523
rect 173605 522478 173623 522512
rect 173657 522478 174623 522512
rect 174657 522478 174674 522512
rect 173605 522436 174674 522478
rect 174801 522507 174813 522541
rect 174847 522507 174859 522541
rect 175574 522523 175644 522724
rect 176314 522722 176382 522837
rect 176314 522688 176331 522722
rect 176365 522688 176382 522722
rect 176314 522671 176382 522688
rect 176678 522758 176748 522773
rect 176678 522724 176695 522758
rect 176729 522724 176748 522758
rect 176678 522523 176748 522724
rect 177418 522722 177486 522837
rect 177418 522688 177435 522722
rect 177469 522688 177486 522722
rect 177418 522671 177486 522688
rect 177782 522758 177852 522773
rect 177782 522724 177799 522758
rect 177833 522724 177852 522758
rect 177782 522523 177852 522724
rect 178522 522722 178590 522837
rect 179309 522792 179827 522851
rect 179953 522852 180011 522946
rect 179953 522818 179965 522852
rect 179999 522818 180011 522852
rect 180045 522885 181114 522946
rect 180045 522851 180063 522885
rect 180097 522851 181063 522885
rect 181097 522851 181114 522885
rect 180045 522837 181114 522851
rect 181149 522885 182218 522946
rect 181149 522851 181167 522885
rect 181201 522851 182167 522885
rect 182201 522851 182218 522885
rect 181149 522837 182218 522851
rect 182253 522885 183322 522946
rect 182253 522851 182271 522885
rect 182305 522851 183271 522885
rect 183305 522851 183322 522885
rect 182253 522837 183322 522851
rect 183357 522885 184426 522946
rect 183357 522851 183375 522885
rect 183409 522851 184375 522885
rect 184409 522851 184426 522885
rect 183357 522837 184426 522851
rect 184461 522885 184979 522946
rect 184461 522851 184479 522885
rect 184513 522851 184927 522885
rect 184961 522851 184979 522885
rect 179953 522801 180011 522818
rect 178522 522688 178539 522722
rect 178573 522688 178590 522722
rect 178522 522671 178590 522688
rect 178886 522758 178956 522773
rect 178886 522724 178903 522758
rect 178937 522724 178956 522758
rect 178886 522523 178956 522724
rect 179309 522722 179551 522792
rect 179309 522688 179387 522722
rect 179421 522688 179497 522722
rect 179531 522688 179551 522722
rect 179585 522724 179605 522758
rect 179639 522724 179715 522758
rect 179749 522724 179827 522758
rect 179585 522654 179827 522724
rect 180362 522722 180430 522837
rect 180362 522688 180379 522722
rect 180413 522688 180430 522722
rect 180362 522671 180430 522688
rect 180726 522758 180796 522773
rect 180726 522724 180743 522758
rect 180777 522724 180796 522758
rect 179309 522614 179827 522654
rect 179309 522580 179327 522614
rect 179361 522580 179775 522614
rect 179809 522580 179827 522614
rect 174801 522436 174859 522507
rect 174893 522512 175962 522523
rect 174893 522478 174911 522512
rect 174945 522478 175911 522512
rect 175945 522478 175962 522512
rect 174893 522436 175962 522478
rect 175997 522512 177066 522523
rect 175997 522478 176015 522512
rect 176049 522478 177015 522512
rect 177049 522478 177066 522512
rect 175997 522436 177066 522478
rect 177101 522512 178170 522523
rect 177101 522478 177119 522512
rect 177153 522478 178119 522512
rect 178153 522478 178170 522512
rect 177101 522436 178170 522478
rect 178205 522512 179274 522523
rect 178205 522478 178223 522512
rect 178257 522478 179223 522512
rect 179257 522478 179274 522512
rect 178205 522436 179274 522478
rect 179309 522512 179827 522580
rect 179309 522478 179327 522512
rect 179361 522478 179775 522512
rect 179809 522478 179827 522512
rect 179309 522436 179827 522478
rect 179953 522634 180011 522669
rect 179953 522600 179965 522634
rect 179999 522600 180011 522634
rect 179953 522541 180011 522600
rect 179953 522507 179965 522541
rect 179999 522507 180011 522541
rect 180726 522523 180796 522724
rect 181466 522722 181534 522837
rect 181466 522688 181483 522722
rect 181517 522688 181534 522722
rect 181466 522671 181534 522688
rect 181830 522758 181900 522773
rect 181830 522724 181847 522758
rect 181881 522724 181900 522758
rect 181830 522523 181900 522724
rect 182570 522722 182638 522837
rect 182570 522688 182587 522722
rect 182621 522688 182638 522722
rect 182570 522671 182638 522688
rect 182934 522758 183004 522773
rect 182934 522724 182951 522758
rect 182985 522724 183004 522758
rect 182934 522523 183004 522724
rect 183674 522722 183742 522837
rect 184461 522792 184979 522851
rect 185105 522852 185163 522946
rect 185105 522818 185117 522852
rect 185151 522818 185163 522852
rect 185197 522885 186266 522946
rect 185197 522851 185215 522885
rect 185249 522851 186215 522885
rect 186249 522851 186266 522885
rect 185197 522837 186266 522851
rect 186301 522885 187003 522946
rect 186301 522851 186319 522885
rect 186353 522851 186951 522885
rect 186985 522851 187003 522885
rect 185105 522801 185163 522818
rect 183674 522688 183691 522722
rect 183725 522688 183742 522722
rect 183674 522671 183742 522688
rect 184038 522758 184108 522773
rect 184038 522724 184055 522758
rect 184089 522724 184108 522758
rect 184038 522523 184108 522724
rect 184461 522722 184703 522792
rect 184461 522688 184539 522722
rect 184573 522688 184649 522722
rect 184683 522688 184703 522722
rect 184737 522724 184757 522758
rect 184791 522724 184867 522758
rect 184901 522724 184979 522758
rect 184737 522654 184979 522724
rect 185514 522722 185582 522837
rect 186301 522792 187003 522851
rect 187221 522883 187463 522946
rect 187221 522849 187239 522883
rect 187273 522849 187411 522883
rect 187445 522849 187463 522883
rect 187221 522796 187463 522849
rect 185514 522688 185531 522722
rect 185565 522688 185582 522722
rect 185514 522671 185582 522688
rect 185878 522758 185948 522773
rect 185878 522724 185895 522758
rect 185929 522724 185948 522758
rect 184461 522614 184979 522654
rect 184461 522580 184479 522614
rect 184513 522580 184927 522614
rect 184961 522580 184979 522614
rect 179953 522436 180011 522507
rect 180045 522512 181114 522523
rect 180045 522478 180063 522512
rect 180097 522478 181063 522512
rect 181097 522478 181114 522512
rect 180045 522436 181114 522478
rect 181149 522512 182218 522523
rect 181149 522478 181167 522512
rect 181201 522478 182167 522512
rect 182201 522478 182218 522512
rect 181149 522436 182218 522478
rect 182253 522512 183322 522523
rect 182253 522478 182271 522512
rect 182305 522478 183271 522512
rect 183305 522478 183322 522512
rect 182253 522436 183322 522478
rect 183357 522512 184426 522523
rect 183357 522478 183375 522512
rect 183409 522478 184375 522512
rect 184409 522478 184426 522512
rect 183357 522436 184426 522478
rect 184461 522512 184979 522580
rect 184461 522478 184479 522512
rect 184513 522478 184927 522512
rect 184961 522478 184979 522512
rect 184461 522436 184979 522478
rect 185105 522634 185163 522669
rect 185105 522600 185117 522634
rect 185151 522600 185163 522634
rect 185105 522541 185163 522600
rect 185105 522507 185117 522541
rect 185151 522507 185163 522541
rect 185878 522523 185948 522724
rect 186301 522722 186631 522792
rect 186301 522688 186379 522722
rect 186413 522688 186478 522722
rect 186512 522688 186577 522722
rect 186611 522688 186631 522722
rect 186665 522724 186685 522758
rect 186719 522724 186788 522758
rect 186822 522724 186891 522758
rect 186925 522724 187003 522758
rect 186665 522654 187003 522724
rect 186301 522614 187003 522654
rect 186301 522580 186319 522614
rect 186353 522580 186951 522614
rect 186985 522580 187003 522614
rect 185105 522436 185163 522507
rect 185197 522512 186266 522523
rect 185197 522478 185215 522512
rect 185249 522478 186215 522512
rect 186249 522478 186266 522512
rect 185197 522436 186266 522478
rect 186301 522512 187003 522580
rect 186301 522478 186319 522512
rect 186353 522478 186951 522512
rect 186985 522478 187003 522512
rect 186301 522436 187003 522478
rect 187221 522728 187271 522762
rect 187305 522728 187325 522762
rect 187221 522654 187325 522728
rect 187359 522722 187463 522796
rect 187359 522688 187379 522722
rect 187413 522688 187463 522722
rect 187221 522607 187463 522654
rect 187221 522573 187239 522607
rect 187273 522573 187411 522607
rect 187445 522573 187463 522607
rect 187221 522512 187463 522573
rect 187221 522478 187239 522512
rect 187273 522478 187411 522512
rect 187445 522478 187463 522512
rect 187221 522436 187463 522478
rect 172208 522402 172237 522436
rect 172271 522402 172329 522436
rect 172363 522402 172421 522436
rect 172455 522402 172513 522436
rect 172547 522402 172605 522436
rect 172639 522402 172697 522436
rect 172731 522402 172789 522436
rect 172823 522402 172881 522436
rect 172915 522402 172973 522436
rect 173007 522402 173065 522436
rect 173099 522402 173157 522436
rect 173191 522402 173249 522436
rect 173283 522402 173341 522436
rect 173375 522402 173433 522436
rect 173467 522402 173525 522436
rect 173559 522402 173617 522436
rect 173651 522402 173709 522436
rect 173743 522402 173801 522436
rect 173835 522402 173893 522436
rect 173927 522402 173985 522436
rect 174019 522402 174077 522436
rect 174111 522402 174169 522436
rect 174203 522402 174261 522436
rect 174295 522402 174353 522436
rect 174387 522402 174445 522436
rect 174479 522402 174537 522436
rect 174571 522402 174629 522436
rect 174663 522402 174721 522436
rect 174755 522402 174813 522436
rect 174847 522402 174905 522436
rect 174939 522402 174997 522436
rect 175031 522402 175089 522436
rect 175123 522402 175181 522436
rect 175215 522402 175273 522436
rect 175307 522402 175365 522436
rect 175399 522402 175457 522436
rect 175491 522402 175549 522436
rect 175583 522402 175641 522436
rect 175675 522402 175733 522436
rect 175767 522402 175825 522436
rect 175859 522402 175917 522436
rect 175951 522402 176009 522436
rect 176043 522402 176101 522436
rect 176135 522402 176193 522436
rect 176227 522402 176285 522436
rect 176319 522402 176377 522436
rect 176411 522402 176469 522436
rect 176503 522402 176561 522436
rect 176595 522402 176653 522436
rect 176687 522402 176745 522436
rect 176779 522402 176837 522436
rect 176871 522402 176929 522436
rect 176963 522402 177021 522436
rect 177055 522402 177113 522436
rect 177147 522402 177205 522436
rect 177239 522402 177297 522436
rect 177331 522402 177389 522436
rect 177423 522402 177481 522436
rect 177515 522402 177573 522436
rect 177607 522402 177665 522436
rect 177699 522402 177757 522436
rect 177791 522402 177849 522436
rect 177883 522402 177941 522436
rect 177975 522402 178033 522436
rect 178067 522402 178125 522436
rect 178159 522402 178217 522436
rect 178251 522402 178309 522436
rect 178343 522402 178401 522436
rect 178435 522402 178493 522436
rect 178527 522402 178585 522436
rect 178619 522402 178677 522436
rect 178711 522402 178769 522436
rect 178803 522402 178861 522436
rect 178895 522402 178953 522436
rect 178987 522402 179045 522436
rect 179079 522402 179137 522436
rect 179171 522402 179229 522436
rect 179263 522402 179321 522436
rect 179355 522402 179413 522436
rect 179447 522402 179505 522436
rect 179539 522402 179597 522436
rect 179631 522402 179689 522436
rect 179723 522402 179781 522436
rect 179815 522402 179873 522436
rect 179907 522402 179965 522436
rect 179999 522402 180057 522436
rect 180091 522402 180149 522436
rect 180183 522402 180241 522436
rect 180275 522402 180333 522436
rect 180367 522402 180425 522436
rect 180459 522402 180517 522436
rect 180551 522402 180609 522436
rect 180643 522402 180701 522436
rect 180735 522402 180793 522436
rect 180827 522402 180885 522436
rect 180919 522402 180977 522436
rect 181011 522402 181069 522436
rect 181103 522402 181161 522436
rect 181195 522402 181253 522436
rect 181287 522402 181345 522436
rect 181379 522402 181437 522436
rect 181471 522402 181529 522436
rect 181563 522402 181621 522436
rect 181655 522402 181713 522436
rect 181747 522402 181805 522436
rect 181839 522402 181897 522436
rect 181931 522402 181989 522436
rect 182023 522402 182081 522436
rect 182115 522402 182173 522436
rect 182207 522402 182265 522436
rect 182299 522402 182357 522436
rect 182391 522402 182449 522436
rect 182483 522402 182541 522436
rect 182575 522402 182633 522436
rect 182667 522402 182725 522436
rect 182759 522402 182817 522436
rect 182851 522402 182909 522436
rect 182943 522402 183001 522436
rect 183035 522402 183093 522436
rect 183127 522402 183185 522436
rect 183219 522402 183277 522436
rect 183311 522402 183369 522436
rect 183403 522402 183461 522436
rect 183495 522402 183553 522436
rect 183587 522402 183645 522436
rect 183679 522402 183737 522436
rect 183771 522402 183829 522436
rect 183863 522402 183921 522436
rect 183955 522402 184013 522436
rect 184047 522402 184105 522436
rect 184139 522402 184197 522436
rect 184231 522402 184289 522436
rect 184323 522402 184381 522436
rect 184415 522402 184473 522436
rect 184507 522402 184565 522436
rect 184599 522402 184657 522436
rect 184691 522402 184749 522436
rect 184783 522402 184841 522436
rect 184875 522402 184933 522436
rect 184967 522402 185025 522436
rect 185059 522402 185117 522436
rect 185151 522402 185209 522436
rect 185243 522402 185301 522436
rect 185335 522402 185393 522436
rect 185427 522402 185485 522436
rect 185519 522402 185577 522436
rect 185611 522402 185669 522436
rect 185703 522402 185761 522436
rect 185795 522402 185853 522436
rect 185887 522402 185945 522436
rect 185979 522402 186037 522436
rect 186071 522402 186129 522436
rect 186163 522402 186221 522436
rect 186255 522402 186313 522436
rect 186347 522402 186405 522436
rect 186439 522402 186497 522436
rect 186531 522402 186589 522436
rect 186623 522402 186681 522436
rect 186715 522402 186773 522436
rect 186807 522402 186865 522436
rect 186899 522402 186957 522436
rect 186991 522402 187049 522436
rect 187083 522402 187141 522436
rect 187175 522402 187233 522436
rect 187267 522402 187325 522436
rect 187359 522402 187417 522436
rect 187451 522402 187480 522436
rect 172225 522360 172467 522402
rect 172225 522326 172243 522360
rect 172277 522326 172415 522360
rect 172449 522326 172467 522360
rect 172225 522265 172467 522326
rect 172501 522360 173570 522402
rect 172501 522326 172519 522360
rect 172553 522326 173519 522360
rect 173553 522326 173570 522360
rect 172501 522315 173570 522326
rect 173605 522360 174674 522402
rect 173605 522326 173623 522360
rect 173657 522326 174623 522360
rect 174657 522326 174674 522360
rect 173605 522315 174674 522326
rect 174709 522360 175778 522402
rect 174709 522326 174727 522360
rect 174761 522326 175727 522360
rect 175761 522326 175778 522360
rect 174709 522315 175778 522326
rect 175813 522360 176882 522402
rect 175813 522326 175831 522360
rect 175865 522326 176831 522360
rect 176865 522326 176882 522360
rect 175813 522315 176882 522326
rect 176917 522360 177251 522402
rect 176917 522326 176935 522360
rect 176969 522326 177199 522360
rect 177233 522326 177251 522360
rect 172225 522231 172243 522265
rect 172277 522231 172415 522265
rect 172449 522231 172467 522265
rect 172225 522184 172467 522231
rect 172225 522116 172275 522150
rect 172309 522116 172329 522150
rect 172225 522042 172329 522116
rect 172363 522110 172467 522184
rect 172363 522076 172383 522110
rect 172417 522076 172467 522110
rect 172818 522150 172886 522167
rect 172818 522116 172835 522150
rect 172869 522116 172886 522150
rect 172225 521989 172467 522042
rect 172818 522001 172886 522116
rect 173182 522114 173252 522315
rect 173182 522080 173199 522114
rect 173233 522080 173252 522114
rect 173182 522065 173252 522080
rect 173922 522150 173990 522167
rect 173922 522116 173939 522150
rect 173973 522116 173990 522150
rect 173922 522001 173990 522116
rect 174286 522114 174356 522315
rect 174286 522080 174303 522114
rect 174337 522080 174356 522114
rect 174286 522065 174356 522080
rect 175026 522150 175094 522167
rect 175026 522116 175043 522150
rect 175077 522116 175094 522150
rect 175026 522001 175094 522116
rect 175390 522114 175460 522315
rect 175390 522080 175407 522114
rect 175441 522080 175460 522114
rect 175390 522065 175460 522080
rect 176130 522150 176198 522167
rect 176130 522116 176147 522150
rect 176181 522116 176198 522150
rect 176130 522001 176198 522116
rect 176494 522114 176564 522315
rect 176917 522258 177251 522326
rect 176917 522224 176935 522258
rect 176969 522224 177199 522258
rect 177233 522224 177251 522258
rect 176917 522184 177251 522224
rect 176494 522080 176511 522114
rect 176545 522080 176564 522114
rect 176494 522065 176564 522080
rect 176917 522116 176937 522150
rect 176971 522116 177067 522150
rect 176917 522046 177067 522116
rect 177101 522114 177251 522184
rect 177377 522331 177435 522402
rect 177377 522297 177389 522331
rect 177423 522297 177435 522331
rect 177469 522360 178538 522402
rect 177469 522326 177487 522360
rect 177521 522326 178487 522360
rect 178521 522326 178538 522360
rect 177469 522315 178538 522326
rect 178573 522360 179642 522402
rect 178573 522326 178591 522360
rect 178625 522326 179591 522360
rect 179625 522326 179642 522360
rect 178573 522315 179642 522326
rect 179677 522360 180746 522402
rect 179677 522326 179695 522360
rect 179729 522326 180695 522360
rect 180729 522326 180746 522360
rect 179677 522315 180746 522326
rect 180781 522360 181850 522402
rect 180781 522326 180799 522360
rect 180833 522326 181799 522360
rect 181833 522326 181850 522360
rect 180781 522315 181850 522326
rect 181885 522360 182403 522402
rect 181885 522326 181903 522360
rect 181937 522326 182351 522360
rect 182385 522326 182403 522360
rect 177377 522238 177435 522297
rect 177377 522204 177389 522238
rect 177423 522204 177435 522238
rect 177377 522169 177435 522204
rect 177101 522080 177197 522114
rect 177231 522080 177251 522114
rect 177786 522150 177854 522167
rect 177786 522116 177803 522150
rect 177837 522116 177854 522150
rect 172225 521955 172243 521989
rect 172277 521955 172415 521989
rect 172449 521955 172467 521989
rect 172225 521892 172467 521955
rect 172501 521987 173570 522001
rect 172501 521953 172519 521987
rect 172553 521953 173519 521987
rect 173553 521953 173570 521987
rect 172501 521892 173570 521953
rect 173605 521987 174674 522001
rect 173605 521953 173623 521987
rect 173657 521953 174623 521987
rect 174657 521953 174674 521987
rect 173605 521892 174674 521953
rect 174709 521987 175778 522001
rect 174709 521953 174727 521987
rect 174761 521953 175727 521987
rect 175761 521953 175778 521987
rect 174709 521892 175778 521953
rect 175813 521987 176882 522001
rect 175813 521953 175831 521987
rect 175865 521953 176831 521987
rect 176865 521953 176882 521987
rect 175813 521892 176882 521953
rect 176917 521994 177251 522046
rect 176917 521960 176935 521994
rect 176969 521960 177199 521994
rect 177233 521960 177251 521994
rect 176917 521892 177251 521960
rect 177377 522020 177435 522037
rect 177377 521986 177389 522020
rect 177423 521986 177435 522020
rect 177786 522001 177854 522116
rect 178150 522114 178220 522315
rect 178150 522080 178167 522114
rect 178201 522080 178220 522114
rect 178150 522065 178220 522080
rect 178890 522150 178958 522167
rect 178890 522116 178907 522150
rect 178941 522116 178958 522150
rect 178890 522001 178958 522116
rect 179254 522114 179324 522315
rect 179254 522080 179271 522114
rect 179305 522080 179324 522114
rect 179254 522065 179324 522080
rect 179994 522150 180062 522167
rect 179994 522116 180011 522150
rect 180045 522116 180062 522150
rect 179994 522001 180062 522116
rect 180358 522114 180428 522315
rect 180358 522080 180375 522114
rect 180409 522080 180428 522114
rect 180358 522065 180428 522080
rect 181098 522150 181166 522167
rect 181098 522116 181115 522150
rect 181149 522116 181166 522150
rect 181098 522001 181166 522116
rect 181462 522114 181532 522315
rect 181885 522258 182403 522326
rect 181885 522224 181903 522258
rect 181937 522224 182351 522258
rect 182385 522224 182403 522258
rect 181885 522184 182403 522224
rect 181462 522080 181479 522114
rect 181513 522080 181532 522114
rect 181462 522065 181532 522080
rect 181885 522116 181963 522150
rect 181997 522116 182073 522150
rect 182107 522116 182127 522150
rect 181885 522046 182127 522116
rect 182161 522114 182403 522184
rect 182529 522331 182587 522402
rect 182529 522297 182541 522331
rect 182575 522297 182587 522331
rect 182621 522360 183690 522402
rect 182621 522326 182639 522360
rect 182673 522326 183639 522360
rect 183673 522326 183690 522360
rect 182621 522315 183690 522326
rect 183725 522360 184794 522402
rect 183725 522326 183743 522360
rect 183777 522326 184743 522360
rect 184777 522326 184794 522360
rect 183725 522315 184794 522326
rect 184829 522360 185898 522402
rect 184829 522326 184847 522360
rect 184881 522326 185847 522360
rect 185881 522326 185898 522360
rect 184829 522315 185898 522326
rect 185933 522360 187002 522402
rect 185933 522326 185951 522360
rect 185985 522326 186951 522360
rect 186985 522326 187002 522360
rect 185933 522315 187002 522326
rect 187221 522360 187463 522402
rect 187221 522326 187239 522360
rect 187273 522326 187411 522360
rect 187445 522326 187463 522360
rect 182529 522238 182587 522297
rect 182529 522204 182541 522238
rect 182575 522204 182587 522238
rect 182529 522169 182587 522204
rect 182161 522080 182181 522114
rect 182215 522080 182291 522114
rect 182325 522080 182403 522114
rect 182938 522150 183006 522167
rect 182938 522116 182955 522150
rect 182989 522116 183006 522150
rect 177377 521892 177435 521986
rect 177469 521987 178538 522001
rect 177469 521953 177487 521987
rect 177521 521953 178487 521987
rect 178521 521953 178538 521987
rect 177469 521892 178538 521953
rect 178573 521987 179642 522001
rect 178573 521953 178591 521987
rect 178625 521953 179591 521987
rect 179625 521953 179642 521987
rect 178573 521892 179642 521953
rect 179677 521987 180746 522001
rect 179677 521953 179695 521987
rect 179729 521953 180695 521987
rect 180729 521953 180746 521987
rect 179677 521892 180746 521953
rect 180781 521987 181850 522001
rect 180781 521953 180799 521987
rect 180833 521953 181799 521987
rect 181833 521953 181850 521987
rect 180781 521892 181850 521953
rect 181885 521987 182403 522046
rect 181885 521953 181903 521987
rect 181937 521953 182351 521987
rect 182385 521953 182403 521987
rect 181885 521892 182403 521953
rect 182529 522020 182587 522037
rect 182529 521986 182541 522020
rect 182575 521986 182587 522020
rect 182938 522001 183006 522116
rect 183302 522114 183372 522315
rect 183302 522080 183319 522114
rect 183353 522080 183372 522114
rect 183302 522065 183372 522080
rect 184042 522150 184110 522167
rect 184042 522116 184059 522150
rect 184093 522116 184110 522150
rect 184042 522001 184110 522116
rect 184406 522114 184476 522315
rect 184406 522080 184423 522114
rect 184457 522080 184476 522114
rect 184406 522065 184476 522080
rect 185146 522150 185214 522167
rect 185146 522116 185163 522150
rect 185197 522116 185214 522150
rect 185146 522001 185214 522116
rect 185510 522114 185580 522315
rect 185510 522080 185527 522114
rect 185561 522080 185580 522114
rect 185510 522065 185580 522080
rect 186250 522150 186318 522167
rect 186250 522116 186267 522150
rect 186301 522116 186318 522150
rect 186250 522001 186318 522116
rect 186614 522114 186684 522315
rect 186614 522080 186631 522114
rect 186665 522080 186684 522114
rect 186614 522065 186684 522080
rect 187221 522265 187463 522326
rect 187221 522231 187239 522265
rect 187273 522231 187411 522265
rect 187445 522231 187463 522265
rect 187221 522184 187463 522231
rect 187221 522110 187325 522184
rect 187221 522076 187271 522110
rect 187305 522076 187325 522110
rect 187359 522116 187379 522150
rect 187413 522116 187463 522150
rect 187359 522042 187463 522116
rect 182529 521892 182587 521986
rect 182621 521987 183690 522001
rect 182621 521953 182639 521987
rect 182673 521953 183639 521987
rect 183673 521953 183690 521987
rect 182621 521892 183690 521953
rect 183725 521987 184794 522001
rect 183725 521953 183743 521987
rect 183777 521953 184743 521987
rect 184777 521953 184794 521987
rect 183725 521892 184794 521953
rect 184829 521987 185898 522001
rect 184829 521953 184847 521987
rect 184881 521953 185847 521987
rect 185881 521953 185898 521987
rect 184829 521892 185898 521953
rect 185933 521987 187002 522001
rect 185933 521953 185951 521987
rect 185985 521953 186951 521987
rect 186985 521953 187002 521987
rect 185933 521892 187002 521953
rect 187221 521989 187463 522042
rect 187221 521955 187239 521989
rect 187273 521955 187411 521989
rect 187445 521955 187463 521989
rect 187221 521892 187463 521955
rect 172208 521858 172237 521892
rect 172271 521858 172329 521892
rect 172363 521858 172421 521892
rect 172455 521858 172513 521892
rect 172547 521858 172605 521892
rect 172639 521858 172697 521892
rect 172731 521858 172789 521892
rect 172823 521858 172881 521892
rect 172915 521858 172973 521892
rect 173007 521858 173065 521892
rect 173099 521858 173157 521892
rect 173191 521858 173249 521892
rect 173283 521858 173341 521892
rect 173375 521858 173433 521892
rect 173467 521858 173525 521892
rect 173559 521858 173617 521892
rect 173651 521858 173709 521892
rect 173743 521858 173801 521892
rect 173835 521858 173893 521892
rect 173927 521858 173985 521892
rect 174019 521858 174077 521892
rect 174111 521858 174169 521892
rect 174203 521858 174261 521892
rect 174295 521858 174353 521892
rect 174387 521858 174445 521892
rect 174479 521858 174537 521892
rect 174571 521858 174629 521892
rect 174663 521858 174721 521892
rect 174755 521858 174813 521892
rect 174847 521858 174905 521892
rect 174939 521858 174997 521892
rect 175031 521858 175089 521892
rect 175123 521858 175181 521892
rect 175215 521858 175273 521892
rect 175307 521858 175365 521892
rect 175399 521858 175457 521892
rect 175491 521858 175549 521892
rect 175583 521858 175641 521892
rect 175675 521858 175733 521892
rect 175767 521858 175825 521892
rect 175859 521858 175917 521892
rect 175951 521858 176009 521892
rect 176043 521858 176101 521892
rect 176135 521858 176193 521892
rect 176227 521858 176285 521892
rect 176319 521858 176377 521892
rect 176411 521858 176469 521892
rect 176503 521858 176561 521892
rect 176595 521858 176653 521892
rect 176687 521858 176745 521892
rect 176779 521858 176837 521892
rect 176871 521858 176929 521892
rect 176963 521858 177021 521892
rect 177055 521858 177113 521892
rect 177147 521858 177205 521892
rect 177239 521858 177297 521892
rect 177331 521858 177389 521892
rect 177423 521858 177481 521892
rect 177515 521858 177573 521892
rect 177607 521858 177665 521892
rect 177699 521858 177757 521892
rect 177791 521858 177849 521892
rect 177883 521858 177941 521892
rect 177975 521858 178033 521892
rect 178067 521858 178125 521892
rect 178159 521858 178217 521892
rect 178251 521858 178309 521892
rect 178343 521858 178401 521892
rect 178435 521858 178493 521892
rect 178527 521858 178585 521892
rect 178619 521858 178677 521892
rect 178711 521858 178769 521892
rect 178803 521858 178861 521892
rect 178895 521858 178953 521892
rect 178987 521858 179045 521892
rect 179079 521858 179137 521892
rect 179171 521858 179229 521892
rect 179263 521858 179321 521892
rect 179355 521858 179413 521892
rect 179447 521858 179505 521892
rect 179539 521858 179597 521892
rect 179631 521858 179689 521892
rect 179723 521858 179781 521892
rect 179815 521858 179873 521892
rect 179907 521858 179965 521892
rect 179999 521858 180057 521892
rect 180091 521858 180149 521892
rect 180183 521858 180241 521892
rect 180275 521858 180333 521892
rect 180367 521858 180425 521892
rect 180459 521858 180517 521892
rect 180551 521858 180609 521892
rect 180643 521858 180701 521892
rect 180735 521858 180793 521892
rect 180827 521858 180885 521892
rect 180919 521858 180977 521892
rect 181011 521858 181069 521892
rect 181103 521858 181161 521892
rect 181195 521858 181253 521892
rect 181287 521858 181345 521892
rect 181379 521858 181437 521892
rect 181471 521858 181529 521892
rect 181563 521858 181621 521892
rect 181655 521858 181713 521892
rect 181747 521858 181805 521892
rect 181839 521858 181897 521892
rect 181931 521858 181989 521892
rect 182023 521858 182081 521892
rect 182115 521858 182173 521892
rect 182207 521858 182265 521892
rect 182299 521858 182357 521892
rect 182391 521858 182449 521892
rect 182483 521858 182541 521892
rect 182575 521858 182633 521892
rect 182667 521858 182725 521892
rect 182759 521858 182817 521892
rect 182851 521858 182909 521892
rect 182943 521858 183001 521892
rect 183035 521858 183093 521892
rect 183127 521858 183185 521892
rect 183219 521858 183277 521892
rect 183311 521858 183369 521892
rect 183403 521858 183461 521892
rect 183495 521858 183553 521892
rect 183587 521858 183645 521892
rect 183679 521858 183737 521892
rect 183771 521858 183829 521892
rect 183863 521858 183921 521892
rect 183955 521858 184013 521892
rect 184047 521858 184105 521892
rect 184139 521858 184197 521892
rect 184231 521858 184289 521892
rect 184323 521858 184381 521892
rect 184415 521858 184473 521892
rect 184507 521858 184565 521892
rect 184599 521858 184657 521892
rect 184691 521858 184749 521892
rect 184783 521858 184841 521892
rect 184875 521858 184933 521892
rect 184967 521858 185025 521892
rect 185059 521858 185117 521892
rect 185151 521858 185209 521892
rect 185243 521858 185301 521892
rect 185335 521858 185393 521892
rect 185427 521858 185485 521892
rect 185519 521858 185577 521892
rect 185611 521858 185669 521892
rect 185703 521858 185761 521892
rect 185795 521858 185853 521892
rect 185887 521858 185945 521892
rect 185979 521858 186037 521892
rect 186071 521858 186129 521892
rect 186163 521858 186221 521892
rect 186255 521858 186313 521892
rect 186347 521858 186405 521892
rect 186439 521858 186497 521892
rect 186531 521858 186589 521892
rect 186623 521858 186681 521892
rect 186715 521858 186773 521892
rect 186807 521858 186865 521892
rect 186899 521858 186957 521892
rect 186991 521858 187049 521892
rect 187083 521858 187141 521892
rect 187175 521858 187233 521892
rect 187267 521858 187325 521892
rect 187359 521858 187417 521892
rect 187451 521858 187480 521892
rect 172225 521795 172467 521858
rect 172225 521761 172243 521795
rect 172277 521761 172415 521795
rect 172449 521761 172467 521795
rect 172225 521708 172467 521761
rect 172501 521797 173570 521858
rect 172501 521763 172519 521797
rect 172553 521763 173519 521797
rect 173553 521763 173570 521797
rect 172501 521749 173570 521763
rect 173605 521797 174674 521858
rect 173605 521763 173623 521797
rect 173657 521763 174623 521797
rect 174657 521763 174674 521797
rect 173605 521749 174674 521763
rect 174801 521764 174859 521858
rect 172225 521634 172329 521708
rect 172225 521600 172275 521634
rect 172309 521600 172329 521634
rect 172363 521640 172383 521674
rect 172417 521640 172467 521674
rect 172363 521566 172467 521640
rect 172818 521634 172886 521749
rect 172818 521600 172835 521634
rect 172869 521600 172886 521634
rect 172818 521583 172886 521600
rect 173182 521670 173252 521685
rect 173182 521636 173199 521670
rect 173233 521636 173252 521670
rect 172225 521519 172467 521566
rect 172225 521485 172243 521519
rect 172277 521485 172415 521519
rect 172449 521485 172467 521519
rect 172225 521424 172467 521485
rect 173182 521435 173252 521636
rect 173922 521634 173990 521749
rect 174801 521730 174813 521764
rect 174847 521730 174859 521764
rect 174893 521797 175962 521858
rect 174893 521763 174911 521797
rect 174945 521763 175911 521797
rect 175945 521763 175962 521797
rect 174893 521749 175962 521763
rect 175997 521797 177066 521858
rect 175997 521763 176015 521797
rect 176049 521763 177015 521797
rect 177049 521763 177066 521797
rect 175997 521749 177066 521763
rect 177101 521797 178170 521858
rect 177101 521763 177119 521797
rect 177153 521763 178119 521797
rect 178153 521763 178170 521797
rect 177101 521749 178170 521763
rect 178205 521797 179274 521858
rect 178205 521763 178223 521797
rect 178257 521763 179223 521797
rect 179257 521763 179274 521797
rect 178205 521749 179274 521763
rect 179309 521797 179827 521858
rect 179309 521763 179327 521797
rect 179361 521763 179775 521797
rect 179809 521763 179827 521797
rect 174801 521713 174859 521730
rect 173922 521600 173939 521634
rect 173973 521600 173990 521634
rect 173922 521583 173990 521600
rect 174286 521670 174356 521685
rect 174286 521636 174303 521670
rect 174337 521636 174356 521670
rect 174286 521435 174356 521636
rect 175210 521634 175278 521749
rect 175210 521600 175227 521634
rect 175261 521600 175278 521634
rect 175210 521583 175278 521600
rect 175574 521670 175644 521685
rect 175574 521636 175591 521670
rect 175625 521636 175644 521670
rect 174801 521546 174859 521581
rect 174801 521512 174813 521546
rect 174847 521512 174859 521546
rect 174801 521453 174859 521512
rect 172225 521390 172243 521424
rect 172277 521390 172415 521424
rect 172449 521390 172467 521424
rect 172225 521348 172467 521390
rect 172501 521424 173570 521435
rect 172501 521390 172519 521424
rect 172553 521390 173519 521424
rect 173553 521390 173570 521424
rect 172501 521348 173570 521390
rect 173605 521424 174674 521435
rect 173605 521390 173623 521424
rect 173657 521390 174623 521424
rect 174657 521390 174674 521424
rect 173605 521348 174674 521390
rect 174801 521419 174813 521453
rect 174847 521419 174859 521453
rect 175574 521435 175644 521636
rect 176314 521634 176382 521749
rect 176314 521600 176331 521634
rect 176365 521600 176382 521634
rect 176314 521583 176382 521600
rect 176678 521670 176748 521685
rect 176678 521636 176695 521670
rect 176729 521636 176748 521670
rect 176678 521435 176748 521636
rect 177418 521634 177486 521749
rect 177418 521600 177435 521634
rect 177469 521600 177486 521634
rect 177418 521583 177486 521600
rect 177782 521670 177852 521685
rect 177782 521636 177799 521670
rect 177833 521636 177852 521670
rect 177782 521435 177852 521636
rect 178522 521634 178590 521749
rect 179309 521704 179827 521763
rect 179953 521764 180011 521858
rect 179953 521730 179965 521764
rect 179999 521730 180011 521764
rect 180045 521797 181114 521858
rect 180045 521763 180063 521797
rect 180097 521763 181063 521797
rect 181097 521763 181114 521797
rect 180045 521749 181114 521763
rect 181149 521797 182218 521858
rect 181149 521763 181167 521797
rect 181201 521763 182167 521797
rect 182201 521763 182218 521797
rect 181149 521749 182218 521763
rect 182253 521797 183322 521858
rect 182253 521763 182271 521797
rect 182305 521763 183271 521797
rect 183305 521763 183322 521797
rect 182253 521749 183322 521763
rect 183357 521797 184426 521858
rect 183357 521763 183375 521797
rect 183409 521763 184375 521797
rect 184409 521763 184426 521797
rect 183357 521749 184426 521763
rect 184461 521797 184979 521858
rect 184461 521763 184479 521797
rect 184513 521763 184927 521797
rect 184961 521763 184979 521797
rect 179953 521713 180011 521730
rect 178522 521600 178539 521634
rect 178573 521600 178590 521634
rect 178522 521583 178590 521600
rect 178886 521670 178956 521685
rect 178886 521636 178903 521670
rect 178937 521636 178956 521670
rect 178886 521435 178956 521636
rect 179309 521634 179551 521704
rect 179309 521600 179387 521634
rect 179421 521600 179497 521634
rect 179531 521600 179551 521634
rect 179585 521636 179605 521670
rect 179639 521636 179715 521670
rect 179749 521636 179827 521670
rect 179585 521566 179827 521636
rect 180362 521634 180430 521749
rect 180362 521600 180379 521634
rect 180413 521600 180430 521634
rect 180362 521583 180430 521600
rect 180726 521670 180796 521685
rect 180726 521636 180743 521670
rect 180777 521636 180796 521670
rect 179309 521526 179827 521566
rect 179309 521492 179327 521526
rect 179361 521492 179775 521526
rect 179809 521492 179827 521526
rect 174801 521348 174859 521419
rect 174893 521424 175962 521435
rect 174893 521390 174911 521424
rect 174945 521390 175911 521424
rect 175945 521390 175962 521424
rect 174893 521348 175962 521390
rect 175997 521424 177066 521435
rect 175997 521390 176015 521424
rect 176049 521390 177015 521424
rect 177049 521390 177066 521424
rect 175997 521348 177066 521390
rect 177101 521424 178170 521435
rect 177101 521390 177119 521424
rect 177153 521390 178119 521424
rect 178153 521390 178170 521424
rect 177101 521348 178170 521390
rect 178205 521424 179274 521435
rect 178205 521390 178223 521424
rect 178257 521390 179223 521424
rect 179257 521390 179274 521424
rect 178205 521348 179274 521390
rect 179309 521424 179827 521492
rect 179309 521390 179327 521424
rect 179361 521390 179775 521424
rect 179809 521390 179827 521424
rect 179309 521348 179827 521390
rect 179953 521546 180011 521581
rect 179953 521512 179965 521546
rect 179999 521512 180011 521546
rect 179953 521453 180011 521512
rect 179953 521419 179965 521453
rect 179999 521419 180011 521453
rect 180726 521435 180796 521636
rect 181466 521634 181534 521749
rect 181466 521600 181483 521634
rect 181517 521600 181534 521634
rect 181466 521583 181534 521600
rect 181830 521670 181900 521685
rect 181830 521636 181847 521670
rect 181881 521636 181900 521670
rect 181830 521435 181900 521636
rect 182570 521634 182638 521749
rect 182570 521600 182587 521634
rect 182621 521600 182638 521634
rect 182570 521583 182638 521600
rect 182934 521670 183004 521685
rect 182934 521636 182951 521670
rect 182985 521636 183004 521670
rect 182934 521435 183004 521636
rect 183674 521634 183742 521749
rect 184461 521704 184979 521763
rect 185105 521764 185163 521858
rect 185105 521730 185117 521764
rect 185151 521730 185163 521764
rect 185197 521797 186266 521858
rect 185197 521763 185215 521797
rect 185249 521763 186215 521797
rect 186249 521763 186266 521797
rect 185197 521749 186266 521763
rect 186301 521797 187003 521858
rect 186301 521763 186319 521797
rect 186353 521763 186951 521797
rect 186985 521763 187003 521797
rect 185105 521713 185163 521730
rect 183674 521600 183691 521634
rect 183725 521600 183742 521634
rect 183674 521583 183742 521600
rect 184038 521670 184108 521685
rect 184038 521636 184055 521670
rect 184089 521636 184108 521670
rect 184038 521435 184108 521636
rect 184461 521634 184703 521704
rect 184461 521600 184539 521634
rect 184573 521600 184649 521634
rect 184683 521600 184703 521634
rect 184737 521636 184757 521670
rect 184791 521636 184867 521670
rect 184901 521636 184979 521670
rect 184737 521566 184979 521636
rect 185514 521634 185582 521749
rect 186301 521704 187003 521763
rect 187221 521795 187463 521858
rect 187221 521761 187239 521795
rect 187273 521761 187411 521795
rect 187445 521761 187463 521795
rect 187221 521708 187463 521761
rect 185514 521600 185531 521634
rect 185565 521600 185582 521634
rect 185514 521583 185582 521600
rect 185878 521670 185948 521685
rect 185878 521636 185895 521670
rect 185929 521636 185948 521670
rect 184461 521526 184979 521566
rect 184461 521492 184479 521526
rect 184513 521492 184927 521526
rect 184961 521492 184979 521526
rect 179953 521348 180011 521419
rect 180045 521424 181114 521435
rect 180045 521390 180063 521424
rect 180097 521390 181063 521424
rect 181097 521390 181114 521424
rect 180045 521348 181114 521390
rect 181149 521424 182218 521435
rect 181149 521390 181167 521424
rect 181201 521390 182167 521424
rect 182201 521390 182218 521424
rect 181149 521348 182218 521390
rect 182253 521424 183322 521435
rect 182253 521390 182271 521424
rect 182305 521390 183271 521424
rect 183305 521390 183322 521424
rect 182253 521348 183322 521390
rect 183357 521424 184426 521435
rect 183357 521390 183375 521424
rect 183409 521390 184375 521424
rect 184409 521390 184426 521424
rect 183357 521348 184426 521390
rect 184461 521424 184979 521492
rect 184461 521390 184479 521424
rect 184513 521390 184927 521424
rect 184961 521390 184979 521424
rect 184461 521348 184979 521390
rect 185105 521546 185163 521581
rect 185105 521512 185117 521546
rect 185151 521512 185163 521546
rect 185105 521453 185163 521512
rect 185105 521419 185117 521453
rect 185151 521419 185163 521453
rect 185878 521435 185948 521636
rect 186301 521634 186631 521704
rect 186301 521600 186379 521634
rect 186413 521600 186478 521634
rect 186512 521600 186577 521634
rect 186611 521600 186631 521634
rect 186665 521636 186685 521670
rect 186719 521636 186788 521670
rect 186822 521636 186891 521670
rect 186925 521636 187003 521670
rect 186665 521566 187003 521636
rect 186301 521526 187003 521566
rect 186301 521492 186319 521526
rect 186353 521492 186951 521526
rect 186985 521492 187003 521526
rect 185105 521348 185163 521419
rect 185197 521424 186266 521435
rect 185197 521390 185215 521424
rect 185249 521390 186215 521424
rect 186249 521390 186266 521424
rect 185197 521348 186266 521390
rect 186301 521424 187003 521492
rect 186301 521390 186319 521424
rect 186353 521390 186951 521424
rect 186985 521390 187003 521424
rect 186301 521348 187003 521390
rect 187221 521640 187271 521674
rect 187305 521640 187325 521674
rect 187221 521566 187325 521640
rect 187359 521634 187463 521708
rect 187359 521600 187379 521634
rect 187413 521600 187463 521634
rect 187221 521519 187463 521566
rect 187221 521485 187239 521519
rect 187273 521485 187411 521519
rect 187445 521485 187463 521519
rect 187221 521424 187463 521485
rect 187221 521390 187239 521424
rect 187273 521390 187411 521424
rect 187445 521390 187463 521424
rect 187221 521348 187463 521390
rect 172208 521314 172237 521348
rect 172271 521314 172329 521348
rect 172363 521314 172421 521348
rect 172455 521314 172513 521348
rect 172547 521314 172605 521348
rect 172639 521314 172697 521348
rect 172731 521314 172789 521348
rect 172823 521314 172881 521348
rect 172915 521314 172973 521348
rect 173007 521314 173065 521348
rect 173099 521314 173157 521348
rect 173191 521314 173249 521348
rect 173283 521314 173341 521348
rect 173375 521314 173433 521348
rect 173467 521314 173525 521348
rect 173559 521314 173617 521348
rect 173651 521314 173709 521348
rect 173743 521314 173801 521348
rect 173835 521314 173893 521348
rect 173927 521314 173985 521348
rect 174019 521314 174077 521348
rect 174111 521314 174169 521348
rect 174203 521314 174261 521348
rect 174295 521314 174353 521348
rect 174387 521314 174445 521348
rect 174479 521314 174537 521348
rect 174571 521314 174629 521348
rect 174663 521314 174721 521348
rect 174755 521314 174813 521348
rect 174847 521314 174905 521348
rect 174939 521314 174997 521348
rect 175031 521314 175089 521348
rect 175123 521314 175181 521348
rect 175215 521314 175273 521348
rect 175307 521314 175365 521348
rect 175399 521314 175457 521348
rect 175491 521314 175549 521348
rect 175583 521314 175641 521348
rect 175675 521314 175733 521348
rect 175767 521314 175825 521348
rect 175859 521314 175917 521348
rect 175951 521314 176009 521348
rect 176043 521314 176101 521348
rect 176135 521314 176193 521348
rect 176227 521314 176285 521348
rect 176319 521314 176377 521348
rect 176411 521314 176469 521348
rect 176503 521314 176561 521348
rect 176595 521314 176653 521348
rect 176687 521314 176745 521348
rect 176779 521314 176837 521348
rect 176871 521314 176929 521348
rect 176963 521314 177021 521348
rect 177055 521314 177113 521348
rect 177147 521314 177205 521348
rect 177239 521314 177297 521348
rect 177331 521314 177389 521348
rect 177423 521314 177481 521348
rect 177515 521314 177573 521348
rect 177607 521314 177665 521348
rect 177699 521314 177757 521348
rect 177791 521314 177849 521348
rect 177883 521314 177941 521348
rect 177975 521314 178033 521348
rect 178067 521314 178125 521348
rect 178159 521314 178217 521348
rect 178251 521314 178309 521348
rect 178343 521314 178401 521348
rect 178435 521314 178493 521348
rect 178527 521314 178585 521348
rect 178619 521314 178677 521348
rect 178711 521314 178769 521348
rect 178803 521314 178861 521348
rect 178895 521314 178953 521348
rect 178987 521314 179045 521348
rect 179079 521314 179137 521348
rect 179171 521314 179229 521348
rect 179263 521314 179321 521348
rect 179355 521314 179413 521348
rect 179447 521314 179505 521348
rect 179539 521314 179597 521348
rect 179631 521314 179689 521348
rect 179723 521314 179781 521348
rect 179815 521314 179873 521348
rect 179907 521314 179965 521348
rect 179999 521314 180057 521348
rect 180091 521314 180149 521348
rect 180183 521314 180241 521348
rect 180275 521314 180333 521348
rect 180367 521314 180425 521348
rect 180459 521314 180517 521348
rect 180551 521314 180609 521348
rect 180643 521314 180701 521348
rect 180735 521314 180793 521348
rect 180827 521314 180885 521348
rect 180919 521314 180977 521348
rect 181011 521314 181069 521348
rect 181103 521314 181161 521348
rect 181195 521314 181253 521348
rect 181287 521314 181345 521348
rect 181379 521314 181437 521348
rect 181471 521314 181529 521348
rect 181563 521314 181621 521348
rect 181655 521314 181713 521348
rect 181747 521314 181805 521348
rect 181839 521314 181897 521348
rect 181931 521314 181989 521348
rect 182023 521314 182081 521348
rect 182115 521314 182173 521348
rect 182207 521314 182265 521348
rect 182299 521314 182357 521348
rect 182391 521314 182449 521348
rect 182483 521314 182541 521348
rect 182575 521314 182633 521348
rect 182667 521314 182725 521348
rect 182759 521314 182817 521348
rect 182851 521314 182909 521348
rect 182943 521314 183001 521348
rect 183035 521314 183093 521348
rect 183127 521314 183185 521348
rect 183219 521314 183277 521348
rect 183311 521314 183369 521348
rect 183403 521314 183461 521348
rect 183495 521314 183553 521348
rect 183587 521314 183645 521348
rect 183679 521314 183737 521348
rect 183771 521314 183829 521348
rect 183863 521314 183921 521348
rect 183955 521314 184013 521348
rect 184047 521314 184105 521348
rect 184139 521314 184197 521348
rect 184231 521314 184289 521348
rect 184323 521314 184381 521348
rect 184415 521314 184473 521348
rect 184507 521314 184565 521348
rect 184599 521314 184657 521348
rect 184691 521314 184749 521348
rect 184783 521314 184841 521348
rect 184875 521314 184933 521348
rect 184967 521314 185025 521348
rect 185059 521314 185117 521348
rect 185151 521314 185209 521348
rect 185243 521314 185301 521348
rect 185335 521314 185393 521348
rect 185427 521314 185485 521348
rect 185519 521314 185577 521348
rect 185611 521314 185669 521348
rect 185703 521314 185761 521348
rect 185795 521314 185853 521348
rect 185887 521314 185945 521348
rect 185979 521314 186037 521348
rect 186071 521314 186129 521348
rect 186163 521314 186221 521348
rect 186255 521314 186313 521348
rect 186347 521314 186405 521348
rect 186439 521314 186497 521348
rect 186531 521314 186589 521348
rect 186623 521314 186681 521348
rect 186715 521314 186773 521348
rect 186807 521314 186865 521348
rect 186899 521314 186957 521348
rect 186991 521314 187049 521348
rect 187083 521314 187141 521348
rect 187175 521314 187233 521348
rect 187267 521314 187325 521348
rect 187359 521314 187417 521348
rect 187451 521314 187480 521348
rect 172225 521272 172467 521314
rect 172225 521238 172243 521272
rect 172277 521238 172415 521272
rect 172449 521238 172467 521272
rect 172225 521177 172467 521238
rect 172501 521272 173570 521314
rect 172501 521238 172519 521272
rect 172553 521238 173519 521272
rect 173553 521238 173570 521272
rect 172501 521227 173570 521238
rect 173605 521272 174674 521314
rect 173605 521238 173623 521272
rect 173657 521238 174623 521272
rect 174657 521238 174674 521272
rect 173605 521227 174674 521238
rect 174709 521272 175778 521314
rect 174709 521238 174727 521272
rect 174761 521238 175727 521272
rect 175761 521238 175778 521272
rect 174709 521227 175778 521238
rect 175813 521272 176882 521314
rect 175813 521238 175831 521272
rect 175865 521238 176831 521272
rect 176865 521238 176882 521272
rect 175813 521227 176882 521238
rect 176917 521272 177251 521314
rect 176917 521238 176935 521272
rect 176969 521238 177199 521272
rect 177233 521238 177251 521272
rect 172225 521143 172243 521177
rect 172277 521143 172415 521177
rect 172449 521143 172467 521177
rect 172225 521096 172467 521143
rect 172225 521028 172275 521062
rect 172309 521028 172329 521062
rect 172225 520954 172329 521028
rect 172363 521022 172467 521096
rect 172363 520988 172383 521022
rect 172417 520988 172467 521022
rect 172818 521062 172886 521079
rect 172818 521028 172835 521062
rect 172869 521028 172886 521062
rect 172225 520901 172467 520954
rect 172818 520913 172886 521028
rect 173182 521026 173252 521227
rect 173182 520992 173199 521026
rect 173233 520992 173252 521026
rect 173182 520977 173252 520992
rect 173922 521062 173990 521079
rect 173922 521028 173939 521062
rect 173973 521028 173990 521062
rect 173922 520913 173990 521028
rect 174286 521026 174356 521227
rect 174286 520992 174303 521026
rect 174337 520992 174356 521026
rect 174286 520977 174356 520992
rect 175026 521062 175094 521079
rect 175026 521028 175043 521062
rect 175077 521028 175094 521062
rect 175026 520913 175094 521028
rect 175390 521026 175460 521227
rect 175390 520992 175407 521026
rect 175441 520992 175460 521026
rect 175390 520977 175460 520992
rect 176130 521062 176198 521079
rect 176130 521028 176147 521062
rect 176181 521028 176198 521062
rect 176130 520913 176198 521028
rect 176494 521026 176564 521227
rect 176917 521170 177251 521238
rect 176917 521136 176935 521170
rect 176969 521136 177199 521170
rect 177233 521136 177251 521170
rect 176917 521096 177251 521136
rect 176494 520992 176511 521026
rect 176545 520992 176564 521026
rect 176494 520977 176564 520992
rect 176917 521028 176937 521062
rect 176971 521028 177067 521062
rect 176917 520958 177067 521028
rect 177101 521026 177251 521096
rect 177377 521243 177435 521314
rect 177377 521209 177389 521243
rect 177423 521209 177435 521243
rect 177469 521272 178538 521314
rect 177469 521238 177487 521272
rect 177521 521238 178487 521272
rect 178521 521238 178538 521272
rect 177469 521227 178538 521238
rect 178573 521272 179642 521314
rect 178573 521238 178591 521272
rect 178625 521238 179591 521272
rect 179625 521238 179642 521272
rect 178573 521227 179642 521238
rect 179677 521272 180746 521314
rect 179677 521238 179695 521272
rect 179729 521238 180695 521272
rect 180729 521238 180746 521272
rect 179677 521227 180746 521238
rect 180781 521272 181850 521314
rect 180781 521238 180799 521272
rect 180833 521238 181799 521272
rect 181833 521238 181850 521272
rect 180781 521227 181850 521238
rect 181885 521272 182403 521314
rect 181885 521238 181903 521272
rect 181937 521238 182351 521272
rect 182385 521238 182403 521272
rect 177377 521150 177435 521209
rect 177377 521116 177389 521150
rect 177423 521116 177435 521150
rect 177377 521081 177435 521116
rect 177101 520992 177197 521026
rect 177231 520992 177251 521026
rect 177786 521062 177854 521079
rect 177786 521028 177803 521062
rect 177837 521028 177854 521062
rect 172225 520867 172243 520901
rect 172277 520867 172415 520901
rect 172449 520867 172467 520901
rect 172225 520804 172467 520867
rect 172501 520899 173570 520913
rect 172501 520865 172519 520899
rect 172553 520865 173519 520899
rect 173553 520865 173570 520899
rect 172501 520804 173570 520865
rect 173605 520899 174674 520913
rect 173605 520865 173623 520899
rect 173657 520865 174623 520899
rect 174657 520865 174674 520899
rect 173605 520804 174674 520865
rect 174709 520899 175778 520913
rect 174709 520865 174727 520899
rect 174761 520865 175727 520899
rect 175761 520865 175778 520899
rect 174709 520804 175778 520865
rect 175813 520899 176882 520913
rect 175813 520865 175831 520899
rect 175865 520865 176831 520899
rect 176865 520865 176882 520899
rect 175813 520804 176882 520865
rect 176917 520906 177251 520958
rect 176917 520872 176935 520906
rect 176969 520872 177199 520906
rect 177233 520872 177251 520906
rect 176917 520804 177251 520872
rect 177377 520932 177435 520949
rect 177377 520898 177389 520932
rect 177423 520898 177435 520932
rect 177786 520913 177854 521028
rect 178150 521026 178220 521227
rect 178150 520992 178167 521026
rect 178201 520992 178220 521026
rect 178150 520977 178220 520992
rect 178890 521062 178958 521079
rect 178890 521028 178907 521062
rect 178941 521028 178958 521062
rect 178890 520913 178958 521028
rect 179254 521026 179324 521227
rect 179254 520992 179271 521026
rect 179305 520992 179324 521026
rect 179254 520977 179324 520992
rect 179994 521062 180062 521079
rect 179994 521028 180011 521062
rect 180045 521028 180062 521062
rect 179994 520913 180062 521028
rect 180358 521026 180428 521227
rect 180358 520992 180375 521026
rect 180409 520992 180428 521026
rect 180358 520977 180428 520992
rect 181098 521062 181166 521079
rect 181098 521028 181115 521062
rect 181149 521028 181166 521062
rect 181098 520913 181166 521028
rect 181462 521026 181532 521227
rect 181885 521170 182403 521238
rect 181885 521136 181903 521170
rect 181937 521136 182351 521170
rect 182385 521136 182403 521170
rect 181885 521096 182403 521136
rect 181462 520992 181479 521026
rect 181513 520992 181532 521026
rect 181462 520977 181532 520992
rect 181885 521028 181963 521062
rect 181997 521028 182073 521062
rect 182107 521028 182127 521062
rect 181885 520958 182127 521028
rect 182161 521026 182403 521096
rect 182529 521243 182587 521314
rect 182529 521209 182541 521243
rect 182575 521209 182587 521243
rect 182621 521272 183690 521314
rect 182621 521238 182639 521272
rect 182673 521238 183639 521272
rect 183673 521238 183690 521272
rect 182621 521227 183690 521238
rect 183725 521272 184794 521314
rect 183725 521238 183743 521272
rect 183777 521238 184743 521272
rect 184777 521238 184794 521272
rect 183725 521227 184794 521238
rect 184829 521272 185898 521314
rect 184829 521238 184847 521272
rect 184881 521238 185847 521272
rect 185881 521238 185898 521272
rect 184829 521227 185898 521238
rect 185933 521272 187002 521314
rect 185933 521238 185951 521272
rect 185985 521238 186951 521272
rect 186985 521238 187002 521272
rect 185933 521227 187002 521238
rect 187221 521272 187463 521314
rect 187221 521238 187239 521272
rect 187273 521238 187411 521272
rect 187445 521238 187463 521272
rect 182529 521150 182587 521209
rect 182529 521116 182541 521150
rect 182575 521116 182587 521150
rect 182529 521081 182587 521116
rect 182161 520992 182181 521026
rect 182215 520992 182291 521026
rect 182325 520992 182403 521026
rect 182938 521062 183006 521079
rect 182938 521028 182955 521062
rect 182989 521028 183006 521062
rect 177377 520804 177435 520898
rect 177469 520899 178538 520913
rect 177469 520865 177487 520899
rect 177521 520865 178487 520899
rect 178521 520865 178538 520899
rect 177469 520804 178538 520865
rect 178573 520899 179642 520913
rect 178573 520865 178591 520899
rect 178625 520865 179591 520899
rect 179625 520865 179642 520899
rect 178573 520804 179642 520865
rect 179677 520899 180746 520913
rect 179677 520865 179695 520899
rect 179729 520865 180695 520899
rect 180729 520865 180746 520899
rect 179677 520804 180746 520865
rect 180781 520899 181850 520913
rect 180781 520865 180799 520899
rect 180833 520865 181799 520899
rect 181833 520865 181850 520899
rect 180781 520804 181850 520865
rect 181885 520899 182403 520958
rect 181885 520865 181903 520899
rect 181937 520865 182351 520899
rect 182385 520865 182403 520899
rect 181885 520804 182403 520865
rect 182529 520932 182587 520949
rect 182529 520898 182541 520932
rect 182575 520898 182587 520932
rect 182938 520913 183006 521028
rect 183302 521026 183372 521227
rect 183302 520992 183319 521026
rect 183353 520992 183372 521026
rect 183302 520977 183372 520992
rect 184042 521062 184110 521079
rect 184042 521028 184059 521062
rect 184093 521028 184110 521062
rect 184042 520913 184110 521028
rect 184406 521026 184476 521227
rect 184406 520992 184423 521026
rect 184457 520992 184476 521026
rect 184406 520977 184476 520992
rect 185146 521062 185214 521079
rect 185146 521028 185163 521062
rect 185197 521028 185214 521062
rect 185146 520913 185214 521028
rect 185510 521026 185580 521227
rect 185510 520992 185527 521026
rect 185561 520992 185580 521026
rect 185510 520977 185580 520992
rect 186250 521062 186318 521079
rect 186250 521028 186267 521062
rect 186301 521028 186318 521062
rect 186250 520913 186318 521028
rect 186614 521026 186684 521227
rect 186614 520992 186631 521026
rect 186665 520992 186684 521026
rect 186614 520977 186684 520992
rect 187221 521177 187463 521238
rect 187221 521143 187239 521177
rect 187273 521143 187411 521177
rect 187445 521143 187463 521177
rect 187221 521096 187463 521143
rect 187221 521022 187325 521096
rect 187221 520988 187271 521022
rect 187305 520988 187325 521022
rect 187359 521028 187379 521062
rect 187413 521028 187463 521062
rect 187359 520954 187463 521028
rect 182529 520804 182587 520898
rect 182621 520899 183690 520913
rect 182621 520865 182639 520899
rect 182673 520865 183639 520899
rect 183673 520865 183690 520899
rect 182621 520804 183690 520865
rect 183725 520899 184794 520913
rect 183725 520865 183743 520899
rect 183777 520865 184743 520899
rect 184777 520865 184794 520899
rect 183725 520804 184794 520865
rect 184829 520899 185898 520913
rect 184829 520865 184847 520899
rect 184881 520865 185847 520899
rect 185881 520865 185898 520899
rect 184829 520804 185898 520865
rect 185933 520899 187002 520913
rect 185933 520865 185951 520899
rect 185985 520865 186951 520899
rect 186985 520865 187002 520899
rect 185933 520804 187002 520865
rect 187221 520901 187463 520954
rect 187221 520867 187239 520901
rect 187273 520867 187411 520901
rect 187445 520867 187463 520901
rect 187221 520804 187463 520867
rect 172208 520770 172237 520804
rect 172271 520770 172329 520804
rect 172363 520770 172421 520804
rect 172455 520770 172513 520804
rect 172547 520770 172605 520804
rect 172639 520770 172697 520804
rect 172731 520770 172789 520804
rect 172823 520770 172881 520804
rect 172915 520770 172973 520804
rect 173007 520770 173065 520804
rect 173099 520770 173157 520804
rect 173191 520770 173249 520804
rect 173283 520770 173341 520804
rect 173375 520770 173433 520804
rect 173467 520770 173525 520804
rect 173559 520770 173617 520804
rect 173651 520770 173709 520804
rect 173743 520770 173801 520804
rect 173835 520770 173893 520804
rect 173927 520770 173985 520804
rect 174019 520770 174077 520804
rect 174111 520770 174169 520804
rect 174203 520770 174261 520804
rect 174295 520770 174353 520804
rect 174387 520770 174445 520804
rect 174479 520770 174537 520804
rect 174571 520770 174629 520804
rect 174663 520770 174721 520804
rect 174755 520770 174813 520804
rect 174847 520770 174905 520804
rect 174939 520770 174997 520804
rect 175031 520770 175089 520804
rect 175123 520770 175181 520804
rect 175215 520770 175273 520804
rect 175307 520770 175365 520804
rect 175399 520770 175457 520804
rect 175491 520770 175549 520804
rect 175583 520770 175641 520804
rect 175675 520770 175733 520804
rect 175767 520770 175825 520804
rect 175859 520770 175917 520804
rect 175951 520770 176009 520804
rect 176043 520770 176101 520804
rect 176135 520770 176193 520804
rect 176227 520770 176285 520804
rect 176319 520770 176377 520804
rect 176411 520770 176469 520804
rect 176503 520770 176561 520804
rect 176595 520770 176653 520804
rect 176687 520770 176745 520804
rect 176779 520770 176837 520804
rect 176871 520770 176929 520804
rect 176963 520770 177021 520804
rect 177055 520770 177113 520804
rect 177147 520770 177205 520804
rect 177239 520770 177297 520804
rect 177331 520770 177389 520804
rect 177423 520770 177481 520804
rect 177515 520770 177573 520804
rect 177607 520770 177665 520804
rect 177699 520770 177757 520804
rect 177791 520770 177849 520804
rect 177883 520770 177941 520804
rect 177975 520770 178033 520804
rect 178067 520770 178125 520804
rect 178159 520770 178217 520804
rect 178251 520770 178309 520804
rect 178343 520770 178401 520804
rect 178435 520770 178493 520804
rect 178527 520770 178585 520804
rect 178619 520770 178677 520804
rect 178711 520770 178769 520804
rect 178803 520770 178861 520804
rect 178895 520770 178953 520804
rect 178987 520770 179045 520804
rect 179079 520770 179137 520804
rect 179171 520770 179229 520804
rect 179263 520770 179321 520804
rect 179355 520770 179413 520804
rect 179447 520770 179505 520804
rect 179539 520770 179597 520804
rect 179631 520770 179689 520804
rect 179723 520770 179781 520804
rect 179815 520770 179873 520804
rect 179907 520770 179965 520804
rect 179999 520770 180057 520804
rect 180091 520770 180149 520804
rect 180183 520770 180241 520804
rect 180275 520770 180333 520804
rect 180367 520770 180425 520804
rect 180459 520770 180517 520804
rect 180551 520770 180609 520804
rect 180643 520770 180701 520804
rect 180735 520770 180793 520804
rect 180827 520770 180885 520804
rect 180919 520770 180977 520804
rect 181011 520770 181069 520804
rect 181103 520770 181161 520804
rect 181195 520770 181253 520804
rect 181287 520770 181345 520804
rect 181379 520770 181437 520804
rect 181471 520770 181529 520804
rect 181563 520770 181621 520804
rect 181655 520770 181713 520804
rect 181747 520770 181805 520804
rect 181839 520770 181897 520804
rect 181931 520770 181989 520804
rect 182023 520770 182081 520804
rect 182115 520770 182173 520804
rect 182207 520770 182265 520804
rect 182299 520770 182357 520804
rect 182391 520770 182449 520804
rect 182483 520770 182541 520804
rect 182575 520770 182633 520804
rect 182667 520770 182725 520804
rect 182759 520770 182817 520804
rect 182851 520770 182909 520804
rect 182943 520770 183001 520804
rect 183035 520770 183093 520804
rect 183127 520770 183185 520804
rect 183219 520770 183277 520804
rect 183311 520770 183369 520804
rect 183403 520770 183461 520804
rect 183495 520770 183553 520804
rect 183587 520770 183645 520804
rect 183679 520770 183737 520804
rect 183771 520770 183829 520804
rect 183863 520770 183921 520804
rect 183955 520770 184013 520804
rect 184047 520770 184105 520804
rect 184139 520770 184197 520804
rect 184231 520770 184289 520804
rect 184323 520770 184381 520804
rect 184415 520770 184473 520804
rect 184507 520770 184565 520804
rect 184599 520770 184657 520804
rect 184691 520770 184749 520804
rect 184783 520770 184841 520804
rect 184875 520770 184933 520804
rect 184967 520770 185025 520804
rect 185059 520770 185117 520804
rect 185151 520770 185209 520804
rect 185243 520770 185301 520804
rect 185335 520770 185393 520804
rect 185427 520770 185485 520804
rect 185519 520770 185577 520804
rect 185611 520770 185669 520804
rect 185703 520770 185761 520804
rect 185795 520770 185853 520804
rect 185887 520770 185945 520804
rect 185979 520770 186037 520804
rect 186071 520770 186129 520804
rect 186163 520770 186221 520804
rect 186255 520770 186313 520804
rect 186347 520770 186405 520804
rect 186439 520770 186497 520804
rect 186531 520770 186589 520804
rect 186623 520770 186681 520804
rect 186715 520770 186773 520804
rect 186807 520770 186865 520804
rect 186899 520770 186957 520804
rect 186991 520770 187049 520804
rect 187083 520770 187141 520804
rect 187175 520770 187233 520804
rect 187267 520770 187325 520804
rect 187359 520770 187417 520804
rect 187451 520770 187480 520804
rect 172225 520707 172467 520770
rect 172225 520673 172243 520707
rect 172277 520673 172415 520707
rect 172449 520673 172467 520707
rect 172225 520620 172467 520673
rect 172501 520709 173570 520770
rect 172501 520675 172519 520709
rect 172553 520675 173519 520709
rect 173553 520675 173570 520709
rect 172501 520661 173570 520675
rect 173605 520709 174674 520770
rect 173605 520675 173623 520709
rect 173657 520675 174623 520709
rect 174657 520675 174674 520709
rect 173605 520661 174674 520675
rect 174801 520676 174859 520770
rect 172225 520546 172329 520620
rect 172225 520512 172275 520546
rect 172309 520512 172329 520546
rect 172363 520552 172383 520586
rect 172417 520552 172467 520586
rect 172363 520478 172467 520552
rect 172818 520546 172886 520661
rect 172818 520512 172835 520546
rect 172869 520512 172886 520546
rect 172818 520495 172886 520512
rect 173182 520582 173252 520597
rect 173182 520548 173199 520582
rect 173233 520548 173252 520582
rect 172225 520431 172467 520478
rect 172225 520397 172243 520431
rect 172277 520397 172415 520431
rect 172449 520397 172467 520431
rect 172225 520336 172467 520397
rect 173182 520347 173252 520548
rect 173922 520546 173990 520661
rect 174801 520642 174813 520676
rect 174847 520642 174859 520676
rect 174893 520709 175962 520770
rect 174893 520675 174911 520709
rect 174945 520675 175911 520709
rect 175945 520675 175962 520709
rect 174893 520661 175962 520675
rect 175997 520709 177066 520770
rect 175997 520675 176015 520709
rect 176049 520675 177015 520709
rect 177049 520675 177066 520709
rect 175997 520661 177066 520675
rect 177101 520709 178170 520770
rect 177101 520675 177119 520709
rect 177153 520675 178119 520709
rect 178153 520675 178170 520709
rect 177101 520661 178170 520675
rect 178205 520709 179274 520770
rect 178205 520675 178223 520709
rect 178257 520675 179223 520709
rect 179257 520675 179274 520709
rect 178205 520661 179274 520675
rect 179309 520709 179827 520770
rect 179309 520675 179327 520709
rect 179361 520675 179775 520709
rect 179809 520675 179827 520709
rect 174801 520625 174859 520642
rect 173922 520512 173939 520546
rect 173973 520512 173990 520546
rect 173922 520495 173990 520512
rect 174286 520582 174356 520597
rect 174286 520548 174303 520582
rect 174337 520548 174356 520582
rect 174286 520347 174356 520548
rect 175210 520546 175278 520661
rect 175210 520512 175227 520546
rect 175261 520512 175278 520546
rect 175210 520495 175278 520512
rect 175574 520582 175644 520597
rect 175574 520548 175591 520582
rect 175625 520548 175644 520582
rect 174801 520458 174859 520493
rect 174801 520424 174813 520458
rect 174847 520424 174859 520458
rect 174801 520365 174859 520424
rect 172225 520302 172243 520336
rect 172277 520302 172415 520336
rect 172449 520302 172467 520336
rect 172225 520260 172467 520302
rect 172501 520336 173570 520347
rect 172501 520302 172519 520336
rect 172553 520302 173519 520336
rect 173553 520302 173570 520336
rect 172501 520260 173570 520302
rect 173605 520336 174674 520347
rect 173605 520302 173623 520336
rect 173657 520302 174623 520336
rect 174657 520302 174674 520336
rect 173605 520260 174674 520302
rect 174801 520331 174813 520365
rect 174847 520331 174859 520365
rect 175574 520347 175644 520548
rect 176314 520546 176382 520661
rect 176314 520512 176331 520546
rect 176365 520512 176382 520546
rect 176314 520495 176382 520512
rect 176678 520582 176748 520597
rect 176678 520548 176695 520582
rect 176729 520548 176748 520582
rect 176678 520347 176748 520548
rect 177418 520546 177486 520661
rect 177418 520512 177435 520546
rect 177469 520512 177486 520546
rect 177418 520495 177486 520512
rect 177782 520582 177852 520597
rect 177782 520548 177799 520582
rect 177833 520548 177852 520582
rect 177782 520347 177852 520548
rect 178522 520546 178590 520661
rect 179309 520616 179827 520675
rect 179953 520676 180011 520770
rect 179953 520642 179965 520676
rect 179999 520642 180011 520676
rect 180045 520709 181114 520770
rect 180045 520675 180063 520709
rect 180097 520675 181063 520709
rect 181097 520675 181114 520709
rect 180045 520661 181114 520675
rect 181149 520709 182218 520770
rect 181149 520675 181167 520709
rect 181201 520675 182167 520709
rect 182201 520675 182218 520709
rect 181149 520661 182218 520675
rect 182253 520709 183322 520770
rect 182253 520675 182271 520709
rect 182305 520675 183271 520709
rect 183305 520675 183322 520709
rect 182253 520661 183322 520675
rect 183357 520709 184426 520770
rect 183357 520675 183375 520709
rect 183409 520675 184375 520709
rect 184409 520675 184426 520709
rect 183357 520661 184426 520675
rect 184461 520709 184979 520770
rect 184461 520675 184479 520709
rect 184513 520675 184927 520709
rect 184961 520675 184979 520709
rect 179953 520625 180011 520642
rect 178522 520512 178539 520546
rect 178573 520512 178590 520546
rect 178522 520495 178590 520512
rect 178886 520582 178956 520597
rect 178886 520548 178903 520582
rect 178937 520548 178956 520582
rect 178886 520347 178956 520548
rect 179309 520546 179551 520616
rect 179309 520512 179387 520546
rect 179421 520512 179497 520546
rect 179531 520512 179551 520546
rect 179585 520548 179605 520582
rect 179639 520548 179715 520582
rect 179749 520548 179827 520582
rect 179585 520478 179827 520548
rect 180362 520546 180430 520661
rect 180362 520512 180379 520546
rect 180413 520512 180430 520546
rect 180362 520495 180430 520512
rect 180726 520582 180796 520597
rect 180726 520548 180743 520582
rect 180777 520548 180796 520582
rect 179309 520438 179827 520478
rect 179309 520404 179327 520438
rect 179361 520404 179775 520438
rect 179809 520404 179827 520438
rect 174801 520260 174859 520331
rect 174893 520336 175962 520347
rect 174893 520302 174911 520336
rect 174945 520302 175911 520336
rect 175945 520302 175962 520336
rect 174893 520260 175962 520302
rect 175997 520336 177066 520347
rect 175997 520302 176015 520336
rect 176049 520302 177015 520336
rect 177049 520302 177066 520336
rect 175997 520260 177066 520302
rect 177101 520336 178170 520347
rect 177101 520302 177119 520336
rect 177153 520302 178119 520336
rect 178153 520302 178170 520336
rect 177101 520260 178170 520302
rect 178205 520336 179274 520347
rect 178205 520302 178223 520336
rect 178257 520302 179223 520336
rect 179257 520302 179274 520336
rect 178205 520260 179274 520302
rect 179309 520336 179827 520404
rect 179309 520302 179327 520336
rect 179361 520302 179775 520336
rect 179809 520302 179827 520336
rect 179309 520260 179827 520302
rect 179953 520458 180011 520493
rect 179953 520424 179965 520458
rect 179999 520424 180011 520458
rect 179953 520365 180011 520424
rect 179953 520331 179965 520365
rect 179999 520331 180011 520365
rect 180726 520347 180796 520548
rect 181466 520546 181534 520661
rect 181466 520512 181483 520546
rect 181517 520512 181534 520546
rect 181466 520495 181534 520512
rect 181830 520582 181900 520597
rect 181830 520548 181847 520582
rect 181881 520548 181900 520582
rect 181830 520347 181900 520548
rect 182570 520546 182638 520661
rect 182570 520512 182587 520546
rect 182621 520512 182638 520546
rect 182570 520495 182638 520512
rect 182934 520582 183004 520597
rect 182934 520548 182951 520582
rect 182985 520548 183004 520582
rect 182934 520347 183004 520548
rect 183674 520546 183742 520661
rect 184461 520616 184979 520675
rect 185105 520676 185163 520770
rect 185105 520642 185117 520676
rect 185151 520642 185163 520676
rect 185197 520709 186266 520770
rect 185197 520675 185215 520709
rect 185249 520675 186215 520709
rect 186249 520675 186266 520709
rect 185197 520661 186266 520675
rect 186301 520709 187003 520770
rect 186301 520675 186319 520709
rect 186353 520675 186951 520709
rect 186985 520675 187003 520709
rect 185105 520625 185163 520642
rect 183674 520512 183691 520546
rect 183725 520512 183742 520546
rect 183674 520495 183742 520512
rect 184038 520582 184108 520597
rect 184038 520548 184055 520582
rect 184089 520548 184108 520582
rect 184038 520347 184108 520548
rect 184461 520546 184703 520616
rect 184461 520512 184539 520546
rect 184573 520512 184649 520546
rect 184683 520512 184703 520546
rect 184737 520548 184757 520582
rect 184791 520548 184867 520582
rect 184901 520548 184979 520582
rect 184737 520478 184979 520548
rect 185514 520546 185582 520661
rect 186301 520616 187003 520675
rect 187221 520707 187463 520770
rect 187221 520673 187239 520707
rect 187273 520673 187411 520707
rect 187445 520673 187463 520707
rect 187221 520620 187463 520673
rect 185514 520512 185531 520546
rect 185565 520512 185582 520546
rect 185514 520495 185582 520512
rect 185878 520582 185948 520597
rect 185878 520548 185895 520582
rect 185929 520548 185948 520582
rect 184461 520438 184979 520478
rect 184461 520404 184479 520438
rect 184513 520404 184927 520438
rect 184961 520404 184979 520438
rect 179953 520260 180011 520331
rect 180045 520336 181114 520347
rect 180045 520302 180063 520336
rect 180097 520302 181063 520336
rect 181097 520302 181114 520336
rect 180045 520260 181114 520302
rect 181149 520336 182218 520347
rect 181149 520302 181167 520336
rect 181201 520302 182167 520336
rect 182201 520302 182218 520336
rect 181149 520260 182218 520302
rect 182253 520336 183322 520347
rect 182253 520302 182271 520336
rect 182305 520302 183271 520336
rect 183305 520302 183322 520336
rect 182253 520260 183322 520302
rect 183357 520336 184426 520347
rect 183357 520302 183375 520336
rect 183409 520302 184375 520336
rect 184409 520302 184426 520336
rect 183357 520260 184426 520302
rect 184461 520336 184979 520404
rect 184461 520302 184479 520336
rect 184513 520302 184927 520336
rect 184961 520302 184979 520336
rect 184461 520260 184979 520302
rect 185105 520458 185163 520493
rect 185105 520424 185117 520458
rect 185151 520424 185163 520458
rect 185105 520365 185163 520424
rect 185105 520331 185117 520365
rect 185151 520331 185163 520365
rect 185878 520347 185948 520548
rect 186301 520546 186631 520616
rect 186301 520512 186379 520546
rect 186413 520512 186478 520546
rect 186512 520512 186577 520546
rect 186611 520512 186631 520546
rect 186665 520548 186685 520582
rect 186719 520548 186788 520582
rect 186822 520548 186891 520582
rect 186925 520548 187003 520582
rect 186665 520478 187003 520548
rect 186301 520438 187003 520478
rect 186301 520404 186319 520438
rect 186353 520404 186951 520438
rect 186985 520404 187003 520438
rect 185105 520260 185163 520331
rect 185197 520336 186266 520347
rect 185197 520302 185215 520336
rect 185249 520302 186215 520336
rect 186249 520302 186266 520336
rect 185197 520260 186266 520302
rect 186301 520336 187003 520404
rect 186301 520302 186319 520336
rect 186353 520302 186951 520336
rect 186985 520302 187003 520336
rect 186301 520260 187003 520302
rect 187221 520552 187271 520586
rect 187305 520552 187325 520586
rect 187221 520478 187325 520552
rect 187359 520546 187463 520620
rect 187359 520512 187379 520546
rect 187413 520512 187463 520546
rect 187221 520431 187463 520478
rect 187221 520397 187239 520431
rect 187273 520397 187411 520431
rect 187445 520397 187463 520431
rect 187221 520336 187463 520397
rect 187221 520302 187239 520336
rect 187273 520302 187411 520336
rect 187445 520302 187463 520336
rect 187221 520260 187463 520302
rect 172208 520226 172237 520260
rect 172271 520226 172329 520260
rect 172363 520226 172421 520260
rect 172455 520226 172513 520260
rect 172547 520226 172605 520260
rect 172639 520226 172697 520260
rect 172731 520226 172789 520260
rect 172823 520226 172881 520260
rect 172915 520226 172973 520260
rect 173007 520226 173065 520260
rect 173099 520226 173157 520260
rect 173191 520226 173249 520260
rect 173283 520226 173341 520260
rect 173375 520226 173433 520260
rect 173467 520226 173525 520260
rect 173559 520226 173617 520260
rect 173651 520226 173709 520260
rect 173743 520226 173801 520260
rect 173835 520226 173893 520260
rect 173927 520226 173985 520260
rect 174019 520226 174077 520260
rect 174111 520226 174169 520260
rect 174203 520226 174261 520260
rect 174295 520226 174353 520260
rect 174387 520226 174445 520260
rect 174479 520226 174537 520260
rect 174571 520226 174629 520260
rect 174663 520226 174721 520260
rect 174755 520226 174813 520260
rect 174847 520226 174905 520260
rect 174939 520226 174997 520260
rect 175031 520226 175089 520260
rect 175123 520226 175181 520260
rect 175215 520226 175273 520260
rect 175307 520226 175365 520260
rect 175399 520226 175457 520260
rect 175491 520226 175549 520260
rect 175583 520226 175641 520260
rect 175675 520226 175733 520260
rect 175767 520226 175825 520260
rect 175859 520226 175917 520260
rect 175951 520226 176009 520260
rect 176043 520226 176101 520260
rect 176135 520226 176193 520260
rect 176227 520226 176285 520260
rect 176319 520226 176377 520260
rect 176411 520226 176469 520260
rect 176503 520226 176561 520260
rect 176595 520226 176653 520260
rect 176687 520226 176745 520260
rect 176779 520226 176837 520260
rect 176871 520226 176929 520260
rect 176963 520226 177021 520260
rect 177055 520226 177113 520260
rect 177147 520226 177205 520260
rect 177239 520226 177297 520260
rect 177331 520226 177389 520260
rect 177423 520226 177481 520260
rect 177515 520226 177573 520260
rect 177607 520226 177665 520260
rect 177699 520226 177757 520260
rect 177791 520226 177849 520260
rect 177883 520226 177941 520260
rect 177975 520226 178033 520260
rect 178067 520226 178125 520260
rect 178159 520226 178217 520260
rect 178251 520226 178309 520260
rect 178343 520226 178401 520260
rect 178435 520226 178493 520260
rect 178527 520226 178585 520260
rect 178619 520226 178677 520260
rect 178711 520226 178769 520260
rect 178803 520226 178861 520260
rect 178895 520226 178953 520260
rect 178987 520226 179045 520260
rect 179079 520226 179137 520260
rect 179171 520226 179229 520260
rect 179263 520226 179321 520260
rect 179355 520226 179413 520260
rect 179447 520226 179505 520260
rect 179539 520226 179597 520260
rect 179631 520226 179689 520260
rect 179723 520226 179781 520260
rect 179815 520226 179873 520260
rect 179907 520226 179965 520260
rect 179999 520226 180057 520260
rect 180091 520226 180149 520260
rect 180183 520226 180241 520260
rect 180275 520226 180333 520260
rect 180367 520226 180425 520260
rect 180459 520226 180517 520260
rect 180551 520226 180609 520260
rect 180643 520226 180701 520260
rect 180735 520226 180793 520260
rect 180827 520226 180885 520260
rect 180919 520226 180977 520260
rect 181011 520226 181069 520260
rect 181103 520226 181161 520260
rect 181195 520226 181253 520260
rect 181287 520226 181345 520260
rect 181379 520226 181437 520260
rect 181471 520226 181529 520260
rect 181563 520226 181621 520260
rect 181655 520226 181713 520260
rect 181747 520226 181805 520260
rect 181839 520226 181897 520260
rect 181931 520226 181989 520260
rect 182023 520226 182081 520260
rect 182115 520226 182173 520260
rect 182207 520226 182265 520260
rect 182299 520226 182357 520260
rect 182391 520226 182449 520260
rect 182483 520226 182541 520260
rect 182575 520226 182633 520260
rect 182667 520226 182725 520260
rect 182759 520226 182817 520260
rect 182851 520226 182909 520260
rect 182943 520226 183001 520260
rect 183035 520226 183093 520260
rect 183127 520226 183185 520260
rect 183219 520226 183277 520260
rect 183311 520226 183369 520260
rect 183403 520226 183461 520260
rect 183495 520226 183553 520260
rect 183587 520226 183645 520260
rect 183679 520226 183737 520260
rect 183771 520226 183829 520260
rect 183863 520226 183921 520260
rect 183955 520226 184013 520260
rect 184047 520226 184105 520260
rect 184139 520226 184197 520260
rect 184231 520226 184289 520260
rect 184323 520226 184381 520260
rect 184415 520226 184473 520260
rect 184507 520226 184565 520260
rect 184599 520226 184657 520260
rect 184691 520226 184749 520260
rect 184783 520226 184841 520260
rect 184875 520226 184933 520260
rect 184967 520226 185025 520260
rect 185059 520226 185117 520260
rect 185151 520226 185209 520260
rect 185243 520226 185301 520260
rect 185335 520226 185393 520260
rect 185427 520226 185485 520260
rect 185519 520226 185577 520260
rect 185611 520226 185669 520260
rect 185703 520226 185761 520260
rect 185795 520226 185853 520260
rect 185887 520226 185945 520260
rect 185979 520226 186037 520260
rect 186071 520226 186129 520260
rect 186163 520226 186221 520260
rect 186255 520226 186313 520260
rect 186347 520226 186405 520260
rect 186439 520226 186497 520260
rect 186531 520226 186589 520260
rect 186623 520226 186681 520260
rect 186715 520226 186773 520260
rect 186807 520226 186865 520260
rect 186899 520226 186957 520260
rect 186991 520226 187049 520260
rect 187083 520226 187141 520260
rect 187175 520226 187233 520260
rect 187267 520226 187325 520260
rect 187359 520226 187417 520260
rect 187451 520226 187480 520260
rect 172225 520184 172467 520226
rect 172225 520150 172243 520184
rect 172277 520150 172415 520184
rect 172449 520150 172467 520184
rect 172225 520089 172467 520150
rect 172501 520184 173570 520226
rect 172501 520150 172519 520184
rect 172553 520150 173519 520184
rect 173553 520150 173570 520184
rect 172501 520139 173570 520150
rect 173605 520184 174674 520226
rect 173605 520150 173623 520184
rect 173657 520150 174623 520184
rect 174657 520150 174674 520184
rect 173605 520139 174674 520150
rect 174709 520184 175778 520226
rect 174709 520150 174727 520184
rect 174761 520150 175727 520184
rect 175761 520150 175778 520184
rect 174709 520139 175778 520150
rect 175813 520184 176882 520226
rect 175813 520150 175831 520184
rect 175865 520150 176831 520184
rect 176865 520150 176882 520184
rect 175813 520139 176882 520150
rect 176917 520184 177251 520226
rect 176917 520150 176935 520184
rect 176969 520150 177199 520184
rect 177233 520150 177251 520184
rect 172225 520055 172243 520089
rect 172277 520055 172415 520089
rect 172449 520055 172467 520089
rect 172225 520008 172467 520055
rect 172225 519940 172275 519974
rect 172309 519940 172329 519974
rect 172225 519866 172329 519940
rect 172363 519934 172467 520008
rect 172363 519900 172383 519934
rect 172417 519900 172467 519934
rect 172818 519974 172886 519991
rect 172818 519940 172835 519974
rect 172869 519940 172886 519974
rect 172225 519813 172467 519866
rect 172818 519825 172886 519940
rect 173182 519938 173252 520139
rect 173182 519904 173199 519938
rect 173233 519904 173252 519938
rect 173182 519889 173252 519904
rect 173922 519974 173990 519991
rect 173922 519940 173939 519974
rect 173973 519940 173990 519974
rect 173922 519825 173990 519940
rect 174286 519938 174356 520139
rect 174286 519904 174303 519938
rect 174337 519904 174356 519938
rect 174286 519889 174356 519904
rect 175026 519974 175094 519991
rect 175026 519940 175043 519974
rect 175077 519940 175094 519974
rect 175026 519825 175094 519940
rect 175390 519938 175460 520139
rect 175390 519904 175407 519938
rect 175441 519904 175460 519938
rect 175390 519889 175460 519904
rect 176130 519974 176198 519991
rect 176130 519940 176147 519974
rect 176181 519940 176198 519974
rect 176130 519825 176198 519940
rect 176494 519938 176564 520139
rect 176917 520082 177251 520150
rect 176917 520048 176935 520082
rect 176969 520048 177199 520082
rect 177233 520048 177251 520082
rect 176917 520008 177251 520048
rect 176494 519904 176511 519938
rect 176545 519904 176564 519938
rect 176494 519889 176564 519904
rect 176917 519940 176937 519974
rect 176971 519940 177067 519974
rect 176917 519870 177067 519940
rect 177101 519938 177251 520008
rect 177377 520155 177435 520226
rect 177377 520121 177389 520155
rect 177423 520121 177435 520155
rect 177469 520184 178538 520226
rect 177469 520150 177487 520184
rect 177521 520150 178487 520184
rect 178521 520150 178538 520184
rect 177469 520139 178538 520150
rect 178573 520184 179642 520226
rect 178573 520150 178591 520184
rect 178625 520150 179591 520184
rect 179625 520150 179642 520184
rect 178573 520139 179642 520150
rect 179677 520184 180746 520226
rect 179677 520150 179695 520184
rect 179729 520150 180695 520184
rect 180729 520150 180746 520184
rect 179677 520139 180746 520150
rect 180781 520184 181850 520226
rect 180781 520150 180799 520184
rect 180833 520150 181799 520184
rect 181833 520150 181850 520184
rect 180781 520139 181850 520150
rect 181885 520184 182403 520226
rect 181885 520150 181903 520184
rect 181937 520150 182351 520184
rect 182385 520150 182403 520184
rect 177377 520062 177435 520121
rect 177377 520028 177389 520062
rect 177423 520028 177435 520062
rect 177377 519993 177435 520028
rect 177101 519904 177197 519938
rect 177231 519904 177251 519938
rect 177786 519974 177854 519991
rect 177786 519940 177803 519974
rect 177837 519940 177854 519974
rect 172225 519779 172243 519813
rect 172277 519779 172415 519813
rect 172449 519779 172467 519813
rect 172225 519716 172467 519779
rect 172501 519811 173570 519825
rect 172501 519777 172519 519811
rect 172553 519777 173519 519811
rect 173553 519777 173570 519811
rect 172501 519716 173570 519777
rect 173605 519811 174674 519825
rect 173605 519777 173623 519811
rect 173657 519777 174623 519811
rect 174657 519777 174674 519811
rect 173605 519716 174674 519777
rect 174709 519811 175778 519825
rect 174709 519777 174727 519811
rect 174761 519777 175727 519811
rect 175761 519777 175778 519811
rect 174709 519716 175778 519777
rect 175813 519811 176882 519825
rect 175813 519777 175831 519811
rect 175865 519777 176831 519811
rect 176865 519777 176882 519811
rect 175813 519716 176882 519777
rect 176917 519818 177251 519870
rect 176917 519784 176935 519818
rect 176969 519784 177199 519818
rect 177233 519784 177251 519818
rect 176917 519716 177251 519784
rect 177377 519844 177435 519861
rect 177377 519810 177389 519844
rect 177423 519810 177435 519844
rect 177786 519825 177854 519940
rect 178150 519938 178220 520139
rect 178150 519904 178167 519938
rect 178201 519904 178220 519938
rect 178150 519889 178220 519904
rect 178890 519974 178958 519991
rect 178890 519940 178907 519974
rect 178941 519940 178958 519974
rect 178890 519825 178958 519940
rect 179254 519938 179324 520139
rect 179254 519904 179271 519938
rect 179305 519904 179324 519938
rect 179254 519889 179324 519904
rect 179994 519974 180062 519991
rect 179994 519940 180011 519974
rect 180045 519940 180062 519974
rect 179994 519825 180062 519940
rect 180358 519938 180428 520139
rect 180358 519904 180375 519938
rect 180409 519904 180428 519938
rect 180358 519889 180428 519904
rect 181098 519974 181166 519991
rect 181098 519940 181115 519974
rect 181149 519940 181166 519974
rect 181098 519825 181166 519940
rect 181462 519938 181532 520139
rect 181885 520082 182403 520150
rect 181885 520048 181903 520082
rect 181937 520048 182351 520082
rect 182385 520048 182403 520082
rect 181885 520008 182403 520048
rect 181462 519904 181479 519938
rect 181513 519904 181532 519938
rect 181462 519889 181532 519904
rect 181885 519940 181963 519974
rect 181997 519940 182073 519974
rect 182107 519940 182127 519974
rect 181885 519870 182127 519940
rect 182161 519938 182403 520008
rect 182529 520155 182587 520226
rect 182529 520121 182541 520155
rect 182575 520121 182587 520155
rect 182621 520184 183690 520226
rect 182621 520150 182639 520184
rect 182673 520150 183639 520184
rect 183673 520150 183690 520184
rect 182621 520139 183690 520150
rect 183725 520184 184794 520226
rect 183725 520150 183743 520184
rect 183777 520150 184743 520184
rect 184777 520150 184794 520184
rect 183725 520139 184794 520150
rect 184829 520184 185898 520226
rect 184829 520150 184847 520184
rect 184881 520150 185847 520184
rect 185881 520150 185898 520184
rect 184829 520139 185898 520150
rect 185933 520184 187002 520226
rect 185933 520150 185951 520184
rect 185985 520150 186951 520184
rect 186985 520150 187002 520184
rect 185933 520139 187002 520150
rect 187221 520184 187463 520226
rect 187221 520150 187239 520184
rect 187273 520150 187411 520184
rect 187445 520150 187463 520184
rect 182529 520062 182587 520121
rect 182529 520028 182541 520062
rect 182575 520028 182587 520062
rect 182529 519993 182587 520028
rect 182161 519904 182181 519938
rect 182215 519904 182291 519938
rect 182325 519904 182403 519938
rect 182938 519974 183006 519991
rect 182938 519940 182955 519974
rect 182989 519940 183006 519974
rect 177377 519716 177435 519810
rect 177469 519811 178538 519825
rect 177469 519777 177487 519811
rect 177521 519777 178487 519811
rect 178521 519777 178538 519811
rect 177469 519716 178538 519777
rect 178573 519811 179642 519825
rect 178573 519777 178591 519811
rect 178625 519777 179591 519811
rect 179625 519777 179642 519811
rect 178573 519716 179642 519777
rect 179677 519811 180746 519825
rect 179677 519777 179695 519811
rect 179729 519777 180695 519811
rect 180729 519777 180746 519811
rect 179677 519716 180746 519777
rect 180781 519811 181850 519825
rect 180781 519777 180799 519811
rect 180833 519777 181799 519811
rect 181833 519777 181850 519811
rect 180781 519716 181850 519777
rect 181885 519811 182403 519870
rect 181885 519777 181903 519811
rect 181937 519777 182351 519811
rect 182385 519777 182403 519811
rect 181885 519716 182403 519777
rect 182529 519844 182587 519861
rect 182529 519810 182541 519844
rect 182575 519810 182587 519844
rect 182938 519825 183006 519940
rect 183302 519938 183372 520139
rect 183302 519904 183319 519938
rect 183353 519904 183372 519938
rect 183302 519889 183372 519904
rect 184042 519974 184110 519991
rect 184042 519940 184059 519974
rect 184093 519940 184110 519974
rect 184042 519825 184110 519940
rect 184406 519938 184476 520139
rect 184406 519904 184423 519938
rect 184457 519904 184476 519938
rect 184406 519889 184476 519904
rect 185146 519974 185214 519991
rect 185146 519940 185163 519974
rect 185197 519940 185214 519974
rect 185146 519825 185214 519940
rect 185510 519938 185580 520139
rect 185510 519904 185527 519938
rect 185561 519904 185580 519938
rect 185510 519889 185580 519904
rect 186250 519974 186318 519991
rect 186250 519940 186267 519974
rect 186301 519940 186318 519974
rect 186250 519825 186318 519940
rect 186614 519938 186684 520139
rect 186614 519904 186631 519938
rect 186665 519904 186684 519938
rect 186614 519889 186684 519904
rect 187221 520089 187463 520150
rect 187221 520055 187239 520089
rect 187273 520055 187411 520089
rect 187445 520055 187463 520089
rect 187221 520008 187463 520055
rect 187221 519934 187325 520008
rect 187221 519900 187271 519934
rect 187305 519900 187325 519934
rect 187359 519940 187379 519974
rect 187413 519940 187463 519974
rect 187359 519866 187463 519940
rect 182529 519716 182587 519810
rect 182621 519811 183690 519825
rect 182621 519777 182639 519811
rect 182673 519777 183639 519811
rect 183673 519777 183690 519811
rect 182621 519716 183690 519777
rect 183725 519811 184794 519825
rect 183725 519777 183743 519811
rect 183777 519777 184743 519811
rect 184777 519777 184794 519811
rect 183725 519716 184794 519777
rect 184829 519811 185898 519825
rect 184829 519777 184847 519811
rect 184881 519777 185847 519811
rect 185881 519777 185898 519811
rect 184829 519716 185898 519777
rect 185933 519811 187002 519825
rect 185933 519777 185951 519811
rect 185985 519777 186951 519811
rect 186985 519777 187002 519811
rect 185933 519716 187002 519777
rect 187221 519813 187463 519866
rect 187221 519779 187239 519813
rect 187273 519779 187411 519813
rect 187445 519779 187463 519813
rect 187221 519716 187463 519779
rect 172208 519682 172237 519716
rect 172271 519682 172329 519716
rect 172363 519682 172421 519716
rect 172455 519682 172513 519716
rect 172547 519682 172605 519716
rect 172639 519682 172697 519716
rect 172731 519682 172789 519716
rect 172823 519682 172881 519716
rect 172915 519682 172973 519716
rect 173007 519682 173065 519716
rect 173099 519682 173157 519716
rect 173191 519682 173249 519716
rect 173283 519682 173341 519716
rect 173375 519682 173433 519716
rect 173467 519682 173525 519716
rect 173559 519682 173617 519716
rect 173651 519682 173709 519716
rect 173743 519682 173801 519716
rect 173835 519682 173893 519716
rect 173927 519682 173985 519716
rect 174019 519682 174077 519716
rect 174111 519682 174169 519716
rect 174203 519682 174261 519716
rect 174295 519682 174353 519716
rect 174387 519682 174445 519716
rect 174479 519682 174537 519716
rect 174571 519682 174629 519716
rect 174663 519682 174721 519716
rect 174755 519682 174813 519716
rect 174847 519682 174905 519716
rect 174939 519682 174997 519716
rect 175031 519682 175089 519716
rect 175123 519682 175181 519716
rect 175215 519682 175273 519716
rect 175307 519682 175365 519716
rect 175399 519682 175457 519716
rect 175491 519682 175549 519716
rect 175583 519682 175641 519716
rect 175675 519682 175733 519716
rect 175767 519682 175825 519716
rect 175859 519682 175917 519716
rect 175951 519682 176009 519716
rect 176043 519682 176101 519716
rect 176135 519682 176193 519716
rect 176227 519682 176285 519716
rect 176319 519682 176377 519716
rect 176411 519682 176469 519716
rect 176503 519682 176561 519716
rect 176595 519682 176653 519716
rect 176687 519682 176745 519716
rect 176779 519682 176837 519716
rect 176871 519682 176929 519716
rect 176963 519682 177021 519716
rect 177055 519682 177113 519716
rect 177147 519682 177205 519716
rect 177239 519682 177297 519716
rect 177331 519682 177389 519716
rect 177423 519682 177481 519716
rect 177515 519682 177573 519716
rect 177607 519682 177665 519716
rect 177699 519682 177757 519716
rect 177791 519682 177849 519716
rect 177883 519682 177941 519716
rect 177975 519682 178033 519716
rect 178067 519682 178125 519716
rect 178159 519682 178217 519716
rect 178251 519682 178309 519716
rect 178343 519682 178401 519716
rect 178435 519682 178493 519716
rect 178527 519682 178585 519716
rect 178619 519682 178677 519716
rect 178711 519682 178769 519716
rect 178803 519682 178861 519716
rect 178895 519682 178953 519716
rect 178987 519682 179045 519716
rect 179079 519682 179137 519716
rect 179171 519682 179229 519716
rect 179263 519682 179321 519716
rect 179355 519682 179413 519716
rect 179447 519682 179505 519716
rect 179539 519682 179597 519716
rect 179631 519682 179689 519716
rect 179723 519682 179781 519716
rect 179815 519682 179873 519716
rect 179907 519682 179965 519716
rect 179999 519682 180057 519716
rect 180091 519682 180149 519716
rect 180183 519682 180241 519716
rect 180275 519682 180333 519716
rect 180367 519682 180425 519716
rect 180459 519682 180517 519716
rect 180551 519682 180609 519716
rect 180643 519682 180701 519716
rect 180735 519682 180793 519716
rect 180827 519682 180885 519716
rect 180919 519682 180977 519716
rect 181011 519682 181069 519716
rect 181103 519682 181161 519716
rect 181195 519682 181253 519716
rect 181287 519682 181345 519716
rect 181379 519682 181437 519716
rect 181471 519682 181529 519716
rect 181563 519682 181621 519716
rect 181655 519682 181713 519716
rect 181747 519682 181805 519716
rect 181839 519682 181897 519716
rect 181931 519682 181989 519716
rect 182023 519682 182081 519716
rect 182115 519682 182173 519716
rect 182207 519682 182265 519716
rect 182299 519682 182357 519716
rect 182391 519682 182449 519716
rect 182483 519682 182541 519716
rect 182575 519682 182633 519716
rect 182667 519682 182725 519716
rect 182759 519682 182817 519716
rect 182851 519682 182909 519716
rect 182943 519682 183001 519716
rect 183035 519682 183093 519716
rect 183127 519682 183185 519716
rect 183219 519682 183277 519716
rect 183311 519682 183369 519716
rect 183403 519682 183461 519716
rect 183495 519682 183553 519716
rect 183587 519682 183645 519716
rect 183679 519682 183737 519716
rect 183771 519682 183829 519716
rect 183863 519682 183921 519716
rect 183955 519682 184013 519716
rect 184047 519682 184105 519716
rect 184139 519682 184197 519716
rect 184231 519682 184289 519716
rect 184323 519682 184381 519716
rect 184415 519682 184473 519716
rect 184507 519682 184565 519716
rect 184599 519682 184657 519716
rect 184691 519682 184749 519716
rect 184783 519682 184841 519716
rect 184875 519682 184933 519716
rect 184967 519682 185025 519716
rect 185059 519682 185117 519716
rect 185151 519682 185209 519716
rect 185243 519682 185301 519716
rect 185335 519682 185393 519716
rect 185427 519682 185485 519716
rect 185519 519682 185577 519716
rect 185611 519682 185669 519716
rect 185703 519682 185761 519716
rect 185795 519682 185853 519716
rect 185887 519682 185945 519716
rect 185979 519682 186037 519716
rect 186071 519682 186129 519716
rect 186163 519682 186221 519716
rect 186255 519682 186313 519716
rect 186347 519682 186405 519716
rect 186439 519682 186497 519716
rect 186531 519682 186589 519716
rect 186623 519682 186681 519716
rect 186715 519682 186773 519716
rect 186807 519682 186865 519716
rect 186899 519682 186957 519716
rect 186991 519682 187049 519716
rect 187083 519682 187141 519716
rect 187175 519682 187233 519716
rect 187267 519682 187325 519716
rect 187359 519682 187417 519716
rect 187451 519682 187480 519716
rect 172225 519619 172467 519682
rect 172225 519585 172243 519619
rect 172277 519585 172415 519619
rect 172449 519585 172467 519619
rect 172225 519532 172467 519585
rect 172501 519621 173570 519682
rect 172501 519587 172519 519621
rect 172553 519587 173519 519621
rect 173553 519587 173570 519621
rect 172501 519573 173570 519587
rect 173605 519621 174674 519682
rect 173605 519587 173623 519621
rect 173657 519587 174623 519621
rect 174657 519587 174674 519621
rect 173605 519573 174674 519587
rect 174801 519588 174859 519682
rect 172225 519458 172329 519532
rect 172225 519424 172275 519458
rect 172309 519424 172329 519458
rect 172363 519464 172383 519498
rect 172417 519464 172467 519498
rect 172363 519390 172467 519464
rect 172818 519458 172886 519573
rect 172818 519424 172835 519458
rect 172869 519424 172886 519458
rect 172818 519407 172886 519424
rect 173182 519494 173252 519509
rect 173182 519460 173199 519494
rect 173233 519460 173252 519494
rect 172225 519343 172467 519390
rect 172225 519309 172243 519343
rect 172277 519309 172415 519343
rect 172449 519309 172467 519343
rect 172225 519248 172467 519309
rect 173182 519259 173252 519460
rect 173922 519458 173990 519573
rect 174801 519554 174813 519588
rect 174847 519554 174859 519588
rect 174893 519621 175962 519682
rect 174893 519587 174911 519621
rect 174945 519587 175911 519621
rect 175945 519587 175962 519621
rect 174893 519573 175962 519587
rect 175997 519621 177066 519682
rect 175997 519587 176015 519621
rect 176049 519587 177015 519621
rect 177049 519587 177066 519621
rect 175997 519573 177066 519587
rect 177101 519621 178170 519682
rect 177101 519587 177119 519621
rect 177153 519587 178119 519621
rect 178153 519587 178170 519621
rect 177101 519573 178170 519587
rect 178205 519621 179274 519682
rect 178205 519587 178223 519621
rect 178257 519587 179223 519621
rect 179257 519587 179274 519621
rect 178205 519573 179274 519587
rect 179309 519621 179827 519682
rect 179309 519587 179327 519621
rect 179361 519587 179775 519621
rect 179809 519587 179827 519621
rect 174801 519537 174859 519554
rect 173922 519424 173939 519458
rect 173973 519424 173990 519458
rect 173922 519407 173990 519424
rect 174286 519494 174356 519509
rect 174286 519460 174303 519494
rect 174337 519460 174356 519494
rect 174286 519259 174356 519460
rect 175210 519458 175278 519573
rect 175210 519424 175227 519458
rect 175261 519424 175278 519458
rect 175210 519407 175278 519424
rect 175574 519494 175644 519509
rect 175574 519460 175591 519494
rect 175625 519460 175644 519494
rect 174801 519370 174859 519405
rect 174801 519336 174813 519370
rect 174847 519336 174859 519370
rect 174801 519277 174859 519336
rect 172225 519214 172243 519248
rect 172277 519214 172415 519248
rect 172449 519214 172467 519248
rect 172225 519172 172467 519214
rect 172501 519248 173570 519259
rect 172501 519214 172519 519248
rect 172553 519214 173519 519248
rect 173553 519214 173570 519248
rect 172501 519172 173570 519214
rect 173605 519248 174674 519259
rect 173605 519214 173623 519248
rect 173657 519214 174623 519248
rect 174657 519214 174674 519248
rect 173605 519172 174674 519214
rect 174801 519243 174813 519277
rect 174847 519243 174859 519277
rect 175574 519259 175644 519460
rect 176314 519458 176382 519573
rect 176314 519424 176331 519458
rect 176365 519424 176382 519458
rect 176314 519407 176382 519424
rect 176678 519494 176748 519509
rect 176678 519460 176695 519494
rect 176729 519460 176748 519494
rect 176678 519259 176748 519460
rect 177418 519458 177486 519573
rect 177418 519424 177435 519458
rect 177469 519424 177486 519458
rect 177418 519407 177486 519424
rect 177782 519494 177852 519509
rect 177782 519460 177799 519494
rect 177833 519460 177852 519494
rect 177782 519259 177852 519460
rect 178522 519458 178590 519573
rect 179309 519528 179827 519587
rect 179953 519588 180011 519682
rect 179953 519554 179965 519588
rect 179999 519554 180011 519588
rect 180045 519621 181114 519682
rect 180045 519587 180063 519621
rect 180097 519587 181063 519621
rect 181097 519587 181114 519621
rect 180045 519573 181114 519587
rect 181149 519621 182218 519682
rect 181149 519587 181167 519621
rect 181201 519587 182167 519621
rect 182201 519587 182218 519621
rect 181149 519573 182218 519587
rect 182253 519621 183322 519682
rect 182253 519587 182271 519621
rect 182305 519587 183271 519621
rect 183305 519587 183322 519621
rect 182253 519573 183322 519587
rect 183357 519621 184426 519682
rect 183357 519587 183375 519621
rect 183409 519587 184375 519621
rect 184409 519587 184426 519621
rect 183357 519573 184426 519587
rect 184461 519621 184979 519682
rect 184461 519587 184479 519621
rect 184513 519587 184927 519621
rect 184961 519587 184979 519621
rect 179953 519537 180011 519554
rect 178522 519424 178539 519458
rect 178573 519424 178590 519458
rect 178522 519407 178590 519424
rect 178886 519494 178956 519509
rect 178886 519460 178903 519494
rect 178937 519460 178956 519494
rect 178886 519259 178956 519460
rect 179309 519458 179551 519528
rect 179309 519424 179387 519458
rect 179421 519424 179497 519458
rect 179531 519424 179551 519458
rect 179585 519460 179605 519494
rect 179639 519460 179715 519494
rect 179749 519460 179827 519494
rect 179585 519390 179827 519460
rect 180362 519458 180430 519573
rect 180362 519424 180379 519458
rect 180413 519424 180430 519458
rect 180362 519407 180430 519424
rect 180726 519494 180796 519509
rect 180726 519460 180743 519494
rect 180777 519460 180796 519494
rect 179309 519350 179827 519390
rect 179309 519316 179327 519350
rect 179361 519316 179775 519350
rect 179809 519316 179827 519350
rect 174801 519172 174859 519243
rect 174893 519248 175962 519259
rect 174893 519214 174911 519248
rect 174945 519214 175911 519248
rect 175945 519214 175962 519248
rect 174893 519172 175962 519214
rect 175997 519248 177066 519259
rect 175997 519214 176015 519248
rect 176049 519214 177015 519248
rect 177049 519214 177066 519248
rect 175997 519172 177066 519214
rect 177101 519248 178170 519259
rect 177101 519214 177119 519248
rect 177153 519214 178119 519248
rect 178153 519214 178170 519248
rect 177101 519172 178170 519214
rect 178205 519248 179274 519259
rect 178205 519214 178223 519248
rect 178257 519214 179223 519248
rect 179257 519214 179274 519248
rect 178205 519172 179274 519214
rect 179309 519248 179827 519316
rect 179309 519214 179327 519248
rect 179361 519214 179775 519248
rect 179809 519214 179827 519248
rect 179309 519172 179827 519214
rect 179953 519370 180011 519405
rect 179953 519336 179965 519370
rect 179999 519336 180011 519370
rect 179953 519277 180011 519336
rect 179953 519243 179965 519277
rect 179999 519243 180011 519277
rect 180726 519259 180796 519460
rect 181466 519458 181534 519573
rect 181466 519424 181483 519458
rect 181517 519424 181534 519458
rect 181466 519407 181534 519424
rect 181830 519494 181900 519509
rect 181830 519460 181847 519494
rect 181881 519460 181900 519494
rect 181830 519259 181900 519460
rect 182570 519458 182638 519573
rect 182570 519424 182587 519458
rect 182621 519424 182638 519458
rect 182570 519407 182638 519424
rect 182934 519494 183004 519509
rect 182934 519460 182951 519494
rect 182985 519460 183004 519494
rect 182934 519259 183004 519460
rect 183674 519458 183742 519573
rect 184461 519528 184979 519587
rect 185105 519588 185163 519682
rect 185105 519554 185117 519588
rect 185151 519554 185163 519588
rect 185197 519621 186266 519682
rect 185197 519587 185215 519621
rect 185249 519587 186215 519621
rect 186249 519587 186266 519621
rect 185197 519573 186266 519587
rect 186301 519621 187003 519682
rect 186301 519587 186319 519621
rect 186353 519587 186951 519621
rect 186985 519587 187003 519621
rect 185105 519537 185163 519554
rect 183674 519424 183691 519458
rect 183725 519424 183742 519458
rect 183674 519407 183742 519424
rect 184038 519494 184108 519509
rect 184038 519460 184055 519494
rect 184089 519460 184108 519494
rect 184038 519259 184108 519460
rect 184461 519458 184703 519528
rect 184461 519424 184539 519458
rect 184573 519424 184649 519458
rect 184683 519424 184703 519458
rect 184737 519460 184757 519494
rect 184791 519460 184867 519494
rect 184901 519460 184979 519494
rect 184737 519390 184979 519460
rect 185514 519458 185582 519573
rect 186301 519528 187003 519587
rect 187221 519619 187463 519682
rect 187221 519585 187239 519619
rect 187273 519585 187411 519619
rect 187445 519585 187463 519619
rect 187221 519532 187463 519585
rect 185514 519424 185531 519458
rect 185565 519424 185582 519458
rect 185514 519407 185582 519424
rect 185878 519494 185948 519509
rect 185878 519460 185895 519494
rect 185929 519460 185948 519494
rect 184461 519350 184979 519390
rect 184461 519316 184479 519350
rect 184513 519316 184927 519350
rect 184961 519316 184979 519350
rect 179953 519172 180011 519243
rect 180045 519248 181114 519259
rect 180045 519214 180063 519248
rect 180097 519214 181063 519248
rect 181097 519214 181114 519248
rect 180045 519172 181114 519214
rect 181149 519248 182218 519259
rect 181149 519214 181167 519248
rect 181201 519214 182167 519248
rect 182201 519214 182218 519248
rect 181149 519172 182218 519214
rect 182253 519248 183322 519259
rect 182253 519214 182271 519248
rect 182305 519214 183271 519248
rect 183305 519214 183322 519248
rect 182253 519172 183322 519214
rect 183357 519248 184426 519259
rect 183357 519214 183375 519248
rect 183409 519214 184375 519248
rect 184409 519214 184426 519248
rect 183357 519172 184426 519214
rect 184461 519248 184979 519316
rect 184461 519214 184479 519248
rect 184513 519214 184927 519248
rect 184961 519214 184979 519248
rect 184461 519172 184979 519214
rect 185105 519370 185163 519405
rect 185105 519336 185117 519370
rect 185151 519336 185163 519370
rect 185105 519277 185163 519336
rect 185105 519243 185117 519277
rect 185151 519243 185163 519277
rect 185878 519259 185948 519460
rect 186301 519458 186631 519528
rect 186301 519424 186379 519458
rect 186413 519424 186478 519458
rect 186512 519424 186577 519458
rect 186611 519424 186631 519458
rect 186665 519460 186685 519494
rect 186719 519460 186788 519494
rect 186822 519460 186891 519494
rect 186925 519460 187003 519494
rect 186665 519390 187003 519460
rect 186301 519350 187003 519390
rect 186301 519316 186319 519350
rect 186353 519316 186951 519350
rect 186985 519316 187003 519350
rect 185105 519172 185163 519243
rect 185197 519248 186266 519259
rect 185197 519214 185215 519248
rect 185249 519214 186215 519248
rect 186249 519214 186266 519248
rect 185197 519172 186266 519214
rect 186301 519248 187003 519316
rect 186301 519214 186319 519248
rect 186353 519214 186951 519248
rect 186985 519214 187003 519248
rect 186301 519172 187003 519214
rect 187221 519464 187271 519498
rect 187305 519464 187325 519498
rect 187221 519390 187325 519464
rect 187359 519458 187463 519532
rect 187359 519424 187379 519458
rect 187413 519424 187463 519458
rect 187221 519343 187463 519390
rect 187221 519309 187239 519343
rect 187273 519309 187411 519343
rect 187445 519309 187463 519343
rect 187221 519248 187463 519309
rect 187221 519214 187239 519248
rect 187273 519214 187411 519248
rect 187445 519214 187463 519248
rect 187221 519172 187463 519214
rect 172208 519138 172237 519172
rect 172271 519138 172329 519172
rect 172363 519138 172421 519172
rect 172455 519138 172513 519172
rect 172547 519138 172605 519172
rect 172639 519138 172697 519172
rect 172731 519138 172789 519172
rect 172823 519138 172881 519172
rect 172915 519138 172973 519172
rect 173007 519138 173065 519172
rect 173099 519138 173157 519172
rect 173191 519138 173249 519172
rect 173283 519138 173341 519172
rect 173375 519138 173433 519172
rect 173467 519138 173525 519172
rect 173559 519138 173617 519172
rect 173651 519138 173709 519172
rect 173743 519138 173801 519172
rect 173835 519138 173893 519172
rect 173927 519138 173985 519172
rect 174019 519138 174077 519172
rect 174111 519138 174169 519172
rect 174203 519138 174261 519172
rect 174295 519138 174353 519172
rect 174387 519138 174445 519172
rect 174479 519138 174537 519172
rect 174571 519138 174629 519172
rect 174663 519138 174721 519172
rect 174755 519138 174813 519172
rect 174847 519138 174905 519172
rect 174939 519138 174997 519172
rect 175031 519138 175089 519172
rect 175123 519138 175181 519172
rect 175215 519138 175273 519172
rect 175307 519138 175365 519172
rect 175399 519138 175457 519172
rect 175491 519138 175549 519172
rect 175583 519138 175641 519172
rect 175675 519138 175733 519172
rect 175767 519138 175825 519172
rect 175859 519138 175917 519172
rect 175951 519138 176009 519172
rect 176043 519138 176101 519172
rect 176135 519138 176193 519172
rect 176227 519138 176285 519172
rect 176319 519138 176377 519172
rect 176411 519138 176469 519172
rect 176503 519138 176561 519172
rect 176595 519138 176653 519172
rect 176687 519138 176745 519172
rect 176779 519138 176837 519172
rect 176871 519138 176929 519172
rect 176963 519138 177021 519172
rect 177055 519138 177113 519172
rect 177147 519138 177205 519172
rect 177239 519138 177297 519172
rect 177331 519138 177389 519172
rect 177423 519138 177481 519172
rect 177515 519138 177573 519172
rect 177607 519138 177665 519172
rect 177699 519138 177757 519172
rect 177791 519138 177849 519172
rect 177883 519138 177941 519172
rect 177975 519138 178033 519172
rect 178067 519138 178125 519172
rect 178159 519138 178217 519172
rect 178251 519138 178309 519172
rect 178343 519138 178401 519172
rect 178435 519138 178493 519172
rect 178527 519138 178585 519172
rect 178619 519138 178677 519172
rect 178711 519138 178769 519172
rect 178803 519138 178861 519172
rect 178895 519138 178953 519172
rect 178987 519138 179045 519172
rect 179079 519138 179137 519172
rect 179171 519138 179229 519172
rect 179263 519138 179321 519172
rect 179355 519138 179413 519172
rect 179447 519138 179505 519172
rect 179539 519138 179597 519172
rect 179631 519138 179689 519172
rect 179723 519138 179781 519172
rect 179815 519138 179873 519172
rect 179907 519138 179965 519172
rect 179999 519138 180057 519172
rect 180091 519138 180149 519172
rect 180183 519138 180241 519172
rect 180275 519138 180333 519172
rect 180367 519138 180425 519172
rect 180459 519138 180517 519172
rect 180551 519138 180609 519172
rect 180643 519138 180701 519172
rect 180735 519138 180793 519172
rect 180827 519138 180885 519172
rect 180919 519138 180977 519172
rect 181011 519138 181069 519172
rect 181103 519138 181161 519172
rect 181195 519138 181253 519172
rect 181287 519138 181345 519172
rect 181379 519138 181437 519172
rect 181471 519138 181529 519172
rect 181563 519138 181621 519172
rect 181655 519138 181713 519172
rect 181747 519138 181805 519172
rect 181839 519138 181897 519172
rect 181931 519138 181989 519172
rect 182023 519138 182081 519172
rect 182115 519138 182173 519172
rect 182207 519138 182265 519172
rect 182299 519138 182357 519172
rect 182391 519138 182449 519172
rect 182483 519138 182541 519172
rect 182575 519138 182633 519172
rect 182667 519138 182725 519172
rect 182759 519138 182817 519172
rect 182851 519138 182909 519172
rect 182943 519138 183001 519172
rect 183035 519138 183093 519172
rect 183127 519138 183185 519172
rect 183219 519138 183277 519172
rect 183311 519138 183369 519172
rect 183403 519138 183461 519172
rect 183495 519138 183553 519172
rect 183587 519138 183645 519172
rect 183679 519138 183737 519172
rect 183771 519138 183829 519172
rect 183863 519138 183921 519172
rect 183955 519138 184013 519172
rect 184047 519138 184105 519172
rect 184139 519138 184197 519172
rect 184231 519138 184289 519172
rect 184323 519138 184381 519172
rect 184415 519138 184473 519172
rect 184507 519138 184565 519172
rect 184599 519138 184657 519172
rect 184691 519138 184749 519172
rect 184783 519138 184841 519172
rect 184875 519138 184933 519172
rect 184967 519138 185025 519172
rect 185059 519138 185117 519172
rect 185151 519138 185209 519172
rect 185243 519138 185301 519172
rect 185335 519138 185393 519172
rect 185427 519138 185485 519172
rect 185519 519138 185577 519172
rect 185611 519138 185669 519172
rect 185703 519138 185761 519172
rect 185795 519138 185853 519172
rect 185887 519138 185945 519172
rect 185979 519138 186037 519172
rect 186071 519138 186129 519172
rect 186163 519138 186221 519172
rect 186255 519138 186313 519172
rect 186347 519138 186405 519172
rect 186439 519138 186497 519172
rect 186531 519138 186589 519172
rect 186623 519138 186681 519172
rect 186715 519138 186773 519172
rect 186807 519138 186865 519172
rect 186899 519138 186957 519172
rect 186991 519138 187049 519172
rect 187083 519138 187141 519172
rect 187175 519138 187233 519172
rect 187267 519138 187325 519172
rect 187359 519138 187417 519172
rect 187451 519138 187480 519172
rect 172225 519096 172467 519138
rect 172225 519062 172243 519096
rect 172277 519062 172415 519096
rect 172449 519062 172467 519096
rect 172225 519001 172467 519062
rect 172501 519096 173570 519138
rect 172501 519062 172519 519096
rect 172553 519062 173519 519096
rect 173553 519062 173570 519096
rect 172501 519051 173570 519062
rect 173605 519096 174674 519138
rect 173605 519062 173623 519096
rect 173657 519062 174623 519096
rect 174657 519062 174674 519096
rect 173605 519051 174674 519062
rect 174709 519096 175778 519138
rect 174709 519062 174727 519096
rect 174761 519062 175727 519096
rect 175761 519062 175778 519096
rect 174709 519051 175778 519062
rect 175813 519096 176882 519138
rect 175813 519062 175831 519096
rect 175865 519062 176831 519096
rect 176865 519062 176882 519096
rect 175813 519051 176882 519062
rect 176917 519096 177251 519138
rect 176917 519062 176935 519096
rect 176969 519062 177199 519096
rect 177233 519062 177251 519096
rect 172225 518967 172243 519001
rect 172277 518967 172415 519001
rect 172449 518967 172467 519001
rect 172225 518920 172467 518967
rect 172225 518852 172275 518886
rect 172309 518852 172329 518886
rect 172225 518778 172329 518852
rect 172363 518846 172467 518920
rect 172363 518812 172383 518846
rect 172417 518812 172467 518846
rect 172818 518886 172886 518903
rect 172818 518852 172835 518886
rect 172869 518852 172886 518886
rect 172225 518725 172467 518778
rect 172818 518737 172886 518852
rect 173182 518850 173252 519051
rect 173182 518816 173199 518850
rect 173233 518816 173252 518850
rect 173182 518801 173252 518816
rect 173922 518886 173990 518903
rect 173922 518852 173939 518886
rect 173973 518852 173990 518886
rect 173922 518737 173990 518852
rect 174286 518850 174356 519051
rect 174286 518816 174303 518850
rect 174337 518816 174356 518850
rect 174286 518801 174356 518816
rect 175026 518886 175094 518903
rect 175026 518852 175043 518886
rect 175077 518852 175094 518886
rect 175026 518737 175094 518852
rect 175390 518850 175460 519051
rect 175390 518816 175407 518850
rect 175441 518816 175460 518850
rect 175390 518801 175460 518816
rect 176130 518886 176198 518903
rect 176130 518852 176147 518886
rect 176181 518852 176198 518886
rect 176130 518737 176198 518852
rect 176494 518850 176564 519051
rect 176917 518994 177251 519062
rect 176917 518960 176935 518994
rect 176969 518960 177199 518994
rect 177233 518960 177251 518994
rect 176917 518920 177251 518960
rect 176494 518816 176511 518850
rect 176545 518816 176564 518850
rect 176494 518801 176564 518816
rect 176917 518852 176937 518886
rect 176971 518852 177067 518886
rect 176917 518782 177067 518852
rect 177101 518850 177251 518920
rect 177377 519067 177435 519138
rect 177377 519033 177389 519067
rect 177423 519033 177435 519067
rect 177469 519096 178538 519138
rect 177469 519062 177487 519096
rect 177521 519062 178487 519096
rect 178521 519062 178538 519096
rect 177469 519051 178538 519062
rect 178573 519096 179642 519138
rect 178573 519062 178591 519096
rect 178625 519062 179591 519096
rect 179625 519062 179642 519096
rect 178573 519051 179642 519062
rect 179677 519096 180746 519138
rect 179677 519062 179695 519096
rect 179729 519062 180695 519096
rect 180729 519062 180746 519096
rect 179677 519051 180746 519062
rect 180781 519096 181850 519138
rect 180781 519062 180799 519096
rect 180833 519062 181799 519096
rect 181833 519062 181850 519096
rect 180781 519051 181850 519062
rect 181885 519096 182403 519138
rect 181885 519062 181903 519096
rect 181937 519062 182351 519096
rect 182385 519062 182403 519096
rect 177377 518974 177435 519033
rect 177377 518940 177389 518974
rect 177423 518940 177435 518974
rect 177377 518905 177435 518940
rect 177101 518816 177197 518850
rect 177231 518816 177251 518850
rect 177786 518886 177854 518903
rect 177786 518852 177803 518886
rect 177837 518852 177854 518886
rect 172225 518691 172243 518725
rect 172277 518691 172415 518725
rect 172449 518691 172467 518725
rect 172225 518628 172467 518691
rect 172501 518723 173570 518737
rect 172501 518689 172519 518723
rect 172553 518689 173519 518723
rect 173553 518689 173570 518723
rect 172501 518628 173570 518689
rect 173605 518723 174674 518737
rect 173605 518689 173623 518723
rect 173657 518689 174623 518723
rect 174657 518689 174674 518723
rect 173605 518628 174674 518689
rect 174709 518723 175778 518737
rect 174709 518689 174727 518723
rect 174761 518689 175727 518723
rect 175761 518689 175778 518723
rect 174709 518628 175778 518689
rect 175813 518723 176882 518737
rect 175813 518689 175831 518723
rect 175865 518689 176831 518723
rect 176865 518689 176882 518723
rect 175813 518628 176882 518689
rect 176917 518730 177251 518782
rect 176917 518696 176935 518730
rect 176969 518696 177199 518730
rect 177233 518696 177251 518730
rect 176917 518628 177251 518696
rect 177377 518756 177435 518773
rect 177377 518722 177389 518756
rect 177423 518722 177435 518756
rect 177786 518737 177854 518852
rect 178150 518850 178220 519051
rect 178150 518816 178167 518850
rect 178201 518816 178220 518850
rect 178150 518801 178220 518816
rect 178890 518886 178958 518903
rect 178890 518852 178907 518886
rect 178941 518852 178958 518886
rect 178890 518737 178958 518852
rect 179254 518850 179324 519051
rect 179254 518816 179271 518850
rect 179305 518816 179324 518850
rect 179254 518801 179324 518816
rect 179994 518886 180062 518903
rect 179994 518852 180011 518886
rect 180045 518852 180062 518886
rect 179994 518737 180062 518852
rect 180358 518850 180428 519051
rect 180358 518816 180375 518850
rect 180409 518816 180428 518850
rect 180358 518801 180428 518816
rect 181098 518886 181166 518903
rect 181098 518852 181115 518886
rect 181149 518852 181166 518886
rect 181098 518737 181166 518852
rect 181462 518850 181532 519051
rect 181885 518994 182403 519062
rect 181885 518960 181903 518994
rect 181937 518960 182351 518994
rect 182385 518960 182403 518994
rect 181885 518920 182403 518960
rect 181462 518816 181479 518850
rect 181513 518816 181532 518850
rect 181462 518801 181532 518816
rect 181885 518852 181963 518886
rect 181997 518852 182073 518886
rect 182107 518852 182127 518886
rect 181885 518782 182127 518852
rect 182161 518850 182403 518920
rect 182529 519067 182587 519138
rect 182529 519033 182541 519067
rect 182575 519033 182587 519067
rect 182621 519096 183690 519138
rect 182621 519062 182639 519096
rect 182673 519062 183639 519096
rect 183673 519062 183690 519096
rect 182621 519051 183690 519062
rect 183725 519096 184794 519138
rect 183725 519062 183743 519096
rect 183777 519062 184743 519096
rect 184777 519062 184794 519096
rect 183725 519051 184794 519062
rect 184829 519096 185898 519138
rect 184829 519062 184847 519096
rect 184881 519062 185847 519096
rect 185881 519062 185898 519096
rect 184829 519051 185898 519062
rect 185933 519096 187002 519138
rect 185933 519062 185951 519096
rect 185985 519062 186951 519096
rect 186985 519062 187002 519096
rect 185933 519051 187002 519062
rect 187221 519096 187463 519138
rect 187221 519062 187239 519096
rect 187273 519062 187411 519096
rect 187445 519062 187463 519096
rect 182529 518974 182587 519033
rect 182529 518940 182541 518974
rect 182575 518940 182587 518974
rect 182529 518905 182587 518940
rect 182161 518816 182181 518850
rect 182215 518816 182291 518850
rect 182325 518816 182403 518850
rect 182938 518886 183006 518903
rect 182938 518852 182955 518886
rect 182989 518852 183006 518886
rect 177377 518628 177435 518722
rect 177469 518723 178538 518737
rect 177469 518689 177487 518723
rect 177521 518689 178487 518723
rect 178521 518689 178538 518723
rect 177469 518628 178538 518689
rect 178573 518723 179642 518737
rect 178573 518689 178591 518723
rect 178625 518689 179591 518723
rect 179625 518689 179642 518723
rect 178573 518628 179642 518689
rect 179677 518723 180746 518737
rect 179677 518689 179695 518723
rect 179729 518689 180695 518723
rect 180729 518689 180746 518723
rect 179677 518628 180746 518689
rect 180781 518723 181850 518737
rect 180781 518689 180799 518723
rect 180833 518689 181799 518723
rect 181833 518689 181850 518723
rect 180781 518628 181850 518689
rect 181885 518723 182403 518782
rect 181885 518689 181903 518723
rect 181937 518689 182351 518723
rect 182385 518689 182403 518723
rect 181885 518628 182403 518689
rect 182529 518756 182587 518773
rect 182529 518722 182541 518756
rect 182575 518722 182587 518756
rect 182938 518737 183006 518852
rect 183302 518850 183372 519051
rect 183302 518816 183319 518850
rect 183353 518816 183372 518850
rect 183302 518801 183372 518816
rect 184042 518886 184110 518903
rect 184042 518852 184059 518886
rect 184093 518852 184110 518886
rect 184042 518737 184110 518852
rect 184406 518850 184476 519051
rect 184406 518816 184423 518850
rect 184457 518816 184476 518850
rect 184406 518801 184476 518816
rect 185146 518886 185214 518903
rect 185146 518852 185163 518886
rect 185197 518852 185214 518886
rect 185146 518737 185214 518852
rect 185510 518850 185580 519051
rect 185510 518816 185527 518850
rect 185561 518816 185580 518850
rect 185510 518801 185580 518816
rect 186250 518886 186318 518903
rect 186250 518852 186267 518886
rect 186301 518852 186318 518886
rect 186250 518737 186318 518852
rect 186614 518850 186684 519051
rect 186614 518816 186631 518850
rect 186665 518816 186684 518850
rect 186614 518801 186684 518816
rect 187221 519001 187463 519062
rect 187221 518967 187239 519001
rect 187273 518967 187411 519001
rect 187445 518967 187463 519001
rect 187221 518920 187463 518967
rect 187221 518846 187325 518920
rect 187221 518812 187271 518846
rect 187305 518812 187325 518846
rect 187359 518852 187379 518886
rect 187413 518852 187463 518886
rect 187359 518778 187463 518852
rect 182529 518628 182587 518722
rect 182621 518723 183690 518737
rect 182621 518689 182639 518723
rect 182673 518689 183639 518723
rect 183673 518689 183690 518723
rect 182621 518628 183690 518689
rect 183725 518723 184794 518737
rect 183725 518689 183743 518723
rect 183777 518689 184743 518723
rect 184777 518689 184794 518723
rect 183725 518628 184794 518689
rect 184829 518723 185898 518737
rect 184829 518689 184847 518723
rect 184881 518689 185847 518723
rect 185881 518689 185898 518723
rect 184829 518628 185898 518689
rect 185933 518723 187002 518737
rect 185933 518689 185951 518723
rect 185985 518689 186951 518723
rect 186985 518689 187002 518723
rect 185933 518628 187002 518689
rect 187221 518725 187463 518778
rect 187221 518691 187239 518725
rect 187273 518691 187411 518725
rect 187445 518691 187463 518725
rect 187221 518628 187463 518691
rect 172208 518594 172237 518628
rect 172271 518594 172329 518628
rect 172363 518594 172421 518628
rect 172455 518594 172513 518628
rect 172547 518594 172605 518628
rect 172639 518594 172697 518628
rect 172731 518594 172789 518628
rect 172823 518594 172881 518628
rect 172915 518594 172973 518628
rect 173007 518594 173065 518628
rect 173099 518594 173157 518628
rect 173191 518594 173249 518628
rect 173283 518594 173341 518628
rect 173375 518594 173433 518628
rect 173467 518594 173525 518628
rect 173559 518594 173617 518628
rect 173651 518594 173709 518628
rect 173743 518594 173801 518628
rect 173835 518594 173893 518628
rect 173927 518594 173985 518628
rect 174019 518594 174077 518628
rect 174111 518594 174169 518628
rect 174203 518594 174261 518628
rect 174295 518594 174353 518628
rect 174387 518594 174445 518628
rect 174479 518594 174537 518628
rect 174571 518594 174629 518628
rect 174663 518594 174721 518628
rect 174755 518594 174813 518628
rect 174847 518594 174905 518628
rect 174939 518594 174997 518628
rect 175031 518594 175089 518628
rect 175123 518594 175181 518628
rect 175215 518594 175273 518628
rect 175307 518594 175365 518628
rect 175399 518594 175457 518628
rect 175491 518594 175549 518628
rect 175583 518594 175641 518628
rect 175675 518594 175733 518628
rect 175767 518594 175825 518628
rect 175859 518594 175917 518628
rect 175951 518594 176009 518628
rect 176043 518594 176101 518628
rect 176135 518594 176193 518628
rect 176227 518594 176285 518628
rect 176319 518594 176377 518628
rect 176411 518594 176469 518628
rect 176503 518594 176561 518628
rect 176595 518594 176653 518628
rect 176687 518594 176745 518628
rect 176779 518594 176837 518628
rect 176871 518594 176929 518628
rect 176963 518594 177021 518628
rect 177055 518594 177113 518628
rect 177147 518594 177205 518628
rect 177239 518594 177297 518628
rect 177331 518594 177389 518628
rect 177423 518594 177481 518628
rect 177515 518594 177573 518628
rect 177607 518594 177665 518628
rect 177699 518594 177757 518628
rect 177791 518594 177849 518628
rect 177883 518594 177941 518628
rect 177975 518594 178033 518628
rect 178067 518594 178125 518628
rect 178159 518594 178217 518628
rect 178251 518594 178309 518628
rect 178343 518594 178401 518628
rect 178435 518594 178493 518628
rect 178527 518594 178585 518628
rect 178619 518594 178677 518628
rect 178711 518594 178769 518628
rect 178803 518594 178861 518628
rect 178895 518594 178953 518628
rect 178987 518594 179045 518628
rect 179079 518594 179137 518628
rect 179171 518594 179229 518628
rect 179263 518594 179321 518628
rect 179355 518594 179413 518628
rect 179447 518594 179505 518628
rect 179539 518594 179597 518628
rect 179631 518594 179689 518628
rect 179723 518594 179781 518628
rect 179815 518594 179873 518628
rect 179907 518594 179965 518628
rect 179999 518594 180057 518628
rect 180091 518594 180149 518628
rect 180183 518594 180241 518628
rect 180275 518594 180333 518628
rect 180367 518594 180425 518628
rect 180459 518594 180517 518628
rect 180551 518594 180609 518628
rect 180643 518594 180701 518628
rect 180735 518594 180793 518628
rect 180827 518594 180885 518628
rect 180919 518594 180977 518628
rect 181011 518594 181069 518628
rect 181103 518594 181161 518628
rect 181195 518594 181253 518628
rect 181287 518594 181345 518628
rect 181379 518594 181437 518628
rect 181471 518594 181529 518628
rect 181563 518594 181621 518628
rect 181655 518594 181713 518628
rect 181747 518594 181805 518628
rect 181839 518594 181897 518628
rect 181931 518594 181989 518628
rect 182023 518594 182081 518628
rect 182115 518594 182173 518628
rect 182207 518594 182265 518628
rect 182299 518594 182357 518628
rect 182391 518594 182449 518628
rect 182483 518594 182541 518628
rect 182575 518594 182633 518628
rect 182667 518594 182725 518628
rect 182759 518594 182817 518628
rect 182851 518594 182909 518628
rect 182943 518594 183001 518628
rect 183035 518594 183093 518628
rect 183127 518594 183185 518628
rect 183219 518594 183277 518628
rect 183311 518594 183369 518628
rect 183403 518594 183461 518628
rect 183495 518594 183553 518628
rect 183587 518594 183645 518628
rect 183679 518594 183737 518628
rect 183771 518594 183829 518628
rect 183863 518594 183921 518628
rect 183955 518594 184013 518628
rect 184047 518594 184105 518628
rect 184139 518594 184197 518628
rect 184231 518594 184289 518628
rect 184323 518594 184381 518628
rect 184415 518594 184473 518628
rect 184507 518594 184565 518628
rect 184599 518594 184657 518628
rect 184691 518594 184749 518628
rect 184783 518594 184841 518628
rect 184875 518594 184933 518628
rect 184967 518594 185025 518628
rect 185059 518594 185117 518628
rect 185151 518594 185209 518628
rect 185243 518594 185301 518628
rect 185335 518594 185393 518628
rect 185427 518594 185485 518628
rect 185519 518594 185577 518628
rect 185611 518594 185669 518628
rect 185703 518594 185761 518628
rect 185795 518594 185853 518628
rect 185887 518594 185945 518628
rect 185979 518594 186037 518628
rect 186071 518594 186129 518628
rect 186163 518594 186221 518628
rect 186255 518594 186313 518628
rect 186347 518594 186405 518628
rect 186439 518594 186497 518628
rect 186531 518594 186589 518628
rect 186623 518594 186681 518628
rect 186715 518594 186773 518628
rect 186807 518594 186865 518628
rect 186899 518594 186957 518628
rect 186991 518594 187049 518628
rect 187083 518594 187141 518628
rect 187175 518594 187233 518628
rect 187267 518594 187325 518628
rect 187359 518594 187417 518628
rect 187451 518594 187480 518628
rect 172225 518531 172467 518594
rect 172225 518497 172243 518531
rect 172277 518497 172415 518531
rect 172449 518497 172467 518531
rect 172225 518444 172467 518497
rect 172501 518533 173570 518594
rect 172501 518499 172519 518533
rect 172553 518499 173519 518533
rect 173553 518499 173570 518533
rect 172501 518485 173570 518499
rect 173605 518533 174674 518594
rect 173605 518499 173623 518533
rect 173657 518499 174623 518533
rect 174657 518499 174674 518533
rect 173605 518485 174674 518499
rect 174801 518500 174859 518594
rect 172225 518370 172329 518444
rect 172225 518336 172275 518370
rect 172309 518336 172329 518370
rect 172363 518376 172383 518410
rect 172417 518376 172467 518410
rect 172363 518302 172467 518376
rect 172818 518370 172886 518485
rect 172818 518336 172835 518370
rect 172869 518336 172886 518370
rect 172818 518319 172886 518336
rect 173182 518406 173252 518421
rect 173182 518372 173199 518406
rect 173233 518372 173252 518406
rect 172225 518255 172467 518302
rect 172225 518221 172243 518255
rect 172277 518221 172415 518255
rect 172449 518221 172467 518255
rect 172225 518160 172467 518221
rect 173182 518171 173252 518372
rect 173922 518370 173990 518485
rect 174801 518466 174813 518500
rect 174847 518466 174859 518500
rect 174893 518533 175962 518594
rect 174893 518499 174911 518533
rect 174945 518499 175911 518533
rect 175945 518499 175962 518533
rect 174893 518485 175962 518499
rect 175997 518533 177066 518594
rect 175997 518499 176015 518533
rect 176049 518499 177015 518533
rect 177049 518499 177066 518533
rect 175997 518485 177066 518499
rect 177101 518533 178170 518594
rect 177101 518499 177119 518533
rect 177153 518499 178119 518533
rect 178153 518499 178170 518533
rect 177101 518485 178170 518499
rect 178205 518533 179274 518594
rect 178205 518499 178223 518533
rect 178257 518499 179223 518533
rect 179257 518499 179274 518533
rect 178205 518485 179274 518499
rect 179309 518533 179827 518594
rect 179309 518499 179327 518533
rect 179361 518499 179775 518533
rect 179809 518499 179827 518533
rect 174801 518449 174859 518466
rect 173922 518336 173939 518370
rect 173973 518336 173990 518370
rect 173922 518319 173990 518336
rect 174286 518406 174356 518421
rect 174286 518372 174303 518406
rect 174337 518372 174356 518406
rect 174286 518171 174356 518372
rect 175210 518370 175278 518485
rect 175210 518336 175227 518370
rect 175261 518336 175278 518370
rect 175210 518319 175278 518336
rect 175574 518406 175644 518421
rect 175574 518372 175591 518406
rect 175625 518372 175644 518406
rect 174801 518282 174859 518317
rect 174801 518248 174813 518282
rect 174847 518248 174859 518282
rect 174801 518189 174859 518248
rect 172225 518126 172243 518160
rect 172277 518126 172415 518160
rect 172449 518126 172467 518160
rect 172225 518084 172467 518126
rect 172501 518160 173570 518171
rect 172501 518126 172519 518160
rect 172553 518126 173519 518160
rect 173553 518126 173570 518160
rect 172501 518084 173570 518126
rect 173605 518160 174674 518171
rect 173605 518126 173623 518160
rect 173657 518126 174623 518160
rect 174657 518126 174674 518160
rect 173605 518084 174674 518126
rect 174801 518155 174813 518189
rect 174847 518155 174859 518189
rect 175574 518171 175644 518372
rect 176314 518370 176382 518485
rect 176314 518336 176331 518370
rect 176365 518336 176382 518370
rect 176314 518319 176382 518336
rect 176678 518406 176748 518421
rect 176678 518372 176695 518406
rect 176729 518372 176748 518406
rect 176678 518171 176748 518372
rect 177418 518370 177486 518485
rect 177418 518336 177435 518370
rect 177469 518336 177486 518370
rect 177418 518319 177486 518336
rect 177782 518406 177852 518421
rect 177782 518372 177799 518406
rect 177833 518372 177852 518406
rect 177782 518171 177852 518372
rect 178522 518370 178590 518485
rect 179309 518440 179827 518499
rect 179953 518500 180011 518594
rect 179953 518466 179965 518500
rect 179999 518466 180011 518500
rect 180045 518533 181114 518594
rect 180045 518499 180063 518533
rect 180097 518499 181063 518533
rect 181097 518499 181114 518533
rect 180045 518485 181114 518499
rect 181149 518533 182218 518594
rect 181149 518499 181167 518533
rect 181201 518499 182167 518533
rect 182201 518499 182218 518533
rect 181149 518485 182218 518499
rect 182253 518533 183322 518594
rect 182253 518499 182271 518533
rect 182305 518499 183271 518533
rect 183305 518499 183322 518533
rect 182253 518485 183322 518499
rect 183357 518533 184426 518594
rect 183357 518499 183375 518533
rect 183409 518499 184375 518533
rect 184409 518499 184426 518533
rect 183357 518485 184426 518499
rect 184461 518533 184979 518594
rect 184461 518499 184479 518533
rect 184513 518499 184927 518533
rect 184961 518499 184979 518533
rect 179953 518449 180011 518466
rect 178522 518336 178539 518370
rect 178573 518336 178590 518370
rect 178522 518319 178590 518336
rect 178886 518406 178956 518421
rect 178886 518372 178903 518406
rect 178937 518372 178956 518406
rect 178886 518171 178956 518372
rect 179309 518370 179551 518440
rect 179309 518336 179387 518370
rect 179421 518336 179497 518370
rect 179531 518336 179551 518370
rect 179585 518372 179605 518406
rect 179639 518372 179715 518406
rect 179749 518372 179827 518406
rect 179585 518302 179827 518372
rect 180362 518370 180430 518485
rect 180362 518336 180379 518370
rect 180413 518336 180430 518370
rect 180362 518319 180430 518336
rect 180726 518406 180796 518421
rect 180726 518372 180743 518406
rect 180777 518372 180796 518406
rect 179309 518262 179827 518302
rect 179309 518228 179327 518262
rect 179361 518228 179775 518262
rect 179809 518228 179827 518262
rect 174801 518084 174859 518155
rect 174893 518160 175962 518171
rect 174893 518126 174911 518160
rect 174945 518126 175911 518160
rect 175945 518126 175962 518160
rect 174893 518084 175962 518126
rect 175997 518160 177066 518171
rect 175997 518126 176015 518160
rect 176049 518126 177015 518160
rect 177049 518126 177066 518160
rect 175997 518084 177066 518126
rect 177101 518160 178170 518171
rect 177101 518126 177119 518160
rect 177153 518126 178119 518160
rect 178153 518126 178170 518160
rect 177101 518084 178170 518126
rect 178205 518160 179274 518171
rect 178205 518126 178223 518160
rect 178257 518126 179223 518160
rect 179257 518126 179274 518160
rect 178205 518084 179274 518126
rect 179309 518160 179827 518228
rect 179309 518126 179327 518160
rect 179361 518126 179775 518160
rect 179809 518126 179827 518160
rect 179309 518084 179827 518126
rect 179953 518282 180011 518317
rect 179953 518248 179965 518282
rect 179999 518248 180011 518282
rect 179953 518189 180011 518248
rect 179953 518155 179965 518189
rect 179999 518155 180011 518189
rect 180726 518171 180796 518372
rect 181466 518370 181534 518485
rect 181466 518336 181483 518370
rect 181517 518336 181534 518370
rect 181466 518319 181534 518336
rect 181830 518406 181900 518421
rect 181830 518372 181847 518406
rect 181881 518372 181900 518406
rect 181830 518171 181900 518372
rect 182570 518370 182638 518485
rect 182570 518336 182587 518370
rect 182621 518336 182638 518370
rect 182570 518319 182638 518336
rect 182934 518406 183004 518421
rect 182934 518372 182951 518406
rect 182985 518372 183004 518406
rect 182934 518171 183004 518372
rect 183674 518370 183742 518485
rect 184461 518440 184979 518499
rect 185105 518500 185163 518594
rect 185105 518466 185117 518500
rect 185151 518466 185163 518500
rect 185197 518533 186266 518594
rect 185197 518499 185215 518533
rect 185249 518499 186215 518533
rect 186249 518499 186266 518533
rect 185197 518485 186266 518499
rect 186301 518533 187003 518594
rect 186301 518499 186319 518533
rect 186353 518499 186951 518533
rect 186985 518499 187003 518533
rect 185105 518449 185163 518466
rect 183674 518336 183691 518370
rect 183725 518336 183742 518370
rect 183674 518319 183742 518336
rect 184038 518406 184108 518421
rect 184038 518372 184055 518406
rect 184089 518372 184108 518406
rect 184038 518171 184108 518372
rect 184461 518370 184703 518440
rect 184461 518336 184539 518370
rect 184573 518336 184649 518370
rect 184683 518336 184703 518370
rect 184737 518372 184757 518406
rect 184791 518372 184867 518406
rect 184901 518372 184979 518406
rect 184737 518302 184979 518372
rect 185514 518370 185582 518485
rect 186301 518440 187003 518499
rect 187221 518531 187463 518594
rect 187221 518497 187239 518531
rect 187273 518497 187411 518531
rect 187445 518497 187463 518531
rect 187221 518444 187463 518497
rect 185514 518336 185531 518370
rect 185565 518336 185582 518370
rect 185514 518319 185582 518336
rect 185878 518406 185948 518421
rect 185878 518372 185895 518406
rect 185929 518372 185948 518406
rect 184461 518262 184979 518302
rect 184461 518228 184479 518262
rect 184513 518228 184927 518262
rect 184961 518228 184979 518262
rect 179953 518084 180011 518155
rect 180045 518160 181114 518171
rect 180045 518126 180063 518160
rect 180097 518126 181063 518160
rect 181097 518126 181114 518160
rect 180045 518084 181114 518126
rect 181149 518160 182218 518171
rect 181149 518126 181167 518160
rect 181201 518126 182167 518160
rect 182201 518126 182218 518160
rect 181149 518084 182218 518126
rect 182253 518160 183322 518171
rect 182253 518126 182271 518160
rect 182305 518126 183271 518160
rect 183305 518126 183322 518160
rect 182253 518084 183322 518126
rect 183357 518160 184426 518171
rect 183357 518126 183375 518160
rect 183409 518126 184375 518160
rect 184409 518126 184426 518160
rect 183357 518084 184426 518126
rect 184461 518160 184979 518228
rect 184461 518126 184479 518160
rect 184513 518126 184927 518160
rect 184961 518126 184979 518160
rect 184461 518084 184979 518126
rect 185105 518282 185163 518317
rect 185105 518248 185117 518282
rect 185151 518248 185163 518282
rect 185105 518189 185163 518248
rect 185105 518155 185117 518189
rect 185151 518155 185163 518189
rect 185878 518171 185948 518372
rect 186301 518370 186631 518440
rect 186301 518336 186379 518370
rect 186413 518336 186478 518370
rect 186512 518336 186577 518370
rect 186611 518336 186631 518370
rect 186665 518372 186685 518406
rect 186719 518372 186788 518406
rect 186822 518372 186891 518406
rect 186925 518372 187003 518406
rect 186665 518302 187003 518372
rect 186301 518262 187003 518302
rect 186301 518228 186319 518262
rect 186353 518228 186951 518262
rect 186985 518228 187003 518262
rect 185105 518084 185163 518155
rect 185197 518160 186266 518171
rect 185197 518126 185215 518160
rect 185249 518126 186215 518160
rect 186249 518126 186266 518160
rect 185197 518084 186266 518126
rect 186301 518160 187003 518228
rect 186301 518126 186319 518160
rect 186353 518126 186951 518160
rect 186985 518126 187003 518160
rect 186301 518084 187003 518126
rect 187221 518376 187271 518410
rect 187305 518376 187325 518410
rect 187221 518302 187325 518376
rect 187359 518370 187463 518444
rect 187359 518336 187379 518370
rect 187413 518336 187463 518370
rect 187221 518255 187463 518302
rect 187221 518221 187239 518255
rect 187273 518221 187411 518255
rect 187445 518221 187463 518255
rect 187221 518160 187463 518221
rect 187221 518126 187239 518160
rect 187273 518126 187411 518160
rect 187445 518126 187463 518160
rect 187221 518084 187463 518126
rect 172208 518050 172237 518084
rect 172271 518050 172329 518084
rect 172363 518050 172421 518084
rect 172455 518050 172513 518084
rect 172547 518050 172605 518084
rect 172639 518050 172697 518084
rect 172731 518050 172789 518084
rect 172823 518050 172881 518084
rect 172915 518050 172973 518084
rect 173007 518050 173065 518084
rect 173099 518050 173157 518084
rect 173191 518050 173249 518084
rect 173283 518050 173341 518084
rect 173375 518050 173433 518084
rect 173467 518050 173525 518084
rect 173559 518050 173617 518084
rect 173651 518050 173709 518084
rect 173743 518050 173801 518084
rect 173835 518050 173893 518084
rect 173927 518050 173985 518084
rect 174019 518050 174077 518084
rect 174111 518050 174169 518084
rect 174203 518050 174261 518084
rect 174295 518050 174353 518084
rect 174387 518050 174445 518084
rect 174479 518050 174537 518084
rect 174571 518050 174629 518084
rect 174663 518050 174721 518084
rect 174755 518050 174813 518084
rect 174847 518050 174905 518084
rect 174939 518050 174997 518084
rect 175031 518050 175089 518084
rect 175123 518050 175181 518084
rect 175215 518050 175273 518084
rect 175307 518050 175365 518084
rect 175399 518050 175457 518084
rect 175491 518050 175549 518084
rect 175583 518050 175641 518084
rect 175675 518050 175733 518084
rect 175767 518050 175825 518084
rect 175859 518050 175917 518084
rect 175951 518050 176009 518084
rect 176043 518050 176101 518084
rect 176135 518050 176193 518084
rect 176227 518050 176285 518084
rect 176319 518050 176377 518084
rect 176411 518050 176469 518084
rect 176503 518050 176561 518084
rect 176595 518050 176653 518084
rect 176687 518050 176745 518084
rect 176779 518050 176837 518084
rect 176871 518050 176929 518084
rect 176963 518050 177021 518084
rect 177055 518050 177113 518084
rect 177147 518050 177205 518084
rect 177239 518050 177297 518084
rect 177331 518050 177389 518084
rect 177423 518050 177481 518084
rect 177515 518050 177573 518084
rect 177607 518050 177665 518084
rect 177699 518050 177757 518084
rect 177791 518050 177849 518084
rect 177883 518050 177941 518084
rect 177975 518050 178033 518084
rect 178067 518050 178125 518084
rect 178159 518050 178217 518084
rect 178251 518050 178309 518084
rect 178343 518050 178401 518084
rect 178435 518050 178493 518084
rect 178527 518050 178585 518084
rect 178619 518050 178677 518084
rect 178711 518050 178769 518084
rect 178803 518050 178861 518084
rect 178895 518050 178953 518084
rect 178987 518050 179045 518084
rect 179079 518050 179137 518084
rect 179171 518050 179229 518084
rect 179263 518050 179321 518084
rect 179355 518050 179413 518084
rect 179447 518050 179505 518084
rect 179539 518050 179597 518084
rect 179631 518050 179689 518084
rect 179723 518050 179781 518084
rect 179815 518050 179873 518084
rect 179907 518050 179965 518084
rect 179999 518050 180057 518084
rect 180091 518050 180149 518084
rect 180183 518050 180241 518084
rect 180275 518050 180333 518084
rect 180367 518050 180425 518084
rect 180459 518050 180517 518084
rect 180551 518050 180609 518084
rect 180643 518050 180701 518084
rect 180735 518050 180793 518084
rect 180827 518050 180885 518084
rect 180919 518050 180977 518084
rect 181011 518050 181069 518084
rect 181103 518050 181161 518084
rect 181195 518050 181253 518084
rect 181287 518050 181345 518084
rect 181379 518050 181437 518084
rect 181471 518050 181529 518084
rect 181563 518050 181621 518084
rect 181655 518050 181713 518084
rect 181747 518050 181805 518084
rect 181839 518050 181897 518084
rect 181931 518050 181989 518084
rect 182023 518050 182081 518084
rect 182115 518050 182173 518084
rect 182207 518050 182265 518084
rect 182299 518050 182357 518084
rect 182391 518050 182449 518084
rect 182483 518050 182541 518084
rect 182575 518050 182633 518084
rect 182667 518050 182725 518084
rect 182759 518050 182817 518084
rect 182851 518050 182909 518084
rect 182943 518050 183001 518084
rect 183035 518050 183093 518084
rect 183127 518050 183185 518084
rect 183219 518050 183277 518084
rect 183311 518050 183369 518084
rect 183403 518050 183461 518084
rect 183495 518050 183553 518084
rect 183587 518050 183645 518084
rect 183679 518050 183737 518084
rect 183771 518050 183829 518084
rect 183863 518050 183921 518084
rect 183955 518050 184013 518084
rect 184047 518050 184105 518084
rect 184139 518050 184197 518084
rect 184231 518050 184289 518084
rect 184323 518050 184381 518084
rect 184415 518050 184473 518084
rect 184507 518050 184565 518084
rect 184599 518050 184657 518084
rect 184691 518050 184749 518084
rect 184783 518050 184841 518084
rect 184875 518050 184933 518084
rect 184967 518050 185025 518084
rect 185059 518050 185117 518084
rect 185151 518050 185209 518084
rect 185243 518050 185301 518084
rect 185335 518050 185393 518084
rect 185427 518050 185485 518084
rect 185519 518050 185577 518084
rect 185611 518050 185669 518084
rect 185703 518050 185761 518084
rect 185795 518050 185853 518084
rect 185887 518050 185945 518084
rect 185979 518050 186037 518084
rect 186071 518050 186129 518084
rect 186163 518050 186221 518084
rect 186255 518050 186313 518084
rect 186347 518050 186405 518084
rect 186439 518050 186497 518084
rect 186531 518050 186589 518084
rect 186623 518050 186681 518084
rect 186715 518050 186773 518084
rect 186807 518050 186865 518084
rect 186899 518050 186957 518084
rect 186991 518050 187049 518084
rect 187083 518050 187141 518084
rect 187175 518050 187233 518084
rect 187267 518050 187325 518084
rect 187359 518050 187417 518084
rect 187451 518050 187480 518084
rect 172225 518008 172467 518050
rect 172225 517974 172243 518008
rect 172277 517974 172415 518008
rect 172449 517974 172467 518008
rect 172225 517913 172467 517974
rect 172501 518008 173570 518050
rect 172501 517974 172519 518008
rect 172553 517974 173519 518008
rect 173553 517974 173570 518008
rect 172501 517963 173570 517974
rect 173605 518008 174674 518050
rect 173605 517974 173623 518008
rect 173657 517974 174623 518008
rect 174657 517974 174674 518008
rect 173605 517963 174674 517974
rect 174709 518008 175778 518050
rect 174709 517974 174727 518008
rect 174761 517974 175727 518008
rect 175761 517974 175778 518008
rect 174709 517963 175778 517974
rect 175813 518008 176882 518050
rect 175813 517974 175831 518008
rect 175865 517974 176831 518008
rect 176865 517974 176882 518008
rect 175813 517963 176882 517974
rect 176917 518008 177251 518050
rect 176917 517974 176935 518008
rect 176969 517974 177199 518008
rect 177233 517974 177251 518008
rect 172225 517879 172243 517913
rect 172277 517879 172415 517913
rect 172449 517879 172467 517913
rect 172225 517832 172467 517879
rect 172225 517764 172275 517798
rect 172309 517764 172329 517798
rect 172225 517690 172329 517764
rect 172363 517758 172467 517832
rect 172363 517724 172383 517758
rect 172417 517724 172467 517758
rect 172818 517798 172886 517815
rect 172818 517764 172835 517798
rect 172869 517764 172886 517798
rect 172225 517637 172467 517690
rect 172818 517649 172886 517764
rect 173182 517762 173252 517963
rect 173182 517728 173199 517762
rect 173233 517728 173252 517762
rect 173182 517713 173252 517728
rect 173922 517798 173990 517815
rect 173922 517764 173939 517798
rect 173973 517764 173990 517798
rect 173922 517649 173990 517764
rect 174286 517762 174356 517963
rect 174286 517728 174303 517762
rect 174337 517728 174356 517762
rect 174286 517713 174356 517728
rect 175026 517798 175094 517815
rect 175026 517764 175043 517798
rect 175077 517764 175094 517798
rect 175026 517649 175094 517764
rect 175390 517762 175460 517963
rect 175390 517728 175407 517762
rect 175441 517728 175460 517762
rect 175390 517713 175460 517728
rect 176130 517798 176198 517815
rect 176130 517764 176147 517798
rect 176181 517764 176198 517798
rect 176130 517649 176198 517764
rect 176494 517762 176564 517963
rect 176917 517906 177251 517974
rect 176917 517872 176935 517906
rect 176969 517872 177199 517906
rect 177233 517872 177251 517906
rect 176917 517832 177251 517872
rect 176494 517728 176511 517762
rect 176545 517728 176564 517762
rect 176494 517713 176564 517728
rect 176917 517764 176937 517798
rect 176971 517764 177067 517798
rect 176917 517694 177067 517764
rect 177101 517762 177251 517832
rect 177377 517979 177435 518050
rect 177377 517945 177389 517979
rect 177423 517945 177435 517979
rect 177469 518008 178538 518050
rect 177469 517974 177487 518008
rect 177521 517974 178487 518008
rect 178521 517974 178538 518008
rect 177469 517963 178538 517974
rect 178573 518008 179642 518050
rect 178573 517974 178591 518008
rect 178625 517974 179591 518008
rect 179625 517974 179642 518008
rect 178573 517963 179642 517974
rect 179677 518008 180746 518050
rect 179677 517974 179695 518008
rect 179729 517974 180695 518008
rect 180729 517974 180746 518008
rect 179677 517963 180746 517974
rect 180781 518008 181850 518050
rect 180781 517974 180799 518008
rect 180833 517974 181799 518008
rect 181833 517974 181850 518008
rect 180781 517963 181850 517974
rect 181885 518008 182403 518050
rect 181885 517974 181903 518008
rect 181937 517974 182351 518008
rect 182385 517974 182403 518008
rect 177377 517886 177435 517945
rect 177377 517852 177389 517886
rect 177423 517852 177435 517886
rect 177377 517817 177435 517852
rect 177101 517728 177197 517762
rect 177231 517728 177251 517762
rect 177786 517798 177854 517815
rect 177786 517764 177803 517798
rect 177837 517764 177854 517798
rect 172225 517603 172243 517637
rect 172277 517603 172415 517637
rect 172449 517603 172467 517637
rect 172225 517540 172467 517603
rect 172501 517635 173570 517649
rect 172501 517601 172519 517635
rect 172553 517601 173519 517635
rect 173553 517601 173570 517635
rect 172501 517540 173570 517601
rect 173605 517635 174674 517649
rect 173605 517601 173623 517635
rect 173657 517601 174623 517635
rect 174657 517601 174674 517635
rect 173605 517540 174674 517601
rect 174709 517635 175778 517649
rect 174709 517601 174727 517635
rect 174761 517601 175727 517635
rect 175761 517601 175778 517635
rect 174709 517540 175778 517601
rect 175813 517635 176882 517649
rect 175813 517601 175831 517635
rect 175865 517601 176831 517635
rect 176865 517601 176882 517635
rect 175813 517540 176882 517601
rect 176917 517642 177251 517694
rect 176917 517608 176935 517642
rect 176969 517608 177199 517642
rect 177233 517608 177251 517642
rect 176917 517540 177251 517608
rect 177377 517668 177435 517685
rect 177377 517634 177389 517668
rect 177423 517634 177435 517668
rect 177786 517649 177854 517764
rect 178150 517762 178220 517963
rect 178150 517728 178167 517762
rect 178201 517728 178220 517762
rect 178150 517713 178220 517728
rect 178890 517798 178958 517815
rect 178890 517764 178907 517798
rect 178941 517764 178958 517798
rect 178890 517649 178958 517764
rect 179254 517762 179324 517963
rect 179254 517728 179271 517762
rect 179305 517728 179324 517762
rect 179254 517713 179324 517728
rect 179994 517798 180062 517815
rect 179994 517764 180011 517798
rect 180045 517764 180062 517798
rect 179994 517649 180062 517764
rect 180358 517762 180428 517963
rect 180358 517728 180375 517762
rect 180409 517728 180428 517762
rect 180358 517713 180428 517728
rect 181098 517798 181166 517815
rect 181098 517764 181115 517798
rect 181149 517764 181166 517798
rect 181098 517649 181166 517764
rect 181462 517762 181532 517963
rect 181885 517906 182403 517974
rect 181885 517872 181903 517906
rect 181937 517872 182351 517906
rect 182385 517872 182403 517906
rect 181885 517832 182403 517872
rect 181462 517728 181479 517762
rect 181513 517728 181532 517762
rect 181462 517713 181532 517728
rect 181885 517764 181963 517798
rect 181997 517764 182073 517798
rect 182107 517764 182127 517798
rect 181885 517694 182127 517764
rect 182161 517762 182403 517832
rect 182529 517979 182587 518050
rect 182529 517945 182541 517979
rect 182575 517945 182587 517979
rect 182621 518008 183690 518050
rect 182621 517974 182639 518008
rect 182673 517974 183639 518008
rect 183673 517974 183690 518008
rect 182621 517963 183690 517974
rect 183725 518008 184794 518050
rect 183725 517974 183743 518008
rect 183777 517974 184743 518008
rect 184777 517974 184794 518008
rect 183725 517963 184794 517974
rect 184829 518008 185898 518050
rect 184829 517974 184847 518008
rect 184881 517974 185847 518008
rect 185881 517974 185898 518008
rect 184829 517963 185898 517974
rect 185933 518008 187002 518050
rect 185933 517974 185951 518008
rect 185985 517974 186951 518008
rect 186985 517974 187002 518008
rect 185933 517963 187002 517974
rect 187221 518008 187463 518050
rect 187221 517974 187239 518008
rect 187273 517974 187411 518008
rect 187445 517974 187463 518008
rect 182529 517886 182587 517945
rect 182529 517852 182541 517886
rect 182575 517852 182587 517886
rect 182529 517817 182587 517852
rect 182161 517728 182181 517762
rect 182215 517728 182291 517762
rect 182325 517728 182403 517762
rect 182938 517798 183006 517815
rect 182938 517764 182955 517798
rect 182989 517764 183006 517798
rect 177377 517540 177435 517634
rect 177469 517635 178538 517649
rect 177469 517601 177487 517635
rect 177521 517601 178487 517635
rect 178521 517601 178538 517635
rect 177469 517540 178538 517601
rect 178573 517635 179642 517649
rect 178573 517601 178591 517635
rect 178625 517601 179591 517635
rect 179625 517601 179642 517635
rect 178573 517540 179642 517601
rect 179677 517635 180746 517649
rect 179677 517601 179695 517635
rect 179729 517601 180695 517635
rect 180729 517601 180746 517635
rect 179677 517540 180746 517601
rect 180781 517635 181850 517649
rect 180781 517601 180799 517635
rect 180833 517601 181799 517635
rect 181833 517601 181850 517635
rect 180781 517540 181850 517601
rect 181885 517635 182403 517694
rect 181885 517601 181903 517635
rect 181937 517601 182351 517635
rect 182385 517601 182403 517635
rect 181885 517540 182403 517601
rect 182529 517668 182587 517685
rect 182529 517634 182541 517668
rect 182575 517634 182587 517668
rect 182938 517649 183006 517764
rect 183302 517762 183372 517963
rect 183302 517728 183319 517762
rect 183353 517728 183372 517762
rect 183302 517713 183372 517728
rect 184042 517798 184110 517815
rect 184042 517764 184059 517798
rect 184093 517764 184110 517798
rect 184042 517649 184110 517764
rect 184406 517762 184476 517963
rect 184406 517728 184423 517762
rect 184457 517728 184476 517762
rect 184406 517713 184476 517728
rect 185146 517798 185214 517815
rect 185146 517764 185163 517798
rect 185197 517764 185214 517798
rect 185146 517649 185214 517764
rect 185510 517762 185580 517963
rect 185510 517728 185527 517762
rect 185561 517728 185580 517762
rect 185510 517713 185580 517728
rect 186250 517798 186318 517815
rect 186250 517764 186267 517798
rect 186301 517764 186318 517798
rect 186250 517649 186318 517764
rect 186614 517762 186684 517963
rect 186614 517728 186631 517762
rect 186665 517728 186684 517762
rect 186614 517713 186684 517728
rect 187221 517913 187463 517974
rect 187221 517879 187239 517913
rect 187273 517879 187411 517913
rect 187445 517879 187463 517913
rect 187221 517832 187463 517879
rect 187221 517758 187325 517832
rect 187221 517724 187271 517758
rect 187305 517724 187325 517758
rect 187359 517764 187379 517798
rect 187413 517764 187463 517798
rect 187359 517690 187463 517764
rect 182529 517540 182587 517634
rect 182621 517635 183690 517649
rect 182621 517601 182639 517635
rect 182673 517601 183639 517635
rect 183673 517601 183690 517635
rect 182621 517540 183690 517601
rect 183725 517635 184794 517649
rect 183725 517601 183743 517635
rect 183777 517601 184743 517635
rect 184777 517601 184794 517635
rect 183725 517540 184794 517601
rect 184829 517635 185898 517649
rect 184829 517601 184847 517635
rect 184881 517601 185847 517635
rect 185881 517601 185898 517635
rect 184829 517540 185898 517601
rect 185933 517635 187002 517649
rect 185933 517601 185951 517635
rect 185985 517601 186951 517635
rect 186985 517601 187002 517635
rect 185933 517540 187002 517601
rect 187221 517637 187463 517690
rect 187221 517603 187239 517637
rect 187273 517603 187411 517637
rect 187445 517603 187463 517637
rect 187221 517540 187463 517603
rect 172208 517506 172237 517540
rect 172271 517506 172329 517540
rect 172363 517506 172421 517540
rect 172455 517506 172513 517540
rect 172547 517506 172605 517540
rect 172639 517506 172697 517540
rect 172731 517506 172789 517540
rect 172823 517506 172881 517540
rect 172915 517506 172973 517540
rect 173007 517506 173065 517540
rect 173099 517506 173157 517540
rect 173191 517506 173249 517540
rect 173283 517506 173341 517540
rect 173375 517506 173433 517540
rect 173467 517506 173525 517540
rect 173559 517506 173617 517540
rect 173651 517506 173709 517540
rect 173743 517506 173801 517540
rect 173835 517506 173893 517540
rect 173927 517506 173985 517540
rect 174019 517506 174077 517540
rect 174111 517506 174169 517540
rect 174203 517506 174261 517540
rect 174295 517506 174353 517540
rect 174387 517506 174445 517540
rect 174479 517506 174537 517540
rect 174571 517506 174629 517540
rect 174663 517506 174721 517540
rect 174755 517506 174813 517540
rect 174847 517506 174905 517540
rect 174939 517506 174997 517540
rect 175031 517506 175089 517540
rect 175123 517506 175181 517540
rect 175215 517506 175273 517540
rect 175307 517506 175365 517540
rect 175399 517506 175457 517540
rect 175491 517506 175549 517540
rect 175583 517506 175641 517540
rect 175675 517506 175733 517540
rect 175767 517506 175825 517540
rect 175859 517506 175917 517540
rect 175951 517506 176009 517540
rect 176043 517506 176101 517540
rect 176135 517506 176193 517540
rect 176227 517506 176285 517540
rect 176319 517506 176377 517540
rect 176411 517506 176469 517540
rect 176503 517506 176561 517540
rect 176595 517506 176653 517540
rect 176687 517506 176745 517540
rect 176779 517506 176837 517540
rect 176871 517506 176929 517540
rect 176963 517506 177021 517540
rect 177055 517506 177113 517540
rect 177147 517506 177205 517540
rect 177239 517506 177297 517540
rect 177331 517506 177389 517540
rect 177423 517506 177481 517540
rect 177515 517506 177573 517540
rect 177607 517506 177665 517540
rect 177699 517506 177757 517540
rect 177791 517506 177849 517540
rect 177883 517506 177941 517540
rect 177975 517506 178033 517540
rect 178067 517506 178125 517540
rect 178159 517506 178217 517540
rect 178251 517506 178309 517540
rect 178343 517506 178401 517540
rect 178435 517506 178493 517540
rect 178527 517506 178585 517540
rect 178619 517506 178677 517540
rect 178711 517506 178769 517540
rect 178803 517506 178861 517540
rect 178895 517506 178953 517540
rect 178987 517506 179045 517540
rect 179079 517506 179137 517540
rect 179171 517506 179229 517540
rect 179263 517506 179321 517540
rect 179355 517506 179413 517540
rect 179447 517506 179505 517540
rect 179539 517506 179597 517540
rect 179631 517506 179689 517540
rect 179723 517506 179781 517540
rect 179815 517506 179873 517540
rect 179907 517506 179965 517540
rect 179999 517506 180057 517540
rect 180091 517506 180149 517540
rect 180183 517506 180241 517540
rect 180275 517506 180333 517540
rect 180367 517506 180425 517540
rect 180459 517506 180517 517540
rect 180551 517506 180609 517540
rect 180643 517506 180701 517540
rect 180735 517506 180793 517540
rect 180827 517506 180885 517540
rect 180919 517506 180977 517540
rect 181011 517506 181069 517540
rect 181103 517506 181161 517540
rect 181195 517506 181253 517540
rect 181287 517506 181345 517540
rect 181379 517506 181437 517540
rect 181471 517506 181529 517540
rect 181563 517506 181621 517540
rect 181655 517506 181713 517540
rect 181747 517506 181805 517540
rect 181839 517506 181897 517540
rect 181931 517506 181989 517540
rect 182023 517506 182081 517540
rect 182115 517506 182173 517540
rect 182207 517506 182265 517540
rect 182299 517506 182357 517540
rect 182391 517506 182449 517540
rect 182483 517506 182541 517540
rect 182575 517506 182633 517540
rect 182667 517506 182725 517540
rect 182759 517506 182817 517540
rect 182851 517506 182909 517540
rect 182943 517506 183001 517540
rect 183035 517506 183093 517540
rect 183127 517506 183185 517540
rect 183219 517506 183277 517540
rect 183311 517506 183369 517540
rect 183403 517506 183461 517540
rect 183495 517506 183553 517540
rect 183587 517506 183645 517540
rect 183679 517506 183737 517540
rect 183771 517506 183829 517540
rect 183863 517506 183921 517540
rect 183955 517506 184013 517540
rect 184047 517506 184105 517540
rect 184139 517506 184197 517540
rect 184231 517506 184289 517540
rect 184323 517506 184381 517540
rect 184415 517506 184473 517540
rect 184507 517506 184565 517540
rect 184599 517506 184657 517540
rect 184691 517506 184749 517540
rect 184783 517506 184841 517540
rect 184875 517506 184933 517540
rect 184967 517506 185025 517540
rect 185059 517506 185117 517540
rect 185151 517506 185209 517540
rect 185243 517506 185301 517540
rect 185335 517506 185393 517540
rect 185427 517506 185485 517540
rect 185519 517506 185577 517540
rect 185611 517506 185669 517540
rect 185703 517506 185761 517540
rect 185795 517506 185853 517540
rect 185887 517506 185945 517540
rect 185979 517506 186037 517540
rect 186071 517506 186129 517540
rect 186163 517506 186221 517540
rect 186255 517506 186313 517540
rect 186347 517506 186405 517540
rect 186439 517506 186497 517540
rect 186531 517506 186589 517540
rect 186623 517506 186681 517540
rect 186715 517506 186773 517540
rect 186807 517506 186865 517540
rect 186899 517506 186957 517540
rect 186991 517506 187049 517540
rect 187083 517506 187141 517540
rect 187175 517506 187233 517540
rect 187267 517506 187325 517540
rect 187359 517506 187417 517540
rect 187451 517506 187480 517540
rect 172225 517443 172467 517506
rect 172225 517409 172243 517443
rect 172277 517409 172415 517443
rect 172449 517409 172467 517443
rect 172225 517356 172467 517409
rect 172501 517445 173570 517506
rect 172501 517411 172519 517445
rect 172553 517411 173519 517445
rect 173553 517411 173570 517445
rect 172501 517397 173570 517411
rect 173605 517445 174674 517506
rect 173605 517411 173623 517445
rect 173657 517411 174623 517445
rect 174657 517411 174674 517445
rect 173605 517397 174674 517411
rect 174801 517412 174859 517506
rect 172225 517282 172329 517356
rect 172225 517248 172275 517282
rect 172309 517248 172329 517282
rect 172363 517288 172383 517322
rect 172417 517288 172467 517322
rect 172363 517214 172467 517288
rect 172818 517282 172886 517397
rect 172818 517248 172835 517282
rect 172869 517248 172886 517282
rect 172818 517231 172886 517248
rect 173182 517318 173252 517333
rect 173182 517284 173199 517318
rect 173233 517284 173252 517318
rect 172225 517167 172467 517214
rect 172225 517133 172243 517167
rect 172277 517133 172415 517167
rect 172449 517133 172467 517167
rect 172225 517072 172467 517133
rect 173182 517083 173252 517284
rect 173922 517282 173990 517397
rect 174801 517378 174813 517412
rect 174847 517378 174859 517412
rect 174893 517445 175962 517506
rect 174893 517411 174911 517445
rect 174945 517411 175911 517445
rect 175945 517411 175962 517445
rect 174893 517397 175962 517411
rect 175997 517445 177066 517506
rect 175997 517411 176015 517445
rect 176049 517411 177015 517445
rect 177049 517411 177066 517445
rect 175997 517397 177066 517411
rect 177101 517445 178170 517506
rect 177101 517411 177119 517445
rect 177153 517411 178119 517445
rect 178153 517411 178170 517445
rect 177101 517397 178170 517411
rect 178205 517445 179274 517506
rect 178205 517411 178223 517445
rect 178257 517411 179223 517445
rect 179257 517411 179274 517445
rect 178205 517397 179274 517411
rect 179309 517445 179827 517506
rect 179309 517411 179327 517445
rect 179361 517411 179775 517445
rect 179809 517411 179827 517445
rect 174801 517361 174859 517378
rect 173922 517248 173939 517282
rect 173973 517248 173990 517282
rect 173922 517231 173990 517248
rect 174286 517318 174356 517333
rect 174286 517284 174303 517318
rect 174337 517284 174356 517318
rect 174286 517083 174356 517284
rect 175210 517282 175278 517397
rect 175210 517248 175227 517282
rect 175261 517248 175278 517282
rect 175210 517231 175278 517248
rect 175574 517318 175644 517333
rect 175574 517284 175591 517318
rect 175625 517284 175644 517318
rect 174801 517194 174859 517229
rect 174801 517160 174813 517194
rect 174847 517160 174859 517194
rect 174801 517101 174859 517160
rect 172225 517038 172243 517072
rect 172277 517038 172415 517072
rect 172449 517038 172467 517072
rect 172225 516996 172467 517038
rect 172501 517072 173570 517083
rect 172501 517038 172519 517072
rect 172553 517038 173519 517072
rect 173553 517038 173570 517072
rect 172501 516996 173570 517038
rect 173605 517072 174674 517083
rect 173605 517038 173623 517072
rect 173657 517038 174623 517072
rect 174657 517038 174674 517072
rect 173605 516996 174674 517038
rect 174801 517067 174813 517101
rect 174847 517067 174859 517101
rect 175574 517083 175644 517284
rect 176314 517282 176382 517397
rect 176314 517248 176331 517282
rect 176365 517248 176382 517282
rect 176314 517231 176382 517248
rect 176678 517318 176748 517333
rect 176678 517284 176695 517318
rect 176729 517284 176748 517318
rect 176678 517083 176748 517284
rect 177418 517282 177486 517397
rect 177418 517248 177435 517282
rect 177469 517248 177486 517282
rect 177418 517231 177486 517248
rect 177782 517318 177852 517333
rect 177782 517284 177799 517318
rect 177833 517284 177852 517318
rect 177782 517083 177852 517284
rect 178522 517282 178590 517397
rect 179309 517352 179827 517411
rect 179953 517412 180011 517506
rect 179953 517378 179965 517412
rect 179999 517378 180011 517412
rect 180045 517445 181114 517506
rect 180045 517411 180063 517445
rect 180097 517411 181063 517445
rect 181097 517411 181114 517445
rect 180045 517397 181114 517411
rect 181149 517445 182218 517506
rect 181149 517411 181167 517445
rect 181201 517411 182167 517445
rect 182201 517411 182218 517445
rect 181149 517397 182218 517411
rect 182253 517445 183322 517506
rect 182253 517411 182271 517445
rect 182305 517411 183271 517445
rect 183305 517411 183322 517445
rect 182253 517397 183322 517411
rect 183357 517445 184426 517506
rect 183357 517411 183375 517445
rect 183409 517411 184375 517445
rect 184409 517411 184426 517445
rect 183357 517397 184426 517411
rect 184461 517445 184979 517506
rect 184461 517411 184479 517445
rect 184513 517411 184927 517445
rect 184961 517411 184979 517445
rect 179953 517361 180011 517378
rect 178522 517248 178539 517282
rect 178573 517248 178590 517282
rect 178522 517231 178590 517248
rect 178886 517318 178956 517333
rect 178886 517284 178903 517318
rect 178937 517284 178956 517318
rect 178886 517083 178956 517284
rect 179309 517282 179551 517352
rect 179309 517248 179387 517282
rect 179421 517248 179497 517282
rect 179531 517248 179551 517282
rect 179585 517284 179605 517318
rect 179639 517284 179715 517318
rect 179749 517284 179827 517318
rect 179585 517214 179827 517284
rect 180362 517282 180430 517397
rect 180362 517248 180379 517282
rect 180413 517248 180430 517282
rect 180362 517231 180430 517248
rect 180726 517318 180796 517333
rect 180726 517284 180743 517318
rect 180777 517284 180796 517318
rect 179309 517174 179827 517214
rect 179309 517140 179327 517174
rect 179361 517140 179775 517174
rect 179809 517140 179827 517174
rect 174801 516996 174859 517067
rect 174893 517072 175962 517083
rect 174893 517038 174911 517072
rect 174945 517038 175911 517072
rect 175945 517038 175962 517072
rect 174893 516996 175962 517038
rect 175997 517072 177066 517083
rect 175997 517038 176015 517072
rect 176049 517038 177015 517072
rect 177049 517038 177066 517072
rect 175997 516996 177066 517038
rect 177101 517072 178170 517083
rect 177101 517038 177119 517072
rect 177153 517038 178119 517072
rect 178153 517038 178170 517072
rect 177101 516996 178170 517038
rect 178205 517072 179274 517083
rect 178205 517038 178223 517072
rect 178257 517038 179223 517072
rect 179257 517038 179274 517072
rect 178205 516996 179274 517038
rect 179309 517072 179827 517140
rect 179309 517038 179327 517072
rect 179361 517038 179775 517072
rect 179809 517038 179827 517072
rect 179309 516996 179827 517038
rect 179953 517194 180011 517229
rect 179953 517160 179965 517194
rect 179999 517160 180011 517194
rect 179953 517101 180011 517160
rect 179953 517067 179965 517101
rect 179999 517067 180011 517101
rect 180726 517083 180796 517284
rect 181466 517282 181534 517397
rect 181466 517248 181483 517282
rect 181517 517248 181534 517282
rect 181466 517231 181534 517248
rect 181830 517318 181900 517333
rect 181830 517284 181847 517318
rect 181881 517284 181900 517318
rect 181830 517083 181900 517284
rect 182570 517282 182638 517397
rect 182570 517248 182587 517282
rect 182621 517248 182638 517282
rect 182570 517231 182638 517248
rect 182934 517318 183004 517333
rect 182934 517284 182951 517318
rect 182985 517284 183004 517318
rect 182934 517083 183004 517284
rect 183674 517282 183742 517397
rect 184461 517352 184979 517411
rect 185105 517412 185163 517506
rect 185105 517378 185117 517412
rect 185151 517378 185163 517412
rect 185197 517445 186266 517506
rect 185197 517411 185215 517445
rect 185249 517411 186215 517445
rect 186249 517411 186266 517445
rect 185197 517397 186266 517411
rect 186301 517445 187003 517506
rect 186301 517411 186319 517445
rect 186353 517411 186951 517445
rect 186985 517411 187003 517445
rect 185105 517361 185163 517378
rect 183674 517248 183691 517282
rect 183725 517248 183742 517282
rect 183674 517231 183742 517248
rect 184038 517318 184108 517333
rect 184038 517284 184055 517318
rect 184089 517284 184108 517318
rect 184038 517083 184108 517284
rect 184461 517282 184703 517352
rect 184461 517248 184539 517282
rect 184573 517248 184649 517282
rect 184683 517248 184703 517282
rect 184737 517284 184757 517318
rect 184791 517284 184867 517318
rect 184901 517284 184979 517318
rect 184737 517214 184979 517284
rect 185514 517282 185582 517397
rect 186301 517352 187003 517411
rect 187221 517443 187463 517506
rect 187221 517409 187239 517443
rect 187273 517409 187411 517443
rect 187445 517409 187463 517443
rect 187221 517356 187463 517409
rect 185514 517248 185531 517282
rect 185565 517248 185582 517282
rect 185514 517231 185582 517248
rect 185878 517318 185948 517333
rect 185878 517284 185895 517318
rect 185929 517284 185948 517318
rect 184461 517174 184979 517214
rect 184461 517140 184479 517174
rect 184513 517140 184927 517174
rect 184961 517140 184979 517174
rect 179953 516996 180011 517067
rect 180045 517072 181114 517083
rect 180045 517038 180063 517072
rect 180097 517038 181063 517072
rect 181097 517038 181114 517072
rect 180045 516996 181114 517038
rect 181149 517072 182218 517083
rect 181149 517038 181167 517072
rect 181201 517038 182167 517072
rect 182201 517038 182218 517072
rect 181149 516996 182218 517038
rect 182253 517072 183322 517083
rect 182253 517038 182271 517072
rect 182305 517038 183271 517072
rect 183305 517038 183322 517072
rect 182253 516996 183322 517038
rect 183357 517072 184426 517083
rect 183357 517038 183375 517072
rect 183409 517038 184375 517072
rect 184409 517038 184426 517072
rect 183357 516996 184426 517038
rect 184461 517072 184979 517140
rect 184461 517038 184479 517072
rect 184513 517038 184927 517072
rect 184961 517038 184979 517072
rect 184461 516996 184979 517038
rect 185105 517194 185163 517229
rect 185105 517160 185117 517194
rect 185151 517160 185163 517194
rect 185105 517101 185163 517160
rect 185105 517067 185117 517101
rect 185151 517067 185163 517101
rect 185878 517083 185948 517284
rect 186301 517282 186631 517352
rect 186301 517248 186379 517282
rect 186413 517248 186478 517282
rect 186512 517248 186577 517282
rect 186611 517248 186631 517282
rect 186665 517284 186685 517318
rect 186719 517284 186788 517318
rect 186822 517284 186891 517318
rect 186925 517284 187003 517318
rect 186665 517214 187003 517284
rect 186301 517174 187003 517214
rect 186301 517140 186319 517174
rect 186353 517140 186951 517174
rect 186985 517140 187003 517174
rect 185105 516996 185163 517067
rect 185197 517072 186266 517083
rect 185197 517038 185215 517072
rect 185249 517038 186215 517072
rect 186249 517038 186266 517072
rect 185197 516996 186266 517038
rect 186301 517072 187003 517140
rect 186301 517038 186319 517072
rect 186353 517038 186951 517072
rect 186985 517038 187003 517072
rect 186301 516996 187003 517038
rect 187221 517288 187271 517322
rect 187305 517288 187325 517322
rect 187221 517214 187325 517288
rect 187359 517282 187463 517356
rect 187359 517248 187379 517282
rect 187413 517248 187463 517282
rect 187221 517167 187463 517214
rect 187221 517133 187239 517167
rect 187273 517133 187411 517167
rect 187445 517133 187463 517167
rect 187221 517072 187463 517133
rect 187221 517038 187239 517072
rect 187273 517038 187411 517072
rect 187445 517038 187463 517072
rect 187221 516996 187463 517038
rect 172208 516962 172237 516996
rect 172271 516962 172329 516996
rect 172363 516962 172421 516996
rect 172455 516962 172513 516996
rect 172547 516962 172605 516996
rect 172639 516962 172697 516996
rect 172731 516962 172789 516996
rect 172823 516962 172881 516996
rect 172915 516962 172973 516996
rect 173007 516962 173065 516996
rect 173099 516962 173157 516996
rect 173191 516962 173249 516996
rect 173283 516962 173341 516996
rect 173375 516962 173433 516996
rect 173467 516962 173525 516996
rect 173559 516962 173617 516996
rect 173651 516962 173709 516996
rect 173743 516962 173801 516996
rect 173835 516962 173893 516996
rect 173927 516962 173985 516996
rect 174019 516962 174077 516996
rect 174111 516962 174169 516996
rect 174203 516962 174261 516996
rect 174295 516962 174353 516996
rect 174387 516962 174445 516996
rect 174479 516962 174537 516996
rect 174571 516962 174629 516996
rect 174663 516962 174721 516996
rect 174755 516962 174813 516996
rect 174847 516962 174905 516996
rect 174939 516962 174997 516996
rect 175031 516962 175089 516996
rect 175123 516962 175181 516996
rect 175215 516962 175273 516996
rect 175307 516962 175365 516996
rect 175399 516962 175457 516996
rect 175491 516962 175549 516996
rect 175583 516962 175641 516996
rect 175675 516962 175733 516996
rect 175767 516962 175825 516996
rect 175859 516962 175917 516996
rect 175951 516962 176009 516996
rect 176043 516962 176101 516996
rect 176135 516962 176193 516996
rect 176227 516962 176285 516996
rect 176319 516962 176377 516996
rect 176411 516962 176469 516996
rect 176503 516962 176561 516996
rect 176595 516962 176653 516996
rect 176687 516962 176745 516996
rect 176779 516962 176837 516996
rect 176871 516962 176929 516996
rect 176963 516962 177021 516996
rect 177055 516962 177113 516996
rect 177147 516962 177205 516996
rect 177239 516962 177297 516996
rect 177331 516962 177389 516996
rect 177423 516962 177481 516996
rect 177515 516962 177573 516996
rect 177607 516962 177665 516996
rect 177699 516962 177757 516996
rect 177791 516962 177849 516996
rect 177883 516962 177941 516996
rect 177975 516962 178033 516996
rect 178067 516962 178125 516996
rect 178159 516962 178217 516996
rect 178251 516962 178309 516996
rect 178343 516962 178401 516996
rect 178435 516962 178493 516996
rect 178527 516962 178585 516996
rect 178619 516962 178677 516996
rect 178711 516962 178769 516996
rect 178803 516962 178861 516996
rect 178895 516962 178953 516996
rect 178987 516962 179045 516996
rect 179079 516962 179137 516996
rect 179171 516962 179229 516996
rect 179263 516962 179321 516996
rect 179355 516962 179413 516996
rect 179447 516962 179505 516996
rect 179539 516962 179597 516996
rect 179631 516962 179689 516996
rect 179723 516962 179781 516996
rect 179815 516962 179873 516996
rect 179907 516962 179965 516996
rect 179999 516962 180057 516996
rect 180091 516962 180149 516996
rect 180183 516962 180241 516996
rect 180275 516962 180333 516996
rect 180367 516962 180425 516996
rect 180459 516962 180517 516996
rect 180551 516962 180609 516996
rect 180643 516962 180701 516996
rect 180735 516962 180793 516996
rect 180827 516962 180885 516996
rect 180919 516962 180977 516996
rect 181011 516962 181069 516996
rect 181103 516962 181161 516996
rect 181195 516962 181253 516996
rect 181287 516962 181345 516996
rect 181379 516962 181437 516996
rect 181471 516962 181529 516996
rect 181563 516962 181621 516996
rect 181655 516962 181713 516996
rect 181747 516962 181805 516996
rect 181839 516962 181897 516996
rect 181931 516962 181989 516996
rect 182023 516962 182081 516996
rect 182115 516962 182173 516996
rect 182207 516962 182265 516996
rect 182299 516962 182357 516996
rect 182391 516962 182449 516996
rect 182483 516962 182541 516996
rect 182575 516962 182633 516996
rect 182667 516962 182725 516996
rect 182759 516962 182817 516996
rect 182851 516962 182909 516996
rect 182943 516962 183001 516996
rect 183035 516962 183093 516996
rect 183127 516962 183185 516996
rect 183219 516962 183277 516996
rect 183311 516962 183369 516996
rect 183403 516962 183461 516996
rect 183495 516962 183553 516996
rect 183587 516962 183645 516996
rect 183679 516962 183737 516996
rect 183771 516962 183829 516996
rect 183863 516962 183921 516996
rect 183955 516962 184013 516996
rect 184047 516962 184105 516996
rect 184139 516962 184197 516996
rect 184231 516962 184289 516996
rect 184323 516962 184381 516996
rect 184415 516962 184473 516996
rect 184507 516962 184565 516996
rect 184599 516962 184657 516996
rect 184691 516962 184749 516996
rect 184783 516962 184841 516996
rect 184875 516962 184933 516996
rect 184967 516962 185025 516996
rect 185059 516962 185117 516996
rect 185151 516962 185209 516996
rect 185243 516962 185301 516996
rect 185335 516962 185393 516996
rect 185427 516962 185485 516996
rect 185519 516962 185577 516996
rect 185611 516962 185669 516996
rect 185703 516962 185761 516996
rect 185795 516962 185853 516996
rect 185887 516962 185945 516996
rect 185979 516962 186037 516996
rect 186071 516962 186129 516996
rect 186163 516962 186221 516996
rect 186255 516962 186313 516996
rect 186347 516962 186405 516996
rect 186439 516962 186497 516996
rect 186531 516962 186589 516996
rect 186623 516962 186681 516996
rect 186715 516962 186773 516996
rect 186807 516962 186865 516996
rect 186899 516962 186957 516996
rect 186991 516962 187049 516996
rect 187083 516962 187141 516996
rect 187175 516962 187233 516996
rect 187267 516962 187325 516996
rect 187359 516962 187417 516996
rect 187451 516962 187480 516996
rect 172225 516920 172467 516962
rect 172225 516886 172243 516920
rect 172277 516886 172415 516920
rect 172449 516886 172467 516920
rect 172225 516825 172467 516886
rect 172501 516920 173570 516962
rect 172501 516886 172519 516920
rect 172553 516886 173519 516920
rect 173553 516886 173570 516920
rect 172501 516875 173570 516886
rect 173605 516920 174674 516962
rect 173605 516886 173623 516920
rect 173657 516886 174623 516920
rect 174657 516886 174674 516920
rect 173605 516875 174674 516886
rect 174709 516920 175778 516962
rect 174709 516886 174727 516920
rect 174761 516886 175727 516920
rect 175761 516886 175778 516920
rect 174709 516875 175778 516886
rect 175813 516920 176882 516962
rect 175813 516886 175831 516920
rect 175865 516886 176831 516920
rect 176865 516886 176882 516920
rect 175813 516875 176882 516886
rect 176917 516920 177251 516962
rect 176917 516886 176935 516920
rect 176969 516886 177199 516920
rect 177233 516886 177251 516920
rect 172225 516791 172243 516825
rect 172277 516791 172415 516825
rect 172449 516791 172467 516825
rect 172225 516744 172467 516791
rect 172225 516676 172275 516710
rect 172309 516676 172329 516710
rect 172225 516602 172329 516676
rect 172363 516670 172467 516744
rect 172363 516636 172383 516670
rect 172417 516636 172467 516670
rect 172818 516710 172886 516727
rect 172818 516676 172835 516710
rect 172869 516676 172886 516710
rect 172225 516549 172467 516602
rect 172818 516561 172886 516676
rect 173182 516674 173252 516875
rect 173182 516640 173199 516674
rect 173233 516640 173252 516674
rect 173182 516625 173252 516640
rect 173922 516710 173990 516727
rect 173922 516676 173939 516710
rect 173973 516676 173990 516710
rect 173922 516561 173990 516676
rect 174286 516674 174356 516875
rect 174286 516640 174303 516674
rect 174337 516640 174356 516674
rect 174286 516625 174356 516640
rect 175026 516710 175094 516727
rect 175026 516676 175043 516710
rect 175077 516676 175094 516710
rect 175026 516561 175094 516676
rect 175390 516674 175460 516875
rect 175390 516640 175407 516674
rect 175441 516640 175460 516674
rect 175390 516625 175460 516640
rect 176130 516710 176198 516727
rect 176130 516676 176147 516710
rect 176181 516676 176198 516710
rect 176130 516561 176198 516676
rect 176494 516674 176564 516875
rect 176917 516818 177251 516886
rect 176917 516784 176935 516818
rect 176969 516784 177199 516818
rect 177233 516784 177251 516818
rect 176917 516744 177251 516784
rect 176494 516640 176511 516674
rect 176545 516640 176564 516674
rect 176494 516625 176564 516640
rect 176917 516676 176937 516710
rect 176971 516676 177067 516710
rect 176917 516606 177067 516676
rect 177101 516674 177251 516744
rect 177377 516891 177435 516962
rect 177377 516857 177389 516891
rect 177423 516857 177435 516891
rect 177469 516920 178538 516962
rect 177469 516886 177487 516920
rect 177521 516886 178487 516920
rect 178521 516886 178538 516920
rect 177469 516875 178538 516886
rect 178573 516920 179642 516962
rect 178573 516886 178591 516920
rect 178625 516886 179591 516920
rect 179625 516886 179642 516920
rect 178573 516875 179642 516886
rect 179677 516920 180746 516962
rect 179677 516886 179695 516920
rect 179729 516886 180695 516920
rect 180729 516886 180746 516920
rect 179677 516875 180746 516886
rect 180781 516920 181850 516962
rect 180781 516886 180799 516920
rect 180833 516886 181799 516920
rect 181833 516886 181850 516920
rect 180781 516875 181850 516886
rect 181885 516920 182403 516962
rect 181885 516886 181903 516920
rect 181937 516886 182351 516920
rect 182385 516886 182403 516920
rect 177377 516798 177435 516857
rect 177377 516764 177389 516798
rect 177423 516764 177435 516798
rect 177377 516729 177435 516764
rect 177101 516640 177197 516674
rect 177231 516640 177251 516674
rect 177786 516710 177854 516727
rect 177786 516676 177803 516710
rect 177837 516676 177854 516710
rect 172225 516515 172243 516549
rect 172277 516515 172415 516549
rect 172449 516515 172467 516549
rect 172225 516452 172467 516515
rect 172501 516547 173570 516561
rect 172501 516513 172519 516547
rect 172553 516513 173519 516547
rect 173553 516513 173570 516547
rect 172501 516452 173570 516513
rect 173605 516547 174674 516561
rect 173605 516513 173623 516547
rect 173657 516513 174623 516547
rect 174657 516513 174674 516547
rect 173605 516452 174674 516513
rect 174709 516547 175778 516561
rect 174709 516513 174727 516547
rect 174761 516513 175727 516547
rect 175761 516513 175778 516547
rect 174709 516452 175778 516513
rect 175813 516547 176882 516561
rect 175813 516513 175831 516547
rect 175865 516513 176831 516547
rect 176865 516513 176882 516547
rect 175813 516452 176882 516513
rect 176917 516554 177251 516606
rect 176917 516520 176935 516554
rect 176969 516520 177199 516554
rect 177233 516520 177251 516554
rect 176917 516452 177251 516520
rect 177377 516580 177435 516597
rect 177377 516546 177389 516580
rect 177423 516546 177435 516580
rect 177786 516561 177854 516676
rect 178150 516674 178220 516875
rect 178150 516640 178167 516674
rect 178201 516640 178220 516674
rect 178150 516625 178220 516640
rect 178890 516710 178958 516727
rect 178890 516676 178907 516710
rect 178941 516676 178958 516710
rect 178890 516561 178958 516676
rect 179254 516674 179324 516875
rect 179254 516640 179271 516674
rect 179305 516640 179324 516674
rect 179254 516625 179324 516640
rect 179994 516710 180062 516727
rect 179994 516676 180011 516710
rect 180045 516676 180062 516710
rect 179994 516561 180062 516676
rect 180358 516674 180428 516875
rect 180358 516640 180375 516674
rect 180409 516640 180428 516674
rect 180358 516625 180428 516640
rect 181098 516710 181166 516727
rect 181098 516676 181115 516710
rect 181149 516676 181166 516710
rect 181098 516561 181166 516676
rect 181462 516674 181532 516875
rect 181885 516818 182403 516886
rect 181885 516784 181903 516818
rect 181937 516784 182351 516818
rect 182385 516784 182403 516818
rect 181885 516744 182403 516784
rect 181462 516640 181479 516674
rect 181513 516640 181532 516674
rect 181462 516625 181532 516640
rect 181885 516676 181963 516710
rect 181997 516676 182073 516710
rect 182107 516676 182127 516710
rect 181885 516606 182127 516676
rect 182161 516674 182403 516744
rect 182529 516891 182587 516962
rect 182529 516857 182541 516891
rect 182575 516857 182587 516891
rect 182621 516920 183690 516962
rect 182621 516886 182639 516920
rect 182673 516886 183639 516920
rect 183673 516886 183690 516920
rect 182621 516875 183690 516886
rect 183725 516920 184794 516962
rect 183725 516886 183743 516920
rect 183777 516886 184743 516920
rect 184777 516886 184794 516920
rect 183725 516875 184794 516886
rect 184829 516920 185898 516962
rect 184829 516886 184847 516920
rect 184881 516886 185847 516920
rect 185881 516886 185898 516920
rect 184829 516875 185898 516886
rect 185933 516920 187002 516962
rect 185933 516886 185951 516920
rect 185985 516886 186951 516920
rect 186985 516886 187002 516920
rect 185933 516875 187002 516886
rect 187221 516920 187463 516962
rect 187221 516886 187239 516920
rect 187273 516886 187411 516920
rect 187445 516886 187463 516920
rect 182529 516798 182587 516857
rect 182529 516764 182541 516798
rect 182575 516764 182587 516798
rect 182529 516729 182587 516764
rect 182161 516640 182181 516674
rect 182215 516640 182291 516674
rect 182325 516640 182403 516674
rect 182938 516710 183006 516727
rect 182938 516676 182955 516710
rect 182989 516676 183006 516710
rect 177377 516452 177435 516546
rect 177469 516547 178538 516561
rect 177469 516513 177487 516547
rect 177521 516513 178487 516547
rect 178521 516513 178538 516547
rect 177469 516452 178538 516513
rect 178573 516547 179642 516561
rect 178573 516513 178591 516547
rect 178625 516513 179591 516547
rect 179625 516513 179642 516547
rect 178573 516452 179642 516513
rect 179677 516547 180746 516561
rect 179677 516513 179695 516547
rect 179729 516513 180695 516547
rect 180729 516513 180746 516547
rect 179677 516452 180746 516513
rect 180781 516547 181850 516561
rect 180781 516513 180799 516547
rect 180833 516513 181799 516547
rect 181833 516513 181850 516547
rect 180781 516452 181850 516513
rect 181885 516547 182403 516606
rect 181885 516513 181903 516547
rect 181937 516513 182351 516547
rect 182385 516513 182403 516547
rect 181885 516452 182403 516513
rect 182529 516580 182587 516597
rect 182529 516546 182541 516580
rect 182575 516546 182587 516580
rect 182938 516561 183006 516676
rect 183302 516674 183372 516875
rect 183302 516640 183319 516674
rect 183353 516640 183372 516674
rect 183302 516625 183372 516640
rect 184042 516710 184110 516727
rect 184042 516676 184059 516710
rect 184093 516676 184110 516710
rect 184042 516561 184110 516676
rect 184406 516674 184476 516875
rect 184406 516640 184423 516674
rect 184457 516640 184476 516674
rect 184406 516625 184476 516640
rect 185146 516710 185214 516727
rect 185146 516676 185163 516710
rect 185197 516676 185214 516710
rect 185146 516561 185214 516676
rect 185510 516674 185580 516875
rect 185510 516640 185527 516674
rect 185561 516640 185580 516674
rect 185510 516625 185580 516640
rect 186250 516710 186318 516727
rect 186250 516676 186267 516710
rect 186301 516676 186318 516710
rect 186250 516561 186318 516676
rect 186614 516674 186684 516875
rect 186614 516640 186631 516674
rect 186665 516640 186684 516674
rect 186614 516625 186684 516640
rect 187221 516825 187463 516886
rect 187221 516791 187239 516825
rect 187273 516791 187411 516825
rect 187445 516791 187463 516825
rect 187221 516744 187463 516791
rect 187221 516670 187325 516744
rect 187221 516636 187271 516670
rect 187305 516636 187325 516670
rect 187359 516676 187379 516710
rect 187413 516676 187463 516710
rect 187359 516602 187463 516676
rect 182529 516452 182587 516546
rect 182621 516547 183690 516561
rect 182621 516513 182639 516547
rect 182673 516513 183639 516547
rect 183673 516513 183690 516547
rect 182621 516452 183690 516513
rect 183725 516547 184794 516561
rect 183725 516513 183743 516547
rect 183777 516513 184743 516547
rect 184777 516513 184794 516547
rect 183725 516452 184794 516513
rect 184829 516547 185898 516561
rect 184829 516513 184847 516547
rect 184881 516513 185847 516547
rect 185881 516513 185898 516547
rect 184829 516452 185898 516513
rect 185933 516547 187002 516561
rect 185933 516513 185951 516547
rect 185985 516513 186951 516547
rect 186985 516513 187002 516547
rect 185933 516452 187002 516513
rect 187221 516549 187463 516602
rect 187221 516515 187239 516549
rect 187273 516515 187411 516549
rect 187445 516515 187463 516549
rect 187221 516452 187463 516515
rect 172208 516418 172237 516452
rect 172271 516418 172329 516452
rect 172363 516418 172421 516452
rect 172455 516418 172513 516452
rect 172547 516418 172605 516452
rect 172639 516418 172697 516452
rect 172731 516418 172789 516452
rect 172823 516418 172881 516452
rect 172915 516418 172973 516452
rect 173007 516418 173065 516452
rect 173099 516418 173157 516452
rect 173191 516418 173249 516452
rect 173283 516418 173341 516452
rect 173375 516418 173433 516452
rect 173467 516418 173525 516452
rect 173559 516418 173617 516452
rect 173651 516418 173709 516452
rect 173743 516418 173801 516452
rect 173835 516418 173893 516452
rect 173927 516418 173985 516452
rect 174019 516418 174077 516452
rect 174111 516418 174169 516452
rect 174203 516418 174261 516452
rect 174295 516418 174353 516452
rect 174387 516418 174445 516452
rect 174479 516418 174537 516452
rect 174571 516418 174629 516452
rect 174663 516418 174721 516452
rect 174755 516418 174813 516452
rect 174847 516418 174905 516452
rect 174939 516418 174997 516452
rect 175031 516418 175089 516452
rect 175123 516418 175181 516452
rect 175215 516418 175273 516452
rect 175307 516418 175365 516452
rect 175399 516418 175457 516452
rect 175491 516418 175549 516452
rect 175583 516418 175641 516452
rect 175675 516418 175733 516452
rect 175767 516418 175825 516452
rect 175859 516418 175917 516452
rect 175951 516418 176009 516452
rect 176043 516418 176101 516452
rect 176135 516418 176193 516452
rect 176227 516418 176285 516452
rect 176319 516418 176377 516452
rect 176411 516418 176469 516452
rect 176503 516418 176561 516452
rect 176595 516418 176653 516452
rect 176687 516418 176745 516452
rect 176779 516418 176837 516452
rect 176871 516418 176929 516452
rect 176963 516418 177021 516452
rect 177055 516418 177113 516452
rect 177147 516418 177205 516452
rect 177239 516418 177297 516452
rect 177331 516418 177389 516452
rect 177423 516418 177481 516452
rect 177515 516418 177573 516452
rect 177607 516418 177665 516452
rect 177699 516418 177757 516452
rect 177791 516418 177849 516452
rect 177883 516418 177941 516452
rect 177975 516418 178033 516452
rect 178067 516418 178125 516452
rect 178159 516418 178217 516452
rect 178251 516418 178309 516452
rect 178343 516418 178401 516452
rect 178435 516418 178493 516452
rect 178527 516418 178585 516452
rect 178619 516418 178677 516452
rect 178711 516418 178769 516452
rect 178803 516418 178861 516452
rect 178895 516418 178953 516452
rect 178987 516418 179045 516452
rect 179079 516418 179137 516452
rect 179171 516418 179229 516452
rect 179263 516418 179321 516452
rect 179355 516418 179413 516452
rect 179447 516418 179505 516452
rect 179539 516418 179597 516452
rect 179631 516418 179689 516452
rect 179723 516418 179781 516452
rect 179815 516418 179873 516452
rect 179907 516418 179965 516452
rect 179999 516418 180057 516452
rect 180091 516418 180149 516452
rect 180183 516418 180241 516452
rect 180275 516418 180333 516452
rect 180367 516418 180425 516452
rect 180459 516418 180517 516452
rect 180551 516418 180609 516452
rect 180643 516418 180701 516452
rect 180735 516418 180793 516452
rect 180827 516418 180885 516452
rect 180919 516418 180977 516452
rect 181011 516418 181069 516452
rect 181103 516418 181161 516452
rect 181195 516418 181253 516452
rect 181287 516418 181345 516452
rect 181379 516418 181437 516452
rect 181471 516418 181529 516452
rect 181563 516418 181621 516452
rect 181655 516418 181713 516452
rect 181747 516418 181805 516452
rect 181839 516418 181897 516452
rect 181931 516418 181989 516452
rect 182023 516418 182081 516452
rect 182115 516418 182173 516452
rect 182207 516418 182265 516452
rect 182299 516418 182357 516452
rect 182391 516418 182449 516452
rect 182483 516418 182541 516452
rect 182575 516418 182633 516452
rect 182667 516418 182725 516452
rect 182759 516418 182817 516452
rect 182851 516418 182909 516452
rect 182943 516418 183001 516452
rect 183035 516418 183093 516452
rect 183127 516418 183185 516452
rect 183219 516418 183277 516452
rect 183311 516418 183369 516452
rect 183403 516418 183461 516452
rect 183495 516418 183553 516452
rect 183587 516418 183645 516452
rect 183679 516418 183737 516452
rect 183771 516418 183829 516452
rect 183863 516418 183921 516452
rect 183955 516418 184013 516452
rect 184047 516418 184105 516452
rect 184139 516418 184197 516452
rect 184231 516418 184289 516452
rect 184323 516418 184381 516452
rect 184415 516418 184473 516452
rect 184507 516418 184565 516452
rect 184599 516418 184657 516452
rect 184691 516418 184749 516452
rect 184783 516418 184841 516452
rect 184875 516418 184933 516452
rect 184967 516418 185025 516452
rect 185059 516418 185117 516452
rect 185151 516418 185209 516452
rect 185243 516418 185301 516452
rect 185335 516418 185393 516452
rect 185427 516418 185485 516452
rect 185519 516418 185577 516452
rect 185611 516418 185669 516452
rect 185703 516418 185761 516452
rect 185795 516418 185853 516452
rect 185887 516418 185945 516452
rect 185979 516418 186037 516452
rect 186071 516418 186129 516452
rect 186163 516418 186221 516452
rect 186255 516418 186313 516452
rect 186347 516418 186405 516452
rect 186439 516418 186497 516452
rect 186531 516418 186589 516452
rect 186623 516418 186681 516452
rect 186715 516418 186773 516452
rect 186807 516418 186865 516452
rect 186899 516418 186957 516452
rect 186991 516418 187049 516452
rect 187083 516418 187141 516452
rect 187175 516418 187233 516452
rect 187267 516418 187325 516452
rect 187359 516418 187417 516452
rect 187451 516418 187480 516452
rect 172225 516355 172467 516418
rect 172225 516321 172243 516355
rect 172277 516321 172415 516355
rect 172449 516321 172467 516355
rect 172225 516268 172467 516321
rect 172501 516357 173570 516418
rect 172501 516323 172519 516357
rect 172553 516323 173519 516357
rect 173553 516323 173570 516357
rect 172501 516309 173570 516323
rect 173605 516357 174674 516418
rect 173605 516323 173623 516357
rect 173657 516323 174623 516357
rect 174657 516323 174674 516357
rect 173605 516309 174674 516323
rect 174801 516324 174859 516418
rect 172225 516194 172329 516268
rect 172225 516160 172275 516194
rect 172309 516160 172329 516194
rect 172363 516200 172383 516234
rect 172417 516200 172467 516234
rect 172363 516126 172467 516200
rect 172818 516194 172886 516309
rect 172818 516160 172835 516194
rect 172869 516160 172886 516194
rect 172818 516143 172886 516160
rect 173182 516230 173252 516245
rect 173182 516196 173199 516230
rect 173233 516196 173252 516230
rect 172225 516079 172467 516126
rect 172225 516045 172243 516079
rect 172277 516045 172415 516079
rect 172449 516045 172467 516079
rect 172225 515984 172467 516045
rect 173182 515995 173252 516196
rect 173922 516194 173990 516309
rect 174801 516290 174813 516324
rect 174847 516290 174859 516324
rect 174893 516357 175962 516418
rect 174893 516323 174911 516357
rect 174945 516323 175911 516357
rect 175945 516323 175962 516357
rect 174893 516309 175962 516323
rect 175997 516357 177066 516418
rect 175997 516323 176015 516357
rect 176049 516323 177015 516357
rect 177049 516323 177066 516357
rect 175997 516309 177066 516323
rect 177101 516357 178170 516418
rect 177101 516323 177119 516357
rect 177153 516323 178119 516357
rect 178153 516323 178170 516357
rect 177101 516309 178170 516323
rect 178205 516357 179274 516418
rect 178205 516323 178223 516357
rect 178257 516323 179223 516357
rect 179257 516323 179274 516357
rect 178205 516309 179274 516323
rect 179309 516357 179827 516418
rect 179309 516323 179327 516357
rect 179361 516323 179775 516357
rect 179809 516323 179827 516357
rect 174801 516273 174859 516290
rect 173922 516160 173939 516194
rect 173973 516160 173990 516194
rect 173922 516143 173990 516160
rect 174286 516230 174356 516245
rect 174286 516196 174303 516230
rect 174337 516196 174356 516230
rect 174286 515995 174356 516196
rect 175210 516194 175278 516309
rect 175210 516160 175227 516194
rect 175261 516160 175278 516194
rect 175210 516143 175278 516160
rect 175574 516230 175644 516245
rect 175574 516196 175591 516230
rect 175625 516196 175644 516230
rect 174801 516106 174859 516141
rect 174801 516072 174813 516106
rect 174847 516072 174859 516106
rect 174801 516013 174859 516072
rect 172225 515950 172243 515984
rect 172277 515950 172415 515984
rect 172449 515950 172467 515984
rect 172225 515908 172467 515950
rect 172501 515984 173570 515995
rect 172501 515950 172519 515984
rect 172553 515950 173519 515984
rect 173553 515950 173570 515984
rect 172501 515908 173570 515950
rect 173605 515984 174674 515995
rect 173605 515950 173623 515984
rect 173657 515950 174623 515984
rect 174657 515950 174674 515984
rect 173605 515908 174674 515950
rect 174801 515979 174813 516013
rect 174847 515979 174859 516013
rect 175574 515995 175644 516196
rect 176314 516194 176382 516309
rect 176314 516160 176331 516194
rect 176365 516160 176382 516194
rect 176314 516143 176382 516160
rect 176678 516230 176748 516245
rect 176678 516196 176695 516230
rect 176729 516196 176748 516230
rect 176678 515995 176748 516196
rect 177418 516194 177486 516309
rect 177418 516160 177435 516194
rect 177469 516160 177486 516194
rect 177418 516143 177486 516160
rect 177782 516230 177852 516245
rect 177782 516196 177799 516230
rect 177833 516196 177852 516230
rect 177782 515995 177852 516196
rect 178522 516194 178590 516309
rect 179309 516264 179827 516323
rect 179953 516324 180011 516418
rect 179953 516290 179965 516324
rect 179999 516290 180011 516324
rect 180045 516357 181114 516418
rect 180045 516323 180063 516357
rect 180097 516323 181063 516357
rect 181097 516323 181114 516357
rect 180045 516309 181114 516323
rect 181149 516357 182218 516418
rect 181149 516323 181167 516357
rect 181201 516323 182167 516357
rect 182201 516323 182218 516357
rect 181149 516309 182218 516323
rect 182253 516357 183322 516418
rect 182253 516323 182271 516357
rect 182305 516323 183271 516357
rect 183305 516323 183322 516357
rect 182253 516309 183322 516323
rect 183357 516357 184426 516418
rect 183357 516323 183375 516357
rect 183409 516323 184375 516357
rect 184409 516323 184426 516357
rect 183357 516309 184426 516323
rect 184461 516357 184979 516418
rect 184461 516323 184479 516357
rect 184513 516323 184927 516357
rect 184961 516323 184979 516357
rect 179953 516273 180011 516290
rect 178522 516160 178539 516194
rect 178573 516160 178590 516194
rect 178522 516143 178590 516160
rect 178886 516230 178956 516245
rect 178886 516196 178903 516230
rect 178937 516196 178956 516230
rect 178886 515995 178956 516196
rect 179309 516194 179551 516264
rect 179309 516160 179387 516194
rect 179421 516160 179497 516194
rect 179531 516160 179551 516194
rect 179585 516196 179605 516230
rect 179639 516196 179715 516230
rect 179749 516196 179827 516230
rect 179585 516126 179827 516196
rect 180362 516194 180430 516309
rect 180362 516160 180379 516194
rect 180413 516160 180430 516194
rect 180362 516143 180430 516160
rect 180726 516230 180796 516245
rect 180726 516196 180743 516230
rect 180777 516196 180796 516230
rect 179309 516086 179827 516126
rect 179309 516052 179327 516086
rect 179361 516052 179775 516086
rect 179809 516052 179827 516086
rect 174801 515908 174859 515979
rect 174893 515984 175962 515995
rect 174893 515950 174911 515984
rect 174945 515950 175911 515984
rect 175945 515950 175962 515984
rect 174893 515908 175962 515950
rect 175997 515984 177066 515995
rect 175997 515950 176015 515984
rect 176049 515950 177015 515984
rect 177049 515950 177066 515984
rect 175997 515908 177066 515950
rect 177101 515984 178170 515995
rect 177101 515950 177119 515984
rect 177153 515950 178119 515984
rect 178153 515950 178170 515984
rect 177101 515908 178170 515950
rect 178205 515984 179274 515995
rect 178205 515950 178223 515984
rect 178257 515950 179223 515984
rect 179257 515950 179274 515984
rect 178205 515908 179274 515950
rect 179309 515984 179827 516052
rect 179309 515950 179327 515984
rect 179361 515950 179775 515984
rect 179809 515950 179827 515984
rect 179309 515908 179827 515950
rect 179953 516106 180011 516141
rect 179953 516072 179965 516106
rect 179999 516072 180011 516106
rect 179953 516013 180011 516072
rect 179953 515979 179965 516013
rect 179999 515979 180011 516013
rect 180726 515995 180796 516196
rect 181466 516194 181534 516309
rect 181466 516160 181483 516194
rect 181517 516160 181534 516194
rect 181466 516143 181534 516160
rect 181830 516230 181900 516245
rect 181830 516196 181847 516230
rect 181881 516196 181900 516230
rect 181830 515995 181900 516196
rect 182570 516194 182638 516309
rect 182570 516160 182587 516194
rect 182621 516160 182638 516194
rect 182570 516143 182638 516160
rect 182934 516230 183004 516245
rect 182934 516196 182951 516230
rect 182985 516196 183004 516230
rect 182934 515995 183004 516196
rect 183674 516194 183742 516309
rect 184461 516264 184979 516323
rect 185105 516324 185163 516418
rect 185105 516290 185117 516324
rect 185151 516290 185163 516324
rect 185197 516357 186266 516418
rect 185197 516323 185215 516357
rect 185249 516323 186215 516357
rect 186249 516323 186266 516357
rect 185197 516309 186266 516323
rect 186301 516357 187003 516418
rect 186301 516323 186319 516357
rect 186353 516323 186951 516357
rect 186985 516323 187003 516357
rect 185105 516273 185163 516290
rect 183674 516160 183691 516194
rect 183725 516160 183742 516194
rect 183674 516143 183742 516160
rect 184038 516230 184108 516245
rect 184038 516196 184055 516230
rect 184089 516196 184108 516230
rect 184038 515995 184108 516196
rect 184461 516194 184703 516264
rect 184461 516160 184539 516194
rect 184573 516160 184649 516194
rect 184683 516160 184703 516194
rect 184737 516196 184757 516230
rect 184791 516196 184867 516230
rect 184901 516196 184979 516230
rect 184737 516126 184979 516196
rect 185514 516194 185582 516309
rect 186301 516264 187003 516323
rect 187221 516355 187463 516418
rect 187221 516321 187239 516355
rect 187273 516321 187411 516355
rect 187445 516321 187463 516355
rect 187221 516268 187463 516321
rect 185514 516160 185531 516194
rect 185565 516160 185582 516194
rect 185514 516143 185582 516160
rect 185878 516230 185948 516245
rect 185878 516196 185895 516230
rect 185929 516196 185948 516230
rect 184461 516086 184979 516126
rect 184461 516052 184479 516086
rect 184513 516052 184927 516086
rect 184961 516052 184979 516086
rect 179953 515908 180011 515979
rect 180045 515984 181114 515995
rect 180045 515950 180063 515984
rect 180097 515950 181063 515984
rect 181097 515950 181114 515984
rect 180045 515908 181114 515950
rect 181149 515984 182218 515995
rect 181149 515950 181167 515984
rect 181201 515950 182167 515984
rect 182201 515950 182218 515984
rect 181149 515908 182218 515950
rect 182253 515984 183322 515995
rect 182253 515950 182271 515984
rect 182305 515950 183271 515984
rect 183305 515950 183322 515984
rect 182253 515908 183322 515950
rect 183357 515984 184426 515995
rect 183357 515950 183375 515984
rect 183409 515950 184375 515984
rect 184409 515950 184426 515984
rect 183357 515908 184426 515950
rect 184461 515984 184979 516052
rect 184461 515950 184479 515984
rect 184513 515950 184927 515984
rect 184961 515950 184979 515984
rect 184461 515908 184979 515950
rect 185105 516106 185163 516141
rect 185105 516072 185117 516106
rect 185151 516072 185163 516106
rect 185105 516013 185163 516072
rect 185105 515979 185117 516013
rect 185151 515979 185163 516013
rect 185878 515995 185948 516196
rect 186301 516194 186631 516264
rect 186301 516160 186379 516194
rect 186413 516160 186478 516194
rect 186512 516160 186577 516194
rect 186611 516160 186631 516194
rect 186665 516196 186685 516230
rect 186719 516196 186788 516230
rect 186822 516196 186891 516230
rect 186925 516196 187003 516230
rect 186665 516126 187003 516196
rect 186301 516086 187003 516126
rect 186301 516052 186319 516086
rect 186353 516052 186951 516086
rect 186985 516052 187003 516086
rect 185105 515908 185163 515979
rect 185197 515984 186266 515995
rect 185197 515950 185215 515984
rect 185249 515950 186215 515984
rect 186249 515950 186266 515984
rect 185197 515908 186266 515950
rect 186301 515984 187003 516052
rect 186301 515950 186319 515984
rect 186353 515950 186951 515984
rect 186985 515950 187003 515984
rect 186301 515908 187003 515950
rect 187221 516200 187271 516234
rect 187305 516200 187325 516234
rect 187221 516126 187325 516200
rect 187359 516194 187463 516268
rect 187359 516160 187379 516194
rect 187413 516160 187463 516194
rect 187221 516079 187463 516126
rect 187221 516045 187239 516079
rect 187273 516045 187411 516079
rect 187445 516045 187463 516079
rect 187221 515984 187463 516045
rect 187221 515950 187239 515984
rect 187273 515950 187411 515984
rect 187445 515950 187463 515984
rect 187221 515908 187463 515950
rect 172208 515874 172237 515908
rect 172271 515874 172329 515908
rect 172363 515874 172421 515908
rect 172455 515874 172513 515908
rect 172547 515874 172605 515908
rect 172639 515874 172697 515908
rect 172731 515874 172789 515908
rect 172823 515874 172881 515908
rect 172915 515874 172973 515908
rect 173007 515874 173065 515908
rect 173099 515874 173157 515908
rect 173191 515874 173249 515908
rect 173283 515874 173341 515908
rect 173375 515874 173433 515908
rect 173467 515874 173525 515908
rect 173559 515874 173617 515908
rect 173651 515874 173709 515908
rect 173743 515874 173801 515908
rect 173835 515874 173893 515908
rect 173927 515874 173985 515908
rect 174019 515874 174077 515908
rect 174111 515874 174169 515908
rect 174203 515874 174261 515908
rect 174295 515874 174353 515908
rect 174387 515874 174445 515908
rect 174479 515874 174537 515908
rect 174571 515874 174629 515908
rect 174663 515874 174721 515908
rect 174755 515874 174813 515908
rect 174847 515874 174905 515908
rect 174939 515874 174997 515908
rect 175031 515874 175089 515908
rect 175123 515874 175181 515908
rect 175215 515874 175273 515908
rect 175307 515874 175365 515908
rect 175399 515874 175457 515908
rect 175491 515874 175549 515908
rect 175583 515874 175641 515908
rect 175675 515874 175733 515908
rect 175767 515874 175825 515908
rect 175859 515874 175917 515908
rect 175951 515874 176009 515908
rect 176043 515874 176101 515908
rect 176135 515874 176193 515908
rect 176227 515874 176285 515908
rect 176319 515874 176377 515908
rect 176411 515874 176469 515908
rect 176503 515874 176561 515908
rect 176595 515874 176653 515908
rect 176687 515874 176745 515908
rect 176779 515874 176837 515908
rect 176871 515874 176929 515908
rect 176963 515874 177021 515908
rect 177055 515874 177113 515908
rect 177147 515874 177205 515908
rect 177239 515874 177297 515908
rect 177331 515874 177389 515908
rect 177423 515874 177481 515908
rect 177515 515874 177573 515908
rect 177607 515874 177665 515908
rect 177699 515874 177757 515908
rect 177791 515874 177849 515908
rect 177883 515874 177941 515908
rect 177975 515874 178033 515908
rect 178067 515874 178125 515908
rect 178159 515874 178217 515908
rect 178251 515874 178309 515908
rect 178343 515874 178401 515908
rect 178435 515874 178493 515908
rect 178527 515874 178585 515908
rect 178619 515874 178677 515908
rect 178711 515874 178769 515908
rect 178803 515874 178861 515908
rect 178895 515874 178953 515908
rect 178987 515874 179045 515908
rect 179079 515874 179137 515908
rect 179171 515874 179229 515908
rect 179263 515874 179321 515908
rect 179355 515874 179413 515908
rect 179447 515874 179505 515908
rect 179539 515874 179597 515908
rect 179631 515874 179689 515908
rect 179723 515874 179781 515908
rect 179815 515874 179873 515908
rect 179907 515874 179965 515908
rect 179999 515874 180057 515908
rect 180091 515874 180149 515908
rect 180183 515874 180241 515908
rect 180275 515874 180333 515908
rect 180367 515874 180425 515908
rect 180459 515874 180517 515908
rect 180551 515874 180609 515908
rect 180643 515874 180701 515908
rect 180735 515874 180793 515908
rect 180827 515874 180885 515908
rect 180919 515874 180977 515908
rect 181011 515874 181069 515908
rect 181103 515874 181161 515908
rect 181195 515874 181253 515908
rect 181287 515874 181345 515908
rect 181379 515874 181437 515908
rect 181471 515874 181529 515908
rect 181563 515874 181621 515908
rect 181655 515874 181713 515908
rect 181747 515874 181805 515908
rect 181839 515874 181897 515908
rect 181931 515874 181989 515908
rect 182023 515874 182081 515908
rect 182115 515874 182173 515908
rect 182207 515874 182265 515908
rect 182299 515874 182357 515908
rect 182391 515874 182449 515908
rect 182483 515874 182541 515908
rect 182575 515874 182633 515908
rect 182667 515874 182725 515908
rect 182759 515874 182817 515908
rect 182851 515874 182909 515908
rect 182943 515874 183001 515908
rect 183035 515874 183093 515908
rect 183127 515874 183185 515908
rect 183219 515874 183277 515908
rect 183311 515874 183369 515908
rect 183403 515874 183461 515908
rect 183495 515874 183553 515908
rect 183587 515874 183645 515908
rect 183679 515874 183737 515908
rect 183771 515874 183829 515908
rect 183863 515874 183921 515908
rect 183955 515874 184013 515908
rect 184047 515874 184105 515908
rect 184139 515874 184197 515908
rect 184231 515874 184289 515908
rect 184323 515874 184381 515908
rect 184415 515874 184473 515908
rect 184507 515874 184565 515908
rect 184599 515874 184657 515908
rect 184691 515874 184749 515908
rect 184783 515874 184841 515908
rect 184875 515874 184933 515908
rect 184967 515874 185025 515908
rect 185059 515874 185117 515908
rect 185151 515874 185209 515908
rect 185243 515874 185301 515908
rect 185335 515874 185393 515908
rect 185427 515874 185485 515908
rect 185519 515874 185577 515908
rect 185611 515874 185669 515908
rect 185703 515874 185761 515908
rect 185795 515874 185853 515908
rect 185887 515874 185945 515908
rect 185979 515874 186037 515908
rect 186071 515874 186129 515908
rect 186163 515874 186221 515908
rect 186255 515874 186313 515908
rect 186347 515874 186405 515908
rect 186439 515874 186497 515908
rect 186531 515874 186589 515908
rect 186623 515874 186681 515908
rect 186715 515874 186773 515908
rect 186807 515874 186865 515908
rect 186899 515874 186957 515908
rect 186991 515874 187049 515908
rect 187083 515874 187141 515908
rect 187175 515874 187233 515908
rect 187267 515874 187325 515908
rect 187359 515874 187417 515908
rect 187451 515874 187480 515908
rect 172225 515832 172467 515874
rect 172225 515798 172243 515832
rect 172277 515798 172415 515832
rect 172449 515798 172467 515832
rect 172225 515737 172467 515798
rect 172225 515703 172243 515737
rect 172277 515703 172415 515737
rect 172449 515703 172467 515737
rect 172225 515656 172467 515703
rect 172501 515832 173203 515874
rect 172501 515798 172519 515832
rect 172553 515798 173151 515832
rect 173185 515798 173203 515832
rect 172501 515730 173203 515798
rect 172501 515696 172519 515730
rect 172553 515696 173151 515730
rect 173185 515696 173203 515730
rect 172501 515656 173203 515696
rect 172225 515588 172275 515622
rect 172309 515588 172329 515622
rect 172225 515514 172329 515588
rect 172363 515582 172467 515656
rect 172363 515548 172383 515582
rect 172417 515548 172467 515582
rect 172501 515588 172579 515622
rect 172613 515588 172678 515622
rect 172712 515588 172777 515622
rect 172811 515588 172831 515622
rect 172501 515518 172831 515588
rect 172865 515586 173203 515656
rect 172865 515552 172885 515586
rect 172919 515552 172988 515586
rect 173022 515552 173091 515586
rect 173125 515552 173203 515586
rect 173421 515824 173483 515840
rect 173421 515790 173439 515824
rect 173473 515790 173483 515824
rect 173421 515702 173483 515790
rect 173517 515832 173579 515874
rect 173517 515798 173525 515832
rect 173559 515798 173579 515832
rect 173517 515764 173579 515798
rect 173517 515730 173525 515764
rect 173559 515730 173579 515764
rect 173517 515714 173579 515730
rect 173613 515806 173665 515840
rect 173613 515772 173617 515806
rect 173651 515797 173665 515806
rect 173613 515763 173621 515772
rect 173655 515763 173665 515797
rect 173699 515832 173750 515874
rect 173699 515798 173707 515832
rect 173741 515798 173750 515832
rect 173699 515782 173750 515798
rect 173785 515824 173837 515840
rect 173785 515790 173793 515824
rect 173827 515790 173837 515824
rect 173613 515748 173665 515763
rect 173785 515756 173837 515790
rect 173785 515748 173793 515756
rect 173613 515722 173793 515748
rect 173827 515722 173837 515756
rect 173613 515714 173837 515722
rect 173421 515668 173439 515702
rect 173473 515680 173483 515702
rect 173785 515688 173837 515714
rect 173871 515818 173928 515874
rect 173871 515784 173879 515818
rect 173913 515784 173928 515818
rect 173871 515750 173928 515784
rect 173871 515716 173879 515750
rect 173913 515716 173928 515750
rect 173871 515700 173928 515716
rect 173973 515832 174675 515874
rect 173973 515798 173991 515832
rect 174025 515798 174623 515832
rect 174657 515798 174675 515832
rect 173973 515730 174675 515798
rect 173473 515668 173627 515680
rect 173421 515646 173627 515668
rect 172225 515461 172467 515514
rect 172225 515427 172243 515461
rect 172277 515427 172415 515461
rect 172449 515427 172467 515461
rect 172225 515364 172467 515427
rect 172501 515459 173203 515518
rect 172501 515425 172519 515459
rect 172553 515425 173151 515459
rect 173185 515425 173203 515459
rect 172501 515364 173203 515425
rect 173421 515464 173455 515646
rect 173489 515596 173559 515612
rect 173523 515562 173559 515596
rect 173593 515596 173627 515646
rect 173785 515654 173793 515688
rect 173827 515664 173837 515688
rect 173973 515696 173991 515730
rect 174025 515696 174623 515730
rect 174657 515696 174675 515730
rect 173827 515654 173936 515664
rect 173973 515656 174675 515696
rect 173785 515630 173936 515654
rect 173593 515562 173635 515596
rect 173669 515562 173703 515596
rect 173737 515562 173771 515596
rect 173805 515562 173821 515596
rect 173489 515534 173559 515562
rect 173489 515500 173525 515534
rect 173855 515528 173936 515630
rect 173489 515498 173559 515500
rect 173606 515494 173936 515528
rect 173973 515588 174051 515622
rect 174085 515588 174150 515622
rect 174184 515588 174249 515622
rect 174283 515588 174303 515622
rect 173973 515518 174303 515588
rect 174337 515586 174675 515656
rect 174801 515803 174859 515874
rect 174801 515769 174813 515803
rect 174847 515769 174859 515803
rect 174893 515832 175962 515874
rect 174893 515798 174911 515832
rect 174945 515798 175911 515832
rect 175945 515798 175962 515832
rect 174893 515787 175962 515798
rect 175997 515832 177066 515874
rect 175997 515798 176015 515832
rect 176049 515798 177015 515832
rect 177049 515798 177066 515832
rect 175997 515787 177066 515798
rect 177101 515832 177343 515874
rect 177101 515798 177119 515832
rect 177153 515798 177291 515832
rect 177325 515798 177343 515832
rect 174801 515710 174859 515769
rect 174801 515676 174813 515710
rect 174847 515676 174859 515710
rect 174801 515641 174859 515676
rect 174337 515552 174357 515586
rect 174391 515552 174460 515586
rect 174494 515552 174563 515586
rect 174597 515552 174675 515586
rect 175210 515622 175278 515639
rect 175210 515588 175227 515622
rect 175261 515588 175278 515622
rect 173606 515466 173665 515494
rect 173421 515448 173481 515464
rect 173421 515414 173439 515448
rect 173473 515414 173481 515448
rect 173421 515398 173481 515414
rect 173515 515444 173570 515460
rect 173515 515410 173525 515444
rect 173559 515410 173570 515444
rect 173606 515432 173622 515466
rect 173656 515432 173665 515466
rect 173785 515466 173837 515494
rect 173606 515416 173665 515432
rect 173699 515444 173750 515460
rect 173515 515364 173570 515410
rect 173699 515410 173708 515444
rect 173742 515410 173750 515444
rect 173785 515432 173794 515466
rect 173828 515432 173837 515466
rect 173785 515416 173837 515432
rect 173871 515444 173927 515460
rect 173699 515364 173750 515410
rect 173871 515410 173880 515444
rect 173914 515410 173927 515444
rect 173871 515364 173927 515410
rect 173973 515459 174675 515518
rect 173973 515425 173991 515459
rect 174025 515425 174623 515459
rect 174657 515425 174675 515459
rect 173973 515364 174675 515425
rect 174801 515492 174859 515509
rect 174801 515458 174813 515492
rect 174847 515458 174859 515492
rect 175210 515473 175278 515588
rect 175574 515586 175644 515787
rect 175574 515552 175591 515586
rect 175625 515552 175644 515586
rect 175574 515537 175644 515552
rect 176314 515622 176382 515639
rect 176314 515588 176331 515622
rect 176365 515588 176382 515622
rect 176314 515473 176382 515588
rect 176678 515586 176748 515787
rect 177101 515737 177343 515798
rect 177101 515703 177119 515737
rect 177153 515703 177291 515737
rect 177325 515703 177343 515737
rect 177101 515656 177343 515703
rect 176678 515552 176695 515586
rect 176729 515552 176748 515586
rect 176678 515537 176748 515552
rect 177101 515588 177151 515622
rect 177185 515588 177205 515622
rect 177101 515514 177205 515588
rect 177239 515582 177343 515656
rect 177377 515803 177435 515874
rect 177377 515769 177389 515803
rect 177423 515769 177435 515803
rect 177469 515832 178538 515874
rect 177469 515798 177487 515832
rect 177521 515798 178487 515832
rect 178521 515798 178538 515832
rect 177469 515787 178538 515798
rect 178573 515832 179642 515874
rect 178573 515798 178591 515832
rect 178625 515798 179591 515832
rect 179625 515798 179642 515832
rect 178573 515787 179642 515798
rect 179677 515832 179919 515874
rect 179677 515798 179695 515832
rect 179729 515798 179867 515832
rect 179901 515798 179919 515832
rect 177377 515710 177435 515769
rect 177377 515676 177389 515710
rect 177423 515676 177435 515710
rect 177377 515641 177435 515676
rect 177239 515548 177259 515582
rect 177293 515548 177343 515582
rect 177786 515622 177854 515639
rect 177786 515588 177803 515622
rect 177837 515588 177854 515622
rect 174801 515364 174859 515458
rect 174893 515459 175962 515473
rect 174893 515425 174911 515459
rect 174945 515425 175911 515459
rect 175945 515425 175962 515459
rect 174893 515364 175962 515425
rect 175997 515459 177066 515473
rect 175997 515425 176015 515459
rect 176049 515425 177015 515459
rect 177049 515425 177066 515459
rect 175997 515364 177066 515425
rect 177101 515461 177343 515514
rect 177101 515427 177119 515461
rect 177153 515427 177291 515461
rect 177325 515427 177343 515461
rect 177101 515364 177343 515427
rect 177377 515492 177435 515509
rect 177377 515458 177389 515492
rect 177423 515458 177435 515492
rect 177786 515473 177854 515588
rect 178150 515586 178220 515787
rect 178150 515552 178167 515586
rect 178201 515552 178220 515586
rect 178150 515537 178220 515552
rect 178890 515622 178958 515639
rect 178890 515588 178907 515622
rect 178941 515588 178958 515622
rect 178890 515473 178958 515588
rect 179254 515586 179324 515787
rect 179677 515737 179919 515798
rect 179677 515703 179695 515737
rect 179729 515703 179867 515737
rect 179901 515703 179919 515737
rect 179677 515656 179919 515703
rect 179254 515552 179271 515586
rect 179305 515552 179324 515586
rect 179254 515537 179324 515552
rect 179677 515588 179727 515622
rect 179761 515588 179781 515622
rect 179677 515514 179781 515588
rect 179815 515582 179919 515656
rect 179953 515803 180011 515874
rect 179953 515769 179965 515803
rect 179999 515769 180011 515803
rect 180045 515832 181114 515874
rect 180045 515798 180063 515832
rect 180097 515798 181063 515832
rect 181097 515798 181114 515832
rect 180045 515787 181114 515798
rect 181149 515832 181851 515874
rect 181149 515798 181167 515832
rect 181201 515798 181799 515832
rect 181833 515798 181851 515832
rect 179953 515710 180011 515769
rect 179953 515676 179965 515710
rect 179999 515676 180011 515710
rect 179953 515641 180011 515676
rect 179815 515548 179835 515582
rect 179869 515548 179919 515582
rect 180362 515622 180430 515639
rect 180362 515588 180379 515622
rect 180413 515588 180430 515622
rect 177377 515364 177435 515458
rect 177469 515459 178538 515473
rect 177469 515425 177487 515459
rect 177521 515425 178487 515459
rect 178521 515425 178538 515459
rect 177469 515364 178538 515425
rect 178573 515459 179642 515473
rect 178573 515425 178591 515459
rect 178625 515425 179591 515459
rect 179625 515425 179642 515459
rect 178573 515364 179642 515425
rect 179677 515461 179919 515514
rect 179677 515427 179695 515461
rect 179729 515427 179867 515461
rect 179901 515427 179919 515461
rect 179677 515364 179919 515427
rect 179953 515492 180011 515509
rect 179953 515458 179965 515492
rect 179999 515458 180011 515492
rect 180362 515473 180430 515588
rect 180726 515586 180796 515787
rect 181149 515730 181851 515798
rect 181149 515696 181167 515730
rect 181201 515696 181799 515730
rect 181833 515696 181851 515730
rect 181149 515656 181851 515696
rect 180726 515552 180743 515586
rect 180777 515552 180796 515586
rect 180726 515537 180796 515552
rect 181149 515588 181227 515622
rect 181261 515588 181326 515622
rect 181360 515588 181425 515622
rect 181459 515588 181479 515622
rect 181149 515518 181479 515588
rect 181513 515586 181851 515656
rect 181513 515552 181533 515586
rect 181567 515552 181636 515586
rect 181670 515552 181739 515586
rect 181773 515552 181851 515586
rect 182069 515824 182123 515840
rect 182069 515806 182087 515824
rect 182069 515772 182081 515806
rect 182121 515790 182123 515824
rect 182115 515772 182123 515790
rect 182069 515743 182123 515772
rect 182069 515709 182087 515743
rect 182121 515709 182123 515743
rect 182157 515824 182223 515874
rect 182157 515790 182173 515824
rect 182207 515790 182223 515824
rect 182157 515756 182223 515790
rect 182157 515722 182173 515756
rect 182207 515722 182223 515756
rect 182259 515824 182295 515840
rect 182293 515790 182295 515824
rect 182259 515756 182295 515790
rect 182293 515722 182295 515756
rect 182069 515659 182123 515709
rect 182259 515688 182295 515722
rect 179953 515364 180011 515458
rect 180045 515459 181114 515473
rect 180045 515425 180063 515459
rect 180097 515425 181063 515459
rect 181097 515425 181114 515459
rect 180045 515364 181114 515425
rect 181149 515459 181851 515518
rect 181149 515425 181167 515459
rect 181201 515425 181799 515459
rect 181833 515425 181851 515459
rect 181149 515364 181851 515425
rect 182069 515499 182105 515659
rect 182160 515654 182295 515688
rect 182529 515803 182587 515874
rect 182529 515769 182541 515803
rect 182575 515769 182587 515803
rect 182621 515832 183690 515874
rect 182621 515798 182639 515832
rect 182673 515798 183639 515832
rect 183673 515798 183690 515832
rect 182621 515787 183690 515798
rect 183725 515832 184794 515874
rect 183725 515798 183743 515832
rect 183777 515798 184743 515832
rect 184777 515798 184794 515832
rect 183725 515787 184794 515798
rect 184829 515832 185071 515874
rect 184829 515798 184847 515832
rect 184881 515798 185019 515832
rect 185053 515798 185071 515832
rect 182529 515710 182587 515769
rect 182529 515676 182541 515710
rect 182575 515676 182587 515710
rect 182160 515625 182194 515654
rect 182529 515641 182587 515676
rect 182139 515609 182194 515625
rect 182938 515622 183006 515639
rect 182173 515575 182194 515609
rect 182139 515559 182194 515575
rect 182160 515508 182194 515559
rect 182239 515602 182307 515618
rect 182239 515596 182265 515602
rect 182239 515562 182257 515596
rect 182299 515568 182307 515602
rect 182291 515562 182307 515568
rect 182239 515544 182307 515562
rect 182938 515588 182955 515622
rect 182989 515588 183006 515622
rect 182069 515470 182121 515499
rect 182160 515474 182293 515508
rect 182069 515436 182087 515470
rect 182259 515453 182293 515474
rect 182069 515398 182121 515436
rect 182157 515406 182173 515440
rect 182207 515406 182223 515440
rect 182157 515364 182223 515406
rect 182259 515398 182293 515419
rect 182529 515492 182587 515509
rect 182529 515458 182541 515492
rect 182575 515458 182587 515492
rect 182938 515473 183006 515588
rect 183302 515586 183372 515787
rect 183302 515552 183319 515586
rect 183353 515552 183372 515586
rect 183302 515537 183372 515552
rect 184042 515622 184110 515639
rect 184042 515588 184059 515622
rect 184093 515588 184110 515622
rect 184042 515473 184110 515588
rect 184406 515586 184476 515787
rect 184829 515737 185071 515798
rect 184829 515703 184847 515737
rect 184881 515703 185019 515737
rect 185053 515703 185071 515737
rect 184829 515656 185071 515703
rect 184406 515552 184423 515586
rect 184457 515552 184476 515586
rect 184406 515537 184476 515552
rect 184829 515588 184879 515622
rect 184913 515588 184933 515622
rect 184829 515514 184933 515588
rect 184967 515582 185071 515656
rect 185105 515803 185163 515874
rect 185105 515769 185117 515803
rect 185151 515769 185163 515803
rect 185197 515832 186266 515874
rect 185197 515798 185215 515832
rect 185249 515798 186215 515832
rect 186249 515798 186266 515832
rect 185197 515787 186266 515798
rect 186393 515824 186455 515840
rect 186393 515790 186411 515824
rect 186445 515790 186455 515824
rect 185105 515710 185163 515769
rect 185105 515676 185117 515710
rect 185151 515676 185163 515710
rect 185105 515641 185163 515676
rect 184967 515548 184987 515582
rect 185021 515548 185071 515582
rect 185514 515622 185582 515639
rect 185514 515588 185531 515622
rect 185565 515588 185582 515622
rect 182529 515364 182587 515458
rect 182621 515459 183690 515473
rect 182621 515425 182639 515459
rect 182673 515425 183639 515459
rect 183673 515425 183690 515459
rect 182621 515364 183690 515425
rect 183725 515459 184794 515473
rect 183725 515425 183743 515459
rect 183777 515425 184743 515459
rect 184777 515425 184794 515459
rect 183725 515364 184794 515425
rect 184829 515461 185071 515514
rect 184829 515427 184847 515461
rect 184881 515427 185019 515461
rect 185053 515427 185071 515461
rect 184829 515364 185071 515427
rect 185105 515492 185163 515509
rect 185105 515458 185117 515492
rect 185151 515458 185163 515492
rect 185514 515473 185582 515588
rect 185878 515586 185948 515787
rect 185878 515552 185895 515586
rect 185929 515552 185948 515586
rect 185878 515537 185948 515552
rect 186393 515702 186455 515790
rect 186489 515832 186551 515874
rect 186489 515798 186497 515832
rect 186531 515798 186551 515832
rect 186489 515764 186551 515798
rect 186489 515730 186497 515764
rect 186531 515730 186551 515764
rect 186489 515714 186551 515730
rect 186585 515806 186637 515840
rect 186585 515772 186589 515806
rect 186623 515797 186637 515806
rect 186585 515763 186593 515772
rect 186627 515763 186637 515797
rect 186671 515832 186722 515874
rect 186671 515798 186679 515832
rect 186713 515798 186722 515832
rect 186671 515782 186722 515798
rect 186757 515824 186809 515840
rect 186757 515790 186765 515824
rect 186799 515790 186809 515824
rect 186585 515748 186637 515763
rect 186757 515756 186809 515790
rect 186757 515748 186765 515756
rect 186585 515722 186765 515748
rect 186799 515722 186809 515756
rect 186585 515714 186809 515722
rect 186393 515668 186411 515702
rect 186445 515680 186455 515702
rect 186757 515688 186809 515714
rect 186843 515818 186900 515874
rect 186843 515784 186851 515818
rect 186885 515784 186900 515818
rect 186843 515750 186900 515784
rect 186843 515716 186851 515750
rect 186885 515716 186900 515750
rect 186843 515700 186900 515716
rect 186945 515832 187187 515874
rect 186945 515798 186963 515832
rect 186997 515798 187135 515832
rect 187169 515798 187187 515832
rect 186945 515737 187187 515798
rect 186945 515703 186963 515737
rect 186997 515703 187135 515737
rect 187169 515703 187187 515737
rect 186445 515668 186599 515680
rect 186393 515646 186599 515668
rect 185105 515364 185163 515458
rect 185197 515459 186266 515473
rect 185197 515425 185215 515459
rect 185249 515425 186215 515459
rect 186249 515425 186266 515459
rect 185197 515364 186266 515425
rect 186393 515464 186427 515646
rect 186461 515596 186531 515612
rect 186495 515562 186531 515596
rect 186565 515596 186599 515646
rect 186757 515654 186765 515688
rect 186799 515664 186809 515688
rect 186799 515654 186908 515664
rect 186945 515656 187187 515703
rect 186757 515630 186908 515654
rect 186565 515562 186607 515596
rect 186641 515562 186675 515596
rect 186709 515562 186743 515596
rect 186777 515562 186793 515596
rect 186461 515534 186531 515562
rect 186461 515500 186497 515534
rect 186827 515528 186908 515630
rect 186461 515498 186531 515500
rect 186578 515494 186908 515528
rect 186945 515588 186995 515622
rect 187029 515588 187049 515622
rect 186945 515514 187049 515588
rect 187083 515582 187187 515656
rect 187083 515548 187103 515582
rect 187137 515548 187187 515582
rect 187221 515832 187463 515874
rect 187221 515798 187239 515832
rect 187273 515798 187411 515832
rect 187445 515798 187463 515832
rect 187221 515737 187463 515798
rect 187221 515703 187239 515737
rect 187273 515703 187411 515737
rect 187445 515703 187463 515737
rect 187221 515656 187463 515703
rect 187221 515582 187325 515656
rect 187221 515548 187271 515582
rect 187305 515548 187325 515582
rect 187359 515588 187379 515622
rect 187413 515588 187463 515622
rect 187359 515514 187463 515588
rect 186578 515466 186637 515494
rect 186393 515448 186453 515464
rect 186393 515414 186411 515448
rect 186445 515414 186453 515448
rect 186393 515398 186453 515414
rect 186487 515444 186542 515460
rect 186487 515410 186497 515444
rect 186531 515410 186542 515444
rect 186578 515432 186594 515466
rect 186628 515432 186637 515466
rect 186757 515466 186809 515494
rect 186578 515416 186637 515432
rect 186671 515444 186722 515460
rect 186487 515364 186542 515410
rect 186671 515410 186680 515444
rect 186714 515410 186722 515444
rect 186757 515432 186766 515466
rect 186800 515432 186809 515466
rect 186945 515461 187187 515514
rect 186757 515416 186809 515432
rect 186843 515444 186899 515460
rect 186671 515364 186722 515410
rect 186843 515410 186852 515444
rect 186886 515410 186899 515444
rect 186843 515364 186899 515410
rect 186945 515427 186963 515461
rect 186997 515427 187135 515461
rect 187169 515427 187187 515461
rect 186945 515364 187187 515427
rect 187221 515461 187463 515514
rect 187221 515427 187239 515461
rect 187273 515427 187411 515461
rect 187445 515427 187463 515461
rect 187221 515364 187463 515427
rect 172208 515330 172237 515364
rect 172271 515330 172329 515364
rect 172363 515330 172421 515364
rect 172455 515330 172513 515364
rect 172547 515330 172605 515364
rect 172639 515330 172697 515364
rect 172731 515330 172789 515364
rect 172823 515330 172881 515364
rect 172915 515330 172973 515364
rect 173007 515330 173065 515364
rect 173099 515330 173157 515364
rect 173191 515330 173249 515364
rect 173283 515330 173341 515364
rect 173375 515330 173433 515364
rect 173467 515330 173525 515364
rect 173559 515330 173617 515364
rect 173651 515330 173709 515364
rect 173743 515330 173801 515364
rect 173835 515330 173893 515364
rect 173927 515330 173985 515364
rect 174019 515330 174077 515364
rect 174111 515330 174169 515364
rect 174203 515330 174261 515364
rect 174295 515330 174353 515364
rect 174387 515330 174445 515364
rect 174479 515330 174537 515364
rect 174571 515330 174629 515364
rect 174663 515330 174721 515364
rect 174755 515330 174813 515364
rect 174847 515330 174905 515364
rect 174939 515330 174997 515364
rect 175031 515330 175089 515364
rect 175123 515330 175181 515364
rect 175215 515330 175273 515364
rect 175307 515330 175365 515364
rect 175399 515330 175457 515364
rect 175491 515330 175549 515364
rect 175583 515330 175641 515364
rect 175675 515330 175733 515364
rect 175767 515330 175825 515364
rect 175859 515330 175917 515364
rect 175951 515330 176009 515364
rect 176043 515330 176101 515364
rect 176135 515330 176193 515364
rect 176227 515330 176285 515364
rect 176319 515330 176377 515364
rect 176411 515330 176469 515364
rect 176503 515330 176561 515364
rect 176595 515330 176653 515364
rect 176687 515330 176745 515364
rect 176779 515330 176837 515364
rect 176871 515330 176929 515364
rect 176963 515330 177021 515364
rect 177055 515330 177113 515364
rect 177147 515330 177205 515364
rect 177239 515330 177297 515364
rect 177331 515330 177389 515364
rect 177423 515330 177481 515364
rect 177515 515330 177573 515364
rect 177607 515330 177665 515364
rect 177699 515330 177757 515364
rect 177791 515330 177849 515364
rect 177883 515330 177941 515364
rect 177975 515330 178033 515364
rect 178067 515330 178125 515364
rect 178159 515330 178217 515364
rect 178251 515330 178309 515364
rect 178343 515330 178401 515364
rect 178435 515330 178493 515364
rect 178527 515330 178585 515364
rect 178619 515330 178677 515364
rect 178711 515330 178769 515364
rect 178803 515330 178861 515364
rect 178895 515330 178953 515364
rect 178987 515330 179045 515364
rect 179079 515330 179137 515364
rect 179171 515330 179229 515364
rect 179263 515330 179321 515364
rect 179355 515330 179413 515364
rect 179447 515330 179505 515364
rect 179539 515330 179597 515364
rect 179631 515330 179689 515364
rect 179723 515330 179781 515364
rect 179815 515330 179873 515364
rect 179907 515330 179965 515364
rect 179999 515330 180057 515364
rect 180091 515330 180149 515364
rect 180183 515330 180241 515364
rect 180275 515330 180333 515364
rect 180367 515330 180425 515364
rect 180459 515330 180517 515364
rect 180551 515330 180609 515364
rect 180643 515330 180701 515364
rect 180735 515330 180793 515364
rect 180827 515330 180885 515364
rect 180919 515330 180977 515364
rect 181011 515330 181069 515364
rect 181103 515330 181161 515364
rect 181195 515330 181253 515364
rect 181287 515330 181345 515364
rect 181379 515330 181437 515364
rect 181471 515330 181529 515364
rect 181563 515330 181621 515364
rect 181655 515330 181713 515364
rect 181747 515330 181805 515364
rect 181839 515330 181897 515364
rect 181931 515330 181989 515364
rect 182023 515330 182081 515364
rect 182115 515330 182173 515364
rect 182207 515330 182265 515364
rect 182299 515330 182357 515364
rect 182391 515330 182449 515364
rect 182483 515330 182541 515364
rect 182575 515330 182633 515364
rect 182667 515330 182725 515364
rect 182759 515330 182817 515364
rect 182851 515330 182909 515364
rect 182943 515330 183001 515364
rect 183035 515330 183093 515364
rect 183127 515330 183185 515364
rect 183219 515330 183277 515364
rect 183311 515330 183369 515364
rect 183403 515330 183461 515364
rect 183495 515330 183553 515364
rect 183587 515330 183645 515364
rect 183679 515330 183737 515364
rect 183771 515330 183829 515364
rect 183863 515330 183921 515364
rect 183955 515330 184013 515364
rect 184047 515330 184105 515364
rect 184139 515330 184197 515364
rect 184231 515330 184289 515364
rect 184323 515330 184381 515364
rect 184415 515330 184473 515364
rect 184507 515330 184565 515364
rect 184599 515330 184657 515364
rect 184691 515330 184749 515364
rect 184783 515330 184841 515364
rect 184875 515330 184933 515364
rect 184967 515330 185025 515364
rect 185059 515330 185117 515364
rect 185151 515330 185209 515364
rect 185243 515330 185301 515364
rect 185335 515330 185393 515364
rect 185427 515330 185485 515364
rect 185519 515330 185577 515364
rect 185611 515330 185669 515364
rect 185703 515330 185761 515364
rect 185795 515330 185853 515364
rect 185887 515330 185945 515364
rect 185979 515330 186037 515364
rect 186071 515330 186129 515364
rect 186163 515330 186221 515364
rect 186255 515330 186313 515364
rect 186347 515330 186405 515364
rect 186439 515330 186497 515364
rect 186531 515330 186589 515364
rect 186623 515330 186681 515364
rect 186715 515330 186773 515364
rect 186807 515330 186865 515364
rect 186899 515330 186957 515364
rect 186991 515330 187049 515364
rect 187083 515330 187141 515364
rect 187175 515330 187233 515364
rect 187267 515330 187325 515364
rect 187359 515330 187417 515364
rect 187451 515330 187480 515364
<< viali >>
rect 164728 541085 164762 541119
rect 165031 541092 165065 541126
rect 165223 541092 165257 541126
rect 165415 541092 165449 541126
rect 165607 541092 165641 541126
rect 165799 541092 165833 541126
rect 165991 541092 166025 541126
rect 166408 541085 166442 541119
rect 164684 540530 164718 541018
rect 164772 540530 164806 541018
rect 164887 540083 164921 540571
rect 164983 540537 165017 541025
rect 165079 540083 165113 540571
rect 165175 540537 165209 541025
rect 165271 540083 165305 540571
rect 165367 540537 165401 541025
rect 165463 540083 165497 540571
rect 165559 540537 165593 541025
rect 165655 540083 165689 540571
rect 165751 540537 165785 541025
rect 165847 540083 165881 540571
rect 165943 540537 165977 541025
rect 166039 540083 166073 540571
rect 166208 540285 166242 540319
rect 166164 540059 166198 540235
rect 166252 540059 166286 540235
rect 166364 540076 166398 540564
rect 166452 540076 166486 540564
rect 166568 540085 166578 540215
rect 166578 540085 166618 540215
rect 166618 540085 166628 540215
rect 164728 539975 164762 540009
rect 164935 539982 164969 540016
rect 165127 539982 165161 540016
rect 165319 539982 165353 540016
rect 165511 539982 165545 540016
rect 165703 539982 165737 540016
rect 165895 539982 165929 540016
rect 166208 539975 166242 540009
rect 166408 539975 166442 540009
rect 168528 541085 168562 541119
rect 168831 541092 168865 541126
rect 169023 541092 169057 541126
rect 169215 541092 169249 541126
rect 169407 541092 169441 541126
rect 169599 541092 169633 541126
rect 169791 541092 169825 541126
rect 170208 541085 170242 541119
rect 168484 540530 168518 541018
rect 168572 540530 168606 541018
rect 168687 540083 168721 540571
rect 168783 540537 168817 541025
rect 168879 540083 168913 540571
rect 168975 540537 169009 541025
rect 169071 540083 169105 540571
rect 169167 540537 169201 541025
rect 169263 540083 169297 540571
rect 169359 540537 169393 541025
rect 169455 540083 169489 540571
rect 169551 540537 169585 541025
rect 169647 540083 169681 540571
rect 169743 540537 169777 541025
rect 169839 540083 169873 540571
rect 170008 540285 170042 540319
rect 169964 540059 169998 540235
rect 170052 540059 170086 540235
rect 170164 540076 170198 540564
rect 170252 540076 170286 540564
rect 170368 540085 170378 540215
rect 170378 540085 170418 540215
rect 170418 540085 170428 540215
rect 168528 539975 168562 540009
rect 168735 539982 168769 540016
rect 168927 539982 168961 540016
rect 169119 539982 169153 540016
rect 169311 539982 169345 540016
rect 169503 539982 169537 540016
rect 169695 539982 169729 540016
rect 170008 539975 170042 540009
rect 170208 539975 170242 540009
rect 172228 541085 172262 541119
rect 172531 541092 172565 541126
rect 172723 541092 172757 541126
rect 172915 541092 172949 541126
rect 173107 541092 173141 541126
rect 173299 541092 173333 541126
rect 173491 541092 173525 541126
rect 173908 541085 173942 541119
rect 172184 540530 172218 541018
rect 172272 540530 172306 541018
rect 172387 540083 172421 540571
rect 172483 540537 172517 541025
rect 172579 540083 172613 540571
rect 172675 540537 172709 541025
rect 172771 540083 172805 540571
rect 172867 540537 172901 541025
rect 172963 540083 172997 540571
rect 173059 540537 173093 541025
rect 173155 540083 173189 540571
rect 173251 540537 173285 541025
rect 173347 540083 173381 540571
rect 173443 540537 173477 541025
rect 173539 540083 173573 540571
rect 173708 540285 173742 540319
rect 173664 540059 173698 540235
rect 173752 540059 173786 540235
rect 173864 540076 173898 540564
rect 173952 540076 173986 540564
rect 174068 540085 174078 540215
rect 174078 540085 174118 540215
rect 174118 540085 174128 540215
rect 172228 539975 172262 540009
rect 172435 539982 172469 540016
rect 172627 539982 172661 540016
rect 172819 539982 172853 540016
rect 173011 539982 173045 540016
rect 173203 539982 173237 540016
rect 173395 539982 173429 540016
rect 173708 539975 173742 540009
rect 173908 539975 173942 540009
rect 175728 541085 175762 541119
rect 176031 541092 176065 541126
rect 176223 541092 176257 541126
rect 176415 541092 176449 541126
rect 176607 541092 176641 541126
rect 176799 541092 176833 541126
rect 176991 541092 177025 541126
rect 177408 541085 177442 541119
rect 175684 540530 175718 541018
rect 175772 540530 175806 541018
rect 175887 540083 175921 540571
rect 175983 540537 176017 541025
rect 176079 540083 176113 540571
rect 176175 540537 176209 541025
rect 176271 540083 176305 540571
rect 176367 540537 176401 541025
rect 176463 540083 176497 540571
rect 176559 540537 176593 541025
rect 176655 540083 176689 540571
rect 176751 540537 176785 541025
rect 176847 540083 176881 540571
rect 176943 540537 176977 541025
rect 177039 540083 177073 540571
rect 177208 540285 177242 540319
rect 177164 540059 177198 540235
rect 177252 540059 177286 540235
rect 177364 540076 177398 540564
rect 177452 540076 177486 540564
rect 177568 540085 177578 540215
rect 177578 540085 177618 540215
rect 177618 540085 177628 540215
rect 175728 539975 175762 540009
rect 175935 539982 175969 540016
rect 176127 539982 176161 540016
rect 176319 539982 176353 540016
rect 176511 539982 176545 540016
rect 176703 539982 176737 540016
rect 176895 539982 176929 540016
rect 177208 539975 177242 540009
rect 177408 539975 177442 540009
rect 179328 541085 179362 541119
rect 179631 541092 179665 541126
rect 179823 541092 179857 541126
rect 180015 541092 180049 541126
rect 180207 541092 180241 541126
rect 180399 541092 180433 541126
rect 180591 541092 180625 541126
rect 181008 541085 181042 541119
rect 179284 540530 179318 541018
rect 179372 540530 179406 541018
rect 179487 540083 179521 540571
rect 179583 540537 179617 541025
rect 179679 540083 179713 540571
rect 179775 540537 179809 541025
rect 179871 540083 179905 540571
rect 179967 540537 180001 541025
rect 180063 540083 180097 540571
rect 180159 540537 180193 541025
rect 180255 540083 180289 540571
rect 180351 540537 180385 541025
rect 180447 540083 180481 540571
rect 180543 540537 180577 541025
rect 180639 540083 180673 540571
rect 180808 540285 180842 540319
rect 180764 540059 180798 540235
rect 180852 540059 180886 540235
rect 180964 540076 180998 540564
rect 181052 540076 181086 540564
rect 181168 540085 181178 540215
rect 181178 540085 181218 540215
rect 181218 540085 181228 540215
rect 179328 539975 179362 540009
rect 179535 539982 179569 540016
rect 179727 539982 179761 540016
rect 179919 539982 179953 540016
rect 180111 539982 180145 540016
rect 180303 539982 180337 540016
rect 180495 539982 180529 540016
rect 180808 539975 180842 540009
rect 181008 539975 181042 540009
rect 182628 541085 182662 541119
rect 182931 541092 182965 541126
rect 183123 541092 183157 541126
rect 183315 541092 183349 541126
rect 183507 541092 183541 541126
rect 183699 541092 183733 541126
rect 183891 541092 183925 541126
rect 184308 541085 184342 541119
rect 182584 540530 182618 541018
rect 182672 540530 182706 541018
rect 182787 540083 182821 540571
rect 182883 540537 182917 541025
rect 182979 540083 183013 540571
rect 183075 540537 183109 541025
rect 183171 540083 183205 540571
rect 183267 540537 183301 541025
rect 183363 540083 183397 540571
rect 183459 540537 183493 541025
rect 183555 540083 183589 540571
rect 183651 540537 183685 541025
rect 183747 540083 183781 540571
rect 183843 540537 183877 541025
rect 183939 540083 183973 540571
rect 184108 540285 184142 540319
rect 184064 540059 184098 540235
rect 184152 540059 184186 540235
rect 184264 540076 184298 540564
rect 184352 540076 184386 540564
rect 184468 540085 184478 540215
rect 184478 540085 184518 540215
rect 184518 540085 184528 540215
rect 182628 539975 182662 540009
rect 182835 539982 182869 540016
rect 183027 539982 183061 540016
rect 183219 539982 183253 540016
rect 183411 539982 183445 540016
rect 183603 539982 183637 540016
rect 183795 539982 183829 540016
rect 184108 539975 184142 540009
rect 184308 539975 184342 540009
rect 185928 541085 185962 541119
rect 186231 541092 186265 541126
rect 186423 541092 186457 541126
rect 186615 541092 186649 541126
rect 186807 541092 186841 541126
rect 186999 541092 187033 541126
rect 187191 541092 187225 541126
rect 187608 541085 187642 541119
rect 185884 540530 185918 541018
rect 185972 540530 186006 541018
rect 186087 540083 186121 540571
rect 186183 540537 186217 541025
rect 186279 540083 186313 540571
rect 186375 540537 186409 541025
rect 186471 540083 186505 540571
rect 186567 540537 186601 541025
rect 186663 540083 186697 540571
rect 186759 540537 186793 541025
rect 186855 540083 186889 540571
rect 186951 540537 186985 541025
rect 187047 540083 187081 540571
rect 187143 540537 187177 541025
rect 187239 540083 187273 540571
rect 187408 540285 187442 540319
rect 187364 540059 187398 540235
rect 187452 540059 187486 540235
rect 187564 540076 187598 540564
rect 187652 540076 187686 540564
rect 187768 540085 187778 540215
rect 187778 540085 187818 540215
rect 187818 540085 187828 540215
rect 185928 539975 185962 540009
rect 186135 539982 186169 540016
rect 186327 539982 186361 540016
rect 186519 539982 186553 540016
rect 186711 539982 186745 540016
rect 186903 539982 186937 540016
rect 187095 539982 187129 540016
rect 187408 539975 187442 540009
rect 187608 539975 187642 540009
rect 189228 541085 189262 541119
rect 189531 541092 189565 541126
rect 189723 541092 189757 541126
rect 189915 541092 189949 541126
rect 190107 541092 190141 541126
rect 190299 541092 190333 541126
rect 190491 541092 190525 541126
rect 190908 541085 190942 541119
rect 189184 540530 189218 541018
rect 189272 540530 189306 541018
rect 189387 540083 189421 540571
rect 189483 540537 189517 541025
rect 189579 540083 189613 540571
rect 189675 540537 189709 541025
rect 189771 540083 189805 540571
rect 189867 540537 189901 541025
rect 189963 540083 189997 540571
rect 190059 540537 190093 541025
rect 190155 540083 190189 540571
rect 190251 540537 190285 541025
rect 190347 540083 190381 540571
rect 190443 540537 190477 541025
rect 190539 540083 190573 540571
rect 190708 540285 190742 540319
rect 190664 540059 190698 540235
rect 190752 540059 190786 540235
rect 190864 540076 190898 540564
rect 190952 540076 190986 540564
rect 191068 540085 191078 540215
rect 191078 540085 191118 540215
rect 191118 540085 191128 540215
rect 189228 539975 189262 540009
rect 189435 539982 189469 540016
rect 189627 539982 189661 540016
rect 189819 539982 189853 540016
rect 190011 539982 190045 540016
rect 190203 539982 190237 540016
rect 190395 539982 190429 540016
rect 190708 539975 190742 540009
rect 190908 539975 190942 540009
rect 191808 540065 191988 540245
rect 162268 538665 162528 538705
rect 158726 538435 158894 538469
rect 159102 538435 159270 538469
rect 159360 538435 159528 538469
rect 159618 538435 159786 538469
rect 159876 538435 160044 538469
rect 160134 538435 160302 538469
rect 160392 538435 160560 538469
rect 160650 538435 160818 538469
rect 160908 538435 161076 538469
rect 161166 538435 161334 538469
rect 161546 538435 161714 538469
rect 161946 538435 162114 538469
rect 162326 538435 162494 538469
rect 158664 538209 158698 538385
rect 158922 538209 158956 538385
rect 159040 538280 159074 538368
rect 159298 538226 159332 538314
rect 159556 538280 159590 538368
rect 159814 538226 159848 538314
rect 160072 538280 160106 538368
rect 160330 538226 160364 538314
rect 160588 538280 160622 538368
rect 160846 538226 160880 538314
rect 161104 538280 161138 538368
rect 161362 538226 161396 538314
rect 161484 538209 161518 538385
rect 161742 538209 161776 538385
rect 161884 538209 161918 538385
rect 162142 538209 162176 538385
rect 162264 538209 162298 538385
rect 162522 538209 162556 538385
rect 158726 538125 158894 538159
rect 159102 538125 159270 538159
rect 159360 538125 159528 538159
rect 159618 538125 159786 538159
rect 159876 538125 160044 538159
rect 160134 538125 160302 538159
rect 160392 538125 160560 538159
rect 160650 538125 160818 538159
rect 160908 538125 161076 538159
rect 161166 538125 161334 538159
rect 161546 538125 161714 538159
rect 161946 538125 162114 538159
rect 162326 538125 162494 538159
rect 164712 539572 164746 539606
rect 165035 539579 165069 539613
rect 165227 539579 165261 539613
rect 165419 539579 165453 539613
rect 165611 539579 165645 539613
rect 165803 539579 165837 539613
rect 165995 539579 166029 539613
rect 166212 539572 166246 539606
rect 166412 539572 166446 539606
rect 164668 538537 164702 539513
rect 164756 538537 164790 539513
rect 164891 538561 164925 539049
rect 164987 539015 165021 539503
rect 165083 538561 165117 539049
rect 165179 539015 165213 539503
rect 165275 538561 165309 539049
rect 165371 539015 165405 539503
rect 165467 538561 165501 539049
rect 165563 539015 165597 539503
rect 165659 538561 165693 539049
rect 165755 539015 165789 539503
rect 165851 538561 165885 539049
rect 165947 539015 165981 539503
rect 166043 538561 166077 539049
rect 166168 538937 166202 539513
rect 166256 538937 166290 539513
rect 166212 538844 166246 538878
rect 166368 538554 166402 539042
rect 166456 538554 166490 539042
rect 166568 539175 166578 539265
rect 166578 539175 166618 539265
rect 164712 538444 164746 538478
rect 164939 538451 164973 538485
rect 165131 538451 165165 538485
rect 165323 538451 165357 538485
rect 165515 538451 165549 538485
rect 165707 538451 165741 538485
rect 165899 538451 165933 538485
rect 166412 538444 166446 538478
rect 168512 539572 168546 539606
rect 168835 539579 168869 539613
rect 169027 539579 169061 539613
rect 169219 539579 169253 539613
rect 169411 539579 169445 539613
rect 169603 539579 169637 539613
rect 169795 539579 169829 539613
rect 170012 539572 170046 539606
rect 170212 539572 170246 539606
rect 168468 538537 168502 539513
rect 168556 538537 168590 539513
rect 168691 538561 168725 539049
rect 168787 539015 168821 539503
rect 168883 538561 168917 539049
rect 168979 539015 169013 539503
rect 169075 538561 169109 539049
rect 169171 539015 169205 539503
rect 169267 538561 169301 539049
rect 169363 539015 169397 539503
rect 169459 538561 169493 539049
rect 169555 539015 169589 539503
rect 169651 538561 169685 539049
rect 169747 539015 169781 539503
rect 169843 538561 169877 539049
rect 169968 538937 170002 539513
rect 170056 538937 170090 539513
rect 170012 538844 170046 538878
rect 170168 538554 170202 539042
rect 170256 538554 170290 539042
rect 170368 539175 170378 539265
rect 170378 539175 170418 539265
rect 168512 538444 168546 538478
rect 168739 538451 168773 538485
rect 168931 538451 168965 538485
rect 169123 538451 169157 538485
rect 169315 538451 169349 538485
rect 169507 538451 169541 538485
rect 169699 538451 169733 538485
rect 170212 538444 170246 538478
rect 172212 539572 172246 539606
rect 172535 539579 172569 539613
rect 172727 539579 172761 539613
rect 172919 539579 172953 539613
rect 173111 539579 173145 539613
rect 173303 539579 173337 539613
rect 173495 539579 173529 539613
rect 173712 539572 173746 539606
rect 173912 539572 173946 539606
rect 172168 538537 172202 539513
rect 172256 538537 172290 539513
rect 172391 538561 172425 539049
rect 172487 539015 172521 539503
rect 172583 538561 172617 539049
rect 172679 539015 172713 539503
rect 172775 538561 172809 539049
rect 172871 539015 172905 539503
rect 172967 538561 173001 539049
rect 173063 539015 173097 539503
rect 173159 538561 173193 539049
rect 173255 539015 173289 539503
rect 173351 538561 173385 539049
rect 173447 539015 173481 539503
rect 173543 538561 173577 539049
rect 173668 538937 173702 539513
rect 173756 538937 173790 539513
rect 173712 538844 173746 538878
rect 173868 538554 173902 539042
rect 173956 538554 173990 539042
rect 174068 539175 174078 539265
rect 174078 539175 174118 539265
rect 172212 538444 172246 538478
rect 172439 538451 172473 538485
rect 172631 538451 172665 538485
rect 172823 538451 172857 538485
rect 173015 538451 173049 538485
rect 173207 538451 173241 538485
rect 173399 538451 173433 538485
rect 173912 538444 173946 538478
rect 175712 539572 175746 539606
rect 176035 539579 176069 539613
rect 176227 539579 176261 539613
rect 176419 539579 176453 539613
rect 176611 539579 176645 539613
rect 176803 539579 176837 539613
rect 176995 539579 177029 539613
rect 177212 539572 177246 539606
rect 177412 539572 177446 539606
rect 175668 538537 175702 539513
rect 175756 538537 175790 539513
rect 175891 538561 175925 539049
rect 175987 539015 176021 539503
rect 176083 538561 176117 539049
rect 176179 539015 176213 539503
rect 176275 538561 176309 539049
rect 176371 539015 176405 539503
rect 176467 538561 176501 539049
rect 176563 539015 176597 539503
rect 176659 538561 176693 539049
rect 176755 539015 176789 539503
rect 176851 538561 176885 539049
rect 176947 539015 176981 539503
rect 177043 538561 177077 539049
rect 177168 538937 177202 539513
rect 177256 538937 177290 539513
rect 177212 538844 177246 538878
rect 177368 538554 177402 539042
rect 177456 538554 177490 539042
rect 177568 539175 177578 539265
rect 177578 539175 177618 539265
rect 175712 538444 175746 538478
rect 175939 538451 175973 538485
rect 176131 538451 176165 538485
rect 176323 538451 176357 538485
rect 176515 538451 176549 538485
rect 176707 538451 176741 538485
rect 176899 538451 176933 538485
rect 177412 538444 177446 538478
rect 179312 539572 179346 539606
rect 179635 539579 179669 539613
rect 179827 539579 179861 539613
rect 180019 539579 180053 539613
rect 180211 539579 180245 539613
rect 180403 539579 180437 539613
rect 180595 539579 180629 539613
rect 180812 539572 180846 539606
rect 181012 539572 181046 539606
rect 179268 538537 179302 539513
rect 179356 538537 179390 539513
rect 179491 538561 179525 539049
rect 179587 539015 179621 539503
rect 179683 538561 179717 539049
rect 179779 539015 179813 539503
rect 179875 538561 179909 539049
rect 179971 539015 180005 539503
rect 180067 538561 180101 539049
rect 180163 539015 180197 539503
rect 180259 538561 180293 539049
rect 180355 539015 180389 539503
rect 180451 538561 180485 539049
rect 180547 539015 180581 539503
rect 180643 538561 180677 539049
rect 180768 538937 180802 539513
rect 180856 538937 180890 539513
rect 180812 538844 180846 538878
rect 180968 538554 181002 539042
rect 181056 538554 181090 539042
rect 181168 539175 181178 539265
rect 181178 539175 181218 539265
rect 179312 538444 179346 538478
rect 179539 538451 179573 538485
rect 179731 538451 179765 538485
rect 179923 538451 179957 538485
rect 180115 538451 180149 538485
rect 180307 538451 180341 538485
rect 180499 538451 180533 538485
rect 181012 538444 181046 538478
rect 182612 539572 182646 539606
rect 182935 539579 182969 539613
rect 183127 539579 183161 539613
rect 183319 539579 183353 539613
rect 183511 539579 183545 539613
rect 183703 539579 183737 539613
rect 183895 539579 183929 539613
rect 184112 539572 184146 539606
rect 184312 539572 184346 539606
rect 182568 538537 182602 539513
rect 182656 538537 182690 539513
rect 182791 538561 182825 539049
rect 182887 539015 182921 539503
rect 182983 538561 183017 539049
rect 183079 539015 183113 539503
rect 183175 538561 183209 539049
rect 183271 539015 183305 539503
rect 183367 538561 183401 539049
rect 183463 539015 183497 539503
rect 183559 538561 183593 539049
rect 183655 539015 183689 539503
rect 183751 538561 183785 539049
rect 183847 539015 183881 539503
rect 183943 538561 183977 539049
rect 184068 538937 184102 539513
rect 184156 538937 184190 539513
rect 184112 538844 184146 538878
rect 184268 538554 184302 539042
rect 184356 538554 184390 539042
rect 184468 539175 184478 539265
rect 184478 539175 184518 539265
rect 182612 538444 182646 538478
rect 182839 538451 182873 538485
rect 183031 538451 183065 538485
rect 183223 538451 183257 538485
rect 183415 538451 183449 538485
rect 183607 538451 183641 538485
rect 183799 538451 183833 538485
rect 184312 538444 184346 538478
rect 185912 539572 185946 539606
rect 186235 539579 186269 539613
rect 186427 539579 186461 539613
rect 186619 539579 186653 539613
rect 186811 539579 186845 539613
rect 187003 539579 187037 539613
rect 187195 539579 187229 539613
rect 187412 539572 187446 539606
rect 187612 539572 187646 539606
rect 185868 538537 185902 539513
rect 185956 538537 185990 539513
rect 186091 538561 186125 539049
rect 186187 539015 186221 539503
rect 186283 538561 186317 539049
rect 186379 539015 186413 539503
rect 186475 538561 186509 539049
rect 186571 539015 186605 539503
rect 186667 538561 186701 539049
rect 186763 539015 186797 539503
rect 186859 538561 186893 539049
rect 186955 539015 186989 539503
rect 187051 538561 187085 539049
rect 187147 539015 187181 539503
rect 187243 538561 187277 539049
rect 187368 538937 187402 539513
rect 187456 538937 187490 539513
rect 187412 538844 187446 538878
rect 187568 538554 187602 539042
rect 187656 538554 187690 539042
rect 187768 539175 187778 539265
rect 187778 539175 187818 539265
rect 185912 538444 185946 538478
rect 186139 538451 186173 538485
rect 186331 538451 186365 538485
rect 186523 538451 186557 538485
rect 186715 538451 186749 538485
rect 186907 538451 186941 538485
rect 187099 538451 187133 538485
rect 187612 538444 187646 538478
rect 189212 539572 189246 539606
rect 189535 539579 189569 539613
rect 189727 539579 189761 539613
rect 189919 539579 189953 539613
rect 190111 539579 190145 539613
rect 190303 539579 190337 539613
rect 190495 539579 190529 539613
rect 190712 539572 190746 539606
rect 190912 539572 190946 539606
rect 189168 538537 189202 539513
rect 189256 538537 189290 539513
rect 189391 538561 189425 539049
rect 189487 539015 189521 539503
rect 189583 538561 189617 539049
rect 189679 539015 189713 539503
rect 189775 538561 189809 539049
rect 189871 539015 189905 539503
rect 189967 538561 190001 539049
rect 190063 539015 190097 539503
rect 190159 538561 190193 539049
rect 190255 539015 190289 539503
rect 190351 538561 190385 539049
rect 190447 539015 190481 539503
rect 190543 538561 190577 539049
rect 190668 538937 190702 539513
rect 190756 538937 190790 539513
rect 190712 538844 190746 538878
rect 190868 538554 190902 539042
rect 190956 538554 190990 539042
rect 191068 539175 191078 539265
rect 191078 539175 191118 539265
rect 189212 538444 189246 538478
rect 189439 538451 189473 538485
rect 189631 538451 189665 538485
rect 189823 538451 189857 538485
rect 190015 538451 190049 538485
rect 190207 538451 190241 538485
rect 190399 538451 190433 538485
rect 190912 538444 190946 538478
rect 161302 537672 161336 537706
rect 161506 537672 161540 537706
rect 161698 537672 161732 537706
rect 161906 537672 161940 537706
rect 162098 537672 162132 537706
rect 162322 537672 162356 537706
rect 161258 537054 161292 537342
rect 161346 537054 161380 537342
rect 161458 537054 161492 537342
rect 161554 537308 161588 537596
rect 161650 537054 161684 537342
rect 161746 537308 161780 537596
rect 161858 537308 161892 537596
rect 161954 537054 161988 537342
rect 162050 537308 162084 537596
rect 162146 537054 162180 537342
rect 162278 537054 162312 537342
rect 162366 537054 162400 537342
rect 161302 536944 161336 536978
rect 161602 536944 161636 536978
rect 162002 536944 162036 536978
rect 162322 536944 162356 536978
rect 157810 536652 157978 536686
rect 158188 536652 158356 536686
rect 158446 536652 158614 536686
rect 158704 536652 158872 536686
rect 158962 536652 159130 536686
rect 159220 536652 159388 536686
rect 159478 536652 159646 536686
rect 159736 536652 159904 536686
rect 159994 536652 160162 536686
rect 160252 536652 160420 536686
rect 160510 536652 160678 536686
rect 160894 536652 161062 536686
rect 161152 536652 161320 536686
rect 161410 536652 161578 536686
rect 161792 536652 161960 536686
rect 162050 536652 162218 536686
rect 162430 536652 162598 536686
rect 157748 536017 157782 536593
rect 158006 536017 158040 536593
rect 158126 536034 158160 536322
rect 158384 536288 158418 536576
rect 158642 536034 158676 536322
rect 158900 536288 158934 536576
rect 159158 536034 159192 536322
rect 159416 536288 159450 536576
rect 159674 536034 159708 536322
rect 159932 536288 159966 536576
rect 160190 536034 160224 536322
rect 160448 536288 160482 536576
rect 160706 536034 160740 536322
rect 160832 536288 160866 536576
rect 161090 536034 161124 536322
rect 161348 536288 161382 536576
rect 161606 536034 161640 536322
rect 161730 536034 161764 536322
rect 161988 536288 162022 536576
rect 162246 536034 162280 536322
rect 162368 536017 162402 536593
rect 162626 536017 162660 536593
rect 157810 535924 157978 535958
rect 158188 535924 158356 535958
rect 158446 535924 158614 535958
rect 158704 535924 158872 535958
rect 158962 535924 159130 535958
rect 159220 535924 159388 535958
rect 159478 535924 159646 535958
rect 159736 535924 159904 535958
rect 159994 535924 160162 535958
rect 160252 535924 160420 535958
rect 160510 535924 160678 535958
rect 160894 535924 161062 535958
rect 161152 535924 161320 535958
rect 161410 535924 161578 535958
rect 161792 535924 161960 535958
rect 162050 535924 162218 535958
rect 162430 535924 162598 535958
rect 164332 537534 164370 537931
rect 164650 537534 164688 537931
rect 164968 537534 165006 537931
rect 165286 537534 165324 537931
rect 165604 537534 165642 537931
rect 165922 537534 165960 537931
rect 166240 537534 166278 537931
rect 166558 537534 166596 537931
rect 164332 536019 164370 536416
rect 164650 536019 164688 536416
rect 164968 536019 165006 536416
rect 165286 536019 165324 536416
rect 165604 536019 165642 536416
rect 165922 536019 165960 536416
rect 166240 536019 166278 536416
rect 166558 536019 166596 536416
rect 168104 537534 168142 537931
rect 168422 537534 168460 537931
rect 168740 537534 168778 537931
rect 169058 537534 169096 537931
rect 168104 536019 168142 536416
rect 168422 536019 168460 536416
rect 168740 536019 168778 536416
rect 169058 536019 169096 536416
rect 171840 537534 171878 537931
rect 172158 537534 172196 537931
rect 171840 536019 171878 536416
rect 172158 536019 172196 536416
rect 175358 537534 175396 537931
rect 175358 536019 175396 536416
rect 178958 537534 178996 537931
rect 178958 536579 178996 536976
rect 182258 537534 182296 537931
rect 182258 536859 182296 537256
rect 185558 537534 185596 537931
rect 185558 536999 185596 537396
rect 188858 537534 188896 537931
rect 188858 536903 188896 537300
rect 162048 535705 162648 535745
rect 164302 535194 164340 535591
rect 164620 535194 164658 535591
rect 164938 535194 164976 535591
rect 165256 535194 165294 535591
rect 165574 535194 165612 535591
rect 165892 535194 165930 535591
rect 166210 535194 166248 535591
rect 166528 535194 166566 535591
rect 164302 533679 164340 534076
rect 164620 533679 164658 534076
rect 164938 533679 164976 534076
rect 165256 533679 165294 534076
rect 165574 533679 165612 534076
rect 165892 533679 165930 534076
rect 166210 533679 166248 534076
rect 166528 533679 166566 534076
rect 172237 530562 172271 530596
rect 172329 530562 172363 530596
rect 172421 530562 172455 530596
rect 172513 530562 172547 530596
rect 172605 530562 172639 530596
rect 172697 530562 172731 530596
rect 172789 530562 172823 530596
rect 172881 530562 172915 530596
rect 172973 530562 173007 530596
rect 173065 530562 173099 530596
rect 173157 530562 173191 530596
rect 173249 530562 173283 530596
rect 173341 530562 173375 530596
rect 173433 530562 173467 530596
rect 173525 530562 173559 530596
rect 173617 530562 173651 530596
rect 173709 530562 173743 530596
rect 173801 530562 173835 530596
rect 173893 530562 173927 530596
rect 173985 530562 174019 530596
rect 174077 530562 174111 530596
rect 174169 530562 174203 530596
rect 174261 530562 174295 530596
rect 174353 530562 174387 530596
rect 174445 530562 174479 530596
rect 174537 530562 174571 530596
rect 174629 530562 174663 530596
rect 174721 530562 174755 530596
rect 174813 530562 174847 530596
rect 174905 530562 174939 530596
rect 174997 530562 175031 530596
rect 175089 530562 175123 530596
rect 175181 530562 175215 530596
rect 175273 530562 175307 530596
rect 175365 530562 175399 530596
rect 175457 530562 175491 530596
rect 175549 530562 175583 530596
rect 175641 530562 175675 530596
rect 175733 530562 175767 530596
rect 175825 530562 175859 530596
rect 175917 530562 175951 530596
rect 176009 530562 176043 530596
rect 176101 530562 176135 530596
rect 176193 530562 176227 530596
rect 176285 530562 176319 530596
rect 176377 530562 176411 530596
rect 176469 530562 176503 530596
rect 176561 530562 176595 530596
rect 176653 530562 176687 530596
rect 176745 530562 176779 530596
rect 176837 530562 176871 530596
rect 176929 530562 176963 530596
rect 177021 530562 177055 530596
rect 177113 530562 177147 530596
rect 177205 530562 177239 530596
rect 177297 530562 177331 530596
rect 177389 530562 177423 530596
rect 177481 530562 177515 530596
rect 177573 530562 177607 530596
rect 177665 530562 177699 530596
rect 177757 530562 177791 530596
rect 177849 530562 177883 530596
rect 177941 530562 177975 530596
rect 178033 530562 178067 530596
rect 178125 530562 178159 530596
rect 178217 530562 178251 530596
rect 178309 530562 178343 530596
rect 178401 530562 178435 530596
rect 178493 530562 178527 530596
rect 178585 530562 178619 530596
rect 178677 530562 178711 530596
rect 178769 530562 178803 530596
rect 178861 530562 178895 530596
rect 178953 530562 178987 530596
rect 179045 530562 179079 530596
rect 179137 530562 179171 530596
rect 179229 530562 179263 530596
rect 179321 530562 179355 530596
rect 179413 530562 179447 530596
rect 179505 530562 179539 530596
rect 179597 530562 179631 530596
rect 179689 530562 179723 530596
rect 179781 530562 179815 530596
rect 179873 530562 179907 530596
rect 179965 530562 179999 530596
rect 180057 530562 180091 530596
rect 180149 530562 180183 530596
rect 180241 530562 180275 530596
rect 180333 530562 180367 530596
rect 180425 530562 180459 530596
rect 180517 530562 180551 530596
rect 180609 530562 180643 530596
rect 180701 530562 180735 530596
rect 180793 530562 180827 530596
rect 180885 530562 180919 530596
rect 180977 530562 181011 530596
rect 181069 530562 181103 530596
rect 181161 530562 181195 530596
rect 181253 530562 181287 530596
rect 181345 530562 181379 530596
rect 181437 530562 181471 530596
rect 181529 530562 181563 530596
rect 181621 530562 181655 530596
rect 181713 530562 181747 530596
rect 181805 530562 181839 530596
rect 181897 530562 181931 530596
rect 181989 530562 182023 530596
rect 182081 530562 182115 530596
rect 182173 530562 182207 530596
rect 182265 530562 182299 530596
rect 182357 530562 182391 530596
rect 182449 530562 182483 530596
rect 182541 530562 182575 530596
rect 182633 530562 182667 530596
rect 182725 530562 182759 530596
rect 182817 530562 182851 530596
rect 182909 530562 182943 530596
rect 183001 530562 183035 530596
rect 183093 530562 183127 530596
rect 183185 530562 183219 530596
rect 183277 530562 183311 530596
rect 183369 530562 183403 530596
rect 183461 530562 183495 530596
rect 183553 530562 183587 530596
rect 183645 530562 183679 530596
rect 183737 530562 183771 530596
rect 183829 530562 183863 530596
rect 183921 530562 183955 530596
rect 184013 530562 184047 530596
rect 184105 530562 184139 530596
rect 184197 530562 184231 530596
rect 184289 530562 184323 530596
rect 184381 530562 184415 530596
rect 184473 530562 184507 530596
rect 184565 530562 184599 530596
rect 184657 530562 184691 530596
rect 184749 530562 184783 530596
rect 184841 530562 184875 530596
rect 184933 530562 184967 530596
rect 185025 530562 185059 530596
rect 185117 530562 185151 530596
rect 185209 530562 185243 530596
rect 185301 530562 185335 530596
rect 185393 530562 185427 530596
rect 185485 530562 185519 530596
rect 185577 530562 185611 530596
rect 185669 530562 185703 530596
rect 185761 530562 185795 530596
rect 185853 530562 185887 530596
rect 185945 530562 185979 530596
rect 186037 530562 186071 530596
rect 186129 530562 186163 530596
rect 186221 530562 186255 530596
rect 186313 530562 186347 530596
rect 186405 530562 186439 530596
rect 186497 530562 186531 530596
rect 186589 530562 186623 530596
rect 186681 530562 186715 530596
rect 186773 530562 186807 530596
rect 186865 530562 186899 530596
rect 186957 530562 186991 530596
rect 187049 530562 187083 530596
rect 187141 530562 187175 530596
rect 187233 530562 187267 530596
rect 187325 530562 187359 530596
rect 187417 530562 187451 530596
rect 172513 530392 172547 530426
rect 172881 530324 172915 530358
rect 174905 530392 174939 530426
rect 175273 530324 175307 530358
rect 175845 530392 175879 530426
rect 175905 530338 175923 530363
rect 175923 530338 175939 530363
rect 175905 530329 175939 530338
rect 175549 530256 175583 530290
rect 176121 530340 176129 530358
rect 176129 530340 176155 530358
rect 176121 530324 176155 530340
rect 176493 530410 176527 530426
rect 176493 530392 176503 530410
rect 176503 530392 176527 530410
rect 176565 530392 176599 530426
rect 176121 530214 176124 530222
rect 176124 530214 176155 530222
rect 176121 530188 176155 530214
rect 176837 530324 176871 530358
rect 176745 530188 176779 530222
rect 177021 530256 177055 530290
rect 177123 530204 177157 530222
rect 177123 530188 177157 530204
rect 177204 530349 177238 530358
rect 177204 530324 177226 530349
rect 177226 530324 177238 530349
rect 177297 530256 177331 530290
rect 177665 530120 177690 530154
rect 177690 530120 177699 530154
rect 178217 530256 178251 530290
rect 178769 530460 178776 530494
rect 178776 530460 178803 530494
rect 178585 530330 178611 530358
rect 178611 530330 178619 530358
rect 178585 530324 178619 530330
rect 179045 530324 179079 530358
rect 178401 530136 178435 530154
rect 178401 530120 178407 530136
rect 178407 530120 178435 530136
rect 179413 530460 179418 530494
rect 179418 530460 179447 530494
rect 179321 530324 179355 530358
rect 180241 530128 180275 530154
rect 180241 530120 180247 530128
rect 180247 530120 180275 530128
rect 180609 530324 180643 530358
rect 180701 530460 180735 530494
rect 180793 530256 180827 530290
rect 181253 530287 181287 530290
rect 181253 530256 181267 530287
rect 181267 530256 181287 530287
rect 181529 530324 181563 530358
rect 181437 530287 181471 530290
rect 181437 530256 181469 530287
rect 181469 530256 181471 530287
rect 181897 530196 181931 530222
rect 181897 530188 181925 530196
rect 181925 530188 181931 530196
rect 182081 530392 182115 530426
rect 182173 530129 182177 530154
rect 182177 530129 182207 530154
rect 182173 530120 182207 530129
rect 183277 530460 183282 530494
rect 183282 530460 183311 530494
rect 183185 530324 183219 530358
rect 185393 530460 185398 530494
rect 185398 530460 185427 530494
rect 185301 530392 185335 530426
rect 187141 530324 187175 530358
rect 172237 530018 172271 530052
rect 172329 530018 172363 530052
rect 172421 530018 172455 530052
rect 172513 530018 172547 530052
rect 172605 530018 172639 530052
rect 172697 530018 172731 530052
rect 172789 530018 172823 530052
rect 172881 530018 172915 530052
rect 172973 530018 173007 530052
rect 173065 530018 173099 530052
rect 173157 530018 173191 530052
rect 173249 530018 173283 530052
rect 173341 530018 173375 530052
rect 173433 530018 173467 530052
rect 173525 530018 173559 530052
rect 173617 530018 173651 530052
rect 173709 530018 173743 530052
rect 173801 530018 173835 530052
rect 173893 530018 173927 530052
rect 173985 530018 174019 530052
rect 174077 530018 174111 530052
rect 174169 530018 174203 530052
rect 174261 530018 174295 530052
rect 174353 530018 174387 530052
rect 174445 530018 174479 530052
rect 174537 530018 174571 530052
rect 174629 530018 174663 530052
rect 174721 530018 174755 530052
rect 174813 530018 174847 530052
rect 174905 530018 174939 530052
rect 174997 530018 175031 530052
rect 175089 530018 175123 530052
rect 175181 530018 175215 530052
rect 175273 530018 175307 530052
rect 175365 530018 175399 530052
rect 175457 530018 175491 530052
rect 175549 530018 175583 530052
rect 175641 530018 175675 530052
rect 175733 530018 175767 530052
rect 175825 530018 175859 530052
rect 175917 530018 175951 530052
rect 176009 530018 176043 530052
rect 176101 530018 176135 530052
rect 176193 530018 176227 530052
rect 176285 530018 176319 530052
rect 176377 530018 176411 530052
rect 176469 530018 176503 530052
rect 176561 530018 176595 530052
rect 176653 530018 176687 530052
rect 176745 530018 176779 530052
rect 176837 530018 176871 530052
rect 176929 530018 176963 530052
rect 177021 530018 177055 530052
rect 177113 530018 177147 530052
rect 177205 530018 177239 530052
rect 177297 530018 177331 530052
rect 177389 530018 177423 530052
rect 177481 530018 177515 530052
rect 177573 530018 177607 530052
rect 177665 530018 177699 530052
rect 177757 530018 177791 530052
rect 177849 530018 177883 530052
rect 177941 530018 177975 530052
rect 178033 530018 178067 530052
rect 178125 530018 178159 530052
rect 178217 530018 178251 530052
rect 178309 530018 178343 530052
rect 178401 530018 178435 530052
rect 178493 530018 178527 530052
rect 178585 530018 178619 530052
rect 178677 530018 178711 530052
rect 178769 530018 178803 530052
rect 178861 530018 178895 530052
rect 178953 530018 178987 530052
rect 179045 530018 179079 530052
rect 179137 530018 179171 530052
rect 179229 530018 179263 530052
rect 179321 530018 179355 530052
rect 179413 530018 179447 530052
rect 179505 530018 179539 530052
rect 179597 530018 179631 530052
rect 179689 530018 179723 530052
rect 179781 530018 179815 530052
rect 179873 530018 179907 530052
rect 179965 530018 179999 530052
rect 180057 530018 180091 530052
rect 180149 530018 180183 530052
rect 180241 530018 180275 530052
rect 180333 530018 180367 530052
rect 180425 530018 180459 530052
rect 180517 530018 180551 530052
rect 180609 530018 180643 530052
rect 180701 530018 180735 530052
rect 180793 530018 180827 530052
rect 180885 530018 180919 530052
rect 180977 530018 181011 530052
rect 181069 530018 181103 530052
rect 181161 530018 181195 530052
rect 181253 530018 181287 530052
rect 181345 530018 181379 530052
rect 181437 530018 181471 530052
rect 181529 530018 181563 530052
rect 181621 530018 181655 530052
rect 181713 530018 181747 530052
rect 181805 530018 181839 530052
rect 181897 530018 181931 530052
rect 181989 530018 182023 530052
rect 182081 530018 182115 530052
rect 182173 530018 182207 530052
rect 182265 530018 182299 530052
rect 182357 530018 182391 530052
rect 182449 530018 182483 530052
rect 182541 530018 182575 530052
rect 182633 530018 182667 530052
rect 182725 530018 182759 530052
rect 182817 530018 182851 530052
rect 182909 530018 182943 530052
rect 183001 530018 183035 530052
rect 183093 530018 183127 530052
rect 183185 530018 183219 530052
rect 183277 530018 183311 530052
rect 183369 530018 183403 530052
rect 183461 530018 183495 530052
rect 183553 530018 183587 530052
rect 183645 530018 183679 530052
rect 183737 530018 183771 530052
rect 183829 530018 183863 530052
rect 183921 530018 183955 530052
rect 184013 530018 184047 530052
rect 184105 530018 184139 530052
rect 184197 530018 184231 530052
rect 184289 530018 184323 530052
rect 184381 530018 184415 530052
rect 184473 530018 184507 530052
rect 184565 530018 184599 530052
rect 184657 530018 184691 530052
rect 184749 530018 184783 530052
rect 184841 530018 184875 530052
rect 184933 530018 184967 530052
rect 185025 530018 185059 530052
rect 185117 530018 185151 530052
rect 185209 530018 185243 530052
rect 185301 530018 185335 530052
rect 185393 530018 185427 530052
rect 185485 530018 185519 530052
rect 185577 530018 185611 530052
rect 185669 530018 185703 530052
rect 185761 530018 185795 530052
rect 185853 530018 185887 530052
rect 185945 530018 185979 530052
rect 186037 530018 186071 530052
rect 186129 530018 186163 530052
rect 186221 530018 186255 530052
rect 186313 530018 186347 530052
rect 186405 530018 186439 530052
rect 186497 530018 186531 530052
rect 186589 530018 186623 530052
rect 186681 530018 186715 530052
rect 186773 530018 186807 530052
rect 186865 530018 186899 530052
rect 186957 530018 186991 530052
rect 187049 530018 187083 530052
rect 187141 530018 187175 530052
rect 187233 530018 187267 530052
rect 187325 530018 187359 530052
rect 187417 530018 187451 530052
rect 174813 529780 174847 529814
rect 175549 529740 175583 529746
rect 175549 529712 175552 529740
rect 175552 529712 175583 529740
rect 175642 529721 175654 529746
rect 175654 529721 175676 529746
rect 175642 529712 175676 529721
rect 175457 529576 175466 529610
rect 175466 529576 175491 529610
rect 175723 529866 175757 529882
rect 175723 529848 175757 529866
rect 175825 529780 175859 529814
rect 176101 529848 176135 529882
rect 176009 529712 176043 529746
rect 176725 529856 176759 529882
rect 176725 529848 176756 529856
rect 176756 529848 176759 529856
rect 176281 529644 176315 529678
rect 176353 529660 176377 529678
rect 176377 529660 176387 529678
rect 176353 529644 176387 529660
rect 176725 529730 176759 529746
rect 176725 529712 176751 529730
rect 176751 529712 176759 529730
rect 177297 529940 177331 529950
rect 177297 529916 177325 529940
rect 177325 529916 177331 529940
rect 176941 529732 176975 529741
rect 176941 529707 176957 529732
rect 176957 529707 176975 529732
rect 177001 529644 177035 529678
rect 177665 529783 177679 529814
rect 177679 529783 177699 529814
rect 177665 529780 177699 529783
rect 177849 529644 177883 529678
rect 177941 529712 177975 529746
rect 178309 529874 178337 529882
rect 178337 529874 178343 529882
rect 178309 529848 178343 529874
rect 178401 529940 178435 529950
rect 178401 529916 178407 529940
rect 178407 529916 178435 529940
rect 178973 529856 179007 529882
rect 178973 529848 178976 529856
rect 178976 529848 179007 529856
rect 178757 529732 178791 529741
rect 178757 529707 178775 529732
rect 178775 529707 178791 529732
rect 178697 529644 178731 529678
rect 178973 529730 179007 529746
rect 178973 529712 178981 529730
rect 178981 529712 179007 529730
rect 179597 529848 179631 529882
rect 179345 529660 179355 529678
rect 179355 529660 179379 529678
rect 179345 529644 179379 529660
rect 179417 529644 179451 529678
rect 179689 529712 179723 529746
rect 179975 529866 180009 529882
rect 179975 529848 180009 529866
rect 179873 529780 179907 529814
rect 180056 529721 180078 529746
rect 180078 529721 180090 529746
rect 180056 529712 180090 529721
rect 180149 529740 180183 529746
rect 180149 529712 180180 529740
rect 180180 529712 180183 529740
rect 180241 529740 180275 529746
rect 180241 529712 180244 529740
rect 180244 529712 180275 529740
rect 180334 529721 180346 529746
rect 180346 529721 180368 529746
rect 180334 529712 180368 529721
rect 180415 529866 180449 529882
rect 180415 529848 180449 529866
rect 180517 529780 180551 529814
rect 180793 529848 180827 529882
rect 180701 529712 180735 529746
rect 181417 529856 181451 529882
rect 181417 529848 181448 529856
rect 181448 529848 181451 529856
rect 180973 529644 181007 529678
rect 181045 529660 181069 529678
rect 181069 529660 181079 529678
rect 181045 529644 181079 529660
rect 181417 529730 181451 529746
rect 181417 529712 181443 529730
rect 181443 529712 181451 529730
rect 181989 529780 182023 529814
rect 181633 529732 181667 529741
rect 181633 529707 181649 529732
rect 181649 529707 181667 529732
rect 181693 529644 181727 529678
rect 182633 529916 182658 529950
rect 182658 529916 182667 529950
rect 183185 529780 183219 529814
rect 172237 529474 172271 529508
rect 172329 529474 172363 529508
rect 172421 529474 172455 529508
rect 172513 529474 172547 529508
rect 172605 529474 172639 529508
rect 172697 529474 172731 529508
rect 172789 529474 172823 529508
rect 172881 529474 172915 529508
rect 172973 529474 173007 529508
rect 173065 529474 173099 529508
rect 173157 529474 173191 529508
rect 173249 529474 173283 529508
rect 173341 529474 173375 529508
rect 173433 529474 173467 529508
rect 173525 529474 173559 529508
rect 173617 529474 173651 529508
rect 173709 529474 173743 529508
rect 173801 529474 173835 529508
rect 173893 529474 173927 529508
rect 173985 529474 174019 529508
rect 174077 529474 174111 529508
rect 174169 529474 174203 529508
rect 174261 529474 174295 529508
rect 174353 529474 174387 529508
rect 174445 529474 174479 529508
rect 174537 529474 174571 529508
rect 174629 529474 174663 529508
rect 174721 529474 174755 529508
rect 174813 529474 174847 529508
rect 174905 529474 174939 529508
rect 174997 529474 175031 529508
rect 175089 529474 175123 529508
rect 175181 529474 175215 529508
rect 175273 529474 175307 529508
rect 175365 529474 175399 529508
rect 175457 529474 175491 529508
rect 175549 529474 175583 529508
rect 175641 529474 175675 529508
rect 175733 529474 175767 529508
rect 175825 529474 175859 529508
rect 175917 529474 175951 529508
rect 176009 529474 176043 529508
rect 176101 529474 176135 529508
rect 176193 529474 176227 529508
rect 176285 529474 176319 529508
rect 176377 529474 176411 529508
rect 176469 529474 176503 529508
rect 176561 529474 176595 529508
rect 176653 529474 176687 529508
rect 176745 529474 176779 529508
rect 176837 529474 176871 529508
rect 176929 529474 176963 529508
rect 177021 529474 177055 529508
rect 177113 529474 177147 529508
rect 177205 529474 177239 529508
rect 177297 529474 177331 529508
rect 177389 529474 177423 529508
rect 177481 529474 177515 529508
rect 177573 529474 177607 529508
rect 177665 529474 177699 529508
rect 177757 529474 177791 529508
rect 177849 529474 177883 529508
rect 177941 529474 177975 529508
rect 178033 529474 178067 529508
rect 178125 529474 178159 529508
rect 178217 529474 178251 529508
rect 178309 529474 178343 529508
rect 178401 529474 178435 529508
rect 178493 529474 178527 529508
rect 178585 529474 178619 529508
rect 178677 529474 178711 529508
rect 178769 529474 178803 529508
rect 178861 529474 178895 529508
rect 178953 529474 178987 529508
rect 179045 529474 179079 529508
rect 179137 529474 179171 529508
rect 179229 529474 179263 529508
rect 179321 529474 179355 529508
rect 179413 529474 179447 529508
rect 179505 529474 179539 529508
rect 179597 529474 179631 529508
rect 179689 529474 179723 529508
rect 179781 529474 179815 529508
rect 179873 529474 179907 529508
rect 179965 529474 179999 529508
rect 180057 529474 180091 529508
rect 180149 529474 180183 529508
rect 180241 529474 180275 529508
rect 180333 529474 180367 529508
rect 180425 529474 180459 529508
rect 180517 529474 180551 529508
rect 180609 529474 180643 529508
rect 180701 529474 180735 529508
rect 180793 529474 180827 529508
rect 180885 529474 180919 529508
rect 180977 529474 181011 529508
rect 181069 529474 181103 529508
rect 181161 529474 181195 529508
rect 181253 529474 181287 529508
rect 181345 529474 181379 529508
rect 181437 529474 181471 529508
rect 181529 529474 181563 529508
rect 181621 529474 181655 529508
rect 181713 529474 181747 529508
rect 181805 529474 181839 529508
rect 181897 529474 181931 529508
rect 181989 529474 182023 529508
rect 182081 529474 182115 529508
rect 182173 529474 182207 529508
rect 182265 529474 182299 529508
rect 182357 529474 182391 529508
rect 182449 529474 182483 529508
rect 182541 529474 182575 529508
rect 182633 529474 182667 529508
rect 182725 529474 182759 529508
rect 182817 529474 182851 529508
rect 182909 529474 182943 529508
rect 183001 529474 183035 529508
rect 183093 529474 183127 529508
rect 183185 529474 183219 529508
rect 183277 529474 183311 529508
rect 183369 529474 183403 529508
rect 183461 529474 183495 529508
rect 183553 529474 183587 529508
rect 183645 529474 183679 529508
rect 183737 529474 183771 529508
rect 183829 529474 183863 529508
rect 183921 529474 183955 529508
rect 184013 529474 184047 529508
rect 184105 529474 184139 529508
rect 184197 529474 184231 529508
rect 184289 529474 184323 529508
rect 184381 529474 184415 529508
rect 184473 529474 184507 529508
rect 184565 529474 184599 529508
rect 184657 529474 184691 529508
rect 184749 529474 184783 529508
rect 184841 529474 184875 529508
rect 184933 529474 184967 529508
rect 185025 529474 185059 529508
rect 185117 529474 185151 529508
rect 185209 529474 185243 529508
rect 185301 529474 185335 529508
rect 185393 529474 185427 529508
rect 185485 529474 185519 529508
rect 185577 529474 185611 529508
rect 185669 529474 185703 529508
rect 185761 529474 185795 529508
rect 185853 529474 185887 529508
rect 185945 529474 185979 529508
rect 186037 529474 186071 529508
rect 186129 529474 186163 529508
rect 186221 529474 186255 529508
rect 186313 529474 186347 529508
rect 186405 529474 186439 529508
rect 186497 529474 186531 529508
rect 186589 529474 186623 529508
rect 186681 529474 186715 529508
rect 186773 529474 186807 529508
rect 186865 529474 186899 529508
rect 186957 529474 186991 529508
rect 187049 529474 187083 529508
rect 187141 529474 187175 529508
rect 187233 529474 187267 529508
rect 187325 529474 187359 529508
rect 187417 529474 187451 529508
rect 175365 529372 175399 529406
rect 175273 529168 175307 529202
rect 175457 529236 175491 529270
rect 177665 529242 177691 529270
rect 177691 529242 177699 529270
rect 177665 529236 177699 529242
rect 175825 529040 175859 529066
rect 175825 529032 175853 529040
rect 175853 529032 175859 529040
rect 176193 529050 176198 529066
rect 176198 529050 176227 529066
rect 176193 529032 176227 529050
rect 177757 529168 177791 529202
rect 177850 529261 177884 529270
rect 177850 529236 177862 529261
rect 177862 529236 177884 529261
rect 178033 529304 178067 529338
rect 177931 529116 177965 529134
rect 177931 529100 177965 529116
rect 178217 529236 178251 529270
rect 178489 529304 178523 529338
rect 178561 529322 178595 529338
rect 178561 529304 178585 529322
rect 178585 529304 178595 529322
rect 178309 529100 178343 529134
rect 178933 529252 178959 529270
rect 178959 529252 178967 529270
rect 178933 529236 178967 529252
rect 179209 529304 179243 529338
rect 179149 529250 179165 529275
rect 179165 529250 179183 529275
rect 179149 529241 179183 529250
rect 178933 529126 178964 529134
rect 178964 529126 178967 529134
rect 178933 529100 178967 529126
rect 179873 529402 179907 529406
rect 179873 529372 179901 529402
rect 179901 529372 179907 529402
rect 179689 529242 179697 529270
rect 179697 529242 179723 529270
rect 179689 529236 179723 529242
rect 179505 529042 179533 529066
rect 179533 529042 179539 529066
rect 179505 529032 179539 529042
rect 180701 529242 180709 529270
rect 180709 529242 180735 529270
rect 180701 529236 180735 529242
rect 182541 529402 182575 529406
rect 182541 529372 182547 529402
rect 182547 529372 182575 529402
rect 181989 529050 181996 529066
rect 181996 529050 182023 529066
rect 181989 529032 182023 529050
rect 182725 529242 182751 529270
rect 182751 529242 182759 529270
rect 182725 529236 182759 529242
rect 172237 528930 172271 528964
rect 172329 528930 172363 528964
rect 172421 528930 172455 528964
rect 172513 528930 172547 528964
rect 172605 528930 172639 528964
rect 172697 528930 172731 528964
rect 172789 528930 172823 528964
rect 172881 528930 172915 528964
rect 172973 528930 173007 528964
rect 173065 528930 173099 528964
rect 173157 528930 173191 528964
rect 173249 528930 173283 528964
rect 173341 528930 173375 528964
rect 173433 528930 173467 528964
rect 173525 528930 173559 528964
rect 173617 528930 173651 528964
rect 173709 528930 173743 528964
rect 173801 528930 173835 528964
rect 173893 528930 173927 528964
rect 173985 528930 174019 528964
rect 174077 528930 174111 528964
rect 174169 528930 174203 528964
rect 174261 528930 174295 528964
rect 174353 528930 174387 528964
rect 174445 528930 174479 528964
rect 174537 528930 174571 528964
rect 174629 528930 174663 528964
rect 174721 528930 174755 528964
rect 174813 528930 174847 528964
rect 174905 528930 174939 528964
rect 174997 528930 175031 528964
rect 175089 528930 175123 528964
rect 175181 528930 175215 528964
rect 175273 528930 175307 528964
rect 175365 528930 175399 528964
rect 175457 528930 175491 528964
rect 175549 528930 175583 528964
rect 175641 528930 175675 528964
rect 175733 528930 175767 528964
rect 175825 528930 175859 528964
rect 175917 528930 175951 528964
rect 176009 528930 176043 528964
rect 176101 528930 176135 528964
rect 176193 528930 176227 528964
rect 176285 528930 176319 528964
rect 176377 528930 176411 528964
rect 176469 528930 176503 528964
rect 176561 528930 176595 528964
rect 176653 528930 176687 528964
rect 176745 528930 176779 528964
rect 176837 528930 176871 528964
rect 176929 528930 176963 528964
rect 177021 528930 177055 528964
rect 177113 528930 177147 528964
rect 177205 528930 177239 528964
rect 177297 528930 177331 528964
rect 177389 528930 177423 528964
rect 177481 528930 177515 528964
rect 177573 528930 177607 528964
rect 177665 528930 177699 528964
rect 177757 528930 177791 528964
rect 177849 528930 177883 528964
rect 177941 528930 177975 528964
rect 178033 528930 178067 528964
rect 178125 528930 178159 528964
rect 178217 528930 178251 528964
rect 178309 528930 178343 528964
rect 178401 528930 178435 528964
rect 178493 528930 178527 528964
rect 178585 528930 178619 528964
rect 178677 528930 178711 528964
rect 178769 528930 178803 528964
rect 178861 528930 178895 528964
rect 178953 528930 178987 528964
rect 179045 528930 179079 528964
rect 179137 528930 179171 528964
rect 179229 528930 179263 528964
rect 179321 528930 179355 528964
rect 179413 528930 179447 528964
rect 179505 528930 179539 528964
rect 179597 528930 179631 528964
rect 179689 528930 179723 528964
rect 179781 528930 179815 528964
rect 179873 528930 179907 528964
rect 179965 528930 179999 528964
rect 180057 528930 180091 528964
rect 180149 528930 180183 528964
rect 180241 528930 180275 528964
rect 180333 528930 180367 528964
rect 180425 528930 180459 528964
rect 180517 528930 180551 528964
rect 180609 528930 180643 528964
rect 180701 528930 180735 528964
rect 180793 528930 180827 528964
rect 180885 528930 180919 528964
rect 180977 528930 181011 528964
rect 181069 528930 181103 528964
rect 181161 528930 181195 528964
rect 181253 528930 181287 528964
rect 181345 528930 181379 528964
rect 181437 528930 181471 528964
rect 181529 528930 181563 528964
rect 181621 528930 181655 528964
rect 181713 528930 181747 528964
rect 181805 528930 181839 528964
rect 181897 528930 181931 528964
rect 181989 528930 182023 528964
rect 182081 528930 182115 528964
rect 182173 528930 182207 528964
rect 182265 528930 182299 528964
rect 182357 528930 182391 528964
rect 182449 528930 182483 528964
rect 182541 528930 182575 528964
rect 182633 528930 182667 528964
rect 182725 528930 182759 528964
rect 182817 528930 182851 528964
rect 182909 528930 182943 528964
rect 183001 528930 183035 528964
rect 183093 528930 183127 528964
rect 183185 528930 183219 528964
rect 183277 528930 183311 528964
rect 183369 528930 183403 528964
rect 183461 528930 183495 528964
rect 183553 528930 183587 528964
rect 183645 528930 183679 528964
rect 183737 528930 183771 528964
rect 183829 528930 183863 528964
rect 183921 528930 183955 528964
rect 184013 528930 184047 528964
rect 184105 528930 184139 528964
rect 184197 528930 184231 528964
rect 184289 528930 184323 528964
rect 184381 528930 184415 528964
rect 184473 528930 184507 528964
rect 184565 528930 184599 528964
rect 184657 528930 184691 528964
rect 184749 528930 184783 528964
rect 184841 528930 184875 528964
rect 184933 528930 184967 528964
rect 185025 528930 185059 528964
rect 185117 528930 185151 528964
rect 185209 528930 185243 528964
rect 185301 528930 185335 528964
rect 185393 528930 185427 528964
rect 185485 528930 185519 528964
rect 185577 528930 185611 528964
rect 185669 528930 185703 528964
rect 185761 528930 185795 528964
rect 185853 528930 185887 528964
rect 185945 528930 185979 528964
rect 186037 528930 186071 528964
rect 186129 528930 186163 528964
rect 186221 528930 186255 528964
rect 186313 528930 186347 528964
rect 186405 528930 186439 528964
rect 186497 528930 186531 528964
rect 186589 528930 186623 528964
rect 186681 528930 186715 528964
rect 186773 528930 186807 528964
rect 186865 528930 186899 528964
rect 186957 528930 186991 528964
rect 187049 528930 187083 528964
rect 187141 528930 187175 528964
rect 187233 528930 187267 528964
rect 187325 528930 187359 528964
rect 187417 528930 187451 528964
rect 176101 528846 176129 528862
rect 176129 528846 176135 528862
rect 176101 528828 176135 528846
rect 175917 528652 175951 528658
rect 175917 528624 175925 528652
rect 175925 528624 175951 528652
rect 176193 528652 176227 528658
rect 176193 528624 176201 528652
rect 176201 528624 176227 528652
rect 176561 528695 176575 528726
rect 176575 528695 176595 528726
rect 176561 528692 176595 528695
rect 176377 528492 176405 528522
rect 176405 528492 176411 528522
rect 176377 528488 176411 528492
rect 176745 528488 176779 528522
rect 176837 528624 176871 528658
rect 177481 528624 177515 528658
rect 177205 528515 177239 528522
rect 177205 528488 177233 528515
rect 177233 528488 177239 528515
rect 178125 528692 178159 528726
rect 179689 528844 179723 528862
rect 179689 528828 179696 528844
rect 179696 528828 179723 528844
rect 180425 528765 180453 528794
rect 180453 528765 180459 528794
rect 180425 528760 180459 528765
rect 178401 528556 178435 528590
rect 180241 528652 180275 528658
rect 180241 528624 180249 528652
rect 180249 528624 180275 528652
rect 180517 528692 180551 528726
rect 180610 528633 180622 528658
rect 180622 528633 180644 528658
rect 180610 528624 180644 528633
rect 180691 528778 180725 528794
rect 180691 528760 180725 528778
rect 180793 528692 180827 528726
rect 181069 528760 181103 528794
rect 180977 528624 181011 528658
rect 181693 528768 181727 528794
rect 181693 528760 181724 528768
rect 181724 528760 181727 528768
rect 181249 528556 181283 528590
rect 181321 528572 181345 528590
rect 181345 528572 181355 528590
rect 181321 528556 181355 528572
rect 181693 528642 181727 528658
rect 181693 528624 181719 528642
rect 181719 528624 181727 528642
rect 182265 528852 182299 528862
rect 182265 528828 182293 528852
rect 182293 528828 182299 528852
rect 181909 528644 181943 528653
rect 181909 528619 181925 528644
rect 181925 528619 181943 528644
rect 181969 528556 182003 528590
rect 172237 528386 172271 528420
rect 172329 528386 172363 528420
rect 172421 528386 172455 528420
rect 172513 528386 172547 528420
rect 172605 528386 172639 528420
rect 172697 528386 172731 528420
rect 172789 528386 172823 528420
rect 172881 528386 172915 528420
rect 172973 528386 173007 528420
rect 173065 528386 173099 528420
rect 173157 528386 173191 528420
rect 173249 528386 173283 528420
rect 173341 528386 173375 528420
rect 173433 528386 173467 528420
rect 173525 528386 173559 528420
rect 173617 528386 173651 528420
rect 173709 528386 173743 528420
rect 173801 528386 173835 528420
rect 173893 528386 173927 528420
rect 173985 528386 174019 528420
rect 174077 528386 174111 528420
rect 174169 528386 174203 528420
rect 174261 528386 174295 528420
rect 174353 528386 174387 528420
rect 174445 528386 174479 528420
rect 174537 528386 174571 528420
rect 174629 528386 174663 528420
rect 174721 528386 174755 528420
rect 174813 528386 174847 528420
rect 174905 528386 174939 528420
rect 174997 528386 175031 528420
rect 175089 528386 175123 528420
rect 175181 528386 175215 528420
rect 175273 528386 175307 528420
rect 175365 528386 175399 528420
rect 175457 528386 175491 528420
rect 175549 528386 175583 528420
rect 175641 528386 175675 528420
rect 175733 528386 175767 528420
rect 175825 528386 175859 528420
rect 175917 528386 175951 528420
rect 176009 528386 176043 528420
rect 176101 528386 176135 528420
rect 176193 528386 176227 528420
rect 176285 528386 176319 528420
rect 176377 528386 176411 528420
rect 176469 528386 176503 528420
rect 176561 528386 176595 528420
rect 176653 528386 176687 528420
rect 176745 528386 176779 528420
rect 176837 528386 176871 528420
rect 176929 528386 176963 528420
rect 177021 528386 177055 528420
rect 177113 528386 177147 528420
rect 177205 528386 177239 528420
rect 177297 528386 177331 528420
rect 177389 528386 177423 528420
rect 177481 528386 177515 528420
rect 177573 528386 177607 528420
rect 177665 528386 177699 528420
rect 177757 528386 177791 528420
rect 177849 528386 177883 528420
rect 177941 528386 177975 528420
rect 178033 528386 178067 528420
rect 178125 528386 178159 528420
rect 178217 528386 178251 528420
rect 178309 528386 178343 528420
rect 178401 528386 178435 528420
rect 178493 528386 178527 528420
rect 178585 528386 178619 528420
rect 178677 528386 178711 528420
rect 178769 528386 178803 528420
rect 178861 528386 178895 528420
rect 178953 528386 178987 528420
rect 179045 528386 179079 528420
rect 179137 528386 179171 528420
rect 179229 528386 179263 528420
rect 179321 528386 179355 528420
rect 179413 528386 179447 528420
rect 179505 528386 179539 528420
rect 179597 528386 179631 528420
rect 179689 528386 179723 528420
rect 179781 528386 179815 528420
rect 179873 528386 179907 528420
rect 179965 528386 179999 528420
rect 180057 528386 180091 528420
rect 180149 528386 180183 528420
rect 180241 528386 180275 528420
rect 180333 528386 180367 528420
rect 180425 528386 180459 528420
rect 180517 528386 180551 528420
rect 180609 528386 180643 528420
rect 180701 528386 180735 528420
rect 180793 528386 180827 528420
rect 180885 528386 180919 528420
rect 180977 528386 181011 528420
rect 181069 528386 181103 528420
rect 181161 528386 181195 528420
rect 181253 528386 181287 528420
rect 181345 528386 181379 528420
rect 181437 528386 181471 528420
rect 181529 528386 181563 528420
rect 181621 528386 181655 528420
rect 181713 528386 181747 528420
rect 181805 528386 181839 528420
rect 181897 528386 181931 528420
rect 181989 528386 182023 528420
rect 182081 528386 182115 528420
rect 182173 528386 182207 528420
rect 182265 528386 182299 528420
rect 182357 528386 182391 528420
rect 182449 528386 182483 528420
rect 182541 528386 182575 528420
rect 182633 528386 182667 528420
rect 182725 528386 182759 528420
rect 182817 528386 182851 528420
rect 182909 528386 182943 528420
rect 183001 528386 183035 528420
rect 183093 528386 183127 528420
rect 183185 528386 183219 528420
rect 183277 528386 183311 528420
rect 183369 528386 183403 528420
rect 183461 528386 183495 528420
rect 183553 528386 183587 528420
rect 183645 528386 183679 528420
rect 183737 528386 183771 528420
rect 183829 528386 183863 528420
rect 183921 528386 183955 528420
rect 184013 528386 184047 528420
rect 184105 528386 184139 528420
rect 184197 528386 184231 528420
rect 184289 528386 184323 528420
rect 184381 528386 184415 528420
rect 184473 528386 184507 528420
rect 184565 528386 184599 528420
rect 184657 528386 184691 528420
rect 184749 528386 184783 528420
rect 184841 528386 184875 528420
rect 184933 528386 184967 528420
rect 185025 528386 185059 528420
rect 185117 528386 185151 528420
rect 185209 528386 185243 528420
rect 185301 528386 185335 528420
rect 185393 528386 185427 528420
rect 185485 528386 185519 528420
rect 185577 528386 185611 528420
rect 185669 528386 185703 528420
rect 185761 528386 185795 528420
rect 185853 528386 185887 528420
rect 185945 528386 185979 528420
rect 186037 528386 186071 528420
rect 186129 528386 186163 528420
rect 186221 528386 186255 528420
rect 186313 528386 186347 528420
rect 186405 528386 186439 528420
rect 186497 528386 186531 528420
rect 186589 528386 186623 528420
rect 186681 528386 186715 528420
rect 186773 528386 186807 528420
rect 186865 528386 186899 528420
rect 186957 528386 186991 528420
rect 187049 528386 187083 528420
rect 187141 528386 187175 528420
rect 187233 528386 187267 528420
rect 187325 528386 187359 528420
rect 187417 528386 187451 528420
rect 176101 528154 176104 528182
rect 176104 528154 176135 528182
rect 176101 528148 176135 528154
rect 176194 528173 176228 528182
rect 176194 528148 176206 528173
rect 176206 528148 176228 528173
rect 176377 528216 176411 528250
rect 176275 528028 176309 528046
rect 176275 528012 176309 528028
rect 176561 528148 176595 528182
rect 176833 528216 176867 528250
rect 176905 528234 176939 528250
rect 176905 528216 176929 528234
rect 176929 528216 176939 528234
rect 176653 528012 176687 528046
rect 177277 528164 177303 528182
rect 177303 528164 177311 528182
rect 177277 528148 177311 528164
rect 177849 528294 177883 528318
rect 177553 528216 177587 528250
rect 177493 528162 177509 528187
rect 177509 528162 177527 528187
rect 177493 528153 177527 528162
rect 177849 528284 177877 528294
rect 177877 528284 177883 528294
rect 177277 528038 177308 528046
rect 177308 528038 177311 528046
rect 177277 528012 177311 528038
rect 178953 528291 178959 528318
rect 178959 528291 178987 528318
rect 178953 528284 178987 528291
rect 178125 528154 178151 528182
rect 178151 528154 178159 528182
rect 178125 528148 178159 528154
rect 177941 528041 177975 528046
rect 177941 528012 177947 528041
rect 177947 528012 177975 528041
rect 179321 528148 179355 528182
rect 179413 528284 179447 528318
rect 180977 528291 180983 528318
rect 180983 528291 181011 528318
rect 180977 528284 181011 528291
rect 179505 528080 179539 528114
rect 181345 528148 181379 528182
rect 181437 528284 181471 528318
rect 181529 528080 181563 528114
rect 172237 527842 172271 527876
rect 172329 527842 172363 527876
rect 172421 527842 172455 527876
rect 172513 527842 172547 527876
rect 172605 527842 172639 527876
rect 172697 527842 172731 527876
rect 172789 527842 172823 527876
rect 172881 527842 172915 527876
rect 172973 527842 173007 527876
rect 173065 527842 173099 527876
rect 173157 527842 173191 527876
rect 173249 527842 173283 527876
rect 173341 527842 173375 527876
rect 173433 527842 173467 527876
rect 173525 527842 173559 527876
rect 173617 527842 173651 527876
rect 173709 527842 173743 527876
rect 173801 527842 173835 527876
rect 173893 527842 173927 527876
rect 173985 527842 174019 527876
rect 174077 527842 174111 527876
rect 174169 527842 174203 527876
rect 174261 527842 174295 527876
rect 174353 527842 174387 527876
rect 174445 527842 174479 527876
rect 174537 527842 174571 527876
rect 174629 527842 174663 527876
rect 174721 527842 174755 527876
rect 174813 527842 174847 527876
rect 174905 527842 174939 527876
rect 174997 527842 175031 527876
rect 175089 527842 175123 527876
rect 175181 527842 175215 527876
rect 175273 527842 175307 527876
rect 175365 527842 175399 527876
rect 175457 527842 175491 527876
rect 175549 527842 175583 527876
rect 175641 527842 175675 527876
rect 175733 527842 175767 527876
rect 175825 527842 175859 527876
rect 175917 527842 175951 527876
rect 176009 527842 176043 527876
rect 176101 527842 176135 527876
rect 176193 527842 176227 527876
rect 176285 527842 176319 527876
rect 176377 527842 176411 527876
rect 176469 527842 176503 527876
rect 176561 527842 176595 527876
rect 176653 527842 176687 527876
rect 176745 527842 176779 527876
rect 176837 527842 176871 527876
rect 176929 527842 176963 527876
rect 177021 527842 177055 527876
rect 177113 527842 177147 527876
rect 177205 527842 177239 527876
rect 177297 527842 177331 527876
rect 177389 527842 177423 527876
rect 177481 527842 177515 527876
rect 177573 527842 177607 527876
rect 177665 527842 177699 527876
rect 177757 527842 177791 527876
rect 177849 527842 177883 527876
rect 177941 527842 177975 527876
rect 178033 527842 178067 527876
rect 178125 527842 178159 527876
rect 178217 527842 178251 527876
rect 178309 527842 178343 527876
rect 178401 527842 178435 527876
rect 178493 527842 178527 527876
rect 178585 527842 178619 527876
rect 178677 527842 178711 527876
rect 178769 527842 178803 527876
rect 178861 527842 178895 527876
rect 178953 527842 178987 527876
rect 179045 527842 179079 527876
rect 179137 527842 179171 527876
rect 179229 527842 179263 527876
rect 179321 527842 179355 527876
rect 179413 527842 179447 527876
rect 179505 527842 179539 527876
rect 179597 527842 179631 527876
rect 179689 527842 179723 527876
rect 179781 527842 179815 527876
rect 179873 527842 179907 527876
rect 179965 527842 179999 527876
rect 180057 527842 180091 527876
rect 180149 527842 180183 527876
rect 180241 527842 180275 527876
rect 180333 527842 180367 527876
rect 180425 527842 180459 527876
rect 180517 527842 180551 527876
rect 180609 527842 180643 527876
rect 180701 527842 180735 527876
rect 180793 527842 180827 527876
rect 180885 527842 180919 527876
rect 180977 527842 181011 527876
rect 181069 527842 181103 527876
rect 181161 527842 181195 527876
rect 181253 527842 181287 527876
rect 181345 527842 181379 527876
rect 181437 527842 181471 527876
rect 181529 527842 181563 527876
rect 181621 527842 181655 527876
rect 181713 527842 181747 527876
rect 181805 527842 181839 527876
rect 181897 527842 181931 527876
rect 181989 527842 182023 527876
rect 182081 527842 182115 527876
rect 182173 527842 182207 527876
rect 182265 527842 182299 527876
rect 182357 527842 182391 527876
rect 182449 527842 182483 527876
rect 182541 527842 182575 527876
rect 182633 527842 182667 527876
rect 182725 527842 182759 527876
rect 182817 527842 182851 527876
rect 182909 527842 182943 527876
rect 183001 527842 183035 527876
rect 183093 527842 183127 527876
rect 183185 527842 183219 527876
rect 183277 527842 183311 527876
rect 183369 527842 183403 527876
rect 183461 527842 183495 527876
rect 183553 527842 183587 527876
rect 183645 527842 183679 527876
rect 183737 527842 183771 527876
rect 183829 527842 183863 527876
rect 183921 527842 183955 527876
rect 184013 527842 184047 527876
rect 184105 527842 184139 527876
rect 184197 527842 184231 527876
rect 184289 527842 184323 527876
rect 184381 527842 184415 527876
rect 184473 527842 184507 527876
rect 184565 527842 184599 527876
rect 184657 527842 184691 527876
rect 184749 527842 184783 527876
rect 184841 527842 184875 527876
rect 184933 527842 184967 527876
rect 185025 527842 185059 527876
rect 185117 527842 185151 527876
rect 185209 527842 185243 527876
rect 185301 527842 185335 527876
rect 185393 527842 185427 527876
rect 185485 527842 185519 527876
rect 185577 527842 185611 527876
rect 185669 527842 185703 527876
rect 185761 527842 185795 527876
rect 185853 527842 185887 527876
rect 185945 527842 185979 527876
rect 186037 527842 186071 527876
rect 186129 527842 186163 527876
rect 186221 527842 186255 527876
rect 186313 527842 186347 527876
rect 186405 527842 186439 527876
rect 186497 527842 186531 527876
rect 186589 527842 186623 527876
rect 186681 527842 186715 527876
rect 186773 527842 186807 527876
rect 186865 527842 186899 527876
rect 186957 527842 186991 527876
rect 187049 527842 187083 527876
rect 187141 527842 187175 527876
rect 187233 527842 187267 527876
rect 187325 527842 187359 527876
rect 187417 527842 187451 527876
rect 176377 527740 176402 527774
rect 176402 527740 176411 527774
rect 177021 527604 177055 527638
rect 178953 527740 178978 527774
rect 178978 527740 178987 527774
rect 179505 527604 179539 527638
rect 172237 527298 172271 527332
rect 172329 527298 172363 527332
rect 172421 527298 172455 527332
rect 172513 527298 172547 527332
rect 172605 527298 172639 527332
rect 172697 527298 172731 527332
rect 172789 527298 172823 527332
rect 172881 527298 172915 527332
rect 172973 527298 173007 527332
rect 173065 527298 173099 527332
rect 173157 527298 173191 527332
rect 173249 527298 173283 527332
rect 173341 527298 173375 527332
rect 173433 527298 173467 527332
rect 173525 527298 173559 527332
rect 173617 527298 173651 527332
rect 173709 527298 173743 527332
rect 173801 527298 173835 527332
rect 173893 527298 173927 527332
rect 173985 527298 174019 527332
rect 174077 527298 174111 527332
rect 174169 527298 174203 527332
rect 174261 527298 174295 527332
rect 174353 527298 174387 527332
rect 174445 527298 174479 527332
rect 174537 527298 174571 527332
rect 174629 527298 174663 527332
rect 174721 527298 174755 527332
rect 174813 527298 174847 527332
rect 174905 527298 174939 527332
rect 174997 527298 175031 527332
rect 175089 527298 175123 527332
rect 175181 527298 175215 527332
rect 175273 527298 175307 527332
rect 175365 527298 175399 527332
rect 175457 527298 175491 527332
rect 175549 527298 175583 527332
rect 175641 527298 175675 527332
rect 175733 527298 175767 527332
rect 175825 527298 175859 527332
rect 175917 527298 175951 527332
rect 176009 527298 176043 527332
rect 176101 527298 176135 527332
rect 176193 527298 176227 527332
rect 176285 527298 176319 527332
rect 176377 527298 176411 527332
rect 176469 527298 176503 527332
rect 176561 527298 176595 527332
rect 176653 527298 176687 527332
rect 176745 527298 176779 527332
rect 176837 527298 176871 527332
rect 176929 527298 176963 527332
rect 177021 527298 177055 527332
rect 177113 527298 177147 527332
rect 177205 527298 177239 527332
rect 177297 527298 177331 527332
rect 177389 527298 177423 527332
rect 177481 527298 177515 527332
rect 177573 527298 177607 527332
rect 177665 527298 177699 527332
rect 177757 527298 177791 527332
rect 177849 527298 177883 527332
rect 177941 527298 177975 527332
rect 178033 527298 178067 527332
rect 178125 527298 178159 527332
rect 178217 527298 178251 527332
rect 178309 527298 178343 527332
rect 178401 527298 178435 527332
rect 178493 527298 178527 527332
rect 178585 527298 178619 527332
rect 178677 527298 178711 527332
rect 178769 527298 178803 527332
rect 178861 527298 178895 527332
rect 178953 527298 178987 527332
rect 179045 527298 179079 527332
rect 179137 527298 179171 527332
rect 179229 527298 179263 527332
rect 179321 527298 179355 527332
rect 179413 527298 179447 527332
rect 179505 527298 179539 527332
rect 179597 527298 179631 527332
rect 179689 527298 179723 527332
rect 179781 527298 179815 527332
rect 179873 527298 179907 527332
rect 179965 527298 179999 527332
rect 180057 527298 180091 527332
rect 180149 527298 180183 527332
rect 180241 527298 180275 527332
rect 180333 527298 180367 527332
rect 180425 527298 180459 527332
rect 180517 527298 180551 527332
rect 180609 527298 180643 527332
rect 180701 527298 180735 527332
rect 180793 527298 180827 527332
rect 180885 527298 180919 527332
rect 180977 527298 181011 527332
rect 181069 527298 181103 527332
rect 181161 527298 181195 527332
rect 181253 527298 181287 527332
rect 181345 527298 181379 527332
rect 181437 527298 181471 527332
rect 181529 527298 181563 527332
rect 181621 527298 181655 527332
rect 181713 527298 181747 527332
rect 181805 527298 181839 527332
rect 181897 527298 181931 527332
rect 181989 527298 182023 527332
rect 182081 527298 182115 527332
rect 182173 527298 182207 527332
rect 182265 527298 182299 527332
rect 182357 527298 182391 527332
rect 182449 527298 182483 527332
rect 182541 527298 182575 527332
rect 182633 527298 182667 527332
rect 182725 527298 182759 527332
rect 182817 527298 182851 527332
rect 182909 527298 182943 527332
rect 183001 527298 183035 527332
rect 183093 527298 183127 527332
rect 183185 527298 183219 527332
rect 183277 527298 183311 527332
rect 183369 527298 183403 527332
rect 183461 527298 183495 527332
rect 183553 527298 183587 527332
rect 183645 527298 183679 527332
rect 183737 527298 183771 527332
rect 183829 527298 183863 527332
rect 183921 527298 183955 527332
rect 184013 527298 184047 527332
rect 184105 527298 184139 527332
rect 184197 527298 184231 527332
rect 184289 527298 184323 527332
rect 184381 527298 184415 527332
rect 184473 527298 184507 527332
rect 184565 527298 184599 527332
rect 184657 527298 184691 527332
rect 184749 527298 184783 527332
rect 184841 527298 184875 527332
rect 184933 527298 184967 527332
rect 185025 527298 185059 527332
rect 185117 527298 185151 527332
rect 185209 527298 185243 527332
rect 185301 527298 185335 527332
rect 185393 527298 185427 527332
rect 185485 527298 185519 527332
rect 185577 527298 185611 527332
rect 185669 527298 185703 527332
rect 185761 527298 185795 527332
rect 185853 527298 185887 527332
rect 185945 527298 185979 527332
rect 186037 527298 186071 527332
rect 186129 527298 186163 527332
rect 186221 527298 186255 527332
rect 186313 527298 186347 527332
rect 186405 527298 186439 527332
rect 186497 527298 186531 527332
rect 186589 527298 186623 527332
rect 186681 527298 186715 527332
rect 186773 527298 186807 527332
rect 186865 527298 186899 527332
rect 186957 527298 186991 527332
rect 187049 527298 187083 527332
rect 187141 527298 187175 527332
rect 187233 527298 187267 527332
rect 187325 527298 187359 527332
rect 187417 527298 187451 527332
rect 172237 526754 172271 526788
rect 172329 526754 172363 526788
rect 172421 526754 172455 526788
rect 172513 526754 172547 526788
rect 172605 526754 172639 526788
rect 172697 526754 172731 526788
rect 172789 526754 172823 526788
rect 172881 526754 172915 526788
rect 172973 526754 173007 526788
rect 173065 526754 173099 526788
rect 173157 526754 173191 526788
rect 173249 526754 173283 526788
rect 173341 526754 173375 526788
rect 173433 526754 173467 526788
rect 173525 526754 173559 526788
rect 173617 526754 173651 526788
rect 173709 526754 173743 526788
rect 173801 526754 173835 526788
rect 173893 526754 173927 526788
rect 173985 526754 174019 526788
rect 174077 526754 174111 526788
rect 174169 526754 174203 526788
rect 174261 526754 174295 526788
rect 174353 526754 174387 526788
rect 174445 526754 174479 526788
rect 174537 526754 174571 526788
rect 174629 526754 174663 526788
rect 174721 526754 174755 526788
rect 174813 526754 174847 526788
rect 174905 526754 174939 526788
rect 174997 526754 175031 526788
rect 175089 526754 175123 526788
rect 175181 526754 175215 526788
rect 175273 526754 175307 526788
rect 175365 526754 175399 526788
rect 175457 526754 175491 526788
rect 175549 526754 175583 526788
rect 175641 526754 175675 526788
rect 175733 526754 175767 526788
rect 175825 526754 175859 526788
rect 175917 526754 175951 526788
rect 176009 526754 176043 526788
rect 176101 526754 176135 526788
rect 176193 526754 176227 526788
rect 176285 526754 176319 526788
rect 176377 526754 176411 526788
rect 176469 526754 176503 526788
rect 176561 526754 176595 526788
rect 176653 526754 176687 526788
rect 176745 526754 176779 526788
rect 176837 526754 176871 526788
rect 176929 526754 176963 526788
rect 177021 526754 177055 526788
rect 177113 526754 177147 526788
rect 177205 526754 177239 526788
rect 177297 526754 177331 526788
rect 177389 526754 177423 526788
rect 177481 526754 177515 526788
rect 177573 526754 177607 526788
rect 177665 526754 177699 526788
rect 177757 526754 177791 526788
rect 177849 526754 177883 526788
rect 177941 526754 177975 526788
rect 178033 526754 178067 526788
rect 178125 526754 178159 526788
rect 178217 526754 178251 526788
rect 178309 526754 178343 526788
rect 178401 526754 178435 526788
rect 178493 526754 178527 526788
rect 178585 526754 178619 526788
rect 178677 526754 178711 526788
rect 178769 526754 178803 526788
rect 178861 526754 178895 526788
rect 178953 526754 178987 526788
rect 179045 526754 179079 526788
rect 179137 526754 179171 526788
rect 179229 526754 179263 526788
rect 179321 526754 179355 526788
rect 179413 526754 179447 526788
rect 179505 526754 179539 526788
rect 179597 526754 179631 526788
rect 179689 526754 179723 526788
rect 179781 526754 179815 526788
rect 179873 526754 179907 526788
rect 179965 526754 179999 526788
rect 180057 526754 180091 526788
rect 180149 526754 180183 526788
rect 180241 526754 180275 526788
rect 180333 526754 180367 526788
rect 180425 526754 180459 526788
rect 180517 526754 180551 526788
rect 180609 526754 180643 526788
rect 180701 526754 180735 526788
rect 180793 526754 180827 526788
rect 180885 526754 180919 526788
rect 180977 526754 181011 526788
rect 181069 526754 181103 526788
rect 181161 526754 181195 526788
rect 181253 526754 181287 526788
rect 181345 526754 181379 526788
rect 181437 526754 181471 526788
rect 181529 526754 181563 526788
rect 181621 526754 181655 526788
rect 181713 526754 181747 526788
rect 181805 526754 181839 526788
rect 181897 526754 181931 526788
rect 181989 526754 182023 526788
rect 182081 526754 182115 526788
rect 182173 526754 182207 526788
rect 182265 526754 182299 526788
rect 182357 526754 182391 526788
rect 182449 526754 182483 526788
rect 182541 526754 182575 526788
rect 182633 526754 182667 526788
rect 182725 526754 182759 526788
rect 182817 526754 182851 526788
rect 182909 526754 182943 526788
rect 183001 526754 183035 526788
rect 183093 526754 183127 526788
rect 183185 526754 183219 526788
rect 183277 526754 183311 526788
rect 183369 526754 183403 526788
rect 183461 526754 183495 526788
rect 183553 526754 183587 526788
rect 183645 526754 183679 526788
rect 183737 526754 183771 526788
rect 183829 526754 183863 526788
rect 183921 526754 183955 526788
rect 184013 526754 184047 526788
rect 184105 526754 184139 526788
rect 184197 526754 184231 526788
rect 184289 526754 184323 526788
rect 184381 526754 184415 526788
rect 184473 526754 184507 526788
rect 184565 526754 184599 526788
rect 184657 526754 184691 526788
rect 184749 526754 184783 526788
rect 184841 526754 184875 526788
rect 184933 526754 184967 526788
rect 185025 526754 185059 526788
rect 185117 526754 185151 526788
rect 185209 526754 185243 526788
rect 185301 526754 185335 526788
rect 185393 526754 185427 526788
rect 185485 526754 185519 526788
rect 185577 526754 185611 526788
rect 185669 526754 185703 526788
rect 185761 526754 185795 526788
rect 185853 526754 185887 526788
rect 185945 526754 185979 526788
rect 186037 526754 186071 526788
rect 186129 526754 186163 526788
rect 186221 526754 186255 526788
rect 186313 526754 186347 526788
rect 186405 526754 186439 526788
rect 186497 526754 186531 526788
rect 186589 526754 186623 526788
rect 186681 526754 186715 526788
rect 186773 526754 186807 526788
rect 186865 526754 186899 526788
rect 186957 526754 186991 526788
rect 187049 526754 187083 526788
rect 187141 526754 187175 526788
rect 187233 526754 187267 526788
rect 187325 526754 187359 526788
rect 187417 526754 187451 526788
rect 172237 526210 172271 526244
rect 172329 526210 172363 526244
rect 172421 526210 172455 526244
rect 172513 526210 172547 526244
rect 172605 526210 172639 526244
rect 172697 526210 172731 526244
rect 172789 526210 172823 526244
rect 172881 526210 172915 526244
rect 172973 526210 173007 526244
rect 173065 526210 173099 526244
rect 173157 526210 173191 526244
rect 173249 526210 173283 526244
rect 173341 526210 173375 526244
rect 173433 526210 173467 526244
rect 173525 526210 173559 526244
rect 173617 526210 173651 526244
rect 173709 526210 173743 526244
rect 173801 526210 173835 526244
rect 173893 526210 173927 526244
rect 173985 526210 174019 526244
rect 174077 526210 174111 526244
rect 174169 526210 174203 526244
rect 174261 526210 174295 526244
rect 174353 526210 174387 526244
rect 174445 526210 174479 526244
rect 174537 526210 174571 526244
rect 174629 526210 174663 526244
rect 174721 526210 174755 526244
rect 174813 526210 174847 526244
rect 174905 526210 174939 526244
rect 174997 526210 175031 526244
rect 175089 526210 175123 526244
rect 175181 526210 175215 526244
rect 175273 526210 175307 526244
rect 175365 526210 175399 526244
rect 175457 526210 175491 526244
rect 175549 526210 175583 526244
rect 175641 526210 175675 526244
rect 175733 526210 175767 526244
rect 175825 526210 175859 526244
rect 175917 526210 175951 526244
rect 176009 526210 176043 526244
rect 176101 526210 176135 526244
rect 176193 526210 176227 526244
rect 176285 526210 176319 526244
rect 176377 526210 176411 526244
rect 176469 526210 176503 526244
rect 176561 526210 176595 526244
rect 176653 526210 176687 526244
rect 176745 526210 176779 526244
rect 176837 526210 176871 526244
rect 176929 526210 176963 526244
rect 177021 526210 177055 526244
rect 177113 526210 177147 526244
rect 177205 526210 177239 526244
rect 177297 526210 177331 526244
rect 177389 526210 177423 526244
rect 177481 526210 177515 526244
rect 177573 526210 177607 526244
rect 177665 526210 177699 526244
rect 177757 526210 177791 526244
rect 177849 526210 177883 526244
rect 177941 526210 177975 526244
rect 178033 526210 178067 526244
rect 178125 526210 178159 526244
rect 178217 526210 178251 526244
rect 178309 526210 178343 526244
rect 178401 526210 178435 526244
rect 178493 526210 178527 526244
rect 178585 526210 178619 526244
rect 178677 526210 178711 526244
rect 178769 526210 178803 526244
rect 178861 526210 178895 526244
rect 178953 526210 178987 526244
rect 179045 526210 179079 526244
rect 179137 526210 179171 526244
rect 179229 526210 179263 526244
rect 179321 526210 179355 526244
rect 179413 526210 179447 526244
rect 179505 526210 179539 526244
rect 179597 526210 179631 526244
rect 179689 526210 179723 526244
rect 179781 526210 179815 526244
rect 179873 526210 179907 526244
rect 179965 526210 179999 526244
rect 180057 526210 180091 526244
rect 180149 526210 180183 526244
rect 180241 526210 180275 526244
rect 180333 526210 180367 526244
rect 180425 526210 180459 526244
rect 180517 526210 180551 526244
rect 180609 526210 180643 526244
rect 180701 526210 180735 526244
rect 180793 526210 180827 526244
rect 180885 526210 180919 526244
rect 180977 526210 181011 526244
rect 181069 526210 181103 526244
rect 181161 526210 181195 526244
rect 181253 526210 181287 526244
rect 181345 526210 181379 526244
rect 181437 526210 181471 526244
rect 181529 526210 181563 526244
rect 181621 526210 181655 526244
rect 181713 526210 181747 526244
rect 181805 526210 181839 526244
rect 181897 526210 181931 526244
rect 181989 526210 182023 526244
rect 182081 526210 182115 526244
rect 182173 526210 182207 526244
rect 182265 526210 182299 526244
rect 182357 526210 182391 526244
rect 182449 526210 182483 526244
rect 182541 526210 182575 526244
rect 182633 526210 182667 526244
rect 182725 526210 182759 526244
rect 182817 526210 182851 526244
rect 182909 526210 182943 526244
rect 183001 526210 183035 526244
rect 183093 526210 183127 526244
rect 183185 526210 183219 526244
rect 183277 526210 183311 526244
rect 183369 526210 183403 526244
rect 183461 526210 183495 526244
rect 183553 526210 183587 526244
rect 183645 526210 183679 526244
rect 183737 526210 183771 526244
rect 183829 526210 183863 526244
rect 183921 526210 183955 526244
rect 184013 526210 184047 526244
rect 184105 526210 184139 526244
rect 184197 526210 184231 526244
rect 184289 526210 184323 526244
rect 184381 526210 184415 526244
rect 184473 526210 184507 526244
rect 184565 526210 184599 526244
rect 184657 526210 184691 526244
rect 184749 526210 184783 526244
rect 184841 526210 184875 526244
rect 184933 526210 184967 526244
rect 185025 526210 185059 526244
rect 185117 526210 185151 526244
rect 185209 526210 185243 526244
rect 185301 526210 185335 526244
rect 185393 526210 185427 526244
rect 185485 526210 185519 526244
rect 185577 526210 185611 526244
rect 185669 526210 185703 526244
rect 185761 526210 185795 526244
rect 185853 526210 185887 526244
rect 185945 526210 185979 526244
rect 186037 526210 186071 526244
rect 186129 526210 186163 526244
rect 186221 526210 186255 526244
rect 186313 526210 186347 526244
rect 186405 526210 186439 526244
rect 186497 526210 186531 526244
rect 186589 526210 186623 526244
rect 186681 526210 186715 526244
rect 186773 526210 186807 526244
rect 186865 526210 186899 526244
rect 186957 526210 186991 526244
rect 187049 526210 187083 526244
rect 187141 526210 187175 526244
rect 187233 526210 187267 526244
rect 187325 526210 187359 526244
rect 187417 526210 187451 526244
rect 172237 525666 172271 525700
rect 172329 525666 172363 525700
rect 172421 525666 172455 525700
rect 172513 525666 172547 525700
rect 172605 525666 172639 525700
rect 172697 525666 172731 525700
rect 172789 525666 172823 525700
rect 172881 525666 172915 525700
rect 172973 525666 173007 525700
rect 173065 525666 173099 525700
rect 173157 525666 173191 525700
rect 173249 525666 173283 525700
rect 173341 525666 173375 525700
rect 173433 525666 173467 525700
rect 173525 525666 173559 525700
rect 173617 525666 173651 525700
rect 173709 525666 173743 525700
rect 173801 525666 173835 525700
rect 173893 525666 173927 525700
rect 173985 525666 174019 525700
rect 174077 525666 174111 525700
rect 174169 525666 174203 525700
rect 174261 525666 174295 525700
rect 174353 525666 174387 525700
rect 174445 525666 174479 525700
rect 174537 525666 174571 525700
rect 174629 525666 174663 525700
rect 174721 525666 174755 525700
rect 174813 525666 174847 525700
rect 174905 525666 174939 525700
rect 174997 525666 175031 525700
rect 175089 525666 175123 525700
rect 175181 525666 175215 525700
rect 175273 525666 175307 525700
rect 175365 525666 175399 525700
rect 175457 525666 175491 525700
rect 175549 525666 175583 525700
rect 175641 525666 175675 525700
rect 175733 525666 175767 525700
rect 175825 525666 175859 525700
rect 175917 525666 175951 525700
rect 176009 525666 176043 525700
rect 176101 525666 176135 525700
rect 176193 525666 176227 525700
rect 176285 525666 176319 525700
rect 176377 525666 176411 525700
rect 176469 525666 176503 525700
rect 176561 525666 176595 525700
rect 176653 525666 176687 525700
rect 176745 525666 176779 525700
rect 176837 525666 176871 525700
rect 176929 525666 176963 525700
rect 177021 525666 177055 525700
rect 177113 525666 177147 525700
rect 177205 525666 177239 525700
rect 177297 525666 177331 525700
rect 177389 525666 177423 525700
rect 177481 525666 177515 525700
rect 177573 525666 177607 525700
rect 177665 525666 177699 525700
rect 177757 525666 177791 525700
rect 177849 525666 177883 525700
rect 177941 525666 177975 525700
rect 178033 525666 178067 525700
rect 178125 525666 178159 525700
rect 178217 525666 178251 525700
rect 178309 525666 178343 525700
rect 178401 525666 178435 525700
rect 178493 525666 178527 525700
rect 178585 525666 178619 525700
rect 178677 525666 178711 525700
rect 178769 525666 178803 525700
rect 178861 525666 178895 525700
rect 178953 525666 178987 525700
rect 179045 525666 179079 525700
rect 179137 525666 179171 525700
rect 179229 525666 179263 525700
rect 179321 525666 179355 525700
rect 179413 525666 179447 525700
rect 179505 525666 179539 525700
rect 179597 525666 179631 525700
rect 179689 525666 179723 525700
rect 179781 525666 179815 525700
rect 179873 525666 179907 525700
rect 179965 525666 179999 525700
rect 180057 525666 180091 525700
rect 180149 525666 180183 525700
rect 180241 525666 180275 525700
rect 180333 525666 180367 525700
rect 180425 525666 180459 525700
rect 180517 525666 180551 525700
rect 180609 525666 180643 525700
rect 180701 525666 180735 525700
rect 180793 525666 180827 525700
rect 180885 525666 180919 525700
rect 180977 525666 181011 525700
rect 181069 525666 181103 525700
rect 181161 525666 181195 525700
rect 181253 525666 181287 525700
rect 181345 525666 181379 525700
rect 181437 525666 181471 525700
rect 181529 525666 181563 525700
rect 181621 525666 181655 525700
rect 181713 525666 181747 525700
rect 181805 525666 181839 525700
rect 181897 525666 181931 525700
rect 181989 525666 182023 525700
rect 182081 525666 182115 525700
rect 182173 525666 182207 525700
rect 182265 525666 182299 525700
rect 182357 525666 182391 525700
rect 182449 525666 182483 525700
rect 182541 525666 182575 525700
rect 182633 525666 182667 525700
rect 182725 525666 182759 525700
rect 182817 525666 182851 525700
rect 182909 525666 182943 525700
rect 183001 525666 183035 525700
rect 183093 525666 183127 525700
rect 183185 525666 183219 525700
rect 183277 525666 183311 525700
rect 183369 525666 183403 525700
rect 183461 525666 183495 525700
rect 183553 525666 183587 525700
rect 183645 525666 183679 525700
rect 183737 525666 183771 525700
rect 183829 525666 183863 525700
rect 183921 525666 183955 525700
rect 184013 525666 184047 525700
rect 184105 525666 184139 525700
rect 184197 525666 184231 525700
rect 184289 525666 184323 525700
rect 184381 525666 184415 525700
rect 184473 525666 184507 525700
rect 184565 525666 184599 525700
rect 184657 525666 184691 525700
rect 184749 525666 184783 525700
rect 184841 525666 184875 525700
rect 184933 525666 184967 525700
rect 185025 525666 185059 525700
rect 185117 525666 185151 525700
rect 185209 525666 185243 525700
rect 185301 525666 185335 525700
rect 185393 525666 185427 525700
rect 185485 525666 185519 525700
rect 185577 525666 185611 525700
rect 185669 525666 185703 525700
rect 185761 525666 185795 525700
rect 185853 525666 185887 525700
rect 185945 525666 185979 525700
rect 186037 525666 186071 525700
rect 186129 525666 186163 525700
rect 186221 525666 186255 525700
rect 186313 525666 186347 525700
rect 186405 525666 186439 525700
rect 186497 525666 186531 525700
rect 186589 525666 186623 525700
rect 186681 525666 186715 525700
rect 186773 525666 186807 525700
rect 186865 525666 186899 525700
rect 186957 525666 186991 525700
rect 187049 525666 187083 525700
rect 187141 525666 187175 525700
rect 187233 525666 187267 525700
rect 187325 525666 187359 525700
rect 187417 525666 187451 525700
rect 172237 525122 172271 525156
rect 172329 525122 172363 525156
rect 172421 525122 172455 525156
rect 172513 525122 172547 525156
rect 172605 525122 172639 525156
rect 172697 525122 172731 525156
rect 172789 525122 172823 525156
rect 172881 525122 172915 525156
rect 172973 525122 173007 525156
rect 173065 525122 173099 525156
rect 173157 525122 173191 525156
rect 173249 525122 173283 525156
rect 173341 525122 173375 525156
rect 173433 525122 173467 525156
rect 173525 525122 173559 525156
rect 173617 525122 173651 525156
rect 173709 525122 173743 525156
rect 173801 525122 173835 525156
rect 173893 525122 173927 525156
rect 173985 525122 174019 525156
rect 174077 525122 174111 525156
rect 174169 525122 174203 525156
rect 174261 525122 174295 525156
rect 174353 525122 174387 525156
rect 174445 525122 174479 525156
rect 174537 525122 174571 525156
rect 174629 525122 174663 525156
rect 174721 525122 174755 525156
rect 174813 525122 174847 525156
rect 174905 525122 174939 525156
rect 174997 525122 175031 525156
rect 175089 525122 175123 525156
rect 175181 525122 175215 525156
rect 175273 525122 175307 525156
rect 175365 525122 175399 525156
rect 175457 525122 175491 525156
rect 175549 525122 175583 525156
rect 175641 525122 175675 525156
rect 175733 525122 175767 525156
rect 175825 525122 175859 525156
rect 175917 525122 175951 525156
rect 176009 525122 176043 525156
rect 176101 525122 176135 525156
rect 176193 525122 176227 525156
rect 176285 525122 176319 525156
rect 176377 525122 176411 525156
rect 176469 525122 176503 525156
rect 176561 525122 176595 525156
rect 176653 525122 176687 525156
rect 176745 525122 176779 525156
rect 176837 525122 176871 525156
rect 176929 525122 176963 525156
rect 177021 525122 177055 525156
rect 177113 525122 177147 525156
rect 177205 525122 177239 525156
rect 177297 525122 177331 525156
rect 177389 525122 177423 525156
rect 177481 525122 177515 525156
rect 177573 525122 177607 525156
rect 177665 525122 177699 525156
rect 177757 525122 177791 525156
rect 177849 525122 177883 525156
rect 177941 525122 177975 525156
rect 178033 525122 178067 525156
rect 178125 525122 178159 525156
rect 178217 525122 178251 525156
rect 178309 525122 178343 525156
rect 178401 525122 178435 525156
rect 178493 525122 178527 525156
rect 178585 525122 178619 525156
rect 178677 525122 178711 525156
rect 178769 525122 178803 525156
rect 178861 525122 178895 525156
rect 178953 525122 178987 525156
rect 179045 525122 179079 525156
rect 179137 525122 179171 525156
rect 179229 525122 179263 525156
rect 179321 525122 179355 525156
rect 179413 525122 179447 525156
rect 179505 525122 179539 525156
rect 179597 525122 179631 525156
rect 179689 525122 179723 525156
rect 179781 525122 179815 525156
rect 179873 525122 179907 525156
rect 179965 525122 179999 525156
rect 180057 525122 180091 525156
rect 180149 525122 180183 525156
rect 180241 525122 180275 525156
rect 180333 525122 180367 525156
rect 180425 525122 180459 525156
rect 180517 525122 180551 525156
rect 180609 525122 180643 525156
rect 180701 525122 180735 525156
rect 180793 525122 180827 525156
rect 180885 525122 180919 525156
rect 180977 525122 181011 525156
rect 181069 525122 181103 525156
rect 181161 525122 181195 525156
rect 181253 525122 181287 525156
rect 181345 525122 181379 525156
rect 181437 525122 181471 525156
rect 181529 525122 181563 525156
rect 181621 525122 181655 525156
rect 181713 525122 181747 525156
rect 181805 525122 181839 525156
rect 181897 525122 181931 525156
rect 181989 525122 182023 525156
rect 182081 525122 182115 525156
rect 182173 525122 182207 525156
rect 182265 525122 182299 525156
rect 182357 525122 182391 525156
rect 182449 525122 182483 525156
rect 182541 525122 182575 525156
rect 182633 525122 182667 525156
rect 182725 525122 182759 525156
rect 182817 525122 182851 525156
rect 182909 525122 182943 525156
rect 183001 525122 183035 525156
rect 183093 525122 183127 525156
rect 183185 525122 183219 525156
rect 183277 525122 183311 525156
rect 183369 525122 183403 525156
rect 183461 525122 183495 525156
rect 183553 525122 183587 525156
rect 183645 525122 183679 525156
rect 183737 525122 183771 525156
rect 183829 525122 183863 525156
rect 183921 525122 183955 525156
rect 184013 525122 184047 525156
rect 184105 525122 184139 525156
rect 184197 525122 184231 525156
rect 184289 525122 184323 525156
rect 184381 525122 184415 525156
rect 184473 525122 184507 525156
rect 184565 525122 184599 525156
rect 184657 525122 184691 525156
rect 184749 525122 184783 525156
rect 184841 525122 184875 525156
rect 184933 525122 184967 525156
rect 185025 525122 185059 525156
rect 185117 525122 185151 525156
rect 185209 525122 185243 525156
rect 185301 525122 185335 525156
rect 185393 525122 185427 525156
rect 185485 525122 185519 525156
rect 185577 525122 185611 525156
rect 185669 525122 185703 525156
rect 185761 525122 185795 525156
rect 185853 525122 185887 525156
rect 185945 525122 185979 525156
rect 186037 525122 186071 525156
rect 186129 525122 186163 525156
rect 186221 525122 186255 525156
rect 186313 525122 186347 525156
rect 186405 525122 186439 525156
rect 186497 525122 186531 525156
rect 186589 525122 186623 525156
rect 186681 525122 186715 525156
rect 186773 525122 186807 525156
rect 186865 525122 186899 525156
rect 186957 525122 186991 525156
rect 187049 525122 187083 525156
rect 187141 525122 187175 525156
rect 187233 525122 187267 525156
rect 187325 525122 187359 525156
rect 187417 525122 187451 525156
rect 172237 524578 172271 524612
rect 172329 524578 172363 524612
rect 172421 524578 172455 524612
rect 172513 524578 172547 524612
rect 172605 524578 172639 524612
rect 172697 524578 172731 524612
rect 172789 524578 172823 524612
rect 172881 524578 172915 524612
rect 172973 524578 173007 524612
rect 173065 524578 173099 524612
rect 173157 524578 173191 524612
rect 173249 524578 173283 524612
rect 173341 524578 173375 524612
rect 173433 524578 173467 524612
rect 173525 524578 173559 524612
rect 173617 524578 173651 524612
rect 173709 524578 173743 524612
rect 173801 524578 173835 524612
rect 173893 524578 173927 524612
rect 173985 524578 174019 524612
rect 174077 524578 174111 524612
rect 174169 524578 174203 524612
rect 174261 524578 174295 524612
rect 174353 524578 174387 524612
rect 174445 524578 174479 524612
rect 174537 524578 174571 524612
rect 174629 524578 174663 524612
rect 174721 524578 174755 524612
rect 174813 524578 174847 524612
rect 174905 524578 174939 524612
rect 174997 524578 175031 524612
rect 175089 524578 175123 524612
rect 175181 524578 175215 524612
rect 175273 524578 175307 524612
rect 175365 524578 175399 524612
rect 175457 524578 175491 524612
rect 175549 524578 175583 524612
rect 175641 524578 175675 524612
rect 175733 524578 175767 524612
rect 175825 524578 175859 524612
rect 175917 524578 175951 524612
rect 176009 524578 176043 524612
rect 176101 524578 176135 524612
rect 176193 524578 176227 524612
rect 176285 524578 176319 524612
rect 176377 524578 176411 524612
rect 176469 524578 176503 524612
rect 176561 524578 176595 524612
rect 176653 524578 176687 524612
rect 176745 524578 176779 524612
rect 176837 524578 176871 524612
rect 176929 524578 176963 524612
rect 177021 524578 177055 524612
rect 177113 524578 177147 524612
rect 177205 524578 177239 524612
rect 177297 524578 177331 524612
rect 177389 524578 177423 524612
rect 177481 524578 177515 524612
rect 177573 524578 177607 524612
rect 177665 524578 177699 524612
rect 177757 524578 177791 524612
rect 177849 524578 177883 524612
rect 177941 524578 177975 524612
rect 178033 524578 178067 524612
rect 178125 524578 178159 524612
rect 178217 524578 178251 524612
rect 178309 524578 178343 524612
rect 178401 524578 178435 524612
rect 178493 524578 178527 524612
rect 178585 524578 178619 524612
rect 178677 524578 178711 524612
rect 178769 524578 178803 524612
rect 178861 524578 178895 524612
rect 178953 524578 178987 524612
rect 179045 524578 179079 524612
rect 179137 524578 179171 524612
rect 179229 524578 179263 524612
rect 179321 524578 179355 524612
rect 179413 524578 179447 524612
rect 179505 524578 179539 524612
rect 179597 524578 179631 524612
rect 179689 524578 179723 524612
rect 179781 524578 179815 524612
rect 179873 524578 179907 524612
rect 179965 524578 179999 524612
rect 180057 524578 180091 524612
rect 180149 524578 180183 524612
rect 180241 524578 180275 524612
rect 180333 524578 180367 524612
rect 180425 524578 180459 524612
rect 180517 524578 180551 524612
rect 180609 524578 180643 524612
rect 180701 524578 180735 524612
rect 180793 524578 180827 524612
rect 180885 524578 180919 524612
rect 180977 524578 181011 524612
rect 181069 524578 181103 524612
rect 181161 524578 181195 524612
rect 181253 524578 181287 524612
rect 181345 524578 181379 524612
rect 181437 524578 181471 524612
rect 181529 524578 181563 524612
rect 181621 524578 181655 524612
rect 181713 524578 181747 524612
rect 181805 524578 181839 524612
rect 181897 524578 181931 524612
rect 181989 524578 182023 524612
rect 182081 524578 182115 524612
rect 182173 524578 182207 524612
rect 182265 524578 182299 524612
rect 182357 524578 182391 524612
rect 182449 524578 182483 524612
rect 182541 524578 182575 524612
rect 182633 524578 182667 524612
rect 182725 524578 182759 524612
rect 182817 524578 182851 524612
rect 182909 524578 182943 524612
rect 183001 524578 183035 524612
rect 183093 524578 183127 524612
rect 183185 524578 183219 524612
rect 183277 524578 183311 524612
rect 183369 524578 183403 524612
rect 183461 524578 183495 524612
rect 183553 524578 183587 524612
rect 183645 524578 183679 524612
rect 183737 524578 183771 524612
rect 183829 524578 183863 524612
rect 183921 524578 183955 524612
rect 184013 524578 184047 524612
rect 184105 524578 184139 524612
rect 184197 524578 184231 524612
rect 184289 524578 184323 524612
rect 184381 524578 184415 524612
rect 184473 524578 184507 524612
rect 184565 524578 184599 524612
rect 184657 524578 184691 524612
rect 184749 524578 184783 524612
rect 184841 524578 184875 524612
rect 184933 524578 184967 524612
rect 185025 524578 185059 524612
rect 185117 524578 185151 524612
rect 185209 524578 185243 524612
rect 185301 524578 185335 524612
rect 185393 524578 185427 524612
rect 185485 524578 185519 524612
rect 185577 524578 185611 524612
rect 185669 524578 185703 524612
rect 185761 524578 185795 524612
rect 185853 524578 185887 524612
rect 185945 524578 185979 524612
rect 186037 524578 186071 524612
rect 186129 524578 186163 524612
rect 186221 524578 186255 524612
rect 186313 524578 186347 524612
rect 186405 524578 186439 524612
rect 186497 524578 186531 524612
rect 186589 524578 186623 524612
rect 186681 524578 186715 524612
rect 186773 524578 186807 524612
rect 186865 524578 186899 524612
rect 186957 524578 186991 524612
rect 187049 524578 187083 524612
rect 187141 524578 187175 524612
rect 187233 524578 187267 524612
rect 187325 524578 187359 524612
rect 187417 524578 187451 524612
rect 172237 524034 172271 524068
rect 172329 524034 172363 524068
rect 172421 524034 172455 524068
rect 172513 524034 172547 524068
rect 172605 524034 172639 524068
rect 172697 524034 172731 524068
rect 172789 524034 172823 524068
rect 172881 524034 172915 524068
rect 172973 524034 173007 524068
rect 173065 524034 173099 524068
rect 173157 524034 173191 524068
rect 173249 524034 173283 524068
rect 173341 524034 173375 524068
rect 173433 524034 173467 524068
rect 173525 524034 173559 524068
rect 173617 524034 173651 524068
rect 173709 524034 173743 524068
rect 173801 524034 173835 524068
rect 173893 524034 173927 524068
rect 173985 524034 174019 524068
rect 174077 524034 174111 524068
rect 174169 524034 174203 524068
rect 174261 524034 174295 524068
rect 174353 524034 174387 524068
rect 174445 524034 174479 524068
rect 174537 524034 174571 524068
rect 174629 524034 174663 524068
rect 174721 524034 174755 524068
rect 174813 524034 174847 524068
rect 174905 524034 174939 524068
rect 174997 524034 175031 524068
rect 175089 524034 175123 524068
rect 175181 524034 175215 524068
rect 175273 524034 175307 524068
rect 175365 524034 175399 524068
rect 175457 524034 175491 524068
rect 175549 524034 175583 524068
rect 175641 524034 175675 524068
rect 175733 524034 175767 524068
rect 175825 524034 175859 524068
rect 175917 524034 175951 524068
rect 176009 524034 176043 524068
rect 176101 524034 176135 524068
rect 176193 524034 176227 524068
rect 176285 524034 176319 524068
rect 176377 524034 176411 524068
rect 176469 524034 176503 524068
rect 176561 524034 176595 524068
rect 176653 524034 176687 524068
rect 176745 524034 176779 524068
rect 176837 524034 176871 524068
rect 176929 524034 176963 524068
rect 177021 524034 177055 524068
rect 177113 524034 177147 524068
rect 177205 524034 177239 524068
rect 177297 524034 177331 524068
rect 177389 524034 177423 524068
rect 177481 524034 177515 524068
rect 177573 524034 177607 524068
rect 177665 524034 177699 524068
rect 177757 524034 177791 524068
rect 177849 524034 177883 524068
rect 177941 524034 177975 524068
rect 178033 524034 178067 524068
rect 178125 524034 178159 524068
rect 178217 524034 178251 524068
rect 178309 524034 178343 524068
rect 178401 524034 178435 524068
rect 178493 524034 178527 524068
rect 178585 524034 178619 524068
rect 178677 524034 178711 524068
rect 178769 524034 178803 524068
rect 178861 524034 178895 524068
rect 178953 524034 178987 524068
rect 179045 524034 179079 524068
rect 179137 524034 179171 524068
rect 179229 524034 179263 524068
rect 179321 524034 179355 524068
rect 179413 524034 179447 524068
rect 179505 524034 179539 524068
rect 179597 524034 179631 524068
rect 179689 524034 179723 524068
rect 179781 524034 179815 524068
rect 179873 524034 179907 524068
rect 179965 524034 179999 524068
rect 180057 524034 180091 524068
rect 180149 524034 180183 524068
rect 180241 524034 180275 524068
rect 180333 524034 180367 524068
rect 180425 524034 180459 524068
rect 180517 524034 180551 524068
rect 180609 524034 180643 524068
rect 180701 524034 180735 524068
rect 180793 524034 180827 524068
rect 180885 524034 180919 524068
rect 180977 524034 181011 524068
rect 181069 524034 181103 524068
rect 181161 524034 181195 524068
rect 181253 524034 181287 524068
rect 181345 524034 181379 524068
rect 181437 524034 181471 524068
rect 181529 524034 181563 524068
rect 181621 524034 181655 524068
rect 181713 524034 181747 524068
rect 181805 524034 181839 524068
rect 181897 524034 181931 524068
rect 181989 524034 182023 524068
rect 182081 524034 182115 524068
rect 182173 524034 182207 524068
rect 182265 524034 182299 524068
rect 182357 524034 182391 524068
rect 182449 524034 182483 524068
rect 182541 524034 182575 524068
rect 182633 524034 182667 524068
rect 182725 524034 182759 524068
rect 182817 524034 182851 524068
rect 182909 524034 182943 524068
rect 183001 524034 183035 524068
rect 183093 524034 183127 524068
rect 183185 524034 183219 524068
rect 183277 524034 183311 524068
rect 183369 524034 183403 524068
rect 183461 524034 183495 524068
rect 183553 524034 183587 524068
rect 183645 524034 183679 524068
rect 183737 524034 183771 524068
rect 183829 524034 183863 524068
rect 183921 524034 183955 524068
rect 184013 524034 184047 524068
rect 184105 524034 184139 524068
rect 184197 524034 184231 524068
rect 184289 524034 184323 524068
rect 184381 524034 184415 524068
rect 184473 524034 184507 524068
rect 184565 524034 184599 524068
rect 184657 524034 184691 524068
rect 184749 524034 184783 524068
rect 184841 524034 184875 524068
rect 184933 524034 184967 524068
rect 185025 524034 185059 524068
rect 185117 524034 185151 524068
rect 185209 524034 185243 524068
rect 185301 524034 185335 524068
rect 185393 524034 185427 524068
rect 185485 524034 185519 524068
rect 185577 524034 185611 524068
rect 185669 524034 185703 524068
rect 185761 524034 185795 524068
rect 185853 524034 185887 524068
rect 185945 524034 185979 524068
rect 186037 524034 186071 524068
rect 186129 524034 186163 524068
rect 186221 524034 186255 524068
rect 186313 524034 186347 524068
rect 186405 524034 186439 524068
rect 186497 524034 186531 524068
rect 186589 524034 186623 524068
rect 186681 524034 186715 524068
rect 186773 524034 186807 524068
rect 186865 524034 186899 524068
rect 186957 524034 186991 524068
rect 187049 524034 187083 524068
rect 187141 524034 187175 524068
rect 187233 524034 187267 524068
rect 187325 524034 187359 524068
rect 187417 524034 187451 524068
rect 172237 523490 172271 523524
rect 172329 523490 172363 523524
rect 172421 523490 172455 523524
rect 172513 523490 172547 523524
rect 172605 523490 172639 523524
rect 172697 523490 172731 523524
rect 172789 523490 172823 523524
rect 172881 523490 172915 523524
rect 172973 523490 173007 523524
rect 173065 523490 173099 523524
rect 173157 523490 173191 523524
rect 173249 523490 173283 523524
rect 173341 523490 173375 523524
rect 173433 523490 173467 523524
rect 173525 523490 173559 523524
rect 173617 523490 173651 523524
rect 173709 523490 173743 523524
rect 173801 523490 173835 523524
rect 173893 523490 173927 523524
rect 173985 523490 174019 523524
rect 174077 523490 174111 523524
rect 174169 523490 174203 523524
rect 174261 523490 174295 523524
rect 174353 523490 174387 523524
rect 174445 523490 174479 523524
rect 174537 523490 174571 523524
rect 174629 523490 174663 523524
rect 174721 523490 174755 523524
rect 174813 523490 174847 523524
rect 174905 523490 174939 523524
rect 174997 523490 175031 523524
rect 175089 523490 175123 523524
rect 175181 523490 175215 523524
rect 175273 523490 175307 523524
rect 175365 523490 175399 523524
rect 175457 523490 175491 523524
rect 175549 523490 175583 523524
rect 175641 523490 175675 523524
rect 175733 523490 175767 523524
rect 175825 523490 175859 523524
rect 175917 523490 175951 523524
rect 176009 523490 176043 523524
rect 176101 523490 176135 523524
rect 176193 523490 176227 523524
rect 176285 523490 176319 523524
rect 176377 523490 176411 523524
rect 176469 523490 176503 523524
rect 176561 523490 176595 523524
rect 176653 523490 176687 523524
rect 176745 523490 176779 523524
rect 176837 523490 176871 523524
rect 176929 523490 176963 523524
rect 177021 523490 177055 523524
rect 177113 523490 177147 523524
rect 177205 523490 177239 523524
rect 177297 523490 177331 523524
rect 177389 523490 177423 523524
rect 177481 523490 177515 523524
rect 177573 523490 177607 523524
rect 177665 523490 177699 523524
rect 177757 523490 177791 523524
rect 177849 523490 177883 523524
rect 177941 523490 177975 523524
rect 178033 523490 178067 523524
rect 178125 523490 178159 523524
rect 178217 523490 178251 523524
rect 178309 523490 178343 523524
rect 178401 523490 178435 523524
rect 178493 523490 178527 523524
rect 178585 523490 178619 523524
rect 178677 523490 178711 523524
rect 178769 523490 178803 523524
rect 178861 523490 178895 523524
rect 178953 523490 178987 523524
rect 179045 523490 179079 523524
rect 179137 523490 179171 523524
rect 179229 523490 179263 523524
rect 179321 523490 179355 523524
rect 179413 523490 179447 523524
rect 179505 523490 179539 523524
rect 179597 523490 179631 523524
rect 179689 523490 179723 523524
rect 179781 523490 179815 523524
rect 179873 523490 179907 523524
rect 179965 523490 179999 523524
rect 180057 523490 180091 523524
rect 180149 523490 180183 523524
rect 180241 523490 180275 523524
rect 180333 523490 180367 523524
rect 180425 523490 180459 523524
rect 180517 523490 180551 523524
rect 180609 523490 180643 523524
rect 180701 523490 180735 523524
rect 180793 523490 180827 523524
rect 180885 523490 180919 523524
rect 180977 523490 181011 523524
rect 181069 523490 181103 523524
rect 181161 523490 181195 523524
rect 181253 523490 181287 523524
rect 181345 523490 181379 523524
rect 181437 523490 181471 523524
rect 181529 523490 181563 523524
rect 181621 523490 181655 523524
rect 181713 523490 181747 523524
rect 181805 523490 181839 523524
rect 181897 523490 181931 523524
rect 181989 523490 182023 523524
rect 182081 523490 182115 523524
rect 182173 523490 182207 523524
rect 182265 523490 182299 523524
rect 182357 523490 182391 523524
rect 182449 523490 182483 523524
rect 182541 523490 182575 523524
rect 182633 523490 182667 523524
rect 182725 523490 182759 523524
rect 182817 523490 182851 523524
rect 182909 523490 182943 523524
rect 183001 523490 183035 523524
rect 183093 523490 183127 523524
rect 183185 523490 183219 523524
rect 183277 523490 183311 523524
rect 183369 523490 183403 523524
rect 183461 523490 183495 523524
rect 183553 523490 183587 523524
rect 183645 523490 183679 523524
rect 183737 523490 183771 523524
rect 183829 523490 183863 523524
rect 183921 523490 183955 523524
rect 184013 523490 184047 523524
rect 184105 523490 184139 523524
rect 184197 523490 184231 523524
rect 184289 523490 184323 523524
rect 184381 523490 184415 523524
rect 184473 523490 184507 523524
rect 184565 523490 184599 523524
rect 184657 523490 184691 523524
rect 184749 523490 184783 523524
rect 184841 523490 184875 523524
rect 184933 523490 184967 523524
rect 185025 523490 185059 523524
rect 185117 523490 185151 523524
rect 185209 523490 185243 523524
rect 185301 523490 185335 523524
rect 185393 523490 185427 523524
rect 185485 523490 185519 523524
rect 185577 523490 185611 523524
rect 185669 523490 185703 523524
rect 185761 523490 185795 523524
rect 185853 523490 185887 523524
rect 185945 523490 185979 523524
rect 186037 523490 186071 523524
rect 186129 523490 186163 523524
rect 186221 523490 186255 523524
rect 186313 523490 186347 523524
rect 186405 523490 186439 523524
rect 186497 523490 186531 523524
rect 186589 523490 186623 523524
rect 186681 523490 186715 523524
rect 186773 523490 186807 523524
rect 186865 523490 186899 523524
rect 186957 523490 186991 523524
rect 187049 523490 187083 523524
rect 187141 523490 187175 523524
rect 187233 523490 187267 523524
rect 187325 523490 187359 523524
rect 187417 523490 187451 523524
rect 172237 522946 172271 522980
rect 172329 522946 172363 522980
rect 172421 522946 172455 522980
rect 172513 522946 172547 522980
rect 172605 522946 172639 522980
rect 172697 522946 172731 522980
rect 172789 522946 172823 522980
rect 172881 522946 172915 522980
rect 172973 522946 173007 522980
rect 173065 522946 173099 522980
rect 173157 522946 173191 522980
rect 173249 522946 173283 522980
rect 173341 522946 173375 522980
rect 173433 522946 173467 522980
rect 173525 522946 173559 522980
rect 173617 522946 173651 522980
rect 173709 522946 173743 522980
rect 173801 522946 173835 522980
rect 173893 522946 173927 522980
rect 173985 522946 174019 522980
rect 174077 522946 174111 522980
rect 174169 522946 174203 522980
rect 174261 522946 174295 522980
rect 174353 522946 174387 522980
rect 174445 522946 174479 522980
rect 174537 522946 174571 522980
rect 174629 522946 174663 522980
rect 174721 522946 174755 522980
rect 174813 522946 174847 522980
rect 174905 522946 174939 522980
rect 174997 522946 175031 522980
rect 175089 522946 175123 522980
rect 175181 522946 175215 522980
rect 175273 522946 175307 522980
rect 175365 522946 175399 522980
rect 175457 522946 175491 522980
rect 175549 522946 175583 522980
rect 175641 522946 175675 522980
rect 175733 522946 175767 522980
rect 175825 522946 175859 522980
rect 175917 522946 175951 522980
rect 176009 522946 176043 522980
rect 176101 522946 176135 522980
rect 176193 522946 176227 522980
rect 176285 522946 176319 522980
rect 176377 522946 176411 522980
rect 176469 522946 176503 522980
rect 176561 522946 176595 522980
rect 176653 522946 176687 522980
rect 176745 522946 176779 522980
rect 176837 522946 176871 522980
rect 176929 522946 176963 522980
rect 177021 522946 177055 522980
rect 177113 522946 177147 522980
rect 177205 522946 177239 522980
rect 177297 522946 177331 522980
rect 177389 522946 177423 522980
rect 177481 522946 177515 522980
rect 177573 522946 177607 522980
rect 177665 522946 177699 522980
rect 177757 522946 177791 522980
rect 177849 522946 177883 522980
rect 177941 522946 177975 522980
rect 178033 522946 178067 522980
rect 178125 522946 178159 522980
rect 178217 522946 178251 522980
rect 178309 522946 178343 522980
rect 178401 522946 178435 522980
rect 178493 522946 178527 522980
rect 178585 522946 178619 522980
rect 178677 522946 178711 522980
rect 178769 522946 178803 522980
rect 178861 522946 178895 522980
rect 178953 522946 178987 522980
rect 179045 522946 179079 522980
rect 179137 522946 179171 522980
rect 179229 522946 179263 522980
rect 179321 522946 179355 522980
rect 179413 522946 179447 522980
rect 179505 522946 179539 522980
rect 179597 522946 179631 522980
rect 179689 522946 179723 522980
rect 179781 522946 179815 522980
rect 179873 522946 179907 522980
rect 179965 522946 179999 522980
rect 180057 522946 180091 522980
rect 180149 522946 180183 522980
rect 180241 522946 180275 522980
rect 180333 522946 180367 522980
rect 180425 522946 180459 522980
rect 180517 522946 180551 522980
rect 180609 522946 180643 522980
rect 180701 522946 180735 522980
rect 180793 522946 180827 522980
rect 180885 522946 180919 522980
rect 180977 522946 181011 522980
rect 181069 522946 181103 522980
rect 181161 522946 181195 522980
rect 181253 522946 181287 522980
rect 181345 522946 181379 522980
rect 181437 522946 181471 522980
rect 181529 522946 181563 522980
rect 181621 522946 181655 522980
rect 181713 522946 181747 522980
rect 181805 522946 181839 522980
rect 181897 522946 181931 522980
rect 181989 522946 182023 522980
rect 182081 522946 182115 522980
rect 182173 522946 182207 522980
rect 182265 522946 182299 522980
rect 182357 522946 182391 522980
rect 182449 522946 182483 522980
rect 182541 522946 182575 522980
rect 182633 522946 182667 522980
rect 182725 522946 182759 522980
rect 182817 522946 182851 522980
rect 182909 522946 182943 522980
rect 183001 522946 183035 522980
rect 183093 522946 183127 522980
rect 183185 522946 183219 522980
rect 183277 522946 183311 522980
rect 183369 522946 183403 522980
rect 183461 522946 183495 522980
rect 183553 522946 183587 522980
rect 183645 522946 183679 522980
rect 183737 522946 183771 522980
rect 183829 522946 183863 522980
rect 183921 522946 183955 522980
rect 184013 522946 184047 522980
rect 184105 522946 184139 522980
rect 184197 522946 184231 522980
rect 184289 522946 184323 522980
rect 184381 522946 184415 522980
rect 184473 522946 184507 522980
rect 184565 522946 184599 522980
rect 184657 522946 184691 522980
rect 184749 522946 184783 522980
rect 184841 522946 184875 522980
rect 184933 522946 184967 522980
rect 185025 522946 185059 522980
rect 185117 522946 185151 522980
rect 185209 522946 185243 522980
rect 185301 522946 185335 522980
rect 185393 522946 185427 522980
rect 185485 522946 185519 522980
rect 185577 522946 185611 522980
rect 185669 522946 185703 522980
rect 185761 522946 185795 522980
rect 185853 522946 185887 522980
rect 185945 522946 185979 522980
rect 186037 522946 186071 522980
rect 186129 522946 186163 522980
rect 186221 522946 186255 522980
rect 186313 522946 186347 522980
rect 186405 522946 186439 522980
rect 186497 522946 186531 522980
rect 186589 522946 186623 522980
rect 186681 522946 186715 522980
rect 186773 522946 186807 522980
rect 186865 522946 186899 522980
rect 186957 522946 186991 522980
rect 187049 522946 187083 522980
rect 187141 522946 187175 522980
rect 187233 522946 187267 522980
rect 187325 522946 187359 522980
rect 187417 522946 187451 522980
rect 172237 522402 172271 522436
rect 172329 522402 172363 522436
rect 172421 522402 172455 522436
rect 172513 522402 172547 522436
rect 172605 522402 172639 522436
rect 172697 522402 172731 522436
rect 172789 522402 172823 522436
rect 172881 522402 172915 522436
rect 172973 522402 173007 522436
rect 173065 522402 173099 522436
rect 173157 522402 173191 522436
rect 173249 522402 173283 522436
rect 173341 522402 173375 522436
rect 173433 522402 173467 522436
rect 173525 522402 173559 522436
rect 173617 522402 173651 522436
rect 173709 522402 173743 522436
rect 173801 522402 173835 522436
rect 173893 522402 173927 522436
rect 173985 522402 174019 522436
rect 174077 522402 174111 522436
rect 174169 522402 174203 522436
rect 174261 522402 174295 522436
rect 174353 522402 174387 522436
rect 174445 522402 174479 522436
rect 174537 522402 174571 522436
rect 174629 522402 174663 522436
rect 174721 522402 174755 522436
rect 174813 522402 174847 522436
rect 174905 522402 174939 522436
rect 174997 522402 175031 522436
rect 175089 522402 175123 522436
rect 175181 522402 175215 522436
rect 175273 522402 175307 522436
rect 175365 522402 175399 522436
rect 175457 522402 175491 522436
rect 175549 522402 175583 522436
rect 175641 522402 175675 522436
rect 175733 522402 175767 522436
rect 175825 522402 175859 522436
rect 175917 522402 175951 522436
rect 176009 522402 176043 522436
rect 176101 522402 176135 522436
rect 176193 522402 176227 522436
rect 176285 522402 176319 522436
rect 176377 522402 176411 522436
rect 176469 522402 176503 522436
rect 176561 522402 176595 522436
rect 176653 522402 176687 522436
rect 176745 522402 176779 522436
rect 176837 522402 176871 522436
rect 176929 522402 176963 522436
rect 177021 522402 177055 522436
rect 177113 522402 177147 522436
rect 177205 522402 177239 522436
rect 177297 522402 177331 522436
rect 177389 522402 177423 522436
rect 177481 522402 177515 522436
rect 177573 522402 177607 522436
rect 177665 522402 177699 522436
rect 177757 522402 177791 522436
rect 177849 522402 177883 522436
rect 177941 522402 177975 522436
rect 178033 522402 178067 522436
rect 178125 522402 178159 522436
rect 178217 522402 178251 522436
rect 178309 522402 178343 522436
rect 178401 522402 178435 522436
rect 178493 522402 178527 522436
rect 178585 522402 178619 522436
rect 178677 522402 178711 522436
rect 178769 522402 178803 522436
rect 178861 522402 178895 522436
rect 178953 522402 178987 522436
rect 179045 522402 179079 522436
rect 179137 522402 179171 522436
rect 179229 522402 179263 522436
rect 179321 522402 179355 522436
rect 179413 522402 179447 522436
rect 179505 522402 179539 522436
rect 179597 522402 179631 522436
rect 179689 522402 179723 522436
rect 179781 522402 179815 522436
rect 179873 522402 179907 522436
rect 179965 522402 179999 522436
rect 180057 522402 180091 522436
rect 180149 522402 180183 522436
rect 180241 522402 180275 522436
rect 180333 522402 180367 522436
rect 180425 522402 180459 522436
rect 180517 522402 180551 522436
rect 180609 522402 180643 522436
rect 180701 522402 180735 522436
rect 180793 522402 180827 522436
rect 180885 522402 180919 522436
rect 180977 522402 181011 522436
rect 181069 522402 181103 522436
rect 181161 522402 181195 522436
rect 181253 522402 181287 522436
rect 181345 522402 181379 522436
rect 181437 522402 181471 522436
rect 181529 522402 181563 522436
rect 181621 522402 181655 522436
rect 181713 522402 181747 522436
rect 181805 522402 181839 522436
rect 181897 522402 181931 522436
rect 181989 522402 182023 522436
rect 182081 522402 182115 522436
rect 182173 522402 182207 522436
rect 182265 522402 182299 522436
rect 182357 522402 182391 522436
rect 182449 522402 182483 522436
rect 182541 522402 182575 522436
rect 182633 522402 182667 522436
rect 182725 522402 182759 522436
rect 182817 522402 182851 522436
rect 182909 522402 182943 522436
rect 183001 522402 183035 522436
rect 183093 522402 183127 522436
rect 183185 522402 183219 522436
rect 183277 522402 183311 522436
rect 183369 522402 183403 522436
rect 183461 522402 183495 522436
rect 183553 522402 183587 522436
rect 183645 522402 183679 522436
rect 183737 522402 183771 522436
rect 183829 522402 183863 522436
rect 183921 522402 183955 522436
rect 184013 522402 184047 522436
rect 184105 522402 184139 522436
rect 184197 522402 184231 522436
rect 184289 522402 184323 522436
rect 184381 522402 184415 522436
rect 184473 522402 184507 522436
rect 184565 522402 184599 522436
rect 184657 522402 184691 522436
rect 184749 522402 184783 522436
rect 184841 522402 184875 522436
rect 184933 522402 184967 522436
rect 185025 522402 185059 522436
rect 185117 522402 185151 522436
rect 185209 522402 185243 522436
rect 185301 522402 185335 522436
rect 185393 522402 185427 522436
rect 185485 522402 185519 522436
rect 185577 522402 185611 522436
rect 185669 522402 185703 522436
rect 185761 522402 185795 522436
rect 185853 522402 185887 522436
rect 185945 522402 185979 522436
rect 186037 522402 186071 522436
rect 186129 522402 186163 522436
rect 186221 522402 186255 522436
rect 186313 522402 186347 522436
rect 186405 522402 186439 522436
rect 186497 522402 186531 522436
rect 186589 522402 186623 522436
rect 186681 522402 186715 522436
rect 186773 522402 186807 522436
rect 186865 522402 186899 522436
rect 186957 522402 186991 522436
rect 187049 522402 187083 522436
rect 187141 522402 187175 522436
rect 187233 522402 187267 522436
rect 187325 522402 187359 522436
rect 187417 522402 187451 522436
rect 172237 521858 172271 521892
rect 172329 521858 172363 521892
rect 172421 521858 172455 521892
rect 172513 521858 172547 521892
rect 172605 521858 172639 521892
rect 172697 521858 172731 521892
rect 172789 521858 172823 521892
rect 172881 521858 172915 521892
rect 172973 521858 173007 521892
rect 173065 521858 173099 521892
rect 173157 521858 173191 521892
rect 173249 521858 173283 521892
rect 173341 521858 173375 521892
rect 173433 521858 173467 521892
rect 173525 521858 173559 521892
rect 173617 521858 173651 521892
rect 173709 521858 173743 521892
rect 173801 521858 173835 521892
rect 173893 521858 173927 521892
rect 173985 521858 174019 521892
rect 174077 521858 174111 521892
rect 174169 521858 174203 521892
rect 174261 521858 174295 521892
rect 174353 521858 174387 521892
rect 174445 521858 174479 521892
rect 174537 521858 174571 521892
rect 174629 521858 174663 521892
rect 174721 521858 174755 521892
rect 174813 521858 174847 521892
rect 174905 521858 174939 521892
rect 174997 521858 175031 521892
rect 175089 521858 175123 521892
rect 175181 521858 175215 521892
rect 175273 521858 175307 521892
rect 175365 521858 175399 521892
rect 175457 521858 175491 521892
rect 175549 521858 175583 521892
rect 175641 521858 175675 521892
rect 175733 521858 175767 521892
rect 175825 521858 175859 521892
rect 175917 521858 175951 521892
rect 176009 521858 176043 521892
rect 176101 521858 176135 521892
rect 176193 521858 176227 521892
rect 176285 521858 176319 521892
rect 176377 521858 176411 521892
rect 176469 521858 176503 521892
rect 176561 521858 176595 521892
rect 176653 521858 176687 521892
rect 176745 521858 176779 521892
rect 176837 521858 176871 521892
rect 176929 521858 176963 521892
rect 177021 521858 177055 521892
rect 177113 521858 177147 521892
rect 177205 521858 177239 521892
rect 177297 521858 177331 521892
rect 177389 521858 177423 521892
rect 177481 521858 177515 521892
rect 177573 521858 177607 521892
rect 177665 521858 177699 521892
rect 177757 521858 177791 521892
rect 177849 521858 177883 521892
rect 177941 521858 177975 521892
rect 178033 521858 178067 521892
rect 178125 521858 178159 521892
rect 178217 521858 178251 521892
rect 178309 521858 178343 521892
rect 178401 521858 178435 521892
rect 178493 521858 178527 521892
rect 178585 521858 178619 521892
rect 178677 521858 178711 521892
rect 178769 521858 178803 521892
rect 178861 521858 178895 521892
rect 178953 521858 178987 521892
rect 179045 521858 179079 521892
rect 179137 521858 179171 521892
rect 179229 521858 179263 521892
rect 179321 521858 179355 521892
rect 179413 521858 179447 521892
rect 179505 521858 179539 521892
rect 179597 521858 179631 521892
rect 179689 521858 179723 521892
rect 179781 521858 179815 521892
rect 179873 521858 179907 521892
rect 179965 521858 179999 521892
rect 180057 521858 180091 521892
rect 180149 521858 180183 521892
rect 180241 521858 180275 521892
rect 180333 521858 180367 521892
rect 180425 521858 180459 521892
rect 180517 521858 180551 521892
rect 180609 521858 180643 521892
rect 180701 521858 180735 521892
rect 180793 521858 180827 521892
rect 180885 521858 180919 521892
rect 180977 521858 181011 521892
rect 181069 521858 181103 521892
rect 181161 521858 181195 521892
rect 181253 521858 181287 521892
rect 181345 521858 181379 521892
rect 181437 521858 181471 521892
rect 181529 521858 181563 521892
rect 181621 521858 181655 521892
rect 181713 521858 181747 521892
rect 181805 521858 181839 521892
rect 181897 521858 181931 521892
rect 181989 521858 182023 521892
rect 182081 521858 182115 521892
rect 182173 521858 182207 521892
rect 182265 521858 182299 521892
rect 182357 521858 182391 521892
rect 182449 521858 182483 521892
rect 182541 521858 182575 521892
rect 182633 521858 182667 521892
rect 182725 521858 182759 521892
rect 182817 521858 182851 521892
rect 182909 521858 182943 521892
rect 183001 521858 183035 521892
rect 183093 521858 183127 521892
rect 183185 521858 183219 521892
rect 183277 521858 183311 521892
rect 183369 521858 183403 521892
rect 183461 521858 183495 521892
rect 183553 521858 183587 521892
rect 183645 521858 183679 521892
rect 183737 521858 183771 521892
rect 183829 521858 183863 521892
rect 183921 521858 183955 521892
rect 184013 521858 184047 521892
rect 184105 521858 184139 521892
rect 184197 521858 184231 521892
rect 184289 521858 184323 521892
rect 184381 521858 184415 521892
rect 184473 521858 184507 521892
rect 184565 521858 184599 521892
rect 184657 521858 184691 521892
rect 184749 521858 184783 521892
rect 184841 521858 184875 521892
rect 184933 521858 184967 521892
rect 185025 521858 185059 521892
rect 185117 521858 185151 521892
rect 185209 521858 185243 521892
rect 185301 521858 185335 521892
rect 185393 521858 185427 521892
rect 185485 521858 185519 521892
rect 185577 521858 185611 521892
rect 185669 521858 185703 521892
rect 185761 521858 185795 521892
rect 185853 521858 185887 521892
rect 185945 521858 185979 521892
rect 186037 521858 186071 521892
rect 186129 521858 186163 521892
rect 186221 521858 186255 521892
rect 186313 521858 186347 521892
rect 186405 521858 186439 521892
rect 186497 521858 186531 521892
rect 186589 521858 186623 521892
rect 186681 521858 186715 521892
rect 186773 521858 186807 521892
rect 186865 521858 186899 521892
rect 186957 521858 186991 521892
rect 187049 521858 187083 521892
rect 187141 521858 187175 521892
rect 187233 521858 187267 521892
rect 187325 521858 187359 521892
rect 187417 521858 187451 521892
rect 172237 521314 172271 521348
rect 172329 521314 172363 521348
rect 172421 521314 172455 521348
rect 172513 521314 172547 521348
rect 172605 521314 172639 521348
rect 172697 521314 172731 521348
rect 172789 521314 172823 521348
rect 172881 521314 172915 521348
rect 172973 521314 173007 521348
rect 173065 521314 173099 521348
rect 173157 521314 173191 521348
rect 173249 521314 173283 521348
rect 173341 521314 173375 521348
rect 173433 521314 173467 521348
rect 173525 521314 173559 521348
rect 173617 521314 173651 521348
rect 173709 521314 173743 521348
rect 173801 521314 173835 521348
rect 173893 521314 173927 521348
rect 173985 521314 174019 521348
rect 174077 521314 174111 521348
rect 174169 521314 174203 521348
rect 174261 521314 174295 521348
rect 174353 521314 174387 521348
rect 174445 521314 174479 521348
rect 174537 521314 174571 521348
rect 174629 521314 174663 521348
rect 174721 521314 174755 521348
rect 174813 521314 174847 521348
rect 174905 521314 174939 521348
rect 174997 521314 175031 521348
rect 175089 521314 175123 521348
rect 175181 521314 175215 521348
rect 175273 521314 175307 521348
rect 175365 521314 175399 521348
rect 175457 521314 175491 521348
rect 175549 521314 175583 521348
rect 175641 521314 175675 521348
rect 175733 521314 175767 521348
rect 175825 521314 175859 521348
rect 175917 521314 175951 521348
rect 176009 521314 176043 521348
rect 176101 521314 176135 521348
rect 176193 521314 176227 521348
rect 176285 521314 176319 521348
rect 176377 521314 176411 521348
rect 176469 521314 176503 521348
rect 176561 521314 176595 521348
rect 176653 521314 176687 521348
rect 176745 521314 176779 521348
rect 176837 521314 176871 521348
rect 176929 521314 176963 521348
rect 177021 521314 177055 521348
rect 177113 521314 177147 521348
rect 177205 521314 177239 521348
rect 177297 521314 177331 521348
rect 177389 521314 177423 521348
rect 177481 521314 177515 521348
rect 177573 521314 177607 521348
rect 177665 521314 177699 521348
rect 177757 521314 177791 521348
rect 177849 521314 177883 521348
rect 177941 521314 177975 521348
rect 178033 521314 178067 521348
rect 178125 521314 178159 521348
rect 178217 521314 178251 521348
rect 178309 521314 178343 521348
rect 178401 521314 178435 521348
rect 178493 521314 178527 521348
rect 178585 521314 178619 521348
rect 178677 521314 178711 521348
rect 178769 521314 178803 521348
rect 178861 521314 178895 521348
rect 178953 521314 178987 521348
rect 179045 521314 179079 521348
rect 179137 521314 179171 521348
rect 179229 521314 179263 521348
rect 179321 521314 179355 521348
rect 179413 521314 179447 521348
rect 179505 521314 179539 521348
rect 179597 521314 179631 521348
rect 179689 521314 179723 521348
rect 179781 521314 179815 521348
rect 179873 521314 179907 521348
rect 179965 521314 179999 521348
rect 180057 521314 180091 521348
rect 180149 521314 180183 521348
rect 180241 521314 180275 521348
rect 180333 521314 180367 521348
rect 180425 521314 180459 521348
rect 180517 521314 180551 521348
rect 180609 521314 180643 521348
rect 180701 521314 180735 521348
rect 180793 521314 180827 521348
rect 180885 521314 180919 521348
rect 180977 521314 181011 521348
rect 181069 521314 181103 521348
rect 181161 521314 181195 521348
rect 181253 521314 181287 521348
rect 181345 521314 181379 521348
rect 181437 521314 181471 521348
rect 181529 521314 181563 521348
rect 181621 521314 181655 521348
rect 181713 521314 181747 521348
rect 181805 521314 181839 521348
rect 181897 521314 181931 521348
rect 181989 521314 182023 521348
rect 182081 521314 182115 521348
rect 182173 521314 182207 521348
rect 182265 521314 182299 521348
rect 182357 521314 182391 521348
rect 182449 521314 182483 521348
rect 182541 521314 182575 521348
rect 182633 521314 182667 521348
rect 182725 521314 182759 521348
rect 182817 521314 182851 521348
rect 182909 521314 182943 521348
rect 183001 521314 183035 521348
rect 183093 521314 183127 521348
rect 183185 521314 183219 521348
rect 183277 521314 183311 521348
rect 183369 521314 183403 521348
rect 183461 521314 183495 521348
rect 183553 521314 183587 521348
rect 183645 521314 183679 521348
rect 183737 521314 183771 521348
rect 183829 521314 183863 521348
rect 183921 521314 183955 521348
rect 184013 521314 184047 521348
rect 184105 521314 184139 521348
rect 184197 521314 184231 521348
rect 184289 521314 184323 521348
rect 184381 521314 184415 521348
rect 184473 521314 184507 521348
rect 184565 521314 184599 521348
rect 184657 521314 184691 521348
rect 184749 521314 184783 521348
rect 184841 521314 184875 521348
rect 184933 521314 184967 521348
rect 185025 521314 185059 521348
rect 185117 521314 185151 521348
rect 185209 521314 185243 521348
rect 185301 521314 185335 521348
rect 185393 521314 185427 521348
rect 185485 521314 185519 521348
rect 185577 521314 185611 521348
rect 185669 521314 185703 521348
rect 185761 521314 185795 521348
rect 185853 521314 185887 521348
rect 185945 521314 185979 521348
rect 186037 521314 186071 521348
rect 186129 521314 186163 521348
rect 186221 521314 186255 521348
rect 186313 521314 186347 521348
rect 186405 521314 186439 521348
rect 186497 521314 186531 521348
rect 186589 521314 186623 521348
rect 186681 521314 186715 521348
rect 186773 521314 186807 521348
rect 186865 521314 186899 521348
rect 186957 521314 186991 521348
rect 187049 521314 187083 521348
rect 187141 521314 187175 521348
rect 187233 521314 187267 521348
rect 187325 521314 187359 521348
rect 187417 521314 187451 521348
rect 172237 520770 172271 520804
rect 172329 520770 172363 520804
rect 172421 520770 172455 520804
rect 172513 520770 172547 520804
rect 172605 520770 172639 520804
rect 172697 520770 172731 520804
rect 172789 520770 172823 520804
rect 172881 520770 172915 520804
rect 172973 520770 173007 520804
rect 173065 520770 173099 520804
rect 173157 520770 173191 520804
rect 173249 520770 173283 520804
rect 173341 520770 173375 520804
rect 173433 520770 173467 520804
rect 173525 520770 173559 520804
rect 173617 520770 173651 520804
rect 173709 520770 173743 520804
rect 173801 520770 173835 520804
rect 173893 520770 173927 520804
rect 173985 520770 174019 520804
rect 174077 520770 174111 520804
rect 174169 520770 174203 520804
rect 174261 520770 174295 520804
rect 174353 520770 174387 520804
rect 174445 520770 174479 520804
rect 174537 520770 174571 520804
rect 174629 520770 174663 520804
rect 174721 520770 174755 520804
rect 174813 520770 174847 520804
rect 174905 520770 174939 520804
rect 174997 520770 175031 520804
rect 175089 520770 175123 520804
rect 175181 520770 175215 520804
rect 175273 520770 175307 520804
rect 175365 520770 175399 520804
rect 175457 520770 175491 520804
rect 175549 520770 175583 520804
rect 175641 520770 175675 520804
rect 175733 520770 175767 520804
rect 175825 520770 175859 520804
rect 175917 520770 175951 520804
rect 176009 520770 176043 520804
rect 176101 520770 176135 520804
rect 176193 520770 176227 520804
rect 176285 520770 176319 520804
rect 176377 520770 176411 520804
rect 176469 520770 176503 520804
rect 176561 520770 176595 520804
rect 176653 520770 176687 520804
rect 176745 520770 176779 520804
rect 176837 520770 176871 520804
rect 176929 520770 176963 520804
rect 177021 520770 177055 520804
rect 177113 520770 177147 520804
rect 177205 520770 177239 520804
rect 177297 520770 177331 520804
rect 177389 520770 177423 520804
rect 177481 520770 177515 520804
rect 177573 520770 177607 520804
rect 177665 520770 177699 520804
rect 177757 520770 177791 520804
rect 177849 520770 177883 520804
rect 177941 520770 177975 520804
rect 178033 520770 178067 520804
rect 178125 520770 178159 520804
rect 178217 520770 178251 520804
rect 178309 520770 178343 520804
rect 178401 520770 178435 520804
rect 178493 520770 178527 520804
rect 178585 520770 178619 520804
rect 178677 520770 178711 520804
rect 178769 520770 178803 520804
rect 178861 520770 178895 520804
rect 178953 520770 178987 520804
rect 179045 520770 179079 520804
rect 179137 520770 179171 520804
rect 179229 520770 179263 520804
rect 179321 520770 179355 520804
rect 179413 520770 179447 520804
rect 179505 520770 179539 520804
rect 179597 520770 179631 520804
rect 179689 520770 179723 520804
rect 179781 520770 179815 520804
rect 179873 520770 179907 520804
rect 179965 520770 179999 520804
rect 180057 520770 180091 520804
rect 180149 520770 180183 520804
rect 180241 520770 180275 520804
rect 180333 520770 180367 520804
rect 180425 520770 180459 520804
rect 180517 520770 180551 520804
rect 180609 520770 180643 520804
rect 180701 520770 180735 520804
rect 180793 520770 180827 520804
rect 180885 520770 180919 520804
rect 180977 520770 181011 520804
rect 181069 520770 181103 520804
rect 181161 520770 181195 520804
rect 181253 520770 181287 520804
rect 181345 520770 181379 520804
rect 181437 520770 181471 520804
rect 181529 520770 181563 520804
rect 181621 520770 181655 520804
rect 181713 520770 181747 520804
rect 181805 520770 181839 520804
rect 181897 520770 181931 520804
rect 181989 520770 182023 520804
rect 182081 520770 182115 520804
rect 182173 520770 182207 520804
rect 182265 520770 182299 520804
rect 182357 520770 182391 520804
rect 182449 520770 182483 520804
rect 182541 520770 182575 520804
rect 182633 520770 182667 520804
rect 182725 520770 182759 520804
rect 182817 520770 182851 520804
rect 182909 520770 182943 520804
rect 183001 520770 183035 520804
rect 183093 520770 183127 520804
rect 183185 520770 183219 520804
rect 183277 520770 183311 520804
rect 183369 520770 183403 520804
rect 183461 520770 183495 520804
rect 183553 520770 183587 520804
rect 183645 520770 183679 520804
rect 183737 520770 183771 520804
rect 183829 520770 183863 520804
rect 183921 520770 183955 520804
rect 184013 520770 184047 520804
rect 184105 520770 184139 520804
rect 184197 520770 184231 520804
rect 184289 520770 184323 520804
rect 184381 520770 184415 520804
rect 184473 520770 184507 520804
rect 184565 520770 184599 520804
rect 184657 520770 184691 520804
rect 184749 520770 184783 520804
rect 184841 520770 184875 520804
rect 184933 520770 184967 520804
rect 185025 520770 185059 520804
rect 185117 520770 185151 520804
rect 185209 520770 185243 520804
rect 185301 520770 185335 520804
rect 185393 520770 185427 520804
rect 185485 520770 185519 520804
rect 185577 520770 185611 520804
rect 185669 520770 185703 520804
rect 185761 520770 185795 520804
rect 185853 520770 185887 520804
rect 185945 520770 185979 520804
rect 186037 520770 186071 520804
rect 186129 520770 186163 520804
rect 186221 520770 186255 520804
rect 186313 520770 186347 520804
rect 186405 520770 186439 520804
rect 186497 520770 186531 520804
rect 186589 520770 186623 520804
rect 186681 520770 186715 520804
rect 186773 520770 186807 520804
rect 186865 520770 186899 520804
rect 186957 520770 186991 520804
rect 187049 520770 187083 520804
rect 187141 520770 187175 520804
rect 187233 520770 187267 520804
rect 187325 520770 187359 520804
rect 187417 520770 187451 520804
rect 172237 520226 172271 520260
rect 172329 520226 172363 520260
rect 172421 520226 172455 520260
rect 172513 520226 172547 520260
rect 172605 520226 172639 520260
rect 172697 520226 172731 520260
rect 172789 520226 172823 520260
rect 172881 520226 172915 520260
rect 172973 520226 173007 520260
rect 173065 520226 173099 520260
rect 173157 520226 173191 520260
rect 173249 520226 173283 520260
rect 173341 520226 173375 520260
rect 173433 520226 173467 520260
rect 173525 520226 173559 520260
rect 173617 520226 173651 520260
rect 173709 520226 173743 520260
rect 173801 520226 173835 520260
rect 173893 520226 173927 520260
rect 173985 520226 174019 520260
rect 174077 520226 174111 520260
rect 174169 520226 174203 520260
rect 174261 520226 174295 520260
rect 174353 520226 174387 520260
rect 174445 520226 174479 520260
rect 174537 520226 174571 520260
rect 174629 520226 174663 520260
rect 174721 520226 174755 520260
rect 174813 520226 174847 520260
rect 174905 520226 174939 520260
rect 174997 520226 175031 520260
rect 175089 520226 175123 520260
rect 175181 520226 175215 520260
rect 175273 520226 175307 520260
rect 175365 520226 175399 520260
rect 175457 520226 175491 520260
rect 175549 520226 175583 520260
rect 175641 520226 175675 520260
rect 175733 520226 175767 520260
rect 175825 520226 175859 520260
rect 175917 520226 175951 520260
rect 176009 520226 176043 520260
rect 176101 520226 176135 520260
rect 176193 520226 176227 520260
rect 176285 520226 176319 520260
rect 176377 520226 176411 520260
rect 176469 520226 176503 520260
rect 176561 520226 176595 520260
rect 176653 520226 176687 520260
rect 176745 520226 176779 520260
rect 176837 520226 176871 520260
rect 176929 520226 176963 520260
rect 177021 520226 177055 520260
rect 177113 520226 177147 520260
rect 177205 520226 177239 520260
rect 177297 520226 177331 520260
rect 177389 520226 177423 520260
rect 177481 520226 177515 520260
rect 177573 520226 177607 520260
rect 177665 520226 177699 520260
rect 177757 520226 177791 520260
rect 177849 520226 177883 520260
rect 177941 520226 177975 520260
rect 178033 520226 178067 520260
rect 178125 520226 178159 520260
rect 178217 520226 178251 520260
rect 178309 520226 178343 520260
rect 178401 520226 178435 520260
rect 178493 520226 178527 520260
rect 178585 520226 178619 520260
rect 178677 520226 178711 520260
rect 178769 520226 178803 520260
rect 178861 520226 178895 520260
rect 178953 520226 178987 520260
rect 179045 520226 179079 520260
rect 179137 520226 179171 520260
rect 179229 520226 179263 520260
rect 179321 520226 179355 520260
rect 179413 520226 179447 520260
rect 179505 520226 179539 520260
rect 179597 520226 179631 520260
rect 179689 520226 179723 520260
rect 179781 520226 179815 520260
rect 179873 520226 179907 520260
rect 179965 520226 179999 520260
rect 180057 520226 180091 520260
rect 180149 520226 180183 520260
rect 180241 520226 180275 520260
rect 180333 520226 180367 520260
rect 180425 520226 180459 520260
rect 180517 520226 180551 520260
rect 180609 520226 180643 520260
rect 180701 520226 180735 520260
rect 180793 520226 180827 520260
rect 180885 520226 180919 520260
rect 180977 520226 181011 520260
rect 181069 520226 181103 520260
rect 181161 520226 181195 520260
rect 181253 520226 181287 520260
rect 181345 520226 181379 520260
rect 181437 520226 181471 520260
rect 181529 520226 181563 520260
rect 181621 520226 181655 520260
rect 181713 520226 181747 520260
rect 181805 520226 181839 520260
rect 181897 520226 181931 520260
rect 181989 520226 182023 520260
rect 182081 520226 182115 520260
rect 182173 520226 182207 520260
rect 182265 520226 182299 520260
rect 182357 520226 182391 520260
rect 182449 520226 182483 520260
rect 182541 520226 182575 520260
rect 182633 520226 182667 520260
rect 182725 520226 182759 520260
rect 182817 520226 182851 520260
rect 182909 520226 182943 520260
rect 183001 520226 183035 520260
rect 183093 520226 183127 520260
rect 183185 520226 183219 520260
rect 183277 520226 183311 520260
rect 183369 520226 183403 520260
rect 183461 520226 183495 520260
rect 183553 520226 183587 520260
rect 183645 520226 183679 520260
rect 183737 520226 183771 520260
rect 183829 520226 183863 520260
rect 183921 520226 183955 520260
rect 184013 520226 184047 520260
rect 184105 520226 184139 520260
rect 184197 520226 184231 520260
rect 184289 520226 184323 520260
rect 184381 520226 184415 520260
rect 184473 520226 184507 520260
rect 184565 520226 184599 520260
rect 184657 520226 184691 520260
rect 184749 520226 184783 520260
rect 184841 520226 184875 520260
rect 184933 520226 184967 520260
rect 185025 520226 185059 520260
rect 185117 520226 185151 520260
rect 185209 520226 185243 520260
rect 185301 520226 185335 520260
rect 185393 520226 185427 520260
rect 185485 520226 185519 520260
rect 185577 520226 185611 520260
rect 185669 520226 185703 520260
rect 185761 520226 185795 520260
rect 185853 520226 185887 520260
rect 185945 520226 185979 520260
rect 186037 520226 186071 520260
rect 186129 520226 186163 520260
rect 186221 520226 186255 520260
rect 186313 520226 186347 520260
rect 186405 520226 186439 520260
rect 186497 520226 186531 520260
rect 186589 520226 186623 520260
rect 186681 520226 186715 520260
rect 186773 520226 186807 520260
rect 186865 520226 186899 520260
rect 186957 520226 186991 520260
rect 187049 520226 187083 520260
rect 187141 520226 187175 520260
rect 187233 520226 187267 520260
rect 187325 520226 187359 520260
rect 187417 520226 187451 520260
rect 172237 519682 172271 519716
rect 172329 519682 172363 519716
rect 172421 519682 172455 519716
rect 172513 519682 172547 519716
rect 172605 519682 172639 519716
rect 172697 519682 172731 519716
rect 172789 519682 172823 519716
rect 172881 519682 172915 519716
rect 172973 519682 173007 519716
rect 173065 519682 173099 519716
rect 173157 519682 173191 519716
rect 173249 519682 173283 519716
rect 173341 519682 173375 519716
rect 173433 519682 173467 519716
rect 173525 519682 173559 519716
rect 173617 519682 173651 519716
rect 173709 519682 173743 519716
rect 173801 519682 173835 519716
rect 173893 519682 173927 519716
rect 173985 519682 174019 519716
rect 174077 519682 174111 519716
rect 174169 519682 174203 519716
rect 174261 519682 174295 519716
rect 174353 519682 174387 519716
rect 174445 519682 174479 519716
rect 174537 519682 174571 519716
rect 174629 519682 174663 519716
rect 174721 519682 174755 519716
rect 174813 519682 174847 519716
rect 174905 519682 174939 519716
rect 174997 519682 175031 519716
rect 175089 519682 175123 519716
rect 175181 519682 175215 519716
rect 175273 519682 175307 519716
rect 175365 519682 175399 519716
rect 175457 519682 175491 519716
rect 175549 519682 175583 519716
rect 175641 519682 175675 519716
rect 175733 519682 175767 519716
rect 175825 519682 175859 519716
rect 175917 519682 175951 519716
rect 176009 519682 176043 519716
rect 176101 519682 176135 519716
rect 176193 519682 176227 519716
rect 176285 519682 176319 519716
rect 176377 519682 176411 519716
rect 176469 519682 176503 519716
rect 176561 519682 176595 519716
rect 176653 519682 176687 519716
rect 176745 519682 176779 519716
rect 176837 519682 176871 519716
rect 176929 519682 176963 519716
rect 177021 519682 177055 519716
rect 177113 519682 177147 519716
rect 177205 519682 177239 519716
rect 177297 519682 177331 519716
rect 177389 519682 177423 519716
rect 177481 519682 177515 519716
rect 177573 519682 177607 519716
rect 177665 519682 177699 519716
rect 177757 519682 177791 519716
rect 177849 519682 177883 519716
rect 177941 519682 177975 519716
rect 178033 519682 178067 519716
rect 178125 519682 178159 519716
rect 178217 519682 178251 519716
rect 178309 519682 178343 519716
rect 178401 519682 178435 519716
rect 178493 519682 178527 519716
rect 178585 519682 178619 519716
rect 178677 519682 178711 519716
rect 178769 519682 178803 519716
rect 178861 519682 178895 519716
rect 178953 519682 178987 519716
rect 179045 519682 179079 519716
rect 179137 519682 179171 519716
rect 179229 519682 179263 519716
rect 179321 519682 179355 519716
rect 179413 519682 179447 519716
rect 179505 519682 179539 519716
rect 179597 519682 179631 519716
rect 179689 519682 179723 519716
rect 179781 519682 179815 519716
rect 179873 519682 179907 519716
rect 179965 519682 179999 519716
rect 180057 519682 180091 519716
rect 180149 519682 180183 519716
rect 180241 519682 180275 519716
rect 180333 519682 180367 519716
rect 180425 519682 180459 519716
rect 180517 519682 180551 519716
rect 180609 519682 180643 519716
rect 180701 519682 180735 519716
rect 180793 519682 180827 519716
rect 180885 519682 180919 519716
rect 180977 519682 181011 519716
rect 181069 519682 181103 519716
rect 181161 519682 181195 519716
rect 181253 519682 181287 519716
rect 181345 519682 181379 519716
rect 181437 519682 181471 519716
rect 181529 519682 181563 519716
rect 181621 519682 181655 519716
rect 181713 519682 181747 519716
rect 181805 519682 181839 519716
rect 181897 519682 181931 519716
rect 181989 519682 182023 519716
rect 182081 519682 182115 519716
rect 182173 519682 182207 519716
rect 182265 519682 182299 519716
rect 182357 519682 182391 519716
rect 182449 519682 182483 519716
rect 182541 519682 182575 519716
rect 182633 519682 182667 519716
rect 182725 519682 182759 519716
rect 182817 519682 182851 519716
rect 182909 519682 182943 519716
rect 183001 519682 183035 519716
rect 183093 519682 183127 519716
rect 183185 519682 183219 519716
rect 183277 519682 183311 519716
rect 183369 519682 183403 519716
rect 183461 519682 183495 519716
rect 183553 519682 183587 519716
rect 183645 519682 183679 519716
rect 183737 519682 183771 519716
rect 183829 519682 183863 519716
rect 183921 519682 183955 519716
rect 184013 519682 184047 519716
rect 184105 519682 184139 519716
rect 184197 519682 184231 519716
rect 184289 519682 184323 519716
rect 184381 519682 184415 519716
rect 184473 519682 184507 519716
rect 184565 519682 184599 519716
rect 184657 519682 184691 519716
rect 184749 519682 184783 519716
rect 184841 519682 184875 519716
rect 184933 519682 184967 519716
rect 185025 519682 185059 519716
rect 185117 519682 185151 519716
rect 185209 519682 185243 519716
rect 185301 519682 185335 519716
rect 185393 519682 185427 519716
rect 185485 519682 185519 519716
rect 185577 519682 185611 519716
rect 185669 519682 185703 519716
rect 185761 519682 185795 519716
rect 185853 519682 185887 519716
rect 185945 519682 185979 519716
rect 186037 519682 186071 519716
rect 186129 519682 186163 519716
rect 186221 519682 186255 519716
rect 186313 519682 186347 519716
rect 186405 519682 186439 519716
rect 186497 519682 186531 519716
rect 186589 519682 186623 519716
rect 186681 519682 186715 519716
rect 186773 519682 186807 519716
rect 186865 519682 186899 519716
rect 186957 519682 186991 519716
rect 187049 519682 187083 519716
rect 187141 519682 187175 519716
rect 187233 519682 187267 519716
rect 187325 519682 187359 519716
rect 187417 519682 187451 519716
rect 172237 519138 172271 519172
rect 172329 519138 172363 519172
rect 172421 519138 172455 519172
rect 172513 519138 172547 519172
rect 172605 519138 172639 519172
rect 172697 519138 172731 519172
rect 172789 519138 172823 519172
rect 172881 519138 172915 519172
rect 172973 519138 173007 519172
rect 173065 519138 173099 519172
rect 173157 519138 173191 519172
rect 173249 519138 173283 519172
rect 173341 519138 173375 519172
rect 173433 519138 173467 519172
rect 173525 519138 173559 519172
rect 173617 519138 173651 519172
rect 173709 519138 173743 519172
rect 173801 519138 173835 519172
rect 173893 519138 173927 519172
rect 173985 519138 174019 519172
rect 174077 519138 174111 519172
rect 174169 519138 174203 519172
rect 174261 519138 174295 519172
rect 174353 519138 174387 519172
rect 174445 519138 174479 519172
rect 174537 519138 174571 519172
rect 174629 519138 174663 519172
rect 174721 519138 174755 519172
rect 174813 519138 174847 519172
rect 174905 519138 174939 519172
rect 174997 519138 175031 519172
rect 175089 519138 175123 519172
rect 175181 519138 175215 519172
rect 175273 519138 175307 519172
rect 175365 519138 175399 519172
rect 175457 519138 175491 519172
rect 175549 519138 175583 519172
rect 175641 519138 175675 519172
rect 175733 519138 175767 519172
rect 175825 519138 175859 519172
rect 175917 519138 175951 519172
rect 176009 519138 176043 519172
rect 176101 519138 176135 519172
rect 176193 519138 176227 519172
rect 176285 519138 176319 519172
rect 176377 519138 176411 519172
rect 176469 519138 176503 519172
rect 176561 519138 176595 519172
rect 176653 519138 176687 519172
rect 176745 519138 176779 519172
rect 176837 519138 176871 519172
rect 176929 519138 176963 519172
rect 177021 519138 177055 519172
rect 177113 519138 177147 519172
rect 177205 519138 177239 519172
rect 177297 519138 177331 519172
rect 177389 519138 177423 519172
rect 177481 519138 177515 519172
rect 177573 519138 177607 519172
rect 177665 519138 177699 519172
rect 177757 519138 177791 519172
rect 177849 519138 177883 519172
rect 177941 519138 177975 519172
rect 178033 519138 178067 519172
rect 178125 519138 178159 519172
rect 178217 519138 178251 519172
rect 178309 519138 178343 519172
rect 178401 519138 178435 519172
rect 178493 519138 178527 519172
rect 178585 519138 178619 519172
rect 178677 519138 178711 519172
rect 178769 519138 178803 519172
rect 178861 519138 178895 519172
rect 178953 519138 178987 519172
rect 179045 519138 179079 519172
rect 179137 519138 179171 519172
rect 179229 519138 179263 519172
rect 179321 519138 179355 519172
rect 179413 519138 179447 519172
rect 179505 519138 179539 519172
rect 179597 519138 179631 519172
rect 179689 519138 179723 519172
rect 179781 519138 179815 519172
rect 179873 519138 179907 519172
rect 179965 519138 179999 519172
rect 180057 519138 180091 519172
rect 180149 519138 180183 519172
rect 180241 519138 180275 519172
rect 180333 519138 180367 519172
rect 180425 519138 180459 519172
rect 180517 519138 180551 519172
rect 180609 519138 180643 519172
rect 180701 519138 180735 519172
rect 180793 519138 180827 519172
rect 180885 519138 180919 519172
rect 180977 519138 181011 519172
rect 181069 519138 181103 519172
rect 181161 519138 181195 519172
rect 181253 519138 181287 519172
rect 181345 519138 181379 519172
rect 181437 519138 181471 519172
rect 181529 519138 181563 519172
rect 181621 519138 181655 519172
rect 181713 519138 181747 519172
rect 181805 519138 181839 519172
rect 181897 519138 181931 519172
rect 181989 519138 182023 519172
rect 182081 519138 182115 519172
rect 182173 519138 182207 519172
rect 182265 519138 182299 519172
rect 182357 519138 182391 519172
rect 182449 519138 182483 519172
rect 182541 519138 182575 519172
rect 182633 519138 182667 519172
rect 182725 519138 182759 519172
rect 182817 519138 182851 519172
rect 182909 519138 182943 519172
rect 183001 519138 183035 519172
rect 183093 519138 183127 519172
rect 183185 519138 183219 519172
rect 183277 519138 183311 519172
rect 183369 519138 183403 519172
rect 183461 519138 183495 519172
rect 183553 519138 183587 519172
rect 183645 519138 183679 519172
rect 183737 519138 183771 519172
rect 183829 519138 183863 519172
rect 183921 519138 183955 519172
rect 184013 519138 184047 519172
rect 184105 519138 184139 519172
rect 184197 519138 184231 519172
rect 184289 519138 184323 519172
rect 184381 519138 184415 519172
rect 184473 519138 184507 519172
rect 184565 519138 184599 519172
rect 184657 519138 184691 519172
rect 184749 519138 184783 519172
rect 184841 519138 184875 519172
rect 184933 519138 184967 519172
rect 185025 519138 185059 519172
rect 185117 519138 185151 519172
rect 185209 519138 185243 519172
rect 185301 519138 185335 519172
rect 185393 519138 185427 519172
rect 185485 519138 185519 519172
rect 185577 519138 185611 519172
rect 185669 519138 185703 519172
rect 185761 519138 185795 519172
rect 185853 519138 185887 519172
rect 185945 519138 185979 519172
rect 186037 519138 186071 519172
rect 186129 519138 186163 519172
rect 186221 519138 186255 519172
rect 186313 519138 186347 519172
rect 186405 519138 186439 519172
rect 186497 519138 186531 519172
rect 186589 519138 186623 519172
rect 186681 519138 186715 519172
rect 186773 519138 186807 519172
rect 186865 519138 186899 519172
rect 186957 519138 186991 519172
rect 187049 519138 187083 519172
rect 187141 519138 187175 519172
rect 187233 519138 187267 519172
rect 187325 519138 187359 519172
rect 187417 519138 187451 519172
rect 172237 518594 172271 518628
rect 172329 518594 172363 518628
rect 172421 518594 172455 518628
rect 172513 518594 172547 518628
rect 172605 518594 172639 518628
rect 172697 518594 172731 518628
rect 172789 518594 172823 518628
rect 172881 518594 172915 518628
rect 172973 518594 173007 518628
rect 173065 518594 173099 518628
rect 173157 518594 173191 518628
rect 173249 518594 173283 518628
rect 173341 518594 173375 518628
rect 173433 518594 173467 518628
rect 173525 518594 173559 518628
rect 173617 518594 173651 518628
rect 173709 518594 173743 518628
rect 173801 518594 173835 518628
rect 173893 518594 173927 518628
rect 173985 518594 174019 518628
rect 174077 518594 174111 518628
rect 174169 518594 174203 518628
rect 174261 518594 174295 518628
rect 174353 518594 174387 518628
rect 174445 518594 174479 518628
rect 174537 518594 174571 518628
rect 174629 518594 174663 518628
rect 174721 518594 174755 518628
rect 174813 518594 174847 518628
rect 174905 518594 174939 518628
rect 174997 518594 175031 518628
rect 175089 518594 175123 518628
rect 175181 518594 175215 518628
rect 175273 518594 175307 518628
rect 175365 518594 175399 518628
rect 175457 518594 175491 518628
rect 175549 518594 175583 518628
rect 175641 518594 175675 518628
rect 175733 518594 175767 518628
rect 175825 518594 175859 518628
rect 175917 518594 175951 518628
rect 176009 518594 176043 518628
rect 176101 518594 176135 518628
rect 176193 518594 176227 518628
rect 176285 518594 176319 518628
rect 176377 518594 176411 518628
rect 176469 518594 176503 518628
rect 176561 518594 176595 518628
rect 176653 518594 176687 518628
rect 176745 518594 176779 518628
rect 176837 518594 176871 518628
rect 176929 518594 176963 518628
rect 177021 518594 177055 518628
rect 177113 518594 177147 518628
rect 177205 518594 177239 518628
rect 177297 518594 177331 518628
rect 177389 518594 177423 518628
rect 177481 518594 177515 518628
rect 177573 518594 177607 518628
rect 177665 518594 177699 518628
rect 177757 518594 177791 518628
rect 177849 518594 177883 518628
rect 177941 518594 177975 518628
rect 178033 518594 178067 518628
rect 178125 518594 178159 518628
rect 178217 518594 178251 518628
rect 178309 518594 178343 518628
rect 178401 518594 178435 518628
rect 178493 518594 178527 518628
rect 178585 518594 178619 518628
rect 178677 518594 178711 518628
rect 178769 518594 178803 518628
rect 178861 518594 178895 518628
rect 178953 518594 178987 518628
rect 179045 518594 179079 518628
rect 179137 518594 179171 518628
rect 179229 518594 179263 518628
rect 179321 518594 179355 518628
rect 179413 518594 179447 518628
rect 179505 518594 179539 518628
rect 179597 518594 179631 518628
rect 179689 518594 179723 518628
rect 179781 518594 179815 518628
rect 179873 518594 179907 518628
rect 179965 518594 179999 518628
rect 180057 518594 180091 518628
rect 180149 518594 180183 518628
rect 180241 518594 180275 518628
rect 180333 518594 180367 518628
rect 180425 518594 180459 518628
rect 180517 518594 180551 518628
rect 180609 518594 180643 518628
rect 180701 518594 180735 518628
rect 180793 518594 180827 518628
rect 180885 518594 180919 518628
rect 180977 518594 181011 518628
rect 181069 518594 181103 518628
rect 181161 518594 181195 518628
rect 181253 518594 181287 518628
rect 181345 518594 181379 518628
rect 181437 518594 181471 518628
rect 181529 518594 181563 518628
rect 181621 518594 181655 518628
rect 181713 518594 181747 518628
rect 181805 518594 181839 518628
rect 181897 518594 181931 518628
rect 181989 518594 182023 518628
rect 182081 518594 182115 518628
rect 182173 518594 182207 518628
rect 182265 518594 182299 518628
rect 182357 518594 182391 518628
rect 182449 518594 182483 518628
rect 182541 518594 182575 518628
rect 182633 518594 182667 518628
rect 182725 518594 182759 518628
rect 182817 518594 182851 518628
rect 182909 518594 182943 518628
rect 183001 518594 183035 518628
rect 183093 518594 183127 518628
rect 183185 518594 183219 518628
rect 183277 518594 183311 518628
rect 183369 518594 183403 518628
rect 183461 518594 183495 518628
rect 183553 518594 183587 518628
rect 183645 518594 183679 518628
rect 183737 518594 183771 518628
rect 183829 518594 183863 518628
rect 183921 518594 183955 518628
rect 184013 518594 184047 518628
rect 184105 518594 184139 518628
rect 184197 518594 184231 518628
rect 184289 518594 184323 518628
rect 184381 518594 184415 518628
rect 184473 518594 184507 518628
rect 184565 518594 184599 518628
rect 184657 518594 184691 518628
rect 184749 518594 184783 518628
rect 184841 518594 184875 518628
rect 184933 518594 184967 518628
rect 185025 518594 185059 518628
rect 185117 518594 185151 518628
rect 185209 518594 185243 518628
rect 185301 518594 185335 518628
rect 185393 518594 185427 518628
rect 185485 518594 185519 518628
rect 185577 518594 185611 518628
rect 185669 518594 185703 518628
rect 185761 518594 185795 518628
rect 185853 518594 185887 518628
rect 185945 518594 185979 518628
rect 186037 518594 186071 518628
rect 186129 518594 186163 518628
rect 186221 518594 186255 518628
rect 186313 518594 186347 518628
rect 186405 518594 186439 518628
rect 186497 518594 186531 518628
rect 186589 518594 186623 518628
rect 186681 518594 186715 518628
rect 186773 518594 186807 518628
rect 186865 518594 186899 518628
rect 186957 518594 186991 518628
rect 187049 518594 187083 518628
rect 187141 518594 187175 518628
rect 187233 518594 187267 518628
rect 187325 518594 187359 518628
rect 187417 518594 187451 518628
rect 172237 518050 172271 518084
rect 172329 518050 172363 518084
rect 172421 518050 172455 518084
rect 172513 518050 172547 518084
rect 172605 518050 172639 518084
rect 172697 518050 172731 518084
rect 172789 518050 172823 518084
rect 172881 518050 172915 518084
rect 172973 518050 173007 518084
rect 173065 518050 173099 518084
rect 173157 518050 173191 518084
rect 173249 518050 173283 518084
rect 173341 518050 173375 518084
rect 173433 518050 173467 518084
rect 173525 518050 173559 518084
rect 173617 518050 173651 518084
rect 173709 518050 173743 518084
rect 173801 518050 173835 518084
rect 173893 518050 173927 518084
rect 173985 518050 174019 518084
rect 174077 518050 174111 518084
rect 174169 518050 174203 518084
rect 174261 518050 174295 518084
rect 174353 518050 174387 518084
rect 174445 518050 174479 518084
rect 174537 518050 174571 518084
rect 174629 518050 174663 518084
rect 174721 518050 174755 518084
rect 174813 518050 174847 518084
rect 174905 518050 174939 518084
rect 174997 518050 175031 518084
rect 175089 518050 175123 518084
rect 175181 518050 175215 518084
rect 175273 518050 175307 518084
rect 175365 518050 175399 518084
rect 175457 518050 175491 518084
rect 175549 518050 175583 518084
rect 175641 518050 175675 518084
rect 175733 518050 175767 518084
rect 175825 518050 175859 518084
rect 175917 518050 175951 518084
rect 176009 518050 176043 518084
rect 176101 518050 176135 518084
rect 176193 518050 176227 518084
rect 176285 518050 176319 518084
rect 176377 518050 176411 518084
rect 176469 518050 176503 518084
rect 176561 518050 176595 518084
rect 176653 518050 176687 518084
rect 176745 518050 176779 518084
rect 176837 518050 176871 518084
rect 176929 518050 176963 518084
rect 177021 518050 177055 518084
rect 177113 518050 177147 518084
rect 177205 518050 177239 518084
rect 177297 518050 177331 518084
rect 177389 518050 177423 518084
rect 177481 518050 177515 518084
rect 177573 518050 177607 518084
rect 177665 518050 177699 518084
rect 177757 518050 177791 518084
rect 177849 518050 177883 518084
rect 177941 518050 177975 518084
rect 178033 518050 178067 518084
rect 178125 518050 178159 518084
rect 178217 518050 178251 518084
rect 178309 518050 178343 518084
rect 178401 518050 178435 518084
rect 178493 518050 178527 518084
rect 178585 518050 178619 518084
rect 178677 518050 178711 518084
rect 178769 518050 178803 518084
rect 178861 518050 178895 518084
rect 178953 518050 178987 518084
rect 179045 518050 179079 518084
rect 179137 518050 179171 518084
rect 179229 518050 179263 518084
rect 179321 518050 179355 518084
rect 179413 518050 179447 518084
rect 179505 518050 179539 518084
rect 179597 518050 179631 518084
rect 179689 518050 179723 518084
rect 179781 518050 179815 518084
rect 179873 518050 179907 518084
rect 179965 518050 179999 518084
rect 180057 518050 180091 518084
rect 180149 518050 180183 518084
rect 180241 518050 180275 518084
rect 180333 518050 180367 518084
rect 180425 518050 180459 518084
rect 180517 518050 180551 518084
rect 180609 518050 180643 518084
rect 180701 518050 180735 518084
rect 180793 518050 180827 518084
rect 180885 518050 180919 518084
rect 180977 518050 181011 518084
rect 181069 518050 181103 518084
rect 181161 518050 181195 518084
rect 181253 518050 181287 518084
rect 181345 518050 181379 518084
rect 181437 518050 181471 518084
rect 181529 518050 181563 518084
rect 181621 518050 181655 518084
rect 181713 518050 181747 518084
rect 181805 518050 181839 518084
rect 181897 518050 181931 518084
rect 181989 518050 182023 518084
rect 182081 518050 182115 518084
rect 182173 518050 182207 518084
rect 182265 518050 182299 518084
rect 182357 518050 182391 518084
rect 182449 518050 182483 518084
rect 182541 518050 182575 518084
rect 182633 518050 182667 518084
rect 182725 518050 182759 518084
rect 182817 518050 182851 518084
rect 182909 518050 182943 518084
rect 183001 518050 183035 518084
rect 183093 518050 183127 518084
rect 183185 518050 183219 518084
rect 183277 518050 183311 518084
rect 183369 518050 183403 518084
rect 183461 518050 183495 518084
rect 183553 518050 183587 518084
rect 183645 518050 183679 518084
rect 183737 518050 183771 518084
rect 183829 518050 183863 518084
rect 183921 518050 183955 518084
rect 184013 518050 184047 518084
rect 184105 518050 184139 518084
rect 184197 518050 184231 518084
rect 184289 518050 184323 518084
rect 184381 518050 184415 518084
rect 184473 518050 184507 518084
rect 184565 518050 184599 518084
rect 184657 518050 184691 518084
rect 184749 518050 184783 518084
rect 184841 518050 184875 518084
rect 184933 518050 184967 518084
rect 185025 518050 185059 518084
rect 185117 518050 185151 518084
rect 185209 518050 185243 518084
rect 185301 518050 185335 518084
rect 185393 518050 185427 518084
rect 185485 518050 185519 518084
rect 185577 518050 185611 518084
rect 185669 518050 185703 518084
rect 185761 518050 185795 518084
rect 185853 518050 185887 518084
rect 185945 518050 185979 518084
rect 186037 518050 186071 518084
rect 186129 518050 186163 518084
rect 186221 518050 186255 518084
rect 186313 518050 186347 518084
rect 186405 518050 186439 518084
rect 186497 518050 186531 518084
rect 186589 518050 186623 518084
rect 186681 518050 186715 518084
rect 186773 518050 186807 518084
rect 186865 518050 186899 518084
rect 186957 518050 186991 518084
rect 187049 518050 187083 518084
rect 187141 518050 187175 518084
rect 187233 518050 187267 518084
rect 187325 518050 187359 518084
rect 187417 518050 187451 518084
rect 172237 517506 172271 517540
rect 172329 517506 172363 517540
rect 172421 517506 172455 517540
rect 172513 517506 172547 517540
rect 172605 517506 172639 517540
rect 172697 517506 172731 517540
rect 172789 517506 172823 517540
rect 172881 517506 172915 517540
rect 172973 517506 173007 517540
rect 173065 517506 173099 517540
rect 173157 517506 173191 517540
rect 173249 517506 173283 517540
rect 173341 517506 173375 517540
rect 173433 517506 173467 517540
rect 173525 517506 173559 517540
rect 173617 517506 173651 517540
rect 173709 517506 173743 517540
rect 173801 517506 173835 517540
rect 173893 517506 173927 517540
rect 173985 517506 174019 517540
rect 174077 517506 174111 517540
rect 174169 517506 174203 517540
rect 174261 517506 174295 517540
rect 174353 517506 174387 517540
rect 174445 517506 174479 517540
rect 174537 517506 174571 517540
rect 174629 517506 174663 517540
rect 174721 517506 174755 517540
rect 174813 517506 174847 517540
rect 174905 517506 174939 517540
rect 174997 517506 175031 517540
rect 175089 517506 175123 517540
rect 175181 517506 175215 517540
rect 175273 517506 175307 517540
rect 175365 517506 175399 517540
rect 175457 517506 175491 517540
rect 175549 517506 175583 517540
rect 175641 517506 175675 517540
rect 175733 517506 175767 517540
rect 175825 517506 175859 517540
rect 175917 517506 175951 517540
rect 176009 517506 176043 517540
rect 176101 517506 176135 517540
rect 176193 517506 176227 517540
rect 176285 517506 176319 517540
rect 176377 517506 176411 517540
rect 176469 517506 176503 517540
rect 176561 517506 176595 517540
rect 176653 517506 176687 517540
rect 176745 517506 176779 517540
rect 176837 517506 176871 517540
rect 176929 517506 176963 517540
rect 177021 517506 177055 517540
rect 177113 517506 177147 517540
rect 177205 517506 177239 517540
rect 177297 517506 177331 517540
rect 177389 517506 177423 517540
rect 177481 517506 177515 517540
rect 177573 517506 177607 517540
rect 177665 517506 177699 517540
rect 177757 517506 177791 517540
rect 177849 517506 177883 517540
rect 177941 517506 177975 517540
rect 178033 517506 178067 517540
rect 178125 517506 178159 517540
rect 178217 517506 178251 517540
rect 178309 517506 178343 517540
rect 178401 517506 178435 517540
rect 178493 517506 178527 517540
rect 178585 517506 178619 517540
rect 178677 517506 178711 517540
rect 178769 517506 178803 517540
rect 178861 517506 178895 517540
rect 178953 517506 178987 517540
rect 179045 517506 179079 517540
rect 179137 517506 179171 517540
rect 179229 517506 179263 517540
rect 179321 517506 179355 517540
rect 179413 517506 179447 517540
rect 179505 517506 179539 517540
rect 179597 517506 179631 517540
rect 179689 517506 179723 517540
rect 179781 517506 179815 517540
rect 179873 517506 179907 517540
rect 179965 517506 179999 517540
rect 180057 517506 180091 517540
rect 180149 517506 180183 517540
rect 180241 517506 180275 517540
rect 180333 517506 180367 517540
rect 180425 517506 180459 517540
rect 180517 517506 180551 517540
rect 180609 517506 180643 517540
rect 180701 517506 180735 517540
rect 180793 517506 180827 517540
rect 180885 517506 180919 517540
rect 180977 517506 181011 517540
rect 181069 517506 181103 517540
rect 181161 517506 181195 517540
rect 181253 517506 181287 517540
rect 181345 517506 181379 517540
rect 181437 517506 181471 517540
rect 181529 517506 181563 517540
rect 181621 517506 181655 517540
rect 181713 517506 181747 517540
rect 181805 517506 181839 517540
rect 181897 517506 181931 517540
rect 181989 517506 182023 517540
rect 182081 517506 182115 517540
rect 182173 517506 182207 517540
rect 182265 517506 182299 517540
rect 182357 517506 182391 517540
rect 182449 517506 182483 517540
rect 182541 517506 182575 517540
rect 182633 517506 182667 517540
rect 182725 517506 182759 517540
rect 182817 517506 182851 517540
rect 182909 517506 182943 517540
rect 183001 517506 183035 517540
rect 183093 517506 183127 517540
rect 183185 517506 183219 517540
rect 183277 517506 183311 517540
rect 183369 517506 183403 517540
rect 183461 517506 183495 517540
rect 183553 517506 183587 517540
rect 183645 517506 183679 517540
rect 183737 517506 183771 517540
rect 183829 517506 183863 517540
rect 183921 517506 183955 517540
rect 184013 517506 184047 517540
rect 184105 517506 184139 517540
rect 184197 517506 184231 517540
rect 184289 517506 184323 517540
rect 184381 517506 184415 517540
rect 184473 517506 184507 517540
rect 184565 517506 184599 517540
rect 184657 517506 184691 517540
rect 184749 517506 184783 517540
rect 184841 517506 184875 517540
rect 184933 517506 184967 517540
rect 185025 517506 185059 517540
rect 185117 517506 185151 517540
rect 185209 517506 185243 517540
rect 185301 517506 185335 517540
rect 185393 517506 185427 517540
rect 185485 517506 185519 517540
rect 185577 517506 185611 517540
rect 185669 517506 185703 517540
rect 185761 517506 185795 517540
rect 185853 517506 185887 517540
rect 185945 517506 185979 517540
rect 186037 517506 186071 517540
rect 186129 517506 186163 517540
rect 186221 517506 186255 517540
rect 186313 517506 186347 517540
rect 186405 517506 186439 517540
rect 186497 517506 186531 517540
rect 186589 517506 186623 517540
rect 186681 517506 186715 517540
rect 186773 517506 186807 517540
rect 186865 517506 186899 517540
rect 186957 517506 186991 517540
rect 187049 517506 187083 517540
rect 187141 517506 187175 517540
rect 187233 517506 187267 517540
rect 187325 517506 187359 517540
rect 187417 517506 187451 517540
rect 172237 516962 172271 516996
rect 172329 516962 172363 516996
rect 172421 516962 172455 516996
rect 172513 516962 172547 516996
rect 172605 516962 172639 516996
rect 172697 516962 172731 516996
rect 172789 516962 172823 516996
rect 172881 516962 172915 516996
rect 172973 516962 173007 516996
rect 173065 516962 173099 516996
rect 173157 516962 173191 516996
rect 173249 516962 173283 516996
rect 173341 516962 173375 516996
rect 173433 516962 173467 516996
rect 173525 516962 173559 516996
rect 173617 516962 173651 516996
rect 173709 516962 173743 516996
rect 173801 516962 173835 516996
rect 173893 516962 173927 516996
rect 173985 516962 174019 516996
rect 174077 516962 174111 516996
rect 174169 516962 174203 516996
rect 174261 516962 174295 516996
rect 174353 516962 174387 516996
rect 174445 516962 174479 516996
rect 174537 516962 174571 516996
rect 174629 516962 174663 516996
rect 174721 516962 174755 516996
rect 174813 516962 174847 516996
rect 174905 516962 174939 516996
rect 174997 516962 175031 516996
rect 175089 516962 175123 516996
rect 175181 516962 175215 516996
rect 175273 516962 175307 516996
rect 175365 516962 175399 516996
rect 175457 516962 175491 516996
rect 175549 516962 175583 516996
rect 175641 516962 175675 516996
rect 175733 516962 175767 516996
rect 175825 516962 175859 516996
rect 175917 516962 175951 516996
rect 176009 516962 176043 516996
rect 176101 516962 176135 516996
rect 176193 516962 176227 516996
rect 176285 516962 176319 516996
rect 176377 516962 176411 516996
rect 176469 516962 176503 516996
rect 176561 516962 176595 516996
rect 176653 516962 176687 516996
rect 176745 516962 176779 516996
rect 176837 516962 176871 516996
rect 176929 516962 176963 516996
rect 177021 516962 177055 516996
rect 177113 516962 177147 516996
rect 177205 516962 177239 516996
rect 177297 516962 177331 516996
rect 177389 516962 177423 516996
rect 177481 516962 177515 516996
rect 177573 516962 177607 516996
rect 177665 516962 177699 516996
rect 177757 516962 177791 516996
rect 177849 516962 177883 516996
rect 177941 516962 177975 516996
rect 178033 516962 178067 516996
rect 178125 516962 178159 516996
rect 178217 516962 178251 516996
rect 178309 516962 178343 516996
rect 178401 516962 178435 516996
rect 178493 516962 178527 516996
rect 178585 516962 178619 516996
rect 178677 516962 178711 516996
rect 178769 516962 178803 516996
rect 178861 516962 178895 516996
rect 178953 516962 178987 516996
rect 179045 516962 179079 516996
rect 179137 516962 179171 516996
rect 179229 516962 179263 516996
rect 179321 516962 179355 516996
rect 179413 516962 179447 516996
rect 179505 516962 179539 516996
rect 179597 516962 179631 516996
rect 179689 516962 179723 516996
rect 179781 516962 179815 516996
rect 179873 516962 179907 516996
rect 179965 516962 179999 516996
rect 180057 516962 180091 516996
rect 180149 516962 180183 516996
rect 180241 516962 180275 516996
rect 180333 516962 180367 516996
rect 180425 516962 180459 516996
rect 180517 516962 180551 516996
rect 180609 516962 180643 516996
rect 180701 516962 180735 516996
rect 180793 516962 180827 516996
rect 180885 516962 180919 516996
rect 180977 516962 181011 516996
rect 181069 516962 181103 516996
rect 181161 516962 181195 516996
rect 181253 516962 181287 516996
rect 181345 516962 181379 516996
rect 181437 516962 181471 516996
rect 181529 516962 181563 516996
rect 181621 516962 181655 516996
rect 181713 516962 181747 516996
rect 181805 516962 181839 516996
rect 181897 516962 181931 516996
rect 181989 516962 182023 516996
rect 182081 516962 182115 516996
rect 182173 516962 182207 516996
rect 182265 516962 182299 516996
rect 182357 516962 182391 516996
rect 182449 516962 182483 516996
rect 182541 516962 182575 516996
rect 182633 516962 182667 516996
rect 182725 516962 182759 516996
rect 182817 516962 182851 516996
rect 182909 516962 182943 516996
rect 183001 516962 183035 516996
rect 183093 516962 183127 516996
rect 183185 516962 183219 516996
rect 183277 516962 183311 516996
rect 183369 516962 183403 516996
rect 183461 516962 183495 516996
rect 183553 516962 183587 516996
rect 183645 516962 183679 516996
rect 183737 516962 183771 516996
rect 183829 516962 183863 516996
rect 183921 516962 183955 516996
rect 184013 516962 184047 516996
rect 184105 516962 184139 516996
rect 184197 516962 184231 516996
rect 184289 516962 184323 516996
rect 184381 516962 184415 516996
rect 184473 516962 184507 516996
rect 184565 516962 184599 516996
rect 184657 516962 184691 516996
rect 184749 516962 184783 516996
rect 184841 516962 184875 516996
rect 184933 516962 184967 516996
rect 185025 516962 185059 516996
rect 185117 516962 185151 516996
rect 185209 516962 185243 516996
rect 185301 516962 185335 516996
rect 185393 516962 185427 516996
rect 185485 516962 185519 516996
rect 185577 516962 185611 516996
rect 185669 516962 185703 516996
rect 185761 516962 185795 516996
rect 185853 516962 185887 516996
rect 185945 516962 185979 516996
rect 186037 516962 186071 516996
rect 186129 516962 186163 516996
rect 186221 516962 186255 516996
rect 186313 516962 186347 516996
rect 186405 516962 186439 516996
rect 186497 516962 186531 516996
rect 186589 516962 186623 516996
rect 186681 516962 186715 516996
rect 186773 516962 186807 516996
rect 186865 516962 186899 516996
rect 186957 516962 186991 516996
rect 187049 516962 187083 516996
rect 187141 516962 187175 516996
rect 187233 516962 187267 516996
rect 187325 516962 187359 516996
rect 187417 516962 187451 516996
rect 172237 516418 172271 516452
rect 172329 516418 172363 516452
rect 172421 516418 172455 516452
rect 172513 516418 172547 516452
rect 172605 516418 172639 516452
rect 172697 516418 172731 516452
rect 172789 516418 172823 516452
rect 172881 516418 172915 516452
rect 172973 516418 173007 516452
rect 173065 516418 173099 516452
rect 173157 516418 173191 516452
rect 173249 516418 173283 516452
rect 173341 516418 173375 516452
rect 173433 516418 173467 516452
rect 173525 516418 173559 516452
rect 173617 516418 173651 516452
rect 173709 516418 173743 516452
rect 173801 516418 173835 516452
rect 173893 516418 173927 516452
rect 173985 516418 174019 516452
rect 174077 516418 174111 516452
rect 174169 516418 174203 516452
rect 174261 516418 174295 516452
rect 174353 516418 174387 516452
rect 174445 516418 174479 516452
rect 174537 516418 174571 516452
rect 174629 516418 174663 516452
rect 174721 516418 174755 516452
rect 174813 516418 174847 516452
rect 174905 516418 174939 516452
rect 174997 516418 175031 516452
rect 175089 516418 175123 516452
rect 175181 516418 175215 516452
rect 175273 516418 175307 516452
rect 175365 516418 175399 516452
rect 175457 516418 175491 516452
rect 175549 516418 175583 516452
rect 175641 516418 175675 516452
rect 175733 516418 175767 516452
rect 175825 516418 175859 516452
rect 175917 516418 175951 516452
rect 176009 516418 176043 516452
rect 176101 516418 176135 516452
rect 176193 516418 176227 516452
rect 176285 516418 176319 516452
rect 176377 516418 176411 516452
rect 176469 516418 176503 516452
rect 176561 516418 176595 516452
rect 176653 516418 176687 516452
rect 176745 516418 176779 516452
rect 176837 516418 176871 516452
rect 176929 516418 176963 516452
rect 177021 516418 177055 516452
rect 177113 516418 177147 516452
rect 177205 516418 177239 516452
rect 177297 516418 177331 516452
rect 177389 516418 177423 516452
rect 177481 516418 177515 516452
rect 177573 516418 177607 516452
rect 177665 516418 177699 516452
rect 177757 516418 177791 516452
rect 177849 516418 177883 516452
rect 177941 516418 177975 516452
rect 178033 516418 178067 516452
rect 178125 516418 178159 516452
rect 178217 516418 178251 516452
rect 178309 516418 178343 516452
rect 178401 516418 178435 516452
rect 178493 516418 178527 516452
rect 178585 516418 178619 516452
rect 178677 516418 178711 516452
rect 178769 516418 178803 516452
rect 178861 516418 178895 516452
rect 178953 516418 178987 516452
rect 179045 516418 179079 516452
rect 179137 516418 179171 516452
rect 179229 516418 179263 516452
rect 179321 516418 179355 516452
rect 179413 516418 179447 516452
rect 179505 516418 179539 516452
rect 179597 516418 179631 516452
rect 179689 516418 179723 516452
rect 179781 516418 179815 516452
rect 179873 516418 179907 516452
rect 179965 516418 179999 516452
rect 180057 516418 180091 516452
rect 180149 516418 180183 516452
rect 180241 516418 180275 516452
rect 180333 516418 180367 516452
rect 180425 516418 180459 516452
rect 180517 516418 180551 516452
rect 180609 516418 180643 516452
rect 180701 516418 180735 516452
rect 180793 516418 180827 516452
rect 180885 516418 180919 516452
rect 180977 516418 181011 516452
rect 181069 516418 181103 516452
rect 181161 516418 181195 516452
rect 181253 516418 181287 516452
rect 181345 516418 181379 516452
rect 181437 516418 181471 516452
rect 181529 516418 181563 516452
rect 181621 516418 181655 516452
rect 181713 516418 181747 516452
rect 181805 516418 181839 516452
rect 181897 516418 181931 516452
rect 181989 516418 182023 516452
rect 182081 516418 182115 516452
rect 182173 516418 182207 516452
rect 182265 516418 182299 516452
rect 182357 516418 182391 516452
rect 182449 516418 182483 516452
rect 182541 516418 182575 516452
rect 182633 516418 182667 516452
rect 182725 516418 182759 516452
rect 182817 516418 182851 516452
rect 182909 516418 182943 516452
rect 183001 516418 183035 516452
rect 183093 516418 183127 516452
rect 183185 516418 183219 516452
rect 183277 516418 183311 516452
rect 183369 516418 183403 516452
rect 183461 516418 183495 516452
rect 183553 516418 183587 516452
rect 183645 516418 183679 516452
rect 183737 516418 183771 516452
rect 183829 516418 183863 516452
rect 183921 516418 183955 516452
rect 184013 516418 184047 516452
rect 184105 516418 184139 516452
rect 184197 516418 184231 516452
rect 184289 516418 184323 516452
rect 184381 516418 184415 516452
rect 184473 516418 184507 516452
rect 184565 516418 184599 516452
rect 184657 516418 184691 516452
rect 184749 516418 184783 516452
rect 184841 516418 184875 516452
rect 184933 516418 184967 516452
rect 185025 516418 185059 516452
rect 185117 516418 185151 516452
rect 185209 516418 185243 516452
rect 185301 516418 185335 516452
rect 185393 516418 185427 516452
rect 185485 516418 185519 516452
rect 185577 516418 185611 516452
rect 185669 516418 185703 516452
rect 185761 516418 185795 516452
rect 185853 516418 185887 516452
rect 185945 516418 185979 516452
rect 186037 516418 186071 516452
rect 186129 516418 186163 516452
rect 186221 516418 186255 516452
rect 186313 516418 186347 516452
rect 186405 516418 186439 516452
rect 186497 516418 186531 516452
rect 186589 516418 186623 516452
rect 186681 516418 186715 516452
rect 186773 516418 186807 516452
rect 186865 516418 186899 516452
rect 186957 516418 186991 516452
rect 187049 516418 187083 516452
rect 187141 516418 187175 516452
rect 187233 516418 187267 516452
rect 187325 516418 187359 516452
rect 187417 516418 187451 516452
rect 172237 515874 172271 515908
rect 172329 515874 172363 515908
rect 172421 515874 172455 515908
rect 172513 515874 172547 515908
rect 172605 515874 172639 515908
rect 172697 515874 172731 515908
rect 172789 515874 172823 515908
rect 172881 515874 172915 515908
rect 172973 515874 173007 515908
rect 173065 515874 173099 515908
rect 173157 515874 173191 515908
rect 173249 515874 173283 515908
rect 173341 515874 173375 515908
rect 173433 515874 173467 515908
rect 173525 515874 173559 515908
rect 173617 515874 173651 515908
rect 173709 515874 173743 515908
rect 173801 515874 173835 515908
rect 173893 515874 173927 515908
rect 173985 515874 174019 515908
rect 174077 515874 174111 515908
rect 174169 515874 174203 515908
rect 174261 515874 174295 515908
rect 174353 515874 174387 515908
rect 174445 515874 174479 515908
rect 174537 515874 174571 515908
rect 174629 515874 174663 515908
rect 174721 515874 174755 515908
rect 174813 515874 174847 515908
rect 174905 515874 174939 515908
rect 174997 515874 175031 515908
rect 175089 515874 175123 515908
rect 175181 515874 175215 515908
rect 175273 515874 175307 515908
rect 175365 515874 175399 515908
rect 175457 515874 175491 515908
rect 175549 515874 175583 515908
rect 175641 515874 175675 515908
rect 175733 515874 175767 515908
rect 175825 515874 175859 515908
rect 175917 515874 175951 515908
rect 176009 515874 176043 515908
rect 176101 515874 176135 515908
rect 176193 515874 176227 515908
rect 176285 515874 176319 515908
rect 176377 515874 176411 515908
rect 176469 515874 176503 515908
rect 176561 515874 176595 515908
rect 176653 515874 176687 515908
rect 176745 515874 176779 515908
rect 176837 515874 176871 515908
rect 176929 515874 176963 515908
rect 177021 515874 177055 515908
rect 177113 515874 177147 515908
rect 177205 515874 177239 515908
rect 177297 515874 177331 515908
rect 177389 515874 177423 515908
rect 177481 515874 177515 515908
rect 177573 515874 177607 515908
rect 177665 515874 177699 515908
rect 177757 515874 177791 515908
rect 177849 515874 177883 515908
rect 177941 515874 177975 515908
rect 178033 515874 178067 515908
rect 178125 515874 178159 515908
rect 178217 515874 178251 515908
rect 178309 515874 178343 515908
rect 178401 515874 178435 515908
rect 178493 515874 178527 515908
rect 178585 515874 178619 515908
rect 178677 515874 178711 515908
rect 178769 515874 178803 515908
rect 178861 515874 178895 515908
rect 178953 515874 178987 515908
rect 179045 515874 179079 515908
rect 179137 515874 179171 515908
rect 179229 515874 179263 515908
rect 179321 515874 179355 515908
rect 179413 515874 179447 515908
rect 179505 515874 179539 515908
rect 179597 515874 179631 515908
rect 179689 515874 179723 515908
rect 179781 515874 179815 515908
rect 179873 515874 179907 515908
rect 179965 515874 179999 515908
rect 180057 515874 180091 515908
rect 180149 515874 180183 515908
rect 180241 515874 180275 515908
rect 180333 515874 180367 515908
rect 180425 515874 180459 515908
rect 180517 515874 180551 515908
rect 180609 515874 180643 515908
rect 180701 515874 180735 515908
rect 180793 515874 180827 515908
rect 180885 515874 180919 515908
rect 180977 515874 181011 515908
rect 181069 515874 181103 515908
rect 181161 515874 181195 515908
rect 181253 515874 181287 515908
rect 181345 515874 181379 515908
rect 181437 515874 181471 515908
rect 181529 515874 181563 515908
rect 181621 515874 181655 515908
rect 181713 515874 181747 515908
rect 181805 515874 181839 515908
rect 181897 515874 181931 515908
rect 181989 515874 182023 515908
rect 182081 515874 182115 515908
rect 182173 515874 182207 515908
rect 182265 515874 182299 515908
rect 182357 515874 182391 515908
rect 182449 515874 182483 515908
rect 182541 515874 182575 515908
rect 182633 515874 182667 515908
rect 182725 515874 182759 515908
rect 182817 515874 182851 515908
rect 182909 515874 182943 515908
rect 183001 515874 183035 515908
rect 183093 515874 183127 515908
rect 183185 515874 183219 515908
rect 183277 515874 183311 515908
rect 183369 515874 183403 515908
rect 183461 515874 183495 515908
rect 183553 515874 183587 515908
rect 183645 515874 183679 515908
rect 183737 515874 183771 515908
rect 183829 515874 183863 515908
rect 183921 515874 183955 515908
rect 184013 515874 184047 515908
rect 184105 515874 184139 515908
rect 184197 515874 184231 515908
rect 184289 515874 184323 515908
rect 184381 515874 184415 515908
rect 184473 515874 184507 515908
rect 184565 515874 184599 515908
rect 184657 515874 184691 515908
rect 184749 515874 184783 515908
rect 184841 515874 184875 515908
rect 184933 515874 184967 515908
rect 185025 515874 185059 515908
rect 185117 515874 185151 515908
rect 185209 515874 185243 515908
rect 185301 515874 185335 515908
rect 185393 515874 185427 515908
rect 185485 515874 185519 515908
rect 185577 515874 185611 515908
rect 185669 515874 185703 515908
rect 185761 515874 185795 515908
rect 185853 515874 185887 515908
rect 185945 515874 185979 515908
rect 186037 515874 186071 515908
rect 186129 515874 186163 515908
rect 186221 515874 186255 515908
rect 186313 515874 186347 515908
rect 186405 515874 186439 515908
rect 186497 515874 186531 515908
rect 186589 515874 186623 515908
rect 186681 515874 186715 515908
rect 186773 515874 186807 515908
rect 186865 515874 186899 515908
rect 186957 515874 186991 515908
rect 187049 515874 187083 515908
rect 187141 515874 187175 515908
rect 187233 515874 187267 515908
rect 187325 515874 187359 515908
rect 187417 515874 187451 515908
rect 173617 515797 173651 515806
rect 173617 515772 173621 515797
rect 173621 515772 173651 515797
rect 173525 515500 173559 515534
rect 182081 515790 182087 515806
rect 182087 515790 182115 515806
rect 182081 515772 182115 515790
rect 182265 515596 182299 515602
rect 182265 515568 182291 515596
rect 182291 515568 182299 515596
rect 186589 515797 186623 515806
rect 186589 515772 186593 515797
rect 186593 515772 186623 515797
rect 186497 515500 186531 515534
rect 172237 515330 172271 515364
rect 172329 515330 172363 515364
rect 172421 515330 172455 515364
rect 172513 515330 172547 515364
rect 172605 515330 172639 515364
rect 172697 515330 172731 515364
rect 172789 515330 172823 515364
rect 172881 515330 172915 515364
rect 172973 515330 173007 515364
rect 173065 515330 173099 515364
rect 173157 515330 173191 515364
rect 173249 515330 173283 515364
rect 173341 515330 173375 515364
rect 173433 515330 173467 515364
rect 173525 515330 173559 515364
rect 173617 515330 173651 515364
rect 173709 515330 173743 515364
rect 173801 515330 173835 515364
rect 173893 515330 173927 515364
rect 173985 515330 174019 515364
rect 174077 515330 174111 515364
rect 174169 515330 174203 515364
rect 174261 515330 174295 515364
rect 174353 515330 174387 515364
rect 174445 515330 174479 515364
rect 174537 515330 174571 515364
rect 174629 515330 174663 515364
rect 174721 515330 174755 515364
rect 174813 515330 174847 515364
rect 174905 515330 174939 515364
rect 174997 515330 175031 515364
rect 175089 515330 175123 515364
rect 175181 515330 175215 515364
rect 175273 515330 175307 515364
rect 175365 515330 175399 515364
rect 175457 515330 175491 515364
rect 175549 515330 175583 515364
rect 175641 515330 175675 515364
rect 175733 515330 175767 515364
rect 175825 515330 175859 515364
rect 175917 515330 175951 515364
rect 176009 515330 176043 515364
rect 176101 515330 176135 515364
rect 176193 515330 176227 515364
rect 176285 515330 176319 515364
rect 176377 515330 176411 515364
rect 176469 515330 176503 515364
rect 176561 515330 176595 515364
rect 176653 515330 176687 515364
rect 176745 515330 176779 515364
rect 176837 515330 176871 515364
rect 176929 515330 176963 515364
rect 177021 515330 177055 515364
rect 177113 515330 177147 515364
rect 177205 515330 177239 515364
rect 177297 515330 177331 515364
rect 177389 515330 177423 515364
rect 177481 515330 177515 515364
rect 177573 515330 177607 515364
rect 177665 515330 177699 515364
rect 177757 515330 177791 515364
rect 177849 515330 177883 515364
rect 177941 515330 177975 515364
rect 178033 515330 178067 515364
rect 178125 515330 178159 515364
rect 178217 515330 178251 515364
rect 178309 515330 178343 515364
rect 178401 515330 178435 515364
rect 178493 515330 178527 515364
rect 178585 515330 178619 515364
rect 178677 515330 178711 515364
rect 178769 515330 178803 515364
rect 178861 515330 178895 515364
rect 178953 515330 178987 515364
rect 179045 515330 179079 515364
rect 179137 515330 179171 515364
rect 179229 515330 179263 515364
rect 179321 515330 179355 515364
rect 179413 515330 179447 515364
rect 179505 515330 179539 515364
rect 179597 515330 179631 515364
rect 179689 515330 179723 515364
rect 179781 515330 179815 515364
rect 179873 515330 179907 515364
rect 179965 515330 179999 515364
rect 180057 515330 180091 515364
rect 180149 515330 180183 515364
rect 180241 515330 180275 515364
rect 180333 515330 180367 515364
rect 180425 515330 180459 515364
rect 180517 515330 180551 515364
rect 180609 515330 180643 515364
rect 180701 515330 180735 515364
rect 180793 515330 180827 515364
rect 180885 515330 180919 515364
rect 180977 515330 181011 515364
rect 181069 515330 181103 515364
rect 181161 515330 181195 515364
rect 181253 515330 181287 515364
rect 181345 515330 181379 515364
rect 181437 515330 181471 515364
rect 181529 515330 181563 515364
rect 181621 515330 181655 515364
rect 181713 515330 181747 515364
rect 181805 515330 181839 515364
rect 181897 515330 181931 515364
rect 181989 515330 182023 515364
rect 182081 515330 182115 515364
rect 182173 515330 182207 515364
rect 182265 515330 182299 515364
rect 182357 515330 182391 515364
rect 182449 515330 182483 515364
rect 182541 515330 182575 515364
rect 182633 515330 182667 515364
rect 182725 515330 182759 515364
rect 182817 515330 182851 515364
rect 182909 515330 182943 515364
rect 183001 515330 183035 515364
rect 183093 515330 183127 515364
rect 183185 515330 183219 515364
rect 183277 515330 183311 515364
rect 183369 515330 183403 515364
rect 183461 515330 183495 515364
rect 183553 515330 183587 515364
rect 183645 515330 183679 515364
rect 183737 515330 183771 515364
rect 183829 515330 183863 515364
rect 183921 515330 183955 515364
rect 184013 515330 184047 515364
rect 184105 515330 184139 515364
rect 184197 515330 184231 515364
rect 184289 515330 184323 515364
rect 184381 515330 184415 515364
rect 184473 515330 184507 515364
rect 184565 515330 184599 515364
rect 184657 515330 184691 515364
rect 184749 515330 184783 515364
rect 184841 515330 184875 515364
rect 184933 515330 184967 515364
rect 185025 515330 185059 515364
rect 185117 515330 185151 515364
rect 185209 515330 185243 515364
rect 185301 515330 185335 515364
rect 185393 515330 185427 515364
rect 185485 515330 185519 515364
rect 185577 515330 185611 515364
rect 185669 515330 185703 515364
rect 185761 515330 185795 515364
rect 185853 515330 185887 515364
rect 185945 515330 185979 515364
rect 186037 515330 186071 515364
rect 186129 515330 186163 515364
rect 186221 515330 186255 515364
rect 186313 515330 186347 515364
rect 186405 515330 186439 515364
rect 186497 515330 186531 515364
rect 186589 515330 186623 515364
rect 186681 515330 186715 515364
rect 186773 515330 186807 515364
rect 186865 515330 186899 515364
rect 186957 515330 186991 515364
rect 187049 515330 187083 515364
rect 187141 515330 187175 515364
rect 187233 515330 187267 515364
rect 187325 515330 187359 515364
rect 187417 515330 187451 515364
<< metal1 >>
rect 17990 699000 18000 701000
rect 20000 699000 20010 701000
rect 69990 699000 70000 701000
rect 72000 699000 72010 701000
rect 121990 699000 122000 701000
rect 124000 699000 124010 701000
rect 18000 687000 20000 699000
rect 70000 691000 72000 699000
rect 122000 695000 124000 699000
rect 122000 693000 156000 695000
rect 70000 689000 152000 691000
rect 18000 685000 148000 687000
rect 2990 682000 3000 684000
rect 5000 682000 11000 684000
rect 9000 533000 11000 682000
rect 146000 628000 148000 685000
rect 145990 626000 146000 628000
rect 148000 626000 148010 628000
rect 150000 549000 152000 689000
rect 154000 553000 156000 693000
rect 153990 551000 154000 553000
rect 156000 551000 156010 553000
rect 150000 547000 179000 549000
rect 145990 544000 146000 546000
rect 148000 544000 163800 546000
rect 177000 544000 179000 547000
rect 163500 542900 163800 544000
rect 178100 542900 178400 544000
rect 153990 538000 154000 540000
rect 156000 538000 156010 540000
rect 163200 538865 163228 538875
rect 163018 538835 163028 538865
rect 158678 538715 163028 538835
rect 158678 538585 158978 538715
rect 158668 538505 158978 538585
rect 158668 538469 158958 538505
rect 158668 538435 158726 538469
rect 158894 538435 158958 538469
rect 158668 538397 158958 538435
rect 158658 538385 158962 538397
rect 158658 538209 158664 538385
rect 158698 538355 158922 538385
rect 158698 538209 158704 538355
rect 158658 538197 158704 538209
rect 158916 538209 158922 538355
rect 158956 538209 158962 538385
rect 159028 538395 159058 538715
rect 161378 538665 161528 538675
rect 161378 538545 161388 538665
rect 161508 538545 161528 538665
rect 161378 538535 161528 538545
rect 159090 538469 159282 538475
rect 159090 538435 159102 538469
rect 159270 538435 159282 538469
rect 159090 538429 159282 538435
rect 159348 538469 159540 538475
rect 159348 538435 159360 538469
rect 159528 538435 159540 538469
rect 159348 538429 159540 538435
rect 159606 538469 159798 538475
rect 159606 538435 159618 538469
rect 159786 538435 159798 538469
rect 159606 538429 159798 538435
rect 159864 538469 160056 538475
rect 159864 538435 159876 538469
rect 160044 538435 160056 538469
rect 159864 538429 160056 538435
rect 160122 538469 160314 538475
rect 160122 538435 160134 538469
rect 160302 538435 160314 538469
rect 160122 538429 160314 538435
rect 160380 538469 160572 538475
rect 160380 538435 160392 538469
rect 160560 538435 160572 538469
rect 160380 538429 160572 538435
rect 160638 538469 160830 538475
rect 160638 538435 160650 538469
rect 160818 538435 160830 538469
rect 160638 538429 160830 538435
rect 160896 538469 161088 538475
rect 160896 538435 160908 538469
rect 161076 538435 161088 538469
rect 160896 538429 161088 538435
rect 161154 538469 161346 538475
rect 161154 538435 161166 538469
rect 161334 538435 161346 538469
rect 161154 538429 161346 538435
rect 161438 538397 161498 538535
rect 161534 538469 161726 538475
rect 161534 538435 161546 538469
rect 161714 538435 161726 538469
rect 161534 538429 161726 538435
rect 161808 538405 161848 538715
rect 162258 538705 162558 538715
rect 162258 538665 162268 538705
rect 162528 538665 162558 538705
rect 163018 538665 163028 538715
rect 163328 538665 163338 538865
rect 161934 538469 162126 538475
rect 161934 538435 161946 538469
rect 162114 538435 162126 538469
rect 161934 538429 162126 538435
rect 162258 538469 162558 538665
rect 163020 538660 163200 538665
rect 162258 538435 162326 538469
rect 162494 538435 162558 538469
rect 161748 538397 161908 538405
rect 162258 538397 162558 538435
rect 159028 538368 161148 538395
rect 159028 538355 159040 538368
rect 159034 538280 159040 538355
rect 159074 538355 159556 538368
rect 159074 538280 159080 538355
rect 159034 538268 159080 538280
rect 159292 538314 159338 538326
rect 159292 538235 159298 538314
rect 158916 538197 158962 538209
rect 159288 538226 159298 538235
rect 159332 538235 159338 538314
rect 159388 538295 159488 538305
rect 159388 538235 159398 538295
rect 159332 538226 159398 538235
rect 159288 538215 159398 538226
rect 159478 538235 159488 538295
rect 159550 538280 159556 538355
rect 159590 538355 160072 538368
rect 159590 538280 159596 538355
rect 159550 538268 159596 538280
rect 159808 538314 159854 538326
rect 159808 538235 159814 538314
rect 159478 538226 159814 538235
rect 159848 538235 159854 538314
rect 160066 538280 160072 538355
rect 160106 538355 160588 538368
rect 160106 538280 160112 538355
rect 160066 538268 160112 538280
rect 160324 538314 160370 538326
rect 160324 538235 160330 538314
rect 159848 538226 160330 538235
rect 160364 538235 160370 538314
rect 160582 538280 160588 538355
rect 160622 538355 161104 538368
rect 160622 538280 160628 538355
rect 160582 538268 160628 538280
rect 160840 538314 160886 538326
rect 160840 538235 160846 538314
rect 160364 538226 160846 538235
rect 160880 538235 160886 538314
rect 161098 538280 161104 538355
rect 161138 538355 161148 538368
rect 161438 538385 161524 538397
rect 161138 538280 161144 538355
rect 161098 538268 161144 538280
rect 161356 538314 161402 538326
rect 161356 538235 161362 538314
rect 160880 538226 161362 538235
rect 161396 538226 161402 538314
rect 159478 538215 161402 538226
rect 159288 538214 161402 538215
rect 159288 538195 161388 538214
rect 161438 538209 161484 538385
rect 161518 538209 161524 538385
rect 161438 538197 161524 538209
rect 161736 538385 161924 538397
rect 161736 538209 161742 538385
rect 161776 538209 161884 538385
rect 161918 538345 161924 538385
rect 162136 538385 162182 538397
rect 161918 538305 161928 538345
rect 161918 538209 161924 538305
rect 161736 538205 161924 538209
rect 161736 538197 161782 538205
rect 161878 538197 161924 538205
rect 162136 538209 162142 538385
rect 162176 538365 162182 538385
rect 162258 538385 162562 538397
rect 162176 538225 162188 538365
rect 162176 538209 162208 538225
rect 162136 538197 162208 538209
rect 162258 538209 162264 538385
rect 162298 538305 162522 538385
rect 162298 538209 162304 538305
rect 162258 538197 162304 538209
rect 162516 538209 162522 538305
rect 162556 538209 162562 538385
rect 162516 538197 162562 538209
rect 161438 538195 161498 538197
rect 158714 538159 158906 538165
rect 158714 538125 158726 538159
rect 158894 538125 158906 538159
rect 159090 538159 159282 538165
rect 159090 538155 159102 538159
rect 158714 538119 158906 538125
rect 159088 538125 159102 538155
rect 159270 538155 159282 538159
rect 159348 538159 159540 538165
rect 159348 538155 159360 538159
rect 159270 538125 159360 538155
rect 159528 538155 159540 538159
rect 159606 538159 159798 538165
rect 159606 538155 159618 538159
rect 159528 538125 159618 538155
rect 159786 538155 159798 538159
rect 159864 538159 160056 538165
rect 159864 538155 159876 538159
rect 159786 538125 159876 538155
rect 160044 538155 160056 538159
rect 160122 538159 160314 538165
rect 160122 538155 160134 538159
rect 160044 538125 160134 538155
rect 160302 538155 160314 538159
rect 160380 538159 160572 538165
rect 160380 538155 160392 538159
rect 160302 538125 160392 538155
rect 160560 538155 160572 538159
rect 160638 538159 160830 538165
rect 160638 538155 160650 538159
rect 160560 538125 160650 538155
rect 160818 538155 160830 538159
rect 160896 538159 161088 538165
rect 160896 538155 160908 538159
rect 160818 538125 160908 538155
rect 161076 538155 161088 538159
rect 161154 538159 161346 538165
rect 161154 538155 161166 538159
rect 161076 538125 161166 538155
rect 161334 538155 161346 538159
rect 161448 538155 161488 538195
rect 162168 538165 162208 538197
rect 161334 538125 161488 538155
rect 161528 538159 162208 538165
rect 161528 538125 161546 538159
rect 161714 538125 161946 538159
rect 162114 538125 162208 538159
rect 159088 538115 161488 538125
rect 161534 538119 161726 538125
rect 161934 538119 162126 538125
rect 154000 537000 156000 538000
rect 161448 537965 161488 538115
rect 162168 537965 162208 538125
rect 162314 538159 162506 538165
rect 162314 538125 162326 538159
rect 162494 538125 162506 538159
rect 162314 538119 162506 538125
rect 163528 538035 163728 542900
rect 178178 541705 178378 542900
rect 164278 541505 188978 541705
rect 164278 540965 164478 541505
rect 164718 541125 164778 541135
rect 165018 541130 166038 541155
rect 165018 541126 166253 541130
rect 164678 541119 164818 541125
rect 164678 541085 164728 541119
rect 164762 541085 164818 541119
rect 165018 541095 165031 541126
rect 165019 541092 165031 541095
rect 165065 541095 165223 541126
rect 165065 541092 165077 541095
rect 165019 541086 165077 541092
rect 165211 541092 165223 541095
rect 165257 541095 165415 541126
rect 165257 541092 165269 541095
rect 165211 541086 165269 541092
rect 165403 541092 165415 541095
rect 165449 541095 165607 541126
rect 165449 541092 165461 541095
rect 165403 541086 165461 541092
rect 165595 541092 165607 541095
rect 165641 541095 165799 541126
rect 165641 541092 165653 541095
rect 165595 541086 165653 541092
rect 165787 541092 165799 541095
rect 165833 541095 165991 541126
rect 165833 541092 165845 541095
rect 165787 541086 165845 541092
rect 165979 541092 165991 541095
rect 166025 541092 166253 541126
rect 165979 541086 166253 541092
rect 164678 541018 164818 541085
rect 166023 541080 166253 541086
rect 164678 540965 164684 541018
rect 164278 540885 164684 540965
rect 164278 540835 164478 540885
rect 164678 540530 164684 540885
rect 164718 540885 164772 541018
rect 164718 540530 164724 540885
rect 164678 540518 164724 540530
rect 164766 540530 164772 540885
rect 164806 540965 164818 541018
rect 164977 541025 165023 541037
rect 165169 541025 165215 541037
rect 165361 541025 165407 541037
rect 165553 541025 165599 541037
rect 165745 541025 165791 541037
rect 165937 541025 165983 541037
rect 164977 540965 164983 541025
rect 164806 540885 164983 540965
rect 164806 540530 164812 540885
rect 164766 540518 164812 540530
rect 164881 540571 164927 540583
rect 164881 540285 164887 540571
rect 164848 540083 164887 540285
rect 164921 540285 164927 540571
rect 164977 540537 164983 540885
rect 165017 540635 165175 541025
rect 165017 540537 165023 540635
rect 164977 540525 165023 540537
rect 165073 540571 165119 540583
rect 165073 540285 165079 540571
rect 164921 540083 165079 540285
rect 165113 540285 165119 540571
rect 165169 540537 165175 540635
rect 165209 540635 165367 541025
rect 165209 540537 165215 540635
rect 165169 540525 165215 540537
rect 165265 540571 165311 540583
rect 165265 540285 165271 540571
rect 165113 540083 165271 540285
rect 165305 540285 165311 540571
rect 165361 540537 165367 540635
rect 165401 540635 165559 541025
rect 165401 540537 165407 540635
rect 165361 540525 165407 540537
rect 165457 540571 165503 540583
rect 165457 540285 165463 540571
rect 165305 540083 165463 540285
rect 165497 540285 165503 540571
rect 165553 540537 165559 540635
rect 165593 540635 165751 541025
rect 165593 540537 165599 540635
rect 165553 540525 165599 540537
rect 165649 540571 165695 540583
rect 165649 540285 165655 540571
rect 165497 540083 165655 540285
rect 165689 540285 165695 540571
rect 165745 540537 165751 540635
rect 165785 540995 165943 541025
rect 165977 540995 166008 541025
rect 165785 540895 165888 540995
rect 165998 540895 166008 540995
rect 165785 540875 165943 540895
rect 165977 540875 166008 540895
rect 165785 540775 165888 540875
rect 165998 540775 166008 540875
rect 166203 540830 166253 541080
rect 166396 541119 166458 541125
rect 166396 541085 166408 541119
rect 166442 541085 166458 541119
rect 166396 541079 166458 541085
rect 166398 541065 166458 541079
rect 168078 540965 168278 541505
rect 168518 541125 168578 541135
rect 168818 541130 169838 541155
rect 168818 541126 170053 541130
rect 168478 541119 168618 541125
rect 168478 541085 168528 541119
rect 168562 541085 168618 541119
rect 168818 541095 168831 541126
rect 168819 541092 168831 541095
rect 168865 541095 169023 541126
rect 168865 541092 168877 541095
rect 168819 541086 168877 541092
rect 169011 541092 169023 541095
rect 169057 541095 169215 541126
rect 169057 541092 169069 541095
rect 169011 541086 169069 541092
rect 169203 541092 169215 541095
rect 169249 541095 169407 541126
rect 169249 541092 169261 541095
rect 169203 541086 169261 541092
rect 169395 541092 169407 541095
rect 169441 541095 169599 541126
rect 169441 541092 169453 541095
rect 169395 541086 169453 541092
rect 169587 541092 169599 541095
rect 169633 541095 169791 541126
rect 169633 541092 169645 541095
rect 169587 541086 169645 541092
rect 169779 541092 169791 541095
rect 169825 541092 170053 541126
rect 169779 541086 170053 541092
rect 168478 541018 168618 541085
rect 169823 541080 170053 541086
rect 168478 540965 168484 541018
rect 166678 540830 167718 540895
rect 168078 540885 168484 540965
rect 168078 540835 168278 540885
rect 165785 540755 165943 540775
rect 165977 540755 166008 540775
rect 165785 540655 165888 540755
rect 165998 540655 166008 540755
rect 165785 540635 165943 540655
rect 165785 540537 165791 540635
rect 165745 540525 165791 540537
rect 165841 540571 165887 540583
rect 165841 540285 165847 540571
rect 165689 540083 165847 540285
rect 165881 540285 165887 540571
rect 165937 540537 165943 540635
rect 165977 540635 166008 540655
rect 166198 540780 167718 540830
rect 165977 540537 165983 540635
rect 165937 540525 165983 540537
rect 166033 540571 166079 540583
rect 166033 540285 166039 540571
rect 165881 540083 166039 540285
rect 166073 540083 166079 540571
rect 166198 540335 166248 540780
rect 166678 540695 167718 540780
rect 166358 540564 166404 540576
rect 166198 540325 166258 540335
rect 166196 540319 166258 540325
rect 166196 540285 166208 540319
rect 166242 540285 166258 540319
rect 166196 540279 166258 540285
rect 166198 540275 166258 540279
rect 166158 540235 166204 540247
rect 166158 540155 166164 540235
rect 164848 540075 166079 540083
rect 164848 540071 164927 540075
rect 165073 540071 165119 540075
rect 165265 540071 165311 540075
rect 165457 540071 165503 540075
rect 165649 540071 165695 540075
rect 165841 540071 165887 540075
rect 166033 540071 166079 540075
rect 164848 540065 164918 540071
rect 164708 540009 164778 540025
rect 164708 539975 164728 540009
rect 164762 539975 164778 540009
rect 164708 539955 164778 539975
rect 164848 539755 164878 540065
rect 166138 540059 166164 540155
rect 166198 540059 166204 540235
rect 166138 540047 166204 540059
rect 166246 540235 166292 540247
rect 166246 540059 166252 540235
rect 166286 540225 166292 540235
rect 166358 540225 166364 540564
rect 166286 540076 166364 540225
rect 166398 540235 166404 540564
rect 166446 540564 166492 540576
rect 166446 540235 166452 540564
rect 166398 540076 166452 540235
rect 166486 540235 166492 540564
rect 166668 540245 166888 540255
rect 166486 540225 166508 540235
rect 166668 540225 166688 540245
rect 166486 540215 166688 540225
rect 166486 540085 166568 540215
rect 166628 540085 166688 540215
rect 166486 540076 166688 540085
rect 166286 540075 166688 540076
rect 166286 540059 166292 540075
rect 166358 540064 166492 540075
rect 166668 540065 166688 540075
rect 166868 540065 166888 540245
rect 166246 540047 166292 540059
rect 164923 540016 164981 540022
rect 164923 540015 164935 540016
rect 164918 539982 164935 540015
rect 164969 540015 164981 540016
rect 165115 540016 165173 540022
rect 165115 540015 165127 540016
rect 164969 539982 165127 540015
rect 165161 540015 165173 540016
rect 165307 540016 165365 540022
rect 165307 540015 165319 540016
rect 165161 539982 165319 540015
rect 165353 540015 165365 540016
rect 165499 540016 165557 540022
rect 165499 540015 165511 540016
rect 165353 539982 165511 540015
rect 165545 540015 165557 540016
rect 165691 540016 165749 540022
rect 165691 540015 165703 540016
rect 165545 539982 165703 540015
rect 165737 540015 165749 540016
rect 165883 540016 165941 540022
rect 165883 540015 165895 540016
rect 165737 539982 165895 540015
rect 165929 539982 165941 540016
rect 164918 539976 165941 539982
rect 164918 539955 165938 539976
rect 161448 537925 161648 537965
rect 161288 537706 161348 537725
rect 161288 537672 161302 537706
rect 161336 537672 161348 537706
rect 161288 537665 161348 537672
rect 161488 537712 161548 537725
rect 161488 537706 161552 537712
rect 161488 537672 161506 537706
rect 161540 537672 161552 537706
rect 161488 537666 161552 537672
rect 161488 537665 161548 537666
rect 161608 537625 161648 537925
rect 162008 537925 162208 537965
rect 162868 537945 162948 537955
rect 161678 537735 161758 537745
rect 161678 537675 161688 537735
rect 161748 537675 161758 537735
rect 161678 537672 161698 537675
rect 161732 537672 161758 537675
rect 161678 537665 161758 537672
rect 161888 537712 161948 537725
rect 161888 537706 161952 537712
rect 161888 537672 161906 537706
rect 161940 537672 161952 537706
rect 161888 537666 161952 537672
rect 161888 537665 161948 537666
rect 161548 537608 161768 537625
rect 162008 537608 162048 537925
rect 162868 537885 162878 537945
rect 162938 537935 162948 537945
rect 163018 537935 163728 538035
rect 162938 537885 163728 537935
rect 162868 537875 162948 537885
rect 163018 537835 163728 537885
rect 164278 539655 164878 539755
rect 164278 537931 164478 539655
rect 164638 539606 164878 539655
rect 164638 539572 164712 539606
rect 164746 539572 164878 539606
rect 164638 539513 164878 539572
rect 165018 539619 166028 539625
rect 165018 539613 166041 539619
rect 165018 539579 165035 539613
rect 165069 539579 165227 539613
rect 165261 539579 165419 539613
rect 165453 539579 165611 539613
rect 165645 539579 165803 539613
rect 165837 539579 165995 539613
rect 166029 539579 166041 539613
rect 165018 539573 166041 539579
rect 165018 539565 166028 539573
rect 166138 539525 166168 540047
rect 166196 540009 166258 540015
rect 166196 539975 166208 540009
rect 166242 539975 166258 540009
rect 166196 539969 166258 539975
rect 166198 539606 166258 539969
rect 166368 540009 166488 540064
rect 166668 540055 166888 540065
rect 166368 539975 166408 540009
rect 166442 539975 166488 540009
rect 166368 539955 166488 539975
rect 166198 539572 166212 539606
rect 166246 539572 166258 539606
rect 166198 539565 166258 539572
rect 166398 539606 166478 539625
rect 166398 539572 166412 539606
rect 166446 539572 166478 539606
rect 166398 539565 166478 539572
rect 164638 539415 164668 539513
rect 164662 538537 164668 539415
rect 164702 539415 164756 539513
rect 164702 538537 164708 539415
rect 164662 538525 164708 538537
rect 164750 538537 164756 539415
rect 164790 539495 164878 539513
rect 164981 539503 165027 539515
rect 164790 539485 164948 539495
rect 164981 539485 164987 539503
rect 164790 539415 164987 539485
rect 164790 538537 164796 539415
rect 164848 539205 164987 539415
rect 164885 539049 164931 539061
rect 164885 538561 164891 539049
rect 164925 538935 164931 539049
rect 164981 539015 164987 539205
rect 165021 539485 165027 539503
rect 165173 539503 165219 539515
rect 165173 539485 165179 539503
rect 165021 539205 165179 539485
rect 165021 539015 165027 539205
rect 164981 539003 165027 539015
rect 165077 539049 165123 539061
rect 165077 538935 165083 539049
rect 164925 538561 165083 538935
rect 165117 538935 165123 539049
rect 165173 539015 165179 539205
rect 165213 539485 165219 539503
rect 165365 539503 165411 539515
rect 165365 539485 165371 539503
rect 165213 539205 165371 539485
rect 165213 539015 165219 539205
rect 165173 539003 165219 539015
rect 165269 539049 165315 539061
rect 165269 538935 165275 539049
rect 165117 538561 165275 538935
rect 165309 538935 165315 539049
rect 165365 539015 165371 539205
rect 165405 539485 165411 539503
rect 165557 539503 165603 539515
rect 165557 539485 165563 539503
rect 165405 539205 165563 539485
rect 165405 539015 165411 539205
rect 165365 539003 165411 539015
rect 165461 539049 165507 539061
rect 165461 538935 165467 539049
rect 165309 538561 165467 538935
rect 165501 538935 165507 539049
rect 165557 539015 165563 539205
rect 165597 539485 165603 539503
rect 165749 539503 165795 539515
rect 165749 539485 165755 539503
rect 165597 539205 165755 539485
rect 165597 539015 165603 539205
rect 165557 539003 165603 539015
rect 165653 539049 165699 539061
rect 165653 538935 165659 539049
rect 165501 538561 165659 538935
rect 165693 538935 165699 539049
rect 165749 539015 165755 539205
rect 165789 539485 165795 539503
rect 165941 539503 165987 539515
rect 165941 539485 165947 539503
rect 165789 539205 165947 539485
rect 165789 539015 165795 539205
rect 165749 539003 165795 539015
rect 165845 539049 165891 539061
rect 165845 538935 165851 539049
rect 165693 538561 165851 538935
rect 165885 538935 165891 539049
rect 165941 539015 165947 539205
rect 165981 539485 165987 539503
rect 166138 539513 166208 539525
rect 165981 539205 165998 539485
rect 166138 539375 166168 539513
rect 165981 539015 165987 539205
rect 165941 539003 165987 539015
rect 166037 539049 166083 539061
rect 166037 538935 166043 539049
rect 165885 538805 166043 538935
rect 165885 538705 165898 538805
rect 166038 538705 166043 538805
rect 165885 538561 166043 538705
rect 166077 538561 166083 539049
rect 166162 539035 166168 539375
rect 164885 538555 166083 538561
rect 164885 538549 164931 538555
rect 165077 538549 165123 538555
rect 165269 538549 165315 538555
rect 165461 538549 165507 538555
rect 165653 538549 165699 538555
rect 165845 538549 165891 538555
rect 166037 538549 166083 538555
rect 166128 538937 166168 539035
rect 166202 538937 166208 539513
rect 166128 538925 166208 538937
rect 166250 539513 166296 539525
rect 166250 538937 166256 539513
rect 166290 539505 166296 539513
rect 166290 539275 166408 539505
rect 166668 539305 166888 539315
rect 166668 539275 166688 539305
rect 166290 539265 166688 539275
rect 166290 539175 166568 539265
rect 166618 539175 166688 539265
rect 166290 539165 166688 539175
rect 166290 539042 166408 539165
rect 166668 539125 166688 539165
rect 166868 539125 166888 539305
rect 166668 539115 166888 539125
rect 166290 538937 166368 539042
rect 166250 538935 166368 538937
rect 166250 538925 166296 538935
rect 164750 538525 164796 538537
rect 164927 538485 164985 538491
rect 165119 538485 165177 538491
rect 165311 538485 165369 538491
rect 165503 538485 165561 538491
rect 165695 538485 165753 538491
rect 165887 538485 165945 538491
rect 166128 538485 166168 538925
rect 166198 538878 166258 538885
rect 166198 538844 166212 538878
rect 166246 538844 166258 538878
rect 166198 538825 166258 538844
rect 166362 538575 166368 538935
rect 164698 538478 164758 538485
rect 164698 538444 164712 538478
rect 164746 538444 164758 538478
rect 164698 538425 164758 538444
rect 164918 538451 164939 538485
rect 164973 538451 165131 538485
rect 165165 538451 165323 538485
rect 165357 538451 165515 538485
rect 165549 538451 165707 538485
rect 165741 538451 165899 538485
rect 165933 538451 166168 538485
rect 164918 538425 166168 538451
rect 166358 538554 166368 538575
rect 166402 538575 166408 539042
rect 166450 539042 166496 539054
rect 166450 538575 166456 539042
rect 166402 538554 166456 538575
rect 166490 538554 166496 539042
rect 166358 538542 166496 538554
rect 166358 538478 166478 538542
rect 166358 538445 166412 538478
rect 166398 538444 166412 538445
rect 166446 538445 166478 538478
rect 166446 538444 166458 538445
rect 166398 538425 166458 538444
rect 166558 537943 167303 537945
rect 164278 537815 164332 537931
rect 162088 537712 162148 537725
rect 162086 537706 162148 537712
rect 162086 537672 162098 537706
rect 162132 537672 162148 537706
rect 162086 537666 162148 537672
rect 162088 537665 162148 537666
rect 162308 537706 162368 537725
rect 162308 537672 162322 537706
rect 162356 537672 162368 537706
rect 162308 537665 162368 537672
rect 161548 537596 161786 537608
rect 161252 537342 161298 537354
rect 161252 537225 161258 537342
rect 161248 537075 161258 537225
rect 161252 537054 161258 537075
rect 161292 537225 161298 537342
rect 161340 537342 161386 537354
rect 161340 537225 161346 537342
rect 161292 537054 161346 537225
rect 161380 537225 161386 537342
rect 161452 537342 161498 537354
rect 161452 537225 161458 537342
rect 161380 537075 161458 537225
rect 161380 537054 161386 537075
rect 161252 537042 161386 537054
rect 161452 537054 161458 537075
rect 161492 537225 161498 537342
rect 161548 537308 161554 537596
rect 161588 537465 161746 537596
rect 161588 537308 161594 537465
rect 161548 537296 161594 537308
rect 161644 537342 161690 537354
rect 161644 537225 161650 537342
rect 161492 537065 161650 537225
rect 161492 537054 161498 537065
rect 161452 537042 161498 537054
rect 161644 537054 161650 537065
rect 161684 537225 161690 537342
rect 161740 537308 161746 537465
rect 161780 537308 161786 537596
rect 161740 537296 161786 537308
rect 161852 537605 161898 537608
rect 162008 537605 162090 537608
rect 161852 537596 162090 537605
rect 161852 537308 161858 537596
rect 161892 537465 162050 537596
rect 161892 537308 161898 537465
rect 161852 537296 161898 537308
rect 161948 537342 161994 537354
rect 161948 537225 161954 537342
rect 161684 537065 161954 537225
rect 161684 537054 161690 537065
rect 161644 537042 161690 537054
rect 154000 536965 156800 537000
rect 161278 536978 161358 537042
rect 154000 536955 156998 536965
rect 154000 536935 157398 536955
rect 161278 536945 161302 536978
rect 161288 536944 161302 536945
rect 161336 536945 161358 536978
rect 161588 536978 161648 536985
rect 161336 536944 161348 536945
rect 154000 536925 157523 536935
rect 161288 536925 161348 536944
rect 161588 536944 161602 536978
rect 161636 536944 161648 536978
rect 161588 536925 161648 536944
rect 154000 536845 157418 536925
rect 157508 536845 157523 536925
rect 154000 536825 157523 536845
rect 161768 536905 161868 537065
rect 161948 537054 161954 537065
rect 161988 537225 161994 537342
rect 162044 537308 162050 537465
rect 162084 537308 162090 537596
rect 164326 537534 164332 537815
rect 164370 537815 164478 537931
rect 164644 537935 164694 537943
rect 164962 537935 165012 537943
rect 164644 537931 165012 537935
rect 164370 537534 164376 537815
rect 164326 537522 164376 537534
rect 164644 537534 164650 537931
rect 164688 537535 164968 537931
rect 164688 537534 164694 537535
rect 164644 537522 164694 537534
rect 164962 537534 164968 537535
rect 165006 537534 165012 537931
rect 164962 537522 165012 537534
rect 165280 537931 165330 537943
rect 165280 537534 165286 537931
rect 165324 537925 165330 537931
rect 165598 537931 165648 537943
rect 165598 537925 165604 537931
rect 165324 537565 165604 537925
rect 165324 537534 165330 537565
rect 165280 537522 165330 537534
rect 165598 537534 165604 537565
rect 165642 537534 165648 537931
rect 165598 537522 165648 537534
rect 165916 537931 165966 537943
rect 165916 537534 165922 537931
rect 165960 537925 165966 537931
rect 166234 537931 166284 537943
rect 166234 537925 166240 537931
rect 165960 537565 166240 537925
rect 165960 537534 165966 537565
rect 165916 537522 165966 537534
rect 166234 537534 166240 537565
rect 166278 537534 166284 537931
rect 166234 537522 166284 537534
rect 166552 537931 167303 537943
rect 166552 537534 166558 537931
rect 166596 537534 167303 537931
rect 166552 537522 167303 537534
rect 166558 537515 167303 537522
rect 162044 537296 162090 537308
rect 162140 537342 162186 537354
rect 162140 537225 162146 537342
rect 161988 537065 162146 537225
rect 161988 537054 161994 537065
rect 161948 537042 161994 537054
rect 162140 537054 162146 537065
rect 162180 537205 162186 537342
rect 162272 537342 162318 537354
rect 162272 537205 162278 537342
rect 162180 537085 162278 537205
rect 162180 537054 162186 537085
rect 162140 537042 162186 537054
rect 162272 537054 162278 537085
rect 162312 537095 162318 537342
rect 162360 537342 162406 537354
rect 162360 537095 162366 537342
rect 162312 537054 162366 537095
rect 162400 537095 162406 537342
rect 163018 537135 163728 537195
rect 162400 537054 162408 537095
rect 162272 537042 162408 537054
rect 161768 536825 161788 536905
rect 161848 536825 161868 536905
rect 154000 536800 157398 536825
rect 161768 536805 161868 536825
rect 161988 536978 162048 536985
rect 161988 536944 162002 536978
rect 162036 536975 162048 536978
rect 162278 536978 162408 537042
rect 162036 536944 162058 536975
rect 161988 536885 162058 536944
rect 162278 536944 162322 536978
rect 162356 536944 162408 536978
rect 162278 536935 162408 536944
rect 162908 537065 163728 537135
rect 162308 536925 162368 536935
rect 162908 536885 162958 537065
rect 163018 536995 163728 537065
rect 161988 536815 162958 536885
rect 156700 536765 157398 536800
rect 156700 536700 156800 536765
rect 157198 536755 157398 536765
rect 162298 536725 162718 536785
rect 162298 536705 162358 536725
rect 157798 536686 157990 536692
rect 157798 536652 157810 536686
rect 157978 536652 157990 536686
rect 157798 536646 157990 536652
rect 158148 536686 162358 536705
rect 162658 536705 162718 536725
rect 163028 536705 163228 536765
rect 158148 536652 158188 536686
rect 158356 536652 158446 536686
rect 158614 536652 158704 536686
rect 158872 536652 158962 536686
rect 159130 536652 159220 536686
rect 159388 536652 159478 536686
rect 159646 536652 159736 536686
rect 159904 536652 159994 536686
rect 160162 536652 160252 536686
rect 160420 536652 160510 536686
rect 160678 536652 160894 536686
rect 161062 536652 161152 536686
rect 161320 536652 161410 536686
rect 161578 536652 161792 536686
rect 161960 536652 162050 536686
rect 162218 536652 162358 536686
rect 158148 536645 162358 536652
rect 162418 536686 162610 536692
rect 162418 536652 162430 536686
rect 162598 536652 162610 536686
rect 162418 536646 162610 536652
rect 162658 536645 163228 536705
rect 157742 536593 157788 536605
rect 157742 536125 157748 536593
rect 157738 536017 157748 536125
rect 157782 536125 157788 536593
rect 158000 536593 158046 536605
rect 158000 536125 158006 536593
rect 157782 536017 158006 536125
rect 158040 536125 158046 536593
rect 161988 536588 162028 536645
rect 158378 536576 158424 536588
rect 158120 536322 158166 536334
rect 158040 536017 158048 536125
rect 158120 536034 158126 536322
rect 158160 536145 158166 536322
rect 158378 536288 158384 536576
rect 158418 536565 158424 536576
rect 158894 536576 158940 536588
rect 158894 536565 158900 536576
rect 158418 536555 158900 536565
rect 158418 536455 158478 536555
rect 158418 536288 158424 536455
rect 158468 536395 158478 536455
rect 158578 536455 158900 536555
rect 158578 536395 158598 536455
rect 158468 536375 158598 536395
rect 158378 536276 158424 536288
rect 158636 536322 158682 536334
rect 158636 536145 158642 536322
rect 158160 536045 158642 536145
rect 158160 536034 158166 536045
rect 158120 536022 158166 536034
rect 158636 536034 158642 536045
rect 158676 536145 158682 536322
rect 158894 536288 158900 536455
rect 158934 536565 158940 536576
rect 159410 536576 159456 536588
rect 159410 536565 159416 536576
rect 158934 536455 159416 536565
rect 158934 536288 158940 536455
rect 158894 536276 158940 536288
rect 159152 536322 159198 536334
rect 159152 536145 159158 536322
rect 158676 536045 159158 536145
rect 158676 536034 158682 536045
rect 158636 536022 158682 536034
rect 159152 536034 159158 536045
rect 159192 536145 159198 536322
rect 159410 536288 159416 536455
rect 159450 536565 159456 536576
rect 159926 536576 159972 536588
rect 159926 536565 159932 536576
rect 159450 536455 159932 536565
rect 159450 536288 159456 536455
rect 159410 536276 159456 536288
rect 159668 536322 159714 536334
rect 159668 536145 159674 536322
rect 159192 536045 159674 536145
rect 159192 536034 159198 536045
rect 159152 536022 159198 536034
rect 159668 536034 159674 536045
rect 159708 536145 159714 536322
rect 159926 536288 159932 536455
rect 159966 536565 159972 536576
rect 160442 536576 160488 536588
rect 160442 536565 160448 536576
rect 159966 536455 160448 536565
rect 159966 536288 159972 536455
rect 159926 536276 159972 536288
rect 160184 536322 160230 536334
rect 160184 536145 160190 536322
rect 159708 536045 160190 536145
rect 159708 536034 159714 536045
rect 159668 536022 159714 536034
rect 160184 536034 160190 536045
rect 160224 536145 160230 536322
rect 160442 536288 160448 536455
rect 160482 536565 160488 536576
rect 160826 536585 160872 536588
rect 161342 536585 161388 536588
rect 160826 536576 161388 536585
rect 160482 536455 160508 536565
rect 160482 536288 160488 536455
rect 160442 536276 160488 536288
rect 160700 536322 160746 536334
rect 160700 536145 160706 536322
rect 160224 536045 160706 536145
rect 160224 536034 160230 536045
rect 160184 536022 160230 536034
rect 160700 536034 160706 536045
rect 160740 536145 160746 536322
rect 160826 536288 160832 536576
rect 160866 536545 161348 536576
rect 160866 536465 161088 536545
rect 161168 536465 161348 536545
rect 160866 536425 161348 536465
rect 160866 536288 160872 536425
rect 160826 536276 160872 536288
rect 161084 536322 161130 536334
rect 161084 536165 161090 536322
rect 160740 536034 160768 536145
rect 161068 536045 161090 536165
rect 160700 536022 160768 536034
rect 161084 536034 161090 536045
rect 161124 536165 161130 536322
rect 161342 536288 161348 536425
rect 161382 536288 161388 536576
rect 161982 536576 162028 536588
rect 161342 536276 161388 536288
rect 161600 536322 161646 536334
rect 161600 536165 161606 536322
rect 161124 536045 161606 536165
rect 161124 536034 161130 536045
rect 161084 536022 161130 536034
rect 161600 536034 161606 536045
rect 161640 536165 161646 536322
rect 161724 536322 161770 536334
rect 161640 536034 161668 536165
rect 161600 536022 161668 536034
rect 161724 536034 161730 536322
rect 161764 536185 161770 536322
rect 161982 536288 161988 536576
rect 162022 536288 162028 536576
rect 162362 536593 162408 536605
rect 161982 536276 162028 536288
rect 162240 536322 162286 536334
rect 162240 536185 162246 536322
rect 161764 536065 162246 536185
rect 161764 536034 161770 536065
rect 161724 536022 161770 536034
rect 162240 536034 162246 536065
rect 162280 536185 162286 536322
rect 162280 536034 162308 536185
rect 162240 536022 162308 536034
rect 157738 535958 158048 536017
rect 157738 535924 157810 535958
rect 157978 535924 158048 535958
rect 157738 535805 158048 535924
rect 158176 535958 158368 535964
rect 158176 535924 158188 535958
rect 158356 535924 158368 535958
rect 158176 535918 158368 535924
rect 158434 535958 158626 535964
rect 158434 535924 158446 535958
rect 158614 535924 158626 535958
rect 158434 535918 158626 535924
rect 158692 535958 158884 535964
rect 158692 535924 158704 535958
rect 158872 535924 158884 535958
rect 158692 535918 158884 535924
rect 158950 535958 159142 535964
rect 158950 535924 158962 535958
rect 159130 535924 159142 535958
rect 158950 535918 159142 535924
rect 159208 535958 159400 535964
rect 159208 535924 159220 535958
rect 159388 535924 159400 535958
rect 159208 535918 159400 535924
rect 159466 535958 159658 535964
rect 159466 535924 159478 535958
rect 159646 535924 159658 535958
rect 159466 535918 159658 535924
rect 159724 535958 159916 535964
rect 159724 535924 159736 535958
rect 159904 535924 159916 535958
rect 159724 535918 159916 535924
rect 159982 535958 160174 535964
rect 159982 535924 159994 535958
rect 160162 535924 160174 535958
rect 159982 535918 160174 535924
rect 160240 535958 160432 535964
rect 160240 535924 160252 535958
rect 160420 535924 160432 535958
rect 160240 535918 160432 535924
rect 160498 535958 160690 535964
rect 160498 535924 160510 535958
rect 160678 535924 160690 535958
rect 160498 535918 160690 535924
rect 160728 535805 160768 536022
rect 160882 535958 161074 535964
rect 160882 535924 160894 535958
rect 161062 535924 161074 535958
rect 160882 535918 161074 535924
rect 161140 535958 161332 535964
rect 161140 535924 161152 535958
rect 161320 535924 161332 535958
rect 161140 535918 161332 535924
rect 161398 535958 161590 535964
rect 161398 535924 161410 535958
rect 161578 535924 161590 535958
rect 161398 535918 161590 535924
rect 161628 535805 161668 536022
rect 161780 535958 161972 535964
rect 161780 535924 161792 535958
rect 161960 535924 161972 535958
rect 161780 535918 161972 535924
rect 162038 535958 162230 535964
rect 162038 535924 162050 535958
rect 162218 535924 162230 535958
rect 162038 535918 162230 535924
rect 162268 535805 162308 536022
rect 162362 536017 162368 536593
rect 162402 536085 162408 536593
rect 162620 536593 162666 536605
rect 162620 536085 162626 536593
rect 162402 536017 162626 536085
rect 162660 536085 162666 536593
rect 162660 536017 162668 536085
rect 162362 536005 162668 536017
rect 162378 535958 162668 536005
rect 162378 535924 162430 535958
rect 162598 535924 162668 535958
rect 162378 535805 162668 535924
rect 157738 535765 162708 535805
rect 157748 535745 162708 535765
rect 157748 535705 162048 535745
rect 162648 535705 162708 535745
rect 157748 535685 162708 535705
rect 160208 535585 160328 535685
rect 160178 535575 160378 535585
rect 160178 535435 160198 535575
rect 160348 535435 160378 535575
rect 160178 535420 160378 535435
rect 163028 533120 163228 536645
rect 163528 536275 163728 536995
rect 164326 536416 164376 536428
rect 163528 536235 164098 536275
rect 163528 535905 163838 536235
rect 164048 535905 164098 536235
rect 164326 536019 164332 536416
rect 164370 536415 164376 536416
rect 164644 536416 164694 536428
rect 164644 536415 164650 536416
rect 164370 536019 164650 536415
rect 164688 536019 164694 536416
rect 164326 536015 164694 536019
rect 164326 536007 164376 536015
rect 164644 536007 164694 536015
rect 164962 536416 165012 536428
rect 164962 536019 164968 536416
rect 165006 536415 165012 536416
rect 165280 536416 165330 536428
rect 165280 536415 165286 536416
rect 165006 536019 165286 536415
rect 165324 536019 165330 536416
rect 164962 536015 165330 536019
rect 164962 536007 165012 536015
rect 165280 536007 165330 536015
rect 165598 536416 165648 536428
rect 165598 536019 165604 536416
rect 165642 536415 165648 536416
rect 165916 536416 165966 536428
rect 165916 536415 165922 536416
rect 165642 536055 165922 536415
rect 165642 536019 165648 536055
rect 165598 536007 165648 536019
rect 165916 536019 165922 536055
rect 165960 536019 165966 536416
rect 165916 536007 165966 536019
rect 166234 536416 166284 536428
rect 166234 536019 166240 536416
rect 166278 536395 166284 536416
rect 166552 536416 166602 536428
rect 166552 536395 166558 536416
rect 166278 536035 166558 536395
rect 166278 536019 166284 536035
rect 166234 536007 166284 536019
rect 166552 536019 166558 536035
rect 166596 536019 166602 536416
rect 166552 536007 166602 536019
rect 166873 536265 167303 537515
rect 166873 536045 166928 536265
rect 167258 536045 167303 536265
rect 166873 535980 167303 536045
rect 163528 535885 164098 535905
rect 163528 535635 163798 535885
rect 163528 535591 164378 535635
rect 163528 535235 164302 535591
rect 163528 535225 163798 535235
rect 164296 535194 164302 535235
rect 164340 535235 164378 535591
rect 164614 535595 164664 535603
rect 164932 535595 164982 535603
rect 164614 535591 164982 535595
rect 164340 535194 164346 535235
rect 164296 535182 164346 535194
rect 164614 535194 164620 535591
rect 164658 535225 164938 535591
rect 164658 535194 164664 535225
rect 164614 535182 164664 535194
rect 164932 535194 164938 535225
rect 164976 535194 164982 535591
rect 164932 535182 164982 535194
rect 165250 535595 165300 535603
rect 165568 535595 165618 535603
rect 165250 535591 165618 535595
rect 165250 535194 165256 535591
rect 165294 535225 165574 535591
rect 165294 535194 165300 535225
rect 165250 535182 165300 535194
rect 165568 535194 165574 535225
rect 165612 535194 165618 535591
rect 165568 535182 165618 535194
rect 165886 535591 165936 535603
rect 165886 535194 165892 535591
rect 165930 535575 165936 535591
rect 166204 535591 166254 535603
rect 166204 535575 166210 535591
rect 165930 535205 166210 535575
rect 165930 535194 165936 535205
rect 165886 535182 165936 535194
rect 166204 535194 166210 535205
rect 166248 535194 166254 535591
rect 166498 535591 167263 535615
rect 166498 535205 166528 535591
rect 166204 535182 166254 535194
rect 166522 535194 166528 535205
rect 166566 535555 167263 535591
rect 166566 535425 166718 535555
rect 166848 535545 167263 535555
rect 166848 535425 166898 535545
rect 166566 535415 166898 535425
rect 167028 535525 167263 535545
rect 167028 535415 167078 535525
rect 166566 535395 167078 535415
rect 167208 535395 167263 535525
rect 166566 535365 167263 535395
rect 166566 535235 166698 535365
rect 166828 535355 167263 535365
rect 166828 535235 166888 535355
rect 166566 535225 166888 535235
rect 167018 535345 167263 535355
rect 167018 535225 167088 535345
rect 166566 535215 167088 535225
rect 167218 535215 167263 535345
rect 166566 535205 167263 535215
rect 166566 535194 166572 535205
rect 166522 535182 166572 535194
rect 164296 534076 164346 534088
rect 164296 533679 164302 534076
rect 164340 534065 164346 534076
rect 164614 534076 164664 534088
rect 164614 534065 164620 534076
rect 164340 533695 164620 534065
rect 164340 533679 164346 533695
rect 164296 533667 164346 533679
rect 164614 533679 164620 533695
rect 164658 534065 164664 534076
rect 164932 534076 164982 534088
rect 164658 533695 164668 534065
rect 164658 533679 164664 533695
rect 164614 533667 164664 533679
rect 164932 533679 164938 534076
rect 164976 534065 164982 534076
rect 165250 534076 165300 534088
rect 165250 534065 165256 534076
rect 164976 533695 165256 534065
rect 164976 533679 164982 533695
rect 164932 533667 164982 533679
rect 165250 533679 165256 533695
rect 165294 533679 165300 534076
rect 165250 533667 165300 533679
rect 165568 534076 165618 534088
rect 165568 533679 165574 534076
rect 165612 534065 165618 534076
rect 165886 534076 165936 534088
rect 165886 534065 165892 534076
rect 165612 533695 165892 534065
rect 165612 533679 165618 533695
rect 165568 533667 165618 533679
rect 165886 533679 165892 533695
rect 165930 533679 165936 534076
rect 165886 533667 165936 533679
rect 166204 534076 166254 534088
rect 166204 533679 166210 534076
rect 166248 534055 166254 534076
rect 166522 534076 166572 534088
rect 166522 534055 166528 534076
rect 166248 533685 166528 534055
rect 166248 533679 166254 533685
rect 166204 533667 166254 533679
rect 166522 533679 166528 533685
rect 166566 533679 166572 534076
rect 166522 533667 166572 533679
rect 163020 533115 163228 533120
rect 163020 533000 163220 533115
rect 9000 531000 163220 533000
rect 167518 532755 167718 540695
rect 168478 540530 168484 540885
rect 168518 540885 168572 541018
rect 168518 540530 168524 540885
rect 168478 540518 168524 540530
rect 168566 540530 168572 540885
rect 168606 540965 168618 541018
rect 168777 541025 168823 541037
rect 168969 541025 169015 541037
rect 169161 541025 169207 541037
rect 169353 541025 169399 541037
rect 169545 541025 169591 541037
rect 169737 541025 169783 541037
rect 168777 540965 168783 541025
rect 168606 540885 168783 540965
rect 168606 540530 168612 540885
rect 168566 540518 168612 540530
rect 168681 540571 168727 540583
rect 168681 540285 168687 540571
rect 168648 540083 168687 540285
rect 168721 540285 168727 540571
rect 168777 540537 168783 540885
rect 168817 540635 168975 541025
rect 168817 540537 168823 540635
rect 168777 540525 168823 540537
rect 168873 540571 168919 540583
rect 168873 540285 168879 540571
rect 168721 540083 168879 540285
rect 168913 540285 168919 540571
rect 168969 540537 168975 540635
rect 169009 540635 169167 541025
rect 169009 540537 169015 540635
rect 168969 540525 169015 540537
rect 169065 540571 169111 540583
rect 169065 540285 169071 540571
rect 168913 540083 169071 540285
rect 169105 540285 169111 540571
rect 169161 540537 169167 540635
rect 169201 540635 169359 541025
rect 169201 540537 169207 540635
rect 169161 540525 169207 540537
rect 169257 540571 169303 540583
rect 169257 540285 169263 540571
rect 169105 540083 169263 540285
rect 169297 540285 169303 540571
rect 169353 540537 169359 540635
rect 169393 540635 169551 541025
rect 169393 540537 169399 540635
rect 169353 540525 169399 540537
rect 169449 540571 169495 540583
rect 169449 540285 169455 540571
rect 169297 540083 169455 540285
rect 169489 540285 169495 540571
rect 169545 540537 169551 540635
rect 169585 540995 169743 541025
rect 169777 540995 169808 541025
rect 169585 540895 169688 540995
rect 169798 540895 169808 540995
rect 169585 540875 169743 540895
rect 169777 540875 169808 540895
rect 169585 540775 169688 540875
rect 169798 540775 169808 540875
rect 170003 540830 170053 541080
rect 170196 541119 170258 541125
rect 170196 541085 170208 541119
rect 170242 541085 170258 541119
rect 170196 541079 170258 541085
rect 170198 541065 170258 541079
rect 171778 540965 171978 541505
rect 172218 541125 172278 541135
rect 172518 541130 173538 541155
rect 172518 541126 173753 541130
rect 172178 541119 172318 541125
rect 172178 541085 172228 541119
rect 172262 541085 172318 541119
rect 172518 541095 172531 541126
rect 172519 541092 172531 541095
rect 172565 541095 172723 541126
rect 172565 541092 172577 541095
rect 172519 541086 172577 541092
rect 172711 541092 172723 541095
rect 172757 541095 172915 541126
rect 172757 541092 172769 541095
rect 172711 541086 172769 541092
rect 172903 541092 172915 541095
rect 172949 541095 173107 541126
rect 172949 541092 172961 541095
rect 172903 541086 172961 541092
rect 173095 541092 173107 541095
rect 173141 541095 173299 541126
rect 173141 541092 173153 541095
rect 173095 541086 173153 541092
rect 173287 541092 173299 541095
rect 173333 541095 173491 541126
rect 173333 541092 173345 541095
rect 173287 541086 173345 541092
rect 173479 541092 173491 541095
rect 173525 541092 173753 541126
rect 173479 541086 173753 541092
rect 172178 541018 172318 541085
rect 173523 541080 173753 541086
rect 172178 540965 172184 541018
rect 170478 540830 171248 540895
rect 171778 540885 172184 540965
rect 171778 540835 171978 540885
rect 169585 540755 169743 540775
rect 169777 540755 169808 540775
rect 169585 540655 169688 540755
rect 169798 540655 169808 540755
rect 169585 540635 169743 540655
rect 169585 540537 169591 540635
rect 169545 540525 169591 540537
rect 169641 540571 169687 540583
rect 169641 540285 169647 540571
rect 169489 540083 169647 540285
rect 169681 540285 169687 540571
rect 169737 540537 169743 540635
rect 169777 540635 169808 540655
rect 169998 540780 171248 540830
rect 169777 540537 169783 540635
rect 169737 540525 169783 540537
rect 169833 540571 169879 540583
rect 169833 540285 169839 540571
rect 169681 540083 169839 540285
rect 169873 540083 169879 540571
rect 169998 540335 170048 540780
rect 170478 540695 171248 540780
rect 170158 540564 170204 540576
rect 169998 540325 170058 540335
rect 169996 540319 170058 540325
rect 169996 540285 170008 540319
rect 170042 540285 170058 540319
rect 169996 540279 170058 540285
rect 169998 540275 170058 540279
rect 169958 540235 170004 540247
rect 169958 540155 169964 540235
rect 168648 540075 169879 540083
rect 168648 540071 168727 540075
rect 168873 540071 168919 540075
rect 169065 540071 169111 540075
rect 169257 540071 169303 540075
rect 169449 540071 169495 540075
rect 169641 540071 169687 540075
rect 169833 540071 169879 540075
rect 168648 540065 168718 540071
rect 168508 540009 168578 540025
rect 168508 539975 168528 540009
rect 168562 539975 168578 540009
rect 168508 539955 168578 539975
rect 168648 539755 168678 540065
rect 169938 540059 169964 540155
rect 169998 540059 170004 540235
rect 169938 540047 170004 540059
rect 170046 540235 170092 540247
rect 170046 540059 170052 540235
rect 170086 540225 170092 540235
rect 170158 540225 170164 540564
rect 170086 540076 170164 540225
rect 170198 540235 170204 540564
rect 170246 540564 170292 540576
rect 170246 540235 170252 540564
rect 170198 540076 170252 540235
rect 170286 540235 170292 540564
rect 170468 540245 170688 540255
rect 170286 540225 170308 540235
rect 170468 540225 170488 540245
rect 170286 540215 170488 540225
rect 170286 540085 170368 540215
rect 170428 540085 170488 540215
rect 170286 540076 170488 540085
rect 170086 540075 170488 540076
rect 170086 540059 170092 540075
rect 170158 540064 170292 540075
rect 170468 540065 170488 540075
rect 170668 540065 170688 540245
rect 170046 540047 170092 540059
rect 168723 540016 168781 540022
rect 168723 540015 168735 540016
rect 168718 539982 168735 540015
rect 168769 540015 168781 540016
rect 168915 540016 168973 540022
rect 168915 540015 168927 540016
rect 168769 539982 168927 540015
rect 168961 540015 168973 540016
rect 169107 540016 169165 540022
rect 169107 540015 169119 540016
rect 168961 539982 169119 540015
rect 169153 540015 169165 540016
rect 169299 540016 169357 540022
rect 169299 540015 169311 540016
rect 169153 539982 169311 540015
rect 169345 540015 169357 540016
rect 169491 540016 169549 540022
rect 169491 540015 169503 540016
rect 169345 539982 169503 540015
rect 169537 540015 169549 540016
rect 169683 540016 169741 540022
rect 169683 540015 169695 540016
rect 169537 539982 169695 540015
rect 169729 539982 169741 540016
rect 168718 539976 169741 539982
rect 168718 539955 169738 539976
rect 168078 539655 168678 539755
rect 168078 537931 168278 539655
rect 168438 539606 168678 539655
rect 168438 539572 168512 539606
rect 168546 539572 168678 539606
rect 168438 539513 168678 539572
rect 168818 539619 169828 539625
rect 168818 539613 169841 539619
rect 168818 539579 168835 539613
rect 168869 539579 169027 539613
rect 169061 539579 169219 539613
rect 169253 539579 169411 539613
rect 169445 539579 169603 539613
rect 169637 539579 169795 539613
rect 169829 539579 169841 539613
rect 168818 539573 169841 539579
rect 168818 539565 169828 539573
rect 169938 539525 169968 540047
rect 169996 540009 170058 540015
rect 169996 539975 170008 540009
rect 170042 539975 170058 540009
rect 169996 539969 170058 539975
rect 169998 539606 170058 539969
rect 170168 540009 170288 540064
rect 170468 540055 170688 540065
rect 170168 539975 170208 540009
rect 170242 539975 170288 540009
rect 170168 539955 170288 539975
rect 169998 539572 170012 539606
rect 170046 539572 170058 539606
rect 169998 539565 170058 539572
rect 170198 539606 170278 539625
rect 170198 539572 170212 539606
rect 170246 539572 170278 539606
rect 170198 539565 170278 539572
rect 168438 539415 168468 539513
rect 168462 538537 168468 539415
rect 168502 539415 168556 539513
rect 168502 538537 168508 539415
rect 168462 538525 168508 538537
rect 168550 538537 168556 539415
rect 168590 539495 168678 539513
rect 168781 539503 168827 539515
rect 168590 539485 168748 539495
rect 168781 539485 168787 539503
rect 168590 539415 168787 539485
rect 168590 538537 168596 539415
rect 168648 539205 168787 539415
rect 168685 539049 168731 539061
rect 168685 538561 168691 539049
rect 168725 538935 168731 539049
rect 168781 539015 168787 539205
rect 168821 539485 168827 539503
rect 168973 539503 169019 539515
rect 168973 539485 168979 539503
rect 168821 539205 168979 539485
rect 168821 539015 168827 539205
rect 168781 539003 168827 539015
rect 168877 539049 168923 539061
rect 168877 538935 168883 539049
rect 168725 538561 168883 538935
rect 168917 538935 168923 539049
rect 168973 539015 168979 539205
rect 169013 539485 169019 539503
rect 169165 539503 169211 539515
rect 169165 539485 169171 539503
rect 169013 539205 169171 539485
rect 169013 539015 169019 539205
rect 168973 539003 169019 539015
rect 169069 539049 169115 539061
rect 169069 538935 169075 539049
rect 168917 538561 169075 538935
rect 169109 538935 169115 539049
rect 169165 539015 169171 539205
rect 169205 539485 169211 539503
rect 169357 539503 169403 539515
rect 169357 539485 169363 539503
rect 169205 539205 169363 539485
rect 169205 539015 169211 539205
rect 169165 539003 169211 539015
rect 169261 539049 169307 539061
rect 169261 538935 169267 539049
rect 169109 538561 169267 538935
rect 169301 538935 169307 539049
rect 169357 539015 169363 539205
rect 169397 539485 169403 539503
rect 169549 539503 169595 539515
rect 169549 539485 169555 539503
rect 169397 539205 169555 539485
rect 169397 539015 169403 539205
rect 169357 539003 169403 539015
rect 169453 539049 169499 539061
rect 169453 538935 169459 539049
rect 169301 538561 169459 538935
rect 169493 538935 169499 539049
rect 169549 539015 169555 539205
rect 169589 539485 169595 539503
rect 169741 539503 169787 539515
rect 169741 539485 169747 539503
rect 169589 539205 169747 539485
rect 169589 539015 169595 539205
rect 169549 539003 169595 539015
rect 169645 539049 169691 539061
rect 169645 538935 169651 539049
rect 169493 538561 169651 538935
rect 169685 538935 169691 539049
rect 169741 539015 169747 539205
rect 169781 539485 169787 539503
rect 169938 539513 170008 539525
rect 169781 539205 169798 539485
rect 169938 539375 169968 539513
rect 169781 539015 169787 539205
rect 169741 539003 169787 539015
rect 169837 539049 169883 539061
rect 169837 538935 169843 539049
rect 169685 538805 169843 538935
rect 169685 538705 169698 538805
rect 169838 538705 169843 538805
rect 169685 538561 169843 538705
rect 169877 538561 169883 539049
rect 169962 539035 169968 539375
rect 168685 538555 169883 538561
rect 168685 538549 168731 538555
rect 168877 538549 168923 538555
rect 169069 538549 169115 538555
rect 169261 538549 169307 538555
rect 169453 538549 169499 538555
rect 169645 538549 169691 538555
rect 169837 538549 169883 538555
rect 169928 538937 169968 539035
rect 170002 538937 170008 539513
rect 169928 538925 170008 538937
rect 170050 539513 170096 539525
rect 170050 538937 170056 539513
rect 170090 539505 170096 539513
rect 170090 539275 170208 539505
rect 170468 539305 170688 539315
rect 170468 539275 170488 539305
rect 170090 539265 170488 539275
rect 170090 539175 170368 539265
rect 170418 539175 170488 539265
rect 170090 539165 170488 539175
rect 170090 539042 170208 539165
rect 170468 539125 170488 539165
rect 170668 539125 170688 539305
rect 170468 539115 170688 539125
rect 170090 538937 170168 539042
rect 170050 538935 170168 538937
rect 170050 538925 170096 538935
rect 168550 538525 168596 538537
rect 168727 538485 168785 538491
rect 168919 538485 168977 538491
rect 169111 538485 169169 538491
rect 169303 538485 169361 538491
rect 169495 538485 169553 538491
rect 169687 538485 169745 538491
rect 169928 538485 169968 538925
rect 169998 538878 170058 538885
rect 169998 538844 170012 538878
rect 170046 538844 170058 538878
rect 169998 538825 170058 538844
rect 170162 538575 170168 538935
rect 168498 538478 168558 538485
rect 168498 538444 168512 538478
rect 168546 538444 168558 538478
rect 168498 538425 168558 538444
rect 168718 538451 168739 538485
rect 168773 538451 168931 538485
rect 168965 538451 169123 538485
rect 169157 538451 169315 538485
rect 169349 538451 169507 538485
rect 169541 538451 169699 538485
rect 169733 538451 169968 538485
rect 168718 538425 169968 538451
rect 170158 538554 170168 538575
rect 170202 538575 170208 539042
rect 170250 539042 170296 539054
rect 170250 538575 170256 539042
rect 170202 538554 170256 538575
rect 170290 538554 170296 539042
rect 170158 538542 170296 538554
rect 170158 538478 170278 538542
rect 170158 538445 170212 538478
rect 170198 538444 170212 538445
rect 170246 538445 170278 538478
rect 170246 538444 170258 538445
rect 170198 538425 170258 538444
rect 168438 537943 168768 537945
rect 169068 537943 169913 537945
rect 168078 537815 168104 537931
rect 168098 537534 168104 537815
rect 168142 537815 168278 537931
rect 168416 537931 168784 537943
rect 168142 537534 168148 537815
rect 168098 537522 168148 537534
rect 168416 537534 168422 537931
rect 168460 537585 168740 537931
rect 168460 537534 168466 537585
rect 168416 537522 168466 537534
rect 168734 537534 168740 537585
rect 168778 537534 168784 537931
rect 168734 537522 168784 537534
rect 169052 537931 169913 537943
rect 169052 537534 169058 537931
rect 169096 537535 169913 537931
rect 169096 537534 169102 537535
rect 169052 537522 169102 537534
rect 168098 536416 168148 536428
rect 168098 536019 168104 536416
rect 168142 536405 168148 536416
rect 168416 536416 168466 536428
rect 168416 536405 168422 536416
rect 168142 536045 168422 536405
rect 168142 536019 168148 536045
rect 168098 536007 168148 536019
rect 168416 536019 168422 536045
rect 168460 536019 168466 536416
rect 168416 536007 168466 536019
rect 168734 536425 168784 536428
rect 169052 536425 169102 536428
rect 168734 536416 169102 536425
rect 168734 536019 168740 536416
rect 168778 536065 169058 536416
rect 168778 536019 168784 536065
rect 168734 536007 168784 536019
rect 169052 536019 169058 536065
rect 169096 536019 169102 536416
rect 169052 536007 169102 536019
rect 169503 536255 169913 537535
rect 169503 535975 169568 536255
rect 169868 535975 169913 536255
rect 169503 535910 169913 535975
rect 171048 533505 171248 540695
rect 172178 540530 172184 540885
rect 172218 540885 172272 541018
rect 172218 540530 172224 540885
rect 172178 540518 172224 540530
rect 172266 540530 172272 540885
rect 172306 540965 172318 541018
rect 172477 541025 172523 541037
rect 172669 541025 172715 541037
rect 172861 541025 172907 541037
rect 173053 541025 173099 541037
rect 173245 541025 173291 541037
rect 173437 541025 173483 541037
rect 172477 540965 172483 541025
rect 172306 540885 172483 540965
rect 172306 540530 172312 540885
rect 172266 540518 172312 540530
rect 172381 540571 172427 540583
rect 172381 540285 172387 540571
rect 172348 540083 172387 540285
rect 172421 540285 172427 540571
rect 172477 540537 172483 540885
rect 172517 540635 172675 541025
rect 172517 540537 172523 540635
rect 172477 540525 172523 540537
rect 172573 540571 172619 540583
rect 172573 540285 172579 540571
rect 172421 540083 172579 540285
rect 172613 540285 172619 540571
rect 172669 540537 172675 540635
rect 172709 540635 172867 541025
rect 172709 540537 172715 540635
rect 172669 540525 172715 540537
rect 172765 540571 172811 540583
rect 172765 540285 172771 540571
rect 172613 540083 172771 540285
rect 172805 540285 172811 540571
rect 172861 540537 172867 540635
rect 172901 540635 173059 541025
rect 172901 540537 172907 540635
rect 172861 540525 172907 540537
rect 172957 540571 173003 540583
rect 172957 540285 172963 540571
rect 172805 540083 172963 540285
rect 172997 540285 173003 540571
rect 173053 540537 173059 540635
rect 173093 540635 173251 541025
rect 173093 540537 173099 540635
rect 173053 540525 173099 540537
rect 173149 540571 173195 540583
rect 173149 540285 173155 540571
rect 172997 540083 173155 540285
rect 173189 540285 173195 540571
rect 173245 540537 173251 540635
rect 173285 540995 173443 541025
rect 173477 540995 173508 541025
rect 173285 540895 173388 540995
rect 173498 540895 173508 540995
rect 173285 540875 173443 540895
rect 173477 540875 173508 540895
rect 173285 540775 173388 540875
rect 173498 540775 173508 540875
rect 173703 540830 173753 541080
rect 173896 541119 173958 541125
rect 173896 541085 173908 541119
rect 173942 541085 173958 541119
rect 173896 541079 173958 541085
rect 173898 541065 173958 541079
rect 175278 540965 175478 541505
rect 175718 541125 175778 541135
rect 176018 541130 177038 541155
rect 176018 541126 177253 541130
rect 175678 541119 175818 541125
rect 175678 541085 175728 541119
rect 175762 541085 175818 541119
rect 176018 541095 176031 541126
rect 176019 541092 176031 541095
rect 176065 541095 176223 541126
rect 176065 541092 176077 541095
rect 176019 541086 176077 541092
rect 176211 541092 176223 541095
rect 176257 541095 176415 541126
rect 176257 541092 176269 541095
rect 176211 541086 176269 541092
rect 176403 541092 176415 541095
rect 176449 541095 176607 541126
rect 176449 541092 176461 541095
rect 176403 541086 176461 541092
rect 176595 541092 176607 541095
rect 176641 541095 176799 541126
rect 176641 541092 176653 541095
rect 176595 541086 176653 541092
rect 176787 541092 176799 541095
rect 176833 541095 176991 541126
rect 176833 541092 176845 541095
rect 176787 541086 176845 541092
rect 176979 541092 176991 541095
rect 177025 541092 177253 541126
rect 176979 541086 177253 541092
rect 175678 541018 175818 541085
rect 177023 541080 177253 541086
rect 175678 540965 175684 541018
rect 174178 540830 174878 540895
rect 175278 540885 175684 540965
rect 175278 540835 175478 540885
rect 173285 540755 173443 540775
rect 173477 540755 173508 540775
rect 173285 540655 173388 540755
rect 173498 540655 173508 540755
rect 173285 540635 173443 540655
rect 173285 540537 173291 540635
rect 173245 540525 173291 540537
rect 173341 540571 173387 540583
rect 173341 540285 173347 540571
rect 173189 540083 173347 540285
rect 173381 540285 173387 540571
rect 173437 540537 173443 540635
rect 173477 540635 173508 540655
rect 173698 540780 174878 540830
rect 173477 540537 173483 540635
rect 173437 540525 173483 540537
rect 173533 540571 173579 540583
rect 173533 540285 173539 540571
rect 173381 540083 173539 540285
rect 173573 540083 173579 540571
rect 173698 540335 173748 540780
rect 174178 540695 174878 540780
rect 173858 540564 173904 540576
rect 173698 540325 173758 540335
rect 173696 540319 173758 540325
rect 173696 540285 173708 540319
rect 173742 540285 173758 540319
rect 173696 540279 173758 540285
rect 173698 540275 173758 540279
rect 173658 540235 173704 540247
rect 173658 540155 173664 540235
rect 172348 540075 173579 540083
rect 172348 540071 172427 540075
rect 172573 540071 172619 540075
rect 172765 540071 172811 540075
rect 172957 540071 173003 540075
rect 173149 540071 173195 540075
rect 173341 540071 173387 540075
rect 173533 540071 173579 540075
rect 172348 540065 172418 540071
rect 172208 540009 172278 540025
rect 172208 539975 172228 540009
rect 172262 539975 172278 540009
rect 172208 539955 172278 539975
rect 172348 539755 172378 540065
rect 173638 540059 173664 540155
rect 173698 540059 173704 540235
rect 173638 540047 173704 540059
rect 173746 540235 173792 540247
rect 173746 540059 173752 540235
rect 173786 540225 173792 540235
rect 173858 540225 173864 540564
rect 173786 540076 173864 540225
rect 173898 540235 173904 540564
rect 173946 540564 173992 540576
rect 173946 540235 173952 540564
rect 173898 540076 173952 540235
rect 173986 540235 173992 540564
rect 174178 540255 174378 540265
rect 173986 540225 174008 540235
rect 174168 540225 174188 540255
rect 173986 540215 174188 540225
rect 173986 540085 174068 540215
rect 174128 540085 174188 540215
rect 173986 540076 174188 540085
rect 173786 540075 174188 540076
rect 174368 540075 174388 540255
rect 173786 540059 173792 540075
rect 173858 540064 173992 540075
rect 173746 540047 173792 540059
rect 172423 540016 172481 540022
rect 172423 540015 172435 540016
rect 172418 539982 172435 540015
rect 172469 540015 172481 540016
rect 172615 540016 172673 540022
rect 172615 540015 172627 540016
rect 172469 539982 172627 540015
rect 172661 540015 172673 540016
rect 172807 540016 172865 540022
rect 172807 540015 172819 540016
rect 172661 539982 172819 540015
rect 172853 540015 172865 540016
rect 172999 540016 173057 540022
rect 172999 540015 173011 540016
rect 172853 539982 173011 540015
rect 173045 540015 173057 540016
rect 173191 540016 173249 540022
rect 173191 540015 173203 540016
rect 173045 539982 173203 540015
rect 173237 540015 173249 540016
rect 173383 540016 173441 540022
rect 173383 540015 173395 540016
rect 173237 539982 173395 540015
rect 173429 539982 173441 540016
rect 172418 539976 173441 539982
rect 172418 539955 173438 539976
rect 171778 539655 172378 539755
rect 171778 537931 171978 539655
rect 172138 539606 172378 539655
rect 172138 539572 172212 539606
rect 172246 539572 172378 539606
rect 172138 539513 172378 539572
rect 172518 539619 173528 539625
rect 172518 539613 173541 539619
rect 172518 539579 172535 539613
rect 172569 539579 172727 539613
rect 172761 539579 172919 539613
rect 172953 539579 173111 539613
rect 173145 539579 173303 539613
rect 173337 539579 173495 539613
rect 173529 539579 173541 539613
rect 172518 539573 173541 539579
rect 172518 539565 173528 539573
rect 173638 539525 173668 540047
rect 173696 540009 173758 540015
rect 173696 539975 173708 540009
rect 173742 539975 173758 540009
rect 173696 539969 173758 539975
rect 173698 539606 173758 539969
rect 173868 540009 173988 540064
rect 174168 540055 174388 540075
rect 173868 539975 173908 540009
rect 173942 539975 173988 540009
rect 173868 539955 173988 539975
rect 173698 539572 173712 539606
rect 173746 539572 173758 539606
rect 173698 539565 173758 539572
rect 173898 539606 173978 539625
rect 173898 539572 173912 539606
rect 173946 539572 173978 539606
rect 173898 539565 173978 539572
rect 172138 539415 172168 539513
rect 172162 538537 172168 539415
rect 172202 539415 172256 539513
rect 172202 538537 172208 539415
rect 172162 538525 172208 538537
rect 172250 538537 172256 539415
rect 172290 539495 172378 539513
rect 172481 539503 172527 539515
rect 172290 539485 172448 539495
rect 172481 539485 172487 539503
rect 172290 539415 172487 539485
rect 172290 538537 172296 539415
rect 172348 539205 172487 539415
rect 172385 539049 172431 539061
rect 172385 538561 172391 539049
rect 172425 538935 172431 539049
rect 172481 539015 172487 539205
rect 172521 539485 172527 539503
rect 172673 539503 172719 539515
rect 172673 539485 172679 539503
rect 172521 539205 172679 539485
rect 172521 539015 172527 539205
rect 172481 539003 172527 539015
rect 172577 539049 172623 539061
rect 172577 538935 172583 539049
rect 172425 538561 172583 538935
rect 172617 538935 172623 539049
rect 172673 539015 172679 539205
rect 172713 539485 172719 539503
rect 172865 539503 172911 539515
rect 172865 539485 172871 539503
rect 172713 539205 172871 539485
rect 172713 539015 172719 539205
rect 172673 539003 172719 539015
rect 172769 539049 172815 539061
rect 172769 538935 172775 539049
rect 172617 538561 172775 538935
rect 172809 538935 172815 539049
rect 172865 539015 172871 539205
rect 172905 539485 172911 539503
rect 173057 539503 173103 539515
rect 173057 539485 173063 539503
rect 172905 539205 173063 539485
rect 172905 539015 172911 539205
rect 172865 539003 172911 539015
rect 172961 539049 173007 539061
rect 172961 538935 172967 539049
rect 172809 538561 172967 538935
rect 173001 538935 173007 539049
rect 173057 539015 173063 539205
rect 173097 539485 173103 539503
rect 173249 539503 173295 539515
rect 173249 539485 173255 539503
rect 173097 539205 173255 539485
rect 173097 539015 173103 539205
rect 173057 539003 173103 539015
rect 173153 539049 173199 539061
rect 173153 538935 173159 539049
rect 173001 538561 173159 538935
rect 173193 538935 173199 539049
rect 173249 539015 173255 539205
rect 173289 539485 173295 539503
rect 173441 539503 173487 539515
rect 173441 539485 173447 539503
rect 173289 539205 173447 539485
rect 173289 539015 173295 539205
rect 173249 539003 173295 539015
rect 173345 539049 173391 539061
rect 173345 538935 173351 539049
rect 173193 538561 173351 538935
rect 173385 538935 173391 539049
rect 173441 539015 173447 539205
rect 173481 539485 173487 539503
rect 173638 539513 173708 539525
rect 173481 539205 173498 539485
rect 173638 539375 173668 539513
rect 173481 539015 173487 539205
rect 173441 539003 173487 539015
rect 173537 539049 173583 539061
rect 173537 538935 173543 539049
rect 173385 538805 173543 538935
rect 173385 538705 173398 538805
rect 173538 538705 173543 538805
rect 173385 538561 173543 538705
rect 173577 538561 173583 539049
rect 173662 539035 173668 539375
rect 172385 538555 173583 538561
rect 172385 538549 172431 538555
rect 172577 538549 172623 538555
rect 172769 538549 172815 538555
rect 172961 538549 173007 538555
rect 173153 538549 173199 538555
rect 173345 538549 173391 538555
rect 173537 538549 173583 538555
rect 173628 538937 173668 539035
rect 173702 538937 173708 539513
rect 173628 538925 173708 538937
rect 173750 539513 173796 539525
rect 173750 538937 173756 539513
rect 173790 539505 173796 539513
rect 173790 539275 173908 539505
rect 174168 539305 174388 539315
rect 174168 539275 174188 539305
rect 173790 539265 174188 539275
rect 173790 539175 174068 539265
rect 174118 539175 174188 539265
rect 173790 539165 174188 539175
rect 173790 539042 173908 539165
rect 174168 539125 174188 539165
rect 174368 539125 174388 539305
rect 174168 539115 174388 539125
rect 173790 538937 173868 539042
rect 173750 538935 173868 538937
rect 173750 538925 173796 538935
rect 172250 538525 172296 538537
rect 172427 538485 172485 538491
rect 172619 538485 172677 538491
rect 172811 538485 172869 538491
rect 173003 538485 173061 538491
rect 173195 538485 173253 538491
rect 173387 538485 173445 538491
rect 173628 538485 173668 538925
rect 173698 538878 173758 538885
rect 173698 538844 173712 538878
rect 173746 538844 173758 538878
rect 173698 538825 173758 538844
rect 173862 538575 173868 538935
rect 172198 538478 172258 538485
rect 172198 538444 172212 538478
rect 172246 538444 172258 538478
rect 172198 538425 172258 538444
rect 172418 538451 172439 538485
rect 172473 538451 172631 538485
rect 172665 538451 172823 538485
rect 172857 538451 173015 538485
rect 173049 538451 173207 538485
rect 173241 538451 173399 538485
rect 173433 538451 173668 538485
rect 172418 538425 173668 538451
rect 173858 538554 173868 538575
rect 173902 538575 173908 539042
rect 173950 539042 173996 539054
rect 173950 538575 173956 539042
rect 173902 538554 173956 538575
rect 173990 538554 173996 539042
rect 173858 538542 173996 538554
rect 173858 538478 173978 538542
rect 173858 538445 173912 538478
rect 173898 538444 173912 538445
rect 173946 538445 173978 538478
rect 173946 538444 173958 538445
rect 173898 538425 173958 538444
rect 171778 537815 171840 537931
rect 171834 537534 171840 537815
rect 171878 537815 171978 537931
rect 172152 537935 172202 537943
rect 172152 537931 172978 537935
rect 171878 537534 171884 537815
rect 171834 537522 171884 537534
rect 172152 537534 172158 537931
rect 172196 537534 172978 537931
rect 172152 537522 172978 537534
rect 172168 537515 172978 537522
rect 171834 536416 171884 536428
rect 171834 536019 171840 536416
rect 171878 536405 171884 536416
rect 172152 536416 172202 536428
rect 172152 536405 172158 536416
rect 171878 536045 172158 536405
rect 171878 536019 171884 536045
rect 171834 536007 171884 536019
rect 172152 536019 172158 536045
rect 172196 536019 172202 536416
rect 172152 536007 172202 536019
rect 172558 536265 172978 537515
rect 172558 535975 172608 536265
rect 172938 535975 172978 536265
rect 172558 535915 172978 535975
rect 174678 533505 174878 540695
rect 175678 540530 175684 540885
rect 175718 540885 175772 541018
rect 175718 540530 175724 540885
rect 175678 540518 175724 540530
rect 175766 540530 175772 540885
rect 175806 540965 175818 541018
rect 175977 541025 176023 541037
rect 176169 541025 176215 541037
rect 176361 541025 176407 541037
rect 176553 541025 176599 541037
rect 176745 541025 176791 541037
rect 176937 541025 176983 541037
rect 175977 540965 175983 541025
rect 175806 540885 175983 540965
rect 175806 540530 175812 540885
rect 175766 540518 175812 540530
rect 175881 540571 175927 540583
rect 175881 540285 175887 540571
rect 175848 540083 175887 540285
rect 175921 540285 175927 540571
rect 175977 540537 175983 540885
rect 176017 540635 176175 541025
rect 176017 540537 176023 540635
rect 175977 540525 176023 540537
rect 176073 540571 176119 540583
rect 176073 540285 176079 540571
rect 175921 540083 176079 540285
rect 176113 540285 176119 540571
rect 176169 540537 176175 540635
rect 176209 540635 176367 541025
rect 176209 540537 176215 540635
rect 176169 540525 176215 540537
rect 176265 540571 176311 540583
rect 176265 540285 176271 540571
rect 176113 540083 176271 540285
rect 176305 540285 176311 540571
rect 176361 540537 176367 540635
rect 176401 540635 176559 541025
rect 176401 540537 176407 540635
rect 176361 540525 176407 540537
rect 176457 540571 176503 540583
rect 176457 540285 176463 540571
rect 176305 540083 176463 540285
rect 176497 540285 176503 540571
rect 176553 540537 176559 540635
rect 176593 540635 176751 541025
rect 176593 540537 176599 540635
rect 176553 540525 176599 540537
rect 176649 540571 176695 540583
rect 176649 540285 176655 540571
rect 176497 540083 176655 540285
rect 176689 540285 176695 540571
rect 176745 540537 176751 540635
rect 176785 540995 176943 541025
rect 176977 540995 177008 541025
rect 176785 540895 176888 540995
rect 176998 540895 177008 540995
rect 176785 540875 176943 540895
rect 176977 540875 177008 540895
rect 176785 540775 176888 540875
rect 176998 540775 177008 540875
rect 177203 540830 177253 541080
rect 177396 541119 177458 541125
rect 177396 541085 177408 541119
rect 177442 541085 177458 541119
rect 177396 541079 177458 541085
rect 177398 541065 177458 541079
rect 178878 540965 179078 541505
rect 179318 541125 179378 541135
rect 179618 541130 180638 541155
rect 179618 541126 180853 541130
rect 179278 541119 179418 541125
rect 179278 541085 179328 541119
rect 179362 541085 179418 541119
rect 179618 541095 179631 541126
rect 179619 541092 179631 541095
rect 179665 541095 179823 541126
rect 179665 541092 179677 541095
rect 179619 541086 179677 541092
rect 179811 541092 179823 541095
rect 179857 541095 180015 541126
rect 179857 541092 179869 541095
rect 179811 541086 179869 541092
rect 180003 541092 180015 541095
rect 180049 541095 180207 541126
rect 180049 541092 180061 541095
rect 180003 541086 180061 541092
rect 180195 541092 180207 541095
rect 180241 541095 180399 541126
rect 180241 541092 180253 541095
rect 180195 541086 180253 541092
rect 180387 541092 180399 541095
rect 180433 541095 180591 541126
rect 180433 541092 180445 541095
rect 180387 541086 180445 541092
rect 180579 541092 180591 541095
rect 180625 541092 180853 541126
rect 180579 541086 180853 541092
rect 179278 541018 179418 541085
rect 180623 541080 180853 541086
rect 179278 540965 179284 541018
rect 177678 540830 178418 540895
rect 178878 540885 179284 540965
rect 178878 540835 179078 540885
rect 176785 540755 176943 540775
rect 176977 540755 177008 540775
rect 176785 540655 176888 540755
rect 176998 540655 177008 540755
rect 176785 540635 176943 540655
rect 176785 540537 176791 540635
rect 176745 540525 176791 540537
rect 176841 540571 176887 540583
rect 176841 540285 176847 540571
rect 176689 540083 176847 540285
rect 176881 540285 176887 540571
rect 176937 540537 176943 540635
rect 176977 540635 177008 540655
rect 177198 540780 178418 540830
rect 176977 540537 176983 540635
rect 176937 540525 176983 540537
rect 177033 540571 177079 540583
rect 177033 540285 177039 540571
rect 176881 540083 177039 540285
rect 177073 540083 177079 540571
rect 177198 540335 177248 540780
rect 177678 540695 178418 540780
rect 177358 540564 177404 540576
rect 177198 540325 177258 540335
rect 177196 540319 177258 540325
rect 177196 540285 177208 540319
rect 177242 540285 177258 540319
rect 177196 540279 177258 540285
rect 177198 540275 177258 540279
rect 177158 540235 177204 540247
rect 177158 540155 177164 540235
rect 175848 540075 177079 540083
rect 175848 540071 175927 540075
rect 176073 540071 176119 540075
rect 176265 540071 176311 540075
rect 176457 540071 176503 540075
rect 176649 540071 176695 540075
rect 176841 540071 176887 540075
rect 177033 540071 177079 540075
rect 175848 540065 175918 540071
rect 175708 540009 175778 540025
rect 175708 539975 175728 540009
rect 175762 539975 175778 540009
rect 175708 539955 175778 539975
rect 175848 539755 175878 540065
rect 177138 540059 177164 540155
rect 177198 540059 177204 540235
rect 177138 540047 177204 540059
rect 177246 540235 177292 540247
rect 177246 540059 177252 540235
rect 177286 540225 177292 540235
rect 177358 540225 177364 540564
rect 177286 540076 177364 540225
rect 177398 540235 177404 540564
rect 177446 540564 177492 540576
rect 177446 540235 177452 540564
rect 177398 540076 177452 540235
rect 177486 540235 177492 540564
rect 177668 540245 177888 540255
rect 177486 540225 177508 540235
rect 177668 540225 177698 540245
rect 177486 540215 177698 540225
rect 177486 540085 177568 540215
rect 177628 540085 177698 540215
rect 177486 540076 177698 540085
rect 177286 540075 177698 540076
rect 177286 540059 177292 540075
rect 177358 540064 177492 540075
rect 177668 540065 177698 540075
rect 177878 540065 177888 540245
rect 177246 540047 177292 540059
rect 175923 540016 175981 540022
rect 175923 540015 175935 540016
rect 175918 539982 175935 540015
rect 175969 540015 175981 540016
rect 176115 540016 176173 540022
rect 176115 540015 176127 540016
rect 175969 539982 176127 540015
rect 176161 540015 176173 540016
rect 176307 540016 176365 540022
rect 176307 540015 176319 540016
rect 176161 539982 176319 540015
rect 176353 540015 176365 540016
rect 176499 540016 176557 540022
rect 176499 540015 176511 540016
rect 176353 539982 176511 540015
rect 176545 540015 176557 540016
rect 176691 540016 176749 540022
rect 176691 540015 176703 540016
rect 176545 539982 176703 540015
rect 176737 540015 176749 540016
rect 176883 540016 176941 540022
rect 176883 540015 176895 540016
rect 176737 539982 176895 540015
rect 176929 539982 176941 540016
rect 175918 539976 176941 539982
rect 175918 539955 176938 539976
rect 175278 539655 175878 539755
rect 175278 537931 175478 539655
rect 175638 539606 175878 539655
rect 175638 539572 175712 539606
rect 175746 539572 175878 539606
rect 175638 539513 175878 539572
rect 176018 539619 177028 539625
rect 176018 539613 177041 539619
rect 176018 539579 176035 539613
rect 176069 539579 176227 539613
rect 176261 539579 176419 539613
rect 176453 539579 176611 539613
rect 176645 539579 176803 539613
rect 176837 539579 176995 539613
rect 177029 539579 177041 539613
rect 176018 539573 177041 539579
rect 176018 539565 177028 539573
rect 177138 539525 177168 540047
rect 177196 540009 177258 540015
rect 177196 539975 177208 540009
rect 177242 539975 177258 540009
rect 177196 539969 177258 539975
rect 177198 539606 177258 539969
rect 177368 540009 177488 540064
rect 177668 540055 177888 540065
rect 177368 539975 177408 540009
rect 177442 539975 177488 540009
rect 177368 539955 177488 539975
rect 177198 539572 177212 539606
rect 177246 539572 177258 539606
rect 177198 539565 177258 539572
rect 177398 539606 177478 539625
rect 177398 539572 177412 539606
rect 177446 539572 177478 539606
rect 177398 539565 177478 539572
rect 175638 539415 175668 539513
rect 175662 538537 175668 539415
rect 175702 539415 175756 539513
rect 175702 538537 175708 539415
rect 175662 538525 175708 538537
rect 175750 538537 175756 539415
rect 175790 539495 175878 539513
rect 175981 539503 176027 539515
rect 175790 539485 175948 539495
rect 175981 539485 175987 539503
rect 175790 539415 175987 539485
rect 175790 538537 175796 539415
rect 175848 539205 175987 539415
rect 175885 539049 175931 539061
rect 175885 538561 175891 539049
rect 175925 538935 175931 539049
rect 175981 539015 175987 539205
rect 176021 539485 176027 539503
rect 176173 539503 176219 539515
rect 176173 539485 176179 539503
rect 176021 539205 176179 539485
rect 176021 539015 176027 539205
rect 175981 539003 176027 539015
rect 176077 539049 176123 539061
rect 176077 538935 176083 539049
rect 175925 538561 176083 538935
rect 176117 538935 176123 539049
rect 176173 539015 176179 539205
rect 176213 539485 176219 539503
rect 176365 539503 176411 539515
rect 176365 539485 176371 539503
rect 176213 539205 176371 539485
rect 176213 539015 176219 539205
rect 176173 539003 176219 539015
rect 176269 539049 176315 539061
rect 176269 538935 176275 539049
rect 176117 538561 176275 538935
rect 176309 538935 176315 539049
rect 176365 539015 176371 539205
rect 176405 539485 176411 539503
rect 176557 539503 176603 539515
rect 176557 539485 176563 539503
rect 176405 539205 176563 539485
rect 176405 539015 176411 539205
rect 176365 539003 176411 539015
rect 176461 539049 176507 539061
rect 176461 538935 176467 539049
rect 176309 538561 176467 538935
rect 176501 538935 176507 539049
rect 176557 539015 176563 539205
rect 176597 539485 176603 539503
rect 176749 539503 176795 539515
rect 176749 539485 176755 539503
rect 176597 539205 176755 539485
rect 176597 539015 176603 539205
rect 176557 539003 176603 539015
rect 176653 539049 176699 539061
rect 176653 538935 176659 539049
rect 176501 538561 176659 538935
rect 176693 538935 176699 539049
rect 176749 539015 176755 539205
rect 176789 539485 176795 539503
rect 176941 539503 176987 539515
rect 176941 539485 176947 539503
rect 176789 539205 176947 539485
rect 176789 539015 176795 539205
rect 176749 539003 176795 539015
rect 176845 539049 176891 539061
rect 176845 538935 176851 539049
rect 176693 538561 176851 538935
rect 176885 538935 176891 539049
rect 176941 539015 176947 539205
rect 176981 539485 176987 539503
rect 177138 539513 177208 539525
rect 176981 539205 176998 539485
rect 177138 539375 177168 539513
rect 176981 539015 176987 539205
rect 176941 539003 176987 539015
rect 177037 539049 177083 539061
rect 177037 538935 177043 539049
rect 176885 538805 177043 538935
rect 176885 538705 176898 538805
rect 177038 538705 177043 538805
rect 176885 538561 177043 538705
rect 177077 538561 177083 539049
rect 177162 539035 177168 539375
rect 175885 538555 177083 538561
rect 175885 538549 175931 538555
rect 176077 538549 176123 538555
rect 176269 538549 176315 538555
rect 176461 538549 176507 538555
rect 176653 538549 176699 538555
rect 176845 538549 176891 538555
rect 177037 538549 177083 538555
rect 177128 538937 177168 539035
rect 177202 538937 177208 539513
rect 177128 538925 177208 538937
rect 177250 539513 177296 539525
rect 177250 538937 177256 539513
rect 177290 539505 177296 539513
rect 177290 539275 177408 539505
rect 177668 539305 177888 539315
rect 177668 539275 177688 539305
rect 177290 539265 177688 539275
rect 177290 539175 177568 539265
rect 177618 539175 177688 539265
rect 177290 539165 177688 539175
rect 177290 539042 177408 539165
rect 177668 539125 177688 539165
rect 177868 539125 177888 539305
rect 177668 539115 177888 539125
rect 177290 538937 177368 539042
rect 177250 538935 177368 538937
rect 177250 538925 177296 538935
rect 175750 538525 175796 538537
rect 175927 538485 175985 538491
rect 176119 538485 176177 538491
rect 176311 538485 176369 538491
rect 176503 538485 176561 538491
rect 176695 538485 176753 538491
rect 176887 538485 176945 538491
rect 177128 538485 177168 538925
rect 177198 538878 177258 538885
rect 177198 538844 177212 538878
rect 177246 538844 177258 538878
rect 177198 538825 177258 538844
rect 177362 538575 177368 538935
rect 175698 538478 175758 538485
rect 175698 538444 175712 538478
rect 175746 538444 175758 538478
rect 175698 538425 175758 538444
rect 175918 538451 175939 538485
rect 175973 538451 176131 538485
rect 176165 538451 176323 538485
rect 176357 538451 176515 538485
rect 176549 538451 176707 538485
rect 176741 538451 176899 538485
rect 176933 538451 177168 538485
rect 175918 538425 177168 538451
rect 177358 538554 177368 538575
rect 177402 538575 177408 539042
rect 177450 539042 177496 539054
rect 177450 538575 177456 539042
rect 177402 538554 177456 538575
rect 177490 538554 177496 539042
rect 177358 538542 177496 538554
rect 177358 538478 177478 538542
rect 177358 538445 177412 538478
rect 177398 538444 177412 538445
rect 177446 538445 177478 538478
rect 177446 538444 177458 538445
rect 177398 538425 177458 538444
rect 175278 537815 175358 537931
rect 175352 537534 175358 537815
rect 175396 537815 175478 537931
rect 175396 537534 175402 537815
rect 175352 537522 175402 537534
rect 175352 536416 175402 536428
rect 175352 536295 175358 536416
rect 175228 536255 175358 536295
rect 175396 536295 175402 536416
rect 175396 536255 175578 536295
rect 175228 535945 175278 536255
rect 175498 535945 175578 536255
rect 175228 535895 175578 535945
rect 171048 533305 173928 533505
rect 174678 533305 176728 533505
rect 173728 532755 173928 533305
rect 167518 532735 172528 532755
rect 167518 532565 172358 532735
rect 172488 532565 172528 532735
rect 167518 532555 172528 532565
rect 173728 532745 174728 532755
rect 173728 532575 174488 532745
rect 174618 532575 174728 532745
rect 173728 532555 174728 532575
rect 176528 532735 176728 533305
rect 176528 532565 176578 532735
rect 176708 532565 176728 532735
rect 176528 532455 176728 532565
rect 178218 532755 178418 540695
rect 179278 540530 179284 540885
rect 179318 540885 179372 541018
rect 179318 540530 179324 540885
rect 179278 540518 179324 540530
rect 179366 540530 179372 540885
rect 179406 540965 179418 541018
rect 179577 541025 179623 541037
rect 179769 541025 179815 541037
rect 179961 541025 180007 541037
rect 180153 541025 180199 541037
rect 180345 541025 180391 541037
rect 180537 541025 180583 541037
rect 179577 540965 179583 541025
rect 179406 540885 179583 540965
rect 179406 540530 179412 540885
rect 179366 540518 179412 540530
rect 179481 540571 179527 540583
rect 179481 540285 179487 540571
rect 179448 540083 179487 540285
rect 179521 540285 179527 540571
rect 179577 540537 179583 540885
rect 179617 540635 179775 541025
rect 179617 540537 179623 540635
rect 179577 540525 179623 540537
rect 179673 540571 179719 540583
rect 179673 540285 179679 540571
rect 179521 540083 179679 540285
rect 179713 540285 179719 540571
rect 179769 540537 179775 540635
rect 179809 540635 179967 541025
rect 179809 540537 179815 540635
rect 179769 540525 179815 540537
rect 179865 540571 179911 540583
rect 179865 540285 179871 540571
rect 179713 540083 179871 540285
rect 179905 540285 179911 540571
rect 179961 540537 179967 540635
rect 180001 540635 180159 541025
rect 180001 540537 180007 540635
rect 179961 540525 180007 540537
rect 180057 540571 180103 540583
rect 180057 540285 180063 540571
rect 179905 540083 180063 540285
rect 180097 540285 180103 540571
rect 180153 540537 180159 540635
rect 180193 540635 180351 541025
rect 180193 540537 180199 540635
rect 180153 540525 180199 540537
rect 180249 540571 180295 540583
rect 180249 540285 180255 540571
rect 180097 540083 180255 540285
rect 180289 540285 180295 540571
rect 180345 540537 180351 540635
rect 180385 540995 180543 541025
rect 180577 540995 180608 541025
rect 180385 540895 180488 540995
rect 180598 540895 180608 540995
rect 180385 540875 180543 540895
rect 180577 540875 180608 540895
rect 180385 540775 180488 540875
rect 180598 540775 180608 540875
rect 180803 540830 180853 541080
rect 180996 541119 181058 541125
rect 180996 541085 181008 541119
rect 181042 541085 181058 541119
rect 180996 541079 181058 541085
rect 180998 541065 181058 541079
rect 182178 540965 182378 541505
rect 182618 541125 182678 541135
rect 182918 541130 183938 541155
rect 182918 541126 184153 541130
rect 182578 541119 182718 541125
rect 182578 541085 182628 541119
rect 182662 541085 182718 541119
rect 182918 541095 182931 541126
rect 182919 541092 182931 541095
rect 182965 541095 183123 541126
rect 182965 541092 182977 541095
rect 182919 541086 182977 541092
rect 183111 541092 183123 541095
rect 183157 541095 183315 541126
rect 183157 541092 183169 541095
rect 183111 541086 183169 541092
rect 183303 541092 183315 541095
rect 183349 541095 183507 541126
rect 183349 541092 183361 541095
rect 183303 541086 183361 541092
rect 183495 541092 183507 541095
rect 183541 541095 183699 541126
rect 183541 541092 183553 541095
rect 183495 541086 183553 541092
rect 183687 541092 183699 541095
rect 183733 541095 183891 541126
rect 183733 541092 183745 541095
rect 183687 541086 183745 541092
rect 183879 541092 183891 541095
rect 183925 541092 184153 541126
rect 183879 541086 184153 541092
rect 182578 541018 182718 541085
rect 183923 541080 184153 541086
rect 182578 540965 182584 541018
rect 181278 540830 181928 540895
rect 182178 540885 182584 540965
rect 182178 540835 182378 540885
rect 180385 540755 180543 540775
rect 180577 540755 180608 540775
rect 180385 540655 180488 540755
rect 180598 540655 180608 540755
rect 180385 540635 180543 540655
rect 180385 540537 180391 540635
rect 180345 540525 180391 540537
rect 180441 540571 180487 540583
rect 180441 540285 180447 540571
rect 180289 540083 180447 540285
rect 180481 540285 180487 540571
rect 180537 540537 180543 540635
rect 180577 540635 180608 540655
rect 180798 540780 181928 540830
rect 180577 540537 180583 540635
rect 180537 540525 180583 540537
rect 180633 540571 180679 540583
rect 180633 540285 180639 540571
rect 180481 540083 180639 540285
rect 180673 540083 180679 540571
rect 180798 540335 180848 540780
rect 181278 540695 181928 540780
rect 180958 540564 181004 540576
rect 180798 540325 180858 540335
rect 180796 540319 180858 540325
rect 180796 540285 180808 540319
rect 180842 540285 180858 540319
rect 180796 540279 180858 540285
rect 180798 540275 180858 540279
rect 180758 540235 180804 540247
rect 180758 540155 180764 540235
rect 179448 540075 180679 540083
rect 179448 540071 179527 540075
rect 179673 540071 179719 540075
rect 179865 540071 179911 540075
rect 180057 540071 180103 540075
rect 180249 540071 180295 540075
rect 180441 540071 180487 540075
rect 180633 540071 180679 540075
rect 179448 540065 179518 540071
rect 179308 540009 179378 540025
rect 179308 539975 179328 540009
rect 179362 539975 179378 540009
rect 179308 539955 179378 539975
rect 179448 539755 179478 540065
rect 180738 540059 180764 540155
rect 180798 540059 180804 540235
rect 180738 540047 180804 540059
rect 180846 540235 180892 540247
rect 180846 540059 180852 540235
rect 180886 540225 180892 540235
rect 180958 540225 180964 540564
rect 180886 540076 180964 540225
rect 180998 540235 181004 540564
rect 181046 540564 181092 540576
rect 181046 540235 181052 540564
rect 180998 540076 181052 540235
rect 181086 540235 181092 540564
rect 181268 540245 181488 540255
rect 181086 540225 181108 540235
rect 181268 540225 181288 540245
rect 181086 540215 181288 540225
rect 181086 540085 181168 540215
rect 181228 540085 181288 540215
rect 181086 540076 181288 540085
rect 180886 540075 181288 540076
rect 180886 540059 180892 540075
rect 180958 540064 181092 540075
rect 181268 540065 181288 540075
rect 181468 540065 181488 540245
rect 180846 540047 180892 540059
rect 179523 540016 179581 540022
rect 179523 540015 179535 540016
rect 179518 539982 179535 540015
rect 179569 540015 179581 540016
rect 179715 540016 179773 540022
rect 179715 540015 179727 540016
rect 179569 539982 179727 540015
rect 179761 540015 179773 540016
rect 179907 540016 179965 540022
rect 179907 540015 179919 540016
rect 179761 539982 179919 540015
rect 179953 540015 179965 540016
rect 180099 540016 180157 540022
rect 180099 540015 180111 540016
rect 179953 539982 180111 540015
rect 180145 540015 180157 540016
rect 180291 540016 180349 540022
rect 180291 540015 180303 540016
rect 180145 539982 180303 540015
rect 180337 540015 180349 540016
rect 180483 540016 180541 540022
rect 180483 540015 180495 540016
rect 180337 539982 180495 540015
rect 180529 539982 180541 540016
rect 179518 539976 180541 539982
rect 179518 539955 180538 539976
rect 178878 539655 179478 539755
rect 178878 537931 179078 539655
rect 179238 539606 179478 539655
rect 179238 539572 179312 539606
rect 179346 539572 179478 539606
rect 179238 539513 179478 539572
rect 179618 539619 180628 539625
rect 179618 539613 180641 539619
rect 179618 539579 179635 539613
rect 179669 539579 179827 539613
rect 179861 539579 180019 539613
rect 180053 539579 180211 539613
rect 180245 539579 180403 539613
rect 180437 539579 180595 539613
rect 180629 539579 180641 539613
rect 179618 539573 180641 539579
rect 179618 539565 180628 539573
rect 180738 539525 180768 540047
rect 180796 540009 180858 540015
rect 180796 539975 180808 540009
rect 180842 539975 180858 540009
rect 180796 539969 180858 539975
rect 180798 539606 180858 539969
rect 180968 540009 181088 540064
rect 181268 540055 181488 540065
rect 180968 539975 181008 540009
rect 181042 539975 181088 540009
rect 180968 539955 181088 539975
rect 180798 539572 180812 539606
rect 180846 539572 180858 539606
rect 180798 539565 180858 539572
rect 180998 539606 181078 539625
rect 180998 539572 181012 539606
rect 181046 539572 181078 539606
rect 180998 539565 181078 539572
rect 179238 539415 179268 539513
rect 179262 538537 179268 539415
rect 179302 539415 179356 539513
rect 179302 538537 179308 539415
rect 179262 538525 179308 538537
rect 179350 538537 179356 539415
rect 179390 539495 179478 539513
rect 179581 539503 179627 539515
rect 179390 539485 179548 539495
rect 179581 539485 179587 539503
rect 179390 539415 179587 539485
rect 179390 538537 179396 539415
rect 179448 539205 179587 539415
rect 179485 539049 179531 539061
rect 179485 538561 179491 539049
rect 179525 538935 179531 539049
rect 179581 539015 179587 539205
rect 179621 539485 179627 539503
rect 179773 539503 179819 539515
rect 179773 539485 179779 539503
rect 179621 539205 179779 539485
rect 179621 539015 179627 539205
rect 179581 539003 179627 539015
rect 179677 539049 179723 539061
rect 179677 538935 179683 539049
rect 179525 538561 179683 538935
rect 179717 538935 179723 539049
rect 179773 539015 179779 539205
rect 179813 539485 179819 539503
rect 179965 539503 180011 539515
rect 179965 539485 179971 539503
rect 179813 539205 179971 539485
rect 179813 539015 179819 539205
rect 179773 539003 179819 539015
rect 179869 539049 179915 539061
rect 179869 538935 179875 539049
rect 179717 538561 179875 538935
rect 179909 538935 179915 539049
rect 179965 539015 179971 539205
rect 180005 539485 180011 539503
rect 180157 539503 180203 539515
rect 180157 539485 180163 539503
rect 180005 539205 180163 539485
rect 180005 539015 180011 539205
rect 179965 539003 180011 539015
rect 180061 539049 180107 539061
rect 180061 538935 180067 539049
rect 179909 538561 180067 538935
rect 180101 538935 180107 539049
rect 180157 539015 180163 539205
rect 180197 539485 180203 539503
rect 180349 539503 180395 539515
rect 180349 539485 180355 539503
rect 180197 539205 180355 539485
rect 180197 539015 180203 539205
rect 180157 539003 180203 539015
rect 180253 539049 180299 539061
rect 180253 538935 180259 539049
rect 180101 538561 180259 538935
rect 180293 538935 180299 539049
rect 180349 539015 180355 539205
rect 180389 539485 180395 539503
rect 180541 539503 180587 539515
rect 180541 539485 180547 539503
rect 180389 539205 180547 539485
rect 180389 539015 180395 539205
rect 180349 539003 180395 539015
rect 180445 539049 180491 539061
rect 180445 538935 180451 539049
rect 180293 538561 180451 538935
rect 180485 538935 180491 539049
rect 180541 539015 180547 539205
rect 180581 539485 180587 539503
rect 180738 539513 180808 539525
rect 180581 539205 180598 539485
rect 180738 539375 180768 539513
rect 180581 539015 180587 539205
rect 180541 539003 180587 539015
rect 180637 539049 180683 539061
rect 180637 538935 180643 539049
rect 180485 538805 180643 538935
rect 180485 538705 180498 538805
rect 180638 538705 180643 538805
rect 180485 538561 180643 538705
rect 180677 538561 180683 539049
rect 180762 539035 180768 539375
rect 179485 538555 180683 538561
rect 179485 538549 179531 538555
rect 179677 538549 179723 538555
rect 179869 538549 179915 538555
rect 180061 538549 180107 538555
rect 180253 538549 180299 538555
rect 180445 538549 180491 538555
rect 180637 538549 180683 538555
rect 180728 538937 180768 539035
rect 180802 538937 180808 539513
rect 180728 538925 180808 538937
rect 180850 539513 180896 539525
rect 180850 538937 180856 539513
rect 180890 539505 180896 539513
rect 180890 539275 181008 539505
rect 181268 539305 181488 539315
rect 181268 539275 181288 539305
rect 180890 539265 181288 539275
rect 180890 539175 181168 539265
rect 181218 539175 181288 539265
rect 180890 539165 181288 539175
rect 180890 539042 181008 539165
rect 181268 539125 181288 539165
rect 181468 539125 181488 539305
rect 181268 539115 181488 539125
rect 180890 538937 180968 539042
rect 180850 538935 180968 538937
rect 180850 538925 180896 538935
rect 179350 538525 179396 538537
rect 179527 538485 179585 538491
rect 179719 538485 179777 538491
rect 179911 538485 179969 538491
rect 180103 538485 180161 538491
rect 180295 538485 180353 538491
rect 180487 538485 180545 538491
rect 180728 538485 180768 538925
rect 180798 538878 180858 538885
rect 180798 538844 180812 538878
rect 180846 538844 180858 538878
rect 180798 538825 180858 538844
rect 180962 538575 180968 538935
rect 179298 538478 179358 538485
rect 179298 538444 179312 538478
rect 179346 538444 179358 538478
rect 179298 538425 179358 538444
rect 179518 538451 179539 538485
rect 179573 538451 179731 538485
rect 179765 538451 179923 538485
rect 179957 538451 180115 538485
rect 180149 538451 180307 538485
rect 180341 538451 180499 538485
rect 180533 538451 180768 538485
rect 179518 538425 180768 538451
rect 180958 538554 180968 538575
rect 181002 538575 181008 539042
rect 181050 539042 181096 539054
rect 181050 538575 181056 539042
rect 181002 538554 181056 538575
rect 181090 538554 181096 539042
rect 180958 538542 181096 538554
rect 180958 538478 181078 538542
rect 180958 538445 181012 538478
rect 180998 538444 181012 538445
rect 181046 538445 181078 538478
rect 181046 538444 181058 538445
rect 180998 538425 181058 538444
rect 178878 537815 178958 537931
rect 178952 537534 178958 537815
rect 178996 537815 179078 537931
rect 178996 537534 179002 537815
rect 178952 537522 179002 537534
rect 178952 536976 179002 536988
rect 178952 536965 178958 536976
rect 178818 536579 178958 536965
rect 178996 536965 179002 536976
rect 178996 536579 179118 536965
rect 178818 536275 179118 536579
rect 178818 535965 178868 536275
rect 179068 535965 179118 536275
rect 178818 535865 179118 535965
rect 181728 533505 181928 540695
rect 182578 540530 182584 540885
rect 182618 540885 182672 541018
rect 182618 540530 182624 540885
rect 182578 540518 182624 540530
rect 182666 540530 182672 540885
rect 182706 540965 182718 541018
rect 182877 541025 182923 541037
rect 183069 541025 183115 541037
rect 183261 541025 183307 541037
rect 183453 541025 183499 541037
rect 183645 541025 183691 541037
rect 183837 541025 183883 541037
rect 182877 540965 182883 541025
rect 182706 540885 182883 540965
rect 182706 540530 182712 540885
rect 182666 540518 182712 540530
rect 182781 540571 182827 540583
rect 182781 540285 182787 540571
rect 182748 540083 182787 540285
rect 182821 540285 182827 540571
rect 182877 540537 182883 540885
rect 182917 540635 183075 541025
rect 182917 540537 182923 540635
rect 182877 540525 182923 540537
rect 182973 540571 183019 540583
rect 182973 540285 182979 540571
rect 182821 540083 182979 540285
rect 183013 540285 183019 540571
rect 183069 540537 183075 540635
rect 183109 540635 183267 541025
rect 183109 540537 183115 540635
rect 183069 540525 183115 540537
rect 183165 540571 183211 540583
rect 183165 540285 183171 540571
rect 183013 540083 183171 540285
rect 183205 540285 183211 540571
rect 183261 540537 183267 540635
rect 183301 540635 183459 541025
rect 183301 540537 183307 540635
rect 183261 540525 183307 540537
rect 183357 540571 183403 540583
rect 183357 540285 183363 540571
rect 183205 540083 183363 540285
rect 183397 540285 183403 540571
rect 183453 540537 183459 540635
rect 183493 540635 183651 541025
rect 183493 540537 183499 540635
rect 183453 540525 183499 540537
rect 183549 540571 183595 540583
rect 183549 540285 183555 540571
rect 183397 540083 183555 540285
rect 183589 540285 183595 540571
rect 183645 540537 183651 540635
rect 183685 540995 183843 541025
rect 183877 540995 183908 541025
rect 183685 540895 183788 540995
rect 183898 540895 183908 540995
rect 183685 540875 183843 540895
rect 183877 540875 183908 540895
rect 183685 540775 183788 540875
rect 183898 540775 183908 540875
rect 184103 540830 184153 541080
rect 184296 541119 184358 541125
rect 184296 541085 184308 541119
rect 184342 541085 184358 541119
rect 184296 541079 184358 541085
rect 184298 541065 184358 541079
rect 185478 540965 185678 541505
rect 185918 541125 185978 541135
rect 186218 541130 187238 541155
rect 186218 541126 187453 541130
rect 185878 541119 186018 541125
rect 185878 541085 185928 541119
rect 185962 541085 186018 541119
rect 186218 541095 186231 541126
rect 186219 541092 186231 541095
rect 186265 541095 186423 541126
rect 186265 541092 186277 541095
rect 186219 541086 186277 541092
rect 186411 541092 186423 541095
rect 186457 541095 186615 541126
rect 186457 541092 186469 541095
rect 186411 541086 186469 541092
rect 186603 541092 186615 541095
rect 186649 541095 186807 541126
rect 186649 541092 186661 541095
rect 186603 541086 186661 541092
rect 186795 541092 186807 541095
rect 186841 541095 186999 541126
rect 186841 541092 186853 541095
rect 186795 541086 186853 541092
rect 186987 541092 186999 541095
rect 187033 541095 187191 541126
rect 187033 541092 187045 541095
rect 186987 541086 187045 541092
rect 187179 541092 187191 541095
rect 187225 541092 187453 541126
rect 187179 541086 187453 541092
rect 185878 541018 186018 541085
rect 187223 541080 187453 541086
rect 185878 540965 185884 541018
rect 184578 540830 185168 540895
rect 185478 540885 185884 540965
rect 185478 540835 185678 540885
rect 183685 540755 183843 540775
rect 183877 540755 183908 540775
rect 183685 540655 183788 540755
rect 183898 540655 183908 540755
rect 183685 540635 183843 540655
rect 183685 540537 183691 540635
rect 183645 540525 183691 540537
rect 183741 540571 183787 540583
rect 183741 540285 183747 540571
rect 183589 540083 183747 540285
rect 183781 540285 183787 540571
rect 183837 540537 183843 540635
rect 183877 540635 183908 540655
rect 184098 540780 185168 540830
rect 183877 540537 183883 540635
rect 183837 540525 183883 540537
rect 183933 540571 183979 540583
rect 183933 540285 183939 540571
rect 183781 540083 183939 540285
rect 183973 540083 183979 540571
rect 184098 540335 184148 540780
rect 184578 540695 185168 540780
rect 184258 540564 184304 540576
rect 184098 540325 184158 540335
rect 184096 540319 184158 540325
rect 184096 540285 184108 540319
rect 184142 540285 184158 540319
rect 184096 540279 184158 540285
rect 184098 540275 184158 540279
rect 184058 540235 184104 540247
rect 184058 540155 184064 540235
rect 182748 540075 183979 540083
rect 182748 540071 182827 540075
rect 182973 540071 183019 540075
rect 183165 540071 183211 540075
rect 183357 540071 183403 540075
rect 183549 540071 183595 540075
rect 183741 540071 183787 540075
rect 183933 540071 183979 540075
rect 182748 540065 182818 540071
rect 182608 540009 182678 540025
rect 182608 539975 182628 540009
rect 182662 539975 182678 540009
rect 182608 539955 182678 539975
rect 182748 539755 182778 540065
rect 184038 540059 184064 540155
rect 184098 540059 184104 540235
rect 184038 540047 184104 540059
rect 184146 540235 184192 540247
rect 184146 540059 184152 540235
rect 184186 540225 184192 540235
rect 184258 540225 184264 540564
rect 184186 540076 184264 540225
rect 184298 540235 184304 540564
rect 184346 540564 184392 540576
rect 184346 540235 184352 540564
rect 184298 540076 184352 540235
rect 184386 540235 184392 540564
rect 184568 540245 184788 540255
rect 184386 540225 184408 540235
rect 184568 540225 184588 540245
rect 184386 540215 184588 540225
rect 184386 540085 184468 540215
rect 184528 540085 184588 540215
rect 184386 540076 184588 540085
rect 184186 540075 184588 540076
rect 184186 540059 184192 540075
rect 184258 540064 184392 540075
rect 184568 540065 184588 540075
rect 184768 540065 184788 540245
rect 184146 540047 184192 540059
rect 182823 540016 182881 540022
rect 182823 540015 182835 540016
rect 182818 539982 182835 540015
rect 182869 540015 182881 540016
rect 183015 540016 183073 540022
rect 183015 540015 183027 540016
rect 182869 539982 183027 540015
rect 183061 540015 183073 540016
rect 183207 540016 183265 540022
rect 183207 540015 183219 540016
rect 183061 539982 183219 540015
rect 183253 540015 183265 540016
rect 183399 540016 183457 540022
rect 183399 540015 183411 540016
rect 183253 539982 183411 540015
rect 183445 540015 183457 540016
rect 183591 540016 183649 540022
rect 183591 540015 183603 540016
rect 183445 539982 183603 540015
rect 183637 540015 183649 540016
rect 183783 540016 183841 540022
rect 183783 540015 183795 540016
rect 183637 539982 183795 540015
rect 183829 539982 183841 540016
rect 182818 539976 183841 539982
rect 182818 539955 183838 539976
rect 182178 539655 182778 539755
rect 182178 537931 182378 539655
rect 182538 539606 182778 539655
rect 182538 539572 182612 539606
rect 182646 539572 182778 539606
rect 182538 539513 182778 539572
rect 182918 539619 183928 539625
rect 182918 539613 183941 539619
rect 182918 539579 182935 539613
rect 182969 539579 183127 539613
rect 183161 539579 183319 539613
rect 183353 539579 183511 539613
rect 183545 539579 183703 539613
rect 183737 539579 183895 539613
rect 183929 539579 183941 539613
rect 182918 539573 183941 539579
rect 182918 539565 183928 539573
rect 184038 539525 184068 540047
rect 184096 540009 184158 540015
rect 184096 539975 184108 540009
rect 184142 539975 184158 540009
rect 184096 539969 184158 539975
rect 184098 539606 184158 539969
rect 184268 540009 184388 540064
rect 184568 540055 184788 540065
rect 184268 539975 184308 540009
rect 184342 539975 184388 540009
rect 184268 539955 184388 539975
rect 184098 539572 184112 539606
rect 184146 539572 184158 539606
rect 184098 539565 184158 539572
rect 184298 539606 184378 539625
rect 184298 539572 184312 539606
rect 184346 539572 184378 539606
rect 184298 539565 184378 539572
rect 182538 539415 182568 539513
rect 182562 538537 182568 539415
rect 182602 539415 182656 539513
rect 182602 538537 182608 539415
rect 182562 538525 182608 538537
rect 182650 538537 182656 539415
rect 182690 539495 182778 539513
rect 182881 539503 182927 539515
rect 182690 539485 182848 539495
rect 182881 539485 182887 539503
rect 182690 539415 182887 539485
rect 182690 538537 182696 539415
rect 182748 539205 182887 539415
rect 182785 539049 182831 539061
rect 182785 538561 182791 539049
rect 182825 538935 182831 539049
rect 182881 539015 182887 539205
rect 182921 539485 182927 539503
rect 183073 539503 183119 539515
rect 183073 539485 183079 539503
rect 182921 539205 183079 539485
rect 182921 539015 182927 539205
rect 182881 539003 182927 539015
rect 182977 539049 183023 539061
rect 182977 538935 182983 539049
rect 182825 538561 182983 538935
rect 183017 538935 183023 539049
rect 183073 539015 183079 539205
rect 183113 539485 183119 539503
rect 183265 539503 183311 539515
rect 183265 539485 183271 539503
rect 183113 539205 183271 539485
rect 183113 539015 183119 539205
rect 183073 539003 183119 539015
rect 183169 539049 183215 539061
rect 183169 538935 183175 539049
rect 183017 538561 183175 538935
rect 183209 538935 183215 539049
rect 183265 539015 183271 539205
rect 183305 539485 183311 539503
rect 183457 539503 183503 539515
rect 183457 539485 183463 539503
rect 183305 539205 183463 539485
rect 183305 539015 183311 539205
rect 183265 539003 183311 539015
rect 183361 539049 183407 539061
rect 183361 538935 183367 539049
rect 183209 538561 183367 538935
rect 183401 538935 183407 539049
rect 183457 539015 183463 539205
rect 183497 539485 183503 539503
rect 183649 539503 183695 539515
rect 183649 539485 183655 539503
rect 183497 539205 183655 539485
rect 183497 539015 183503 539205
rect 183457 539003 183503 539015
rect 183553 539049 183599 539061
rect 183553 538935 183559 539049
rect 183401 538561 183559 538935
rect 183593 538935 183599 539049
rect 183649 539015 183655 539205
rect 183689 539485 183695 539503
rect 183841 539503 183887 539515
rect 183841 539485 183847 539503
rect 183689 539205 183847 539485
rect 183689 539015 183695 539205
rect 183649 539003 183695 539015
rect 183745 539049 183791 539061
rect 183745 538935 183751 539049
rect 183593 538561 183751 538935
rect 183785 538935 183791 539049
rect 183841 539015 183847 539205
rect 183881 539485 183887 539503
rect 184038 539513 184108 539525
rect 183881 539205 183898 539485
rect 184038 539375 184068 539513
rect 183881 539015 183887 539205
rect 183841 539003 183887 539015
rect 183937 539049 183983 539061
rect 183937 538935 183943 539049
rect 183785 538805 183943 538935
rect 183785 538705 183798 538805
rect 183938 538705 183943 538805
rect 183785 538561 183943 538705
rect 183977 538561 183983 539049
rect 184062 539035 184068 539375
rect 182785 538555 183983 538561
rect 182785 538549 182831 538555
rect 182977 538549 183023 538555
rect 183169 538549 183215 538555
rect 183361 538549 183407 538555
rect 183553 538549 183599 538555
rect 183745 538549 183791 538555
rect 183937 538549 183983 538555
rect 184028 538937 184068 539035
rect 184102 538937 184108 539513
rect 184028 538925 184108 538937
rect 184150 539513 184196 539525
rect 184150 538937 184156 539513
rect 184190 539505 184196 539513
rect 184190 539275 184308 539505
rect 184568 539305 184788 539315
rect 184568 539275 184588 539305
rect 184190 539265 184588 539275
rect 184190 539175 184468 539265
rect 184518 539175 184588 539265
rect 184190 539165 184588 539175
rect 184190 539042 184308 539165
rect 184568 539125 184588 539165
rect 184768 539125 184788 539305
rect 184568 539115 184788 539125
rect 184190 538937 184268 539042
rect 184150 538935 184268 538937
rect 184150 538925 184196 538935
rect 182650 538525 182696 538537
rect 182827 538485 182885 538491
rect 183019 538485 183077 538491
rect 183211 538485 183269 538491
rect 183403 538485 183461 538491
rect 183595 538485 183653 538491
rect 183787 538485 183845 538491
rect 184028 538485 184068 538925
rect 184098 538878 184158 538885
rect 184098 538844 184112 538878
rect 184146 538844 184158 538878
rect 184098 538825 184158 538844
rect 184262 538575 184268 538935
rect 182598 538478 182658 538485
rect 182598 538444 182612 538478
rect 182646 538444 182658 538478
rect 182598 538425 182658 538444
rect 182818 538451 182839 538485
rect 182873 538451 183031 538485
rect 183065 538451 183223 538485
rect 183257 538451 183415 538485
rect 183449 538451 183607 538485
rect 183641 538451 183799 538485
rect 183833 538451 184068 538485
rect 182818 538425 184068 538451
rect 184258 538554 184268 538575
rect 184302 538575 184308 539042
rect 184350 539042 184396 539054
rect 184350 538575 184356 539042
rect 184302 538554 184356 538575
rect 184390 538554 184396 539042
rect 184258 538542 184396 538554
rect 184258 538478 184378 538542
rect 184258 538445 184312 538478
rect 184298 538444 184312 538445
rect 184346 538445 184378 538478
rect 184346 538444 184358 538445
rect 184298 538425 184358 538444
rect 182178 537815 182258 537931
rect 182252 537534 182258 537815
rect 182296 537815 182378 537931
rect 182296 537534 182302 537815
rect 182252 537522 182302 537534
rect 182252 537256 182302 537268
rect 182252 537085 182258 537256
rect 182128 536859 182258 537085
rect 182296 537085 182302 537256
rect 182296 536859 182428 537085
rect 182128 536285 182428 536859
rect 182128 536025 182188 536285
rect 182388 536025 182428 536285
rect 182128 535985 182428 536025
rect 184968 533555 185168 540695
rect 185878 540530 185884 540885
rect 185918 540885 185972 541018
rect 185918 540530 185924 540885
rect 185878 540518 185924 540530
rect 185966 540530 185972 540885
rect 186006 540965 186018 541018
rect 186177 541025 186223 541037
rect 186369 541025 186415 541037
rect 186561 541025 186607 541037
rect 186753 541025 186799 541037
rect 186945 541025 186991 541037
rect 187137 541025 187183 541037
rect 186177 540965 186183 541025
rect 186006 540885 186183 540965
rect 186006 540530 186012 540885
rect 185966 540518 186012 540530
rect 186081 540571 186127 540583
rect 186081 540285 186087 540571
rect 186048 540083 186087 540285
rect 186121 540285 186127 540571
rect 186177 540537 186183 540885
rect 186217 540635 186375 541025
rect 186217 540537 186223 540635
rect 186177 540525 186223 540537
rect 186273 540571 186319 540583
rect 186273 540285 186279 540571
rect 186121 540083 186279 540285
rect 186313 540285 186319 540571
rect 186369 540537 186375 540635
rect 186409 540635 186567 541025
rect 186409 540537 186415 540635
rect 186369 540525 186415 540537
rect 186465 540571 186511 540583
rect 186465 540285 186471 540571
rect 186313 540083 186471 540285
rect 186505 540285 186511 540571
rect 186561 540537 186567 540635
rect 186601 540635 186759 541025
rect 186601 540537 186607 540635
rect 186561 540525 186607 540537
rect 186657 540571 186703 540583
rect 186657 540285 186663 540571
rect 186505 540083 186663 540285
rect 186697 540285 186703 540571
rect 186753 540537 186759 540635
rect 186793 540635 186951 541025
rect 186793 540537 186799 540635
rect 186753 540525 186799 540537
rect 186849 540571 186895 540583
rect 186849 540285 186855 540571
rect 186697 540083 186855 540285
rect 186889 540285 186895 540571
rect 186945 540537 186951 540635
rect 186985 540995 187143 541025
rect 187177 540995 187208 541025
rect 186985 540895 187088 540995
rect 187198 540895 187208 540995
rect 186985 540875 187143 540895
rect 187177 540875 187208 540895
rect 186985 540775 187088 540875
rect 187198 540775 187208 540875
rect 187403 540830 187453 541080
rect 187596 541119 187658 541125
rect 187596 541085 187608 541119
rect 187642 541085 187658 541119
rect 187596 541079 187658 541085
rect 187598 541065 187658 541079
rect 188778 540965 188978 541505
rect 189218 541125 189278 541135
rect 189518 541130 190538 541155
rect 189518 541126 190753 541130
rect 189178 541119 189318 541125
rect 189178 541085 189228 541119
rect 189262 541085 189318 541119
rect 189518 541095 189531 541126
rect 189519 541092 189531 541095
rect 189565 541095 189723 541126
rect 189565 541092 189577 541095
rect 189519 541086 189577 541092
rect 189711 541092 189723 541095
rect 189757 541095 189915 541126
rect 189757 541092 189769 541095
rect 189711 541086 189769 541092
rect 189903 541092 189915 541095
rect 189949 541095 190107 541126
rect 189949 541092 189961 541095
rect 189903 541086 189961 541092
rect 190095 541092 190107 541095
rect 190141 541095 190299 541126
rect 190141 541092 190153 541095
rect 190095 541086 190153 541092
rect 190287 541092 190299 541095
rect 190333 541095 190491 541126
rect 190333 541092 190345 541095
rect 190287 541086 190345 541092
rect 190479 541092 190491 541095
rect 190525 541092 190753 541126
rect 190479 541086 190753 541092
rect 189178 541018 189318 541085
rect 190523 541080 190753 541086
rect 189178 540965 189184 541018
rect 187878 540830 188398 540895
rect 188778 540885 189184 540965
rect 188778 540835 188978 540885
rect 186985 540755 187143 540775
rect 187177 540755 187208 540775
rect 186985 540655 187088 540755
rect 187198 540655 187208 540755
rect 186985 540635 187143 540655
rect 186985 540537 186991 540635
rect 186945 540525 186991 540537
rect 187041 540571 187087 540583
rect 187041 540285 187047 540571
rect 186889 540083 187047 540285
rect 187081 540285 187087 540571
rect 187137 540537 187143 540635
rect 187177 540635 187208 540655
rect 187398 540780 188398 540830
rect 187177 540537 187183 540635
rect 187137 540525 187183 540537
rect 187233 540571 187279 540583
rect 187233 540285 187239 540571
rect 187081 540083 187239 540285
rect 187273 540083 187279 540571
rect 187398 540335 187448 540780
rect 187878 540695 188398 540780
rect 187558 540564 187604 540576
rect 187398 540325 187458 540335
rect 187396 540319 187458 540325
rect 187396 540285 187408 540319
rect 187442 540285 187458 540319
rect 187396 540279 187458 540285
rect 187398 540275 187458 540279
rect 187358 540235 187404 540247
rect 187358 540155 187364 540235
rect 186048 540075 187279 540083
rect 186048 540071 186127 540075
rect 186273 540071 186319 540075
rect 186465 540071 186511 540075
rect 186657 540071 186703 540075
rect 186849 540071 186895 540075
rect 187041 540071 187087 540075
rect 187233 540071 187279 540075
rect 186048 540065 186118 540071
rect 185908 540009 185978 540025
rect 185908 539975 185928 540009
rect 185962 539975 185978 540009
rect 185908 539955 185978 539975
rect 186048 539755 186078 540065
rect 187338 540059 187364 540155
rect 187398 540059 187404 540235
rect 187338 540047 187404 540059
rect 187446 540235 187492 540247
rect 187446 540059 187452 540235
rect 187486 540225 187492 540235
rect 187558 540225 187564 540564
rect 187486 540076 187564 540225
rect 187598 540235 187604 540564
rect 187646 540564 187692 540576
rect 187646 540235 187652 540564
rect 187598 540076 187652 540235
rect 187686 540235 187692 540564
rect 187868 540245 188088 540255
rect 187686 540225 187708 540235
rect 187868 540225 187898 540245
rect 187686 540215 187898 540225
rect 187686 540085 187768 540215
rect 187828 540085 187898 540215
rect 187686 540076 187898 540085
rect 187486 540075 187898 540076
rect 187486 540059 187492 540075
rect 187558 540064 187692 540075
rect 187868 540065 187898 540075
rect 188078 540065 188088 540245
rect 187446 540047 187492 540059
rect 186123 540016 186181 540022
rect 186123 540015 186135 540016
rect 186118 539982 186135 540015
rect 186169 540015 186181 540016
rect 186315 540016 186373 540022
rect 186315 540015 186327 540016
rect 186169 539982 186327 540015
rect 186361 540015 186373 540016
rect 186507 540016 186565 540022
rect 186507 540015 186519 540016
rect 186361 539982 186519 540015
rect 186553 540015 186565 540016
rect 186699 540016 186757 540022
rect 186699 540015 186711 540016
rect 186553 539982 186711 540015
rect 186745 540015 186757 540016
rect 186891 540016 186949 540022
rect 186891 540015 186903 540016
rect 186745 539982 186903 540015
rect 186937 540015 186949 540016
rect 187083 540016 187141 540022
rect 187083 540015 187095 540016
rect 186937 539982 187095 540015
rect 187129 539982 187141 540016
rect 186118 539976 187141 539982
rect 186118 539955 187138 539976
rect 185478 539655 186078 539755
rect 185478 537931 185678 539655
rect 185838 539606 186078 539655
rect 185838 539572 185912 539606
rect 185946 539572 186078 539606
rect 185838 539513 186078 539572
rect 186218 539619 187228 539625
rect 186218 539613 187241 539619
rect 186218 539579 186235 539613
rect 186269 539579 186427 539613
rect 186461 539579 186619 539613
rect 186653 539579 186811 539613
rect 186845 539579 187003 539613
rect 187037 539579 187195 539613
rect 187229 539579 187241 539613
rect 186218 539573 187241 539579
rect 186218 539565 187228 539573
rect 187338 539525 187368 540047
rect 187396 540009 187458 540015
rect 187396 539975 187408 540009
rect 187442 539975 187458 540009
rect 187396 539969 187458 539975
rect 187398 539606 187458 539969
rect 187568 540009 187688 540064
rect 187868 540055 188088 540065
rect 187568 539975 187608 540009
rect 187642 539975 187688 540009
rect 187568 539955 187688 539975
rect 187398 539572 187412 539606
rect 187446 539572 187458 539606
rect 187398 539565 187458 539572
rect 187598 539606 187678 539625
rect 187598 539572 187612 539606
rect 187646 539572 187678 539606
rect 187598 539565 187678 539572
rect 185838 539415 185868 539513
rect 185862 538537 185868 539415
rect 185902 539415 185956 539513
rect 185902 538537 185908 539415
rect 185862 538525 185908 538537
rect 185950 538537 185956 539415
rect 185990 539495 186078 539513
rect 186181 539503 186227 539515
rect 185990 539485 186148 539495
rect 186181 539485 186187 539503
rect 185990 539415 186187 539485
rect 185990 538537 185996 539415
rect 186048 539205 186187 539415
rect 186085 539049 186131 539061
rect 186085 538561 186091 539049
rect 186125 538935 186131 539049
rect 186181 539015 186187 539205
rect 186221 539485 186227 539503
rect 186373 539503 186419 539515
rect 186373 539485 186379 539503
rect 186221 539205 186379 539485
rect 186221 539015 186227 539205
rect 186181 539003 186227 539015
rect 186277 539049 186323 539061
rect 186277 538935 186283 539049
rect 186125 538561 186283 538935
rect 186317 538935 186323 539049
rect 186373 539015 186379 539205
rect 186413 539485 186419 539503
rect 186565 539503 186611 539515
rect 186565 539485 186571 539503
rect 186413 539205 186571 539485
rect 186413 539015 186419 539205
rect 186373 539003 186419 539015
rect 186469 539049 186515 539061
rect 186469 538935 186475 539049
rect 186317 538561 186475 538935
rect 186509 538935 186515 539049
rect 186565 539015 186571 539205
rect 186605 539485 186611 539503
rect 186757 539503 186803 539515
rect 186757 539485 186763 539503
rect 186605 539205 186763 539485
rect 186605 539015 186611 539205
rect 186565 539003 186611 539015
rect 186661 539049 186707 539061
rect 186661 538935 186667 539049
rect 186509 538561 186667 538935
rect 186701 538935 186707 539049
rect 186757 539015 186763 539205
rect 186797 539485 186803 539503
rect 186949 539503 186995 539515
rect 186949 539485 186955 539503
rect 186797 539205 186955 539485
rect 186797 539015 186803 539205
rect 186757 539003 186803 539015
rect 186853 539049 186899 539061
rect 186853 538935 186859 539049
rect 186701 538561 186859 538935
rect 186893 538935 186899 539049
rect 186949 539015 186955 539205
rect 186989 539485 186995 539503
rect 187141 539503 187187 539515
rect 187141 539485 187147 539503
rect 186989 539205 187147 539485
rect 186989 539015 186995 539205
rect 186949 539003 186995 539015
rect 187045 539049 187091 539061
rect 187045 538935 187051 539049
rect 186893 538561 187051 538935
rect 187085 538935 187091 539049
rect 187141 539015 187147 539205
rect 187181 539485 187187 539503
rect 187338 539513 187408 539525
rect 187181 539205 187198 539485
rect 187338 539375 187368 539513
rect 187181 539015 187187 539205
rect 187141 539003 187187 539015
rect 187237 539049 187283 539061
rect 187237 538935 187243 539049
rect 187085 538805 187243 538935
rect 187085 538705 187098 538805
rect 187238 538705 187243 538805
rect 187085 538561 187243 538705
rect 187277 538561 187283 539049
rect 187362 539035 187368 539375
rect 186085 538555 187283 538561
rect 186085 538549 186131 538555
rect 186277 538549 186323 538555
rect 186469 538549 186515 538555
rect 186661 538549 186707 538555
rect 186853 538549 186899 538555
rect 187045 538549 187091 538555
rect 187237 538549 187283 538555
rect 187328 538937 187368 539035
rect 187402 538937 187408 539513
rect 187328 538925 187408 538937
rect 187450 539513 187496 539525
rect 187450 538937 187456 539513
rect 187490 539505 187496 539513
rect 187490 539275 187608 539505
rect 187868 539305 188088 539315
rect 187868 539275 187888 539305
rect 187490 539265 187888 539275
rect 187490 539175 187768 539265
rect 187818 539175 187888 539265
rect 187490 539165 187888 539175
rect 187490 539042 187608 539165
rect 187868 539125 187888 539165
rect 188068 539125 188088 539305
rect 187868 539115 188088 539125
rect 187490 538937 187568 539042
rect 187450 538935 187568 538937
rect 187450 538925 187496 538935
rect 185950 538525 185996 538537
rect 186127 538485 186185 538491
rect 186319 538485 186377 538491
rect 186511 538485 186569 538491
rect 186703 538485 186761 538491
rect 186895 538485 186953 538491
rect 187087 538485 187145 538491
rect 187328 538485 187368 538925
rect 187398 538878 187458 538885
rect 187398 538844 187412 538878
rect 187446 538844 187458 538878
rect 187398 538825 187458 538844
rect 187562 538575 187568 538935
rect 185898 538478 185958 538485
rect 185898 538444 185912 538478
rect 185946 538444 185958 538478
rect 185898 538425 185958 538444
rect 186118 538451 186139 538485
rect 186173 538451 186331 538485
rect 186365 538451 186523 538485
rect 186557 538451 186715 538485
rect 186749 538451 186907 538485
rect 186941 538451 187099 538485
rect 187133 538451 187368 538485
rect 186118 538425 187368 538451
rect 187558 538554 187568 538575
rect 187602 538575 187608 539042
rect 187650 539042 187696 539054
rect 187650 538575 187656 539042
rect 187602 538554 187656 538575
rect 187690 538554 187696 539042
rect 187558 538542 187696 538554
rect 187558 538478 187678 538542
rect 187558 538445 187612 538478
rect 187598 538444 187612 538445
rect 187646 538445 187678 538478
rect 187646 538444 187658 538445
rect 187598 538425 187658 538444
rect 185478 537815 185558 537931
rect 185552 537534 185558 537815
rect 185596 537815 185678 537931
rect 185596 537534 185602 537815
rect 185552 537522 185602 537534
rect 185552 537396 185602 537408
rect 185552 537205 185558 537396
rect 185428 536999 185558 537205
rect 185596 537205 185602 537396
rect 185596 536999 185728 537205
rect 185428 536265 185728 536999
rect 185428 536145 185488 536265
rect 185698 536145 185728 536265
rect 185428 536105 185728 536145
rect 180828 533305 181928 533505
rect 182928 533355 185168 533555
rect 178218 532735 178928 532755
rect 178218 532565 178698 532735
rect 178828 532565 178928 532735
rect 178218 532555 178928 532565
rect 180828 532735 181028 533305
rect 180828 532565 180868 532735
rect 180998 532565 181028 532735
rect 180828 532455 181028 532565
rect 182928 532735 183128 533355
rect 184968 533305 185168 533355
rect 188198 533255 188398 540695
rect 189178 540530 189184 540885
rect 189218 540885 189272 541018
rect 189218 540530 189224 540885
rect 189178 540518 189224 540530
rect 189266 540530 189272 540885
rect 189306 540965 189318 541018
rect 189477 541025 189523 541037
rect 189669 541025 189715 541037
rect 189861 541025 189907 541037
rect 190053 541025 190099 541037
rect 190245 541025 190291 541037
rect 190437 541025 190483 541037
rect 189477 540965 189483 541025
rect 189306 540885 189483 540965
rect 189306 540530 189312 540885
rect 189266 540518 189312 540530
rect 189381 540571 189427 540583
rect 189381 540285 189387 540571
rect 189348 540083 189387 540285
rect 189421 540285 189427 540571
rect 189477 540537 189483 540885
rect 189517 540635 189675 541025
rect 189517 540537 189523 540635
rect 189477 540525 189523 540537
rect 189573 540571 189619 540583
rect 189573 540285 189579 540571
rect 189421 540083 189579 540285
rect 189613 540285 189619 540571
rect 189669 540537 189675 540635
rect 189709 540635 189867 541025
rect 189709 540537 189715 540635
rect 189669 540525 189715 540537
rect 189765 540571 189811 540583
rect 189765 540285 189771 540571
rect 189613 540083 189771 540285
rect 189805 540285 189811 540571
rect 189861 540537 189867 540635
rect 189901 540635 190059 541025
rect 189901 540537 189907 540635
rect 189861 540525 189907 540537
rect 189957 540571 190003 540583
rect 189957 540285 189963 540571
rect 189805 540083 189963 540285
rect 189997 540285 190003 540571
rect 190053 540537 190059 540635
rect 190093 540635 190251 541025
rect 190093 540537 190099 540635
rect 190053 540525 190099 540537
rect 190149 540571 190195 540583
rect 190149 540285 190155 540571
rect 189997 540083 190155 540285
rect 190189 540285 190195 540571
rect 190245 540537 190251 540635
rect 190285 540995 190443 541025
rect 190477 540995 190508 541025
rect 190285 540895 190388 540995
rect 190498 540895 190508 540995
rect 190285 540875 190443 540895
rect 190477 540875 190508 540895
rect 190285 540775 190388 540875
rect 190498 540775 190508 540875
rect 190703 540830 190753 541080
rect 190896 541119 190958 541125
rect 190896 541085 190908 541119
rect 190942 541085 190958 541119
rect 190896 541079 190958 541085
rect 190898 541065 190958 541079
rect 191178 540830 191678 540895
rect 190285 540755 190443 540775
rect 190477 540755 190508 540775
rect 190285 540655 190388 540755
rect 190498 540655 190508 540755
rect 190285 540635 190443 540655
rect 190285 540537 190291 540635
rect 190245 540525 190291 540537
rect 190341 540571 190387 540583
rect 190341 540285 190347 540571
rect 190189 540083 190347 540285
rect 190381 540285 190387 540571
rect 190437 540537 190443 540635
rect 190477 540635 190508 540655
rect 190698 540780 191678 540830
rect 190477 540537 190483 540635
rect 190437 540525 190483 540537
rect 190533 540571 190579 540583
rect 190533 540285 190539 540571
rect 190381 540083 190539 540285
rect 190573 540083 190579 540571
rect 190698 540335 190748 540780
rect 191178 540695 191678 540780
rect 190858 540564 190904 540576
rect 190698 540325 190758 540335
rect 190696 540319 190758 540325
rect 190696 540285 190708 540319
rect 190742 540285 190758 540319
rect 190696 540279 190758 540285
rect 190698 540275 190758 540279
rect 190658 540235 190704 540247
rect 190658 540155 190664 540235
rect 189348 540075 190579 540083
rect 189348 540071 189427 540075
rect 189573 540071 189619 540075
rect 189765 540071 189811 540075
rect 189957 540071 190003 540075
rect 190149 540071 190195 540075
rect 190341 540071 190387 540075
rect 190533 540071 190579 540075
rect 189348 540065 189418 540071
rect 189208 540009 189278 540025
rect 189208 539975 189228 540009
rect 189262 539975 189278 540009
rect 189208 539955 189278 539975
rect 189348 539755 189378 540065
rect 190638 540059 190664 540155
rect 190698 540059 190704 540235
rect 190638 540047 190704 540059
rect 190746 540235 190792 540247
rect 190746 540059 190752 540235
rect 190786 540225 190792 540235
rect 190858 540225 190864 540564
rect 190786 540076 190864 540225
rect 190898 540235 190904 540564
rect 190946 540564 190992 540576
rect 190946 540235 190952 540564
rect 190898 540076 190952 540235
rect 190986 540235 190992 540564
rect 191168 540245 191388 540255
rect 190986 540225 191008 540235
rect 191168 540225 191188 540245
rect 190986 540215 191188 540225
rect 190986 540085 191068 540215
rect 191128 540085 191188 540215
rect 190986 540076 191188 540085
rect 190786 540075 191188 540076
rect 190786 540059 190792 540075
rect 190858 540064 190992 540075
rect 191168 540065 191188 540075
rect 191368 540065 191388 540245
rect 190746 540047 190792 540059
rect 189423 540016 189481 540022
rect 189423 540015 189435 540016
rect 189418 539982 189435 540015
rect 189469 540015 189481 540016
rect 189615 540016 189673 540022
rect 189615 540015 189627 540016
rect 189469 539982 189627 540015
rect 189661 540015 189673 540016
rect 189807 540016 189865 540022
rect 189807 540015 189819 540016
rect 189661 539982 189819 540015
rect 189853 540015 189865 540016
rect 189999 540016 190057 540022
rect 189999 540015 190011 540016
rect 189853 539982 190011 540015
rect 190045 540015 190057 540016
rect 190191 540016 190249 540022
rect 190191 540015 190203 540016
rect 190045 539982 190203 540015
rect 190237 540015 190249 540016
rect 190383 540016 190441 540022
rect 190383 540015 190395 540016
rect 190237 539982 190395 540015
rect 190429 539982 190441 540016
rect 189418 539976 190441 539982
rect 189418 539955 190438 539976
rect 188778 539655 189378 539755
rect 188778 537931 188978 539655
rect 189138 539606 189378 539655
rect 189138 539572 189212 539606
rect 189246 539572 189378 539606
rect 189138 539513 189378 539572
rect 189518 539619 190528 539625
rect 189518 539613 190541 539619
rect 189518 539579 189535 539613
rect 189569 539579 189727 539613
rect 189761 539579 189919 539613
rect 189953 539579 190111 539613
rect 190145 539579 190303 539613
rect 190337 539579 190495 539613
rect 190529 539579 190541 539613
rect 189518 539573 190541 539579
rect 189518 539565 190528 539573
rect 190638 539525 190668 540047
rect 190696 540009 190758 540015
rect 190696 539975 190708 540009
rect 190742 539975 190758 540009
rect 190696 539969 190758 539975
rect 190698 539606 190758 539969
rect 190868 540009 190988 540064
rect 191168 540055 191388 540065
rect 190868 539975 190908 540009
rect 190942 539975 190988 540009
rect 190868 539955 190988 539975
rect 190698 539572 190712 539606
rect 190746 539572 190758 539606
rect 190698 539565 190758 539572
rect 190898 539606 190978 539625
rect 190898 539572 190912 539606
rect 190946 539572 190978 539606
rect 190898 539565 190978 539572
rect 189138 539415 189168 539513
rect 189162 538537 189168 539415
rect 189202 539415 189256 539513
rect 189202 538537 189208 539415
rect 189162 538525 189208 538537
rect 189250 538537 189256 539415
rect 189290 539495 189378 539513
rect 189481 539503 189527 539515
rect 189290 539485 189448 539495
rect 189481 539485 189487 539503
rect 189290 539415 189487 539485
rect 189290 538537 189296 539415
rect 189348 539205 189487 539415
rect 189385 539049 189431 539061
rect 189385 538561 189391 539049
rect 189425 538935 189431 539049
rect 189481 539015 189487 539205
rect 189521 539485 189527 539503
rect 189673 539503 189719 539515
rect 189673 539485 189679 539503
rect 189521 539205 189679 539485
rect 189521 539015 189527 539205
rect 189481 539003 189527 539015
rect 189577 539049 189623 539061
rect 189577 538935 189583 539049
rect 189425 538561 189583 538935
rect 189617 538935 189623 539049
rect 189673 539015 189679 539205
rect 189713 539485 189719 539503
rect 189865 539503 189911 539515
rect 189865 539485 189871 539503
rect 189713 539205 189871 539485
rect 189713 539015 189719 539205
rect 189673 539003 189719 539015
rect 189769 539049 189815 539061
rect 189769 538935 189775 539049
rect 189617 538561 189775 538935
rect 189809 538935 189815 539049
rect 189865 539015 189871 539205
rect 189905 539485 189911 539503
rect 190057 539503 190103 539515
rect 190057 539485 190063 539503
rect 189905 539205 190063 539485
rect 189905 539015 189911 539205
rect 189865 539003 189911 539015
rect 189961 539049 190007 539061
rect 189961 538935 189967 539049
rect 189809 538561 189967 538935
rect 190001 538935 190007 539049
rect 190057 539015 190063 539205
rect 190097 539485 190103 539503
rect 190249 539503 190295 539515
rect 190249 539485 190255 539503
rect 190097 539205 190255 539485
rect 190097 539015 190103 539205
rect 190057 539003 190103 539015
rect 190153 539049 190199 539061
rect 190153 538935 190159 539049
rect 190001 538561 190159 538935
rect 190193 538935 190199 539049
rect 190249 539015 190255 539205
rect 190289 539485 190295 539503
rect 190441 539503 190487 539515
rect 190441 539485 190447 539503
rect 190289 539205 190447 539485
rect 190289 539015 190295 539205
rect 190249 539003 190295 539015
rect 190345 539049 190391 539061
rect 190345 538935 190351 539049
rect 190193 538561 190351 538935
rect 190385 538935 190391 539049
rect 190441 539015 190447 539205
rect 190481 539485 190487 539503
rect 190638 539513 190708 539525
rect 190481 539205 190498 539485
rect 190638 539375 190668 539513
rect 190481 539015 190487 539205
rect 190441 539003 190487 539015
rect 190537 539049 190583 539061
rect 190537 538935 190543 539049
rect 190385 538805 190543 538935
rect 190385 538705 190398 538805
rect 190538 538705 190543 538805
rect 190385 538561 190543 538705
rect 190577 538561 190583 539049
rect 190662 539035 190668 539375
rect 189385 538555 190583 538561
rect 189385 538549 189431 538555
rect 189577 538549 189623 538555
rect 189769 538549 189815 538555
rect 189961 538549 190007 538555
rect 190153 538549 190199 538555
rect 190345 538549 190391 538555
rect 190537 538549 190583 538555
rect 190628 538937 190668 539035
rect 190702 538937 190708 539513
rect 190628 538925 190708 538937
rect 190750 539513 190796 539525
rect 190750 538937 190756 539513
rect 190790 539505 190796 539513
rect 190790 539275 190908 539505
rect 191188 539315 191388 539325
rect 191168 539275 191198 539315
rect 190790 539265 191198 539275
rect 190790 539175 191068 539265
rect 191118 539175 191198 539265
rect 190790 539165 191198 539175
rect 190790 539042 190908 539165
rect 191168 539135 191198 539165
rect 191378 539135 191388 539315
rect 191168 539115 191388 539135
rect 190790 538937 190868 539042
rect 190750 538935 190868 538937
rect 190750 538925 190796 538935
rect 189250 538525 189296 538537
rect 189427 538485 189485 538491
rect 189619 538485 189677 538491
rect 189811 538485 189869 538491
rect 190003 538485 190061 538491
rect 190195 538485 190253 538491
rect 190387 538485 190445 538491
rect 190628 538485 190668 538925
rect 190698 538878 190758 538885
rect 190698 538844 190712 538878
rect 190746 538844 190758 538878
rect 190698 538825 190758 538844
rect 190862 538575 190868 538935
rect 189198 538478 189258 538485
rect 189198 538444 189212 538478
rect 189246 538444 189258 538478
rect 189198 538425 189258 538444
rect 189418 538451 189439 538485
rect 189473 538451 189631 538485
rect 189665 538451 189823 538485
rect 189857 538451 190015 538485
rect 190049 538451 190207 538485
rect 190241 538451 190399 538485
rect 190433 538451 190668 538485
rect 189418 538425 190668 538451
rect 190858 538554 190868 538575
rect 190902 538575 190908 539042
rect 190950 539042 190996 539054
rect 190950 538575 190956 539042
rect 190902 538554 190956 538575
rect 190990 538554 190996 539042
rect 190858 538542 190996 538554
rect 190858 538478 190978 538542
rect 190858 538445 190912 538478
rect 190898 538444 190912 538445
rect 190946 538445 190978 538478
rect 190946 538444 190958 538445
rect 190898 538425 190958 538444
rect 188778 537815 188858 537931
rect 188852 537534 188858 537815
rect 188896 537815 188978 537931
rect 188896 537534 188902 537815
rect 188852 537522 188902 537534
rect 188852 537300 188902 537312
rect 188852 537105 188858 537300
rect 188728 536903 188858 537105
rect 188896 537105 188902 537300
rect 188896 536903 189028 537105
rect 188728 536275 189028 536903
rect 188728 536035 188778 536275
rect 188998 536035 189028 536275
rect 188728 536005 189028 536035
rect 182928 532565 182958 532735
rect 183088 532565 183128 532735
rect 182928 532455 183128 532565
rect 185028 533055 188398 533255
rect 185028 532775 185228 533055
rect 185028 532605 185058 532775
rect 185188 532605 185228 532775
rect 191478 532755 191678 540695
rect 193000 540260 195000 542000
rect 192620 540255 195000 540260
rect 191748 540245 195000 540255
rect 191748 540065 191808 540245
rect 191988 540065 195000 540245
rect 191748 540055 192228 540065
rect 192428 540055 195000 540065
rect 192620 540050 195000 540055
rect 193000 540000 195000 540050
rect 192620 539315 195000 539320
rect 191808 539305 195000 539315
rect 191808 539125 191818 539305
rect 191998 539125 195000 539305
rect 191808 539115 195000 539125
rect 192620 539110 195000 539115
rect 193000 537320 195000 539110
rect 185028 532555 185228 532605
rect 187128 532735 191678 532755
rect 187128 532595 187168 532735
rect 187268 532595 191678 532735
rect 187128 532555 191678 532595
rect 172208 530605 187480 530627
rect 172208 530596 174623 530605
rect 172208 530562 172237 530596
rect 172271 530562 172329 530596
rect 172363 530562 172421 530596
rect 172455 530562 172513 530596
rect 172547 530562 172605 530596
rect 172639 530562 172697 530596
rect 172731 530562 172789 530596
rect 172823 530562 172881 530596
rect 172915 530562 172973 530596
rect 173007 530562 173065 530596
rect 173099 530562 173157 530596
rect 173191 530562 173249 530596
rect 173283 530562 173341 530596
rect 173375 530562 173433 530596
rect 173467 530562 173525 530596
rect 173559 530562 173617 530596
rect 173651 530562 173709 530596
rect 173743 530562 173801 530596
rect 173835 530562 173893 530596
rect 173927 530562 173985 530596
rect 174019 530562 174077 530596
rect 174111 530562 174169 530596
rect 174203 530562 174261 530596
rect 174295 530562 174353 530596
rect 174387 530562 174445 530596
rect 174479 530562 174537 530596
rect 174571 530562 174623 530596
rect 172208 530553 174623 530562
rect 174675 530553 174687 530605
rect 174739 530596 174751 530605
rect 174803 530596 174815 530605
rect 174803 530562 174813 530596
rect 174739 530553 174751 530562
rect 174803 530553 174815 530562
rect 174867 530553 174879 530605
rect 174931 530596 178441 530605
rect 174939 530562 174997 530596
rect 175031 530562 175089 530596
rect 175123 530562 175181 530596
rect 175215 530562 175273 530596
rect 175307 530562 175365 530596
rect 175399 530562 175457 530596
rect 175491 530562 175549 530596
rect 175583 530562 175641 530596
rect 175675 530562 175733 530596
rect 175767 530562 175825 530596
rect 175859 530562 175917 530596
rect 175951 530562 176009 530596
rect 176043 530562 176101 530596
rect 176135 530562 176193 530596
rect 176227 530562 176285 530596
rect 176319 530562 176377 530596
rect 176411 530562 176469 530596
rect 176503 530562 176561 530596
rect 176595 530562 176653 530596
rect 176687 530562 176745 530596
rect 176779 530562 176837 530596
rect 176871 530562 176929 530596
rect 176963 530562 177021 530596
rect 177055 530562 177113 530596
rect 177147 530562 177205 530596
rect 177239 530562 177297 530596
rect 177331 530562 177389 530596
rect 177423 530562 177481 530596
rect 177515 530562 177573 530596
rect 177607 530562 177665 530596
rect 177699 530562 177757 530596
rect 177791 530562 177849 530596
rect 177883 530562 177941 530596
rect 177975 530562 178033 530596
rect 178067 530562 178125 530596
rect 178159 530562 178217 530596
rect 178251 530562 178309 530596
rect 178343 530562 178401 530596
rect 178435 530562 178441 530596
rect 174931 530553 178441 530562
rect 178493 530596 178505 530605
rect 178493 530553 178505 530562
rect 178557 530553 178569 530605
rect 178621 530553 178633 530605
rect 178685 530596 178697 530605
rect 178749 530596 182259 530605
rect 178749 530562 178769 530596
rect 178803 530562 178861 530596
rect 178895 530562 178953 530596
rect 178987 530562 179045 530596
rect 179079 530562 179137 530596
rect 179171 530562 179229 530596
rect 179263 530562 179321 530596
rect 179355 530562 179413 530596
rect 179447 530562 179505 530596
rect 179539 530562 179597 530596
rect 179631 530562 179689 530596
rect 179723 530562 179781 530596
rect 179815 530562 179873 530596
rect 179907 530562 179965 530596
rect 179999 530562 180057 530596
rect 180091 530562 180149 530596
rect 180183 530562 180241 530596
rect 180275 530562 180333 530596
rect 180367 530562 180425 530596
rect 180459 530562 180517 530596
rect 180551 530562 180609 530596
rect 180643 530562 180701 530596
rect 180735 530562 180793 530596
rect 180827 530562 180885 530596
rect 180919 530562 180977 530596
rect 181011 530562 181069 530596
rect 181103 530562 181161 530596
rect 181195 530562 181253 530596
rect 181287 530562 181345 530596
rect 181379 530562 181437 530596
rect 181471 530562 181529 530596
rect 181563 530562 181621 530596
rect 181655 530562 181713 530596
rect 181747 530562 181805 530596
rect 181839 530562 181897 530596
rect 181931 530562 181989 530596
rect 182023 530562 182081 530596
rect 182115 530562 182173 530596
rect 182207 530562 182259 530596
rect 178685 530553 178697 530562
rect 178749 530553 182259 530562
rect 182311 530553 182323 530605
rect 182375 530596 182387 530605
rect 182439 530596 182451 530605
rect 182439 530562 182449 530596
rect 182375 530553 182387 530562
rect 182439 530553 182451 530562
rect 182503 530553 182515 530605
rect 182567 530596 186077 530605
rect 182575 530562 182633 530596
rect 182667 530562 182725 530596
rect 182759 530562 182817 530596
rect 182851 530562 182909 530596
rect 182943 530562 183001 530596
rect 183035 530562 183093 530596
rect 183127 530562 183185 530596
rect 183219 530562 183277 530596
rect 183311 530562 183369 530596
rect 183403 530562 183461 530596
rect 183495 530562 183553 530596
rect 183587 530562 183645 530596
rect 183679 530562 183737 530596
rect 183771 530562 183829 530596
rect 183863 530562 183921 530596
rect 183955 530562 184013 530596
rect 184047 530562 184105 530596
rect 184139 530562 184197 530596
rect 184231 530562 184289 530596
rect 184323 530562 184381 530596
rect 184415 530562 184473 530596
rect 184507 530562 184565 530596
rect 184599 530562 184657 530596
rect 184691 530562 184749 530596
rect 184783 530562 184841 530596
rect 184875 530562 184933 530596
rect 184967 530562 185025 530596
rect 185059 530562 185117 530596
rect 185151 530562 185209 530596
rect 185243 530562 185301 530596
rect 185335 530562 185393 530596
rect 185427 530562 185485 530596
rect 185519 530562 185577 530596
rect 185611 530562 185669 530596
rect 185703 530562 185761 530596
rect 185795 530562 185853 530596
rect 185887 530562 185945 530596
rect 185979 530562 186037 530596
rect 186071 530562 186077 530596
rect 182567 530553 186077 530562
rect 186129 530596 186141 530605
rect 186129 530553 186141 530562
rect 186193 530553 186205 530605
rect 186257 530553 186269 530605
rect 186321 530596 186333 530605
rect 186385 530596 187480 530605
rect 186385 530562 186405 530596
rect 186439 530562 186497 530596
rect 186531 530562 186589 530596
rect 186623 530562 186681 530596
rect 186715 530562 186773 530596
rect 186807 530562 186865 530596
rect 186899 530562 186957 530596
rect 186991 530562 187049 530596
rect 187083 530562 187141 530596
rect 187175 530562 187233 530596
rect 187267 530562 187325 530596
rect 187359 530562 187417 530596
rect 187451 530562 187480 530596
rect 186321 530553 186333 530562
rect 186385 530553 187480 530562
rect 172208 530531 187480 530553
rect 176822 530491 176828 530503
rect 176656 530463 176828 530491
rect 172406 530383 172412 530435
rect 172464 530423 172470 530435
rect 172501 530426 172559 530432
rect 172501 530423 172513 530426
rect 172464 530395 172513 530423
rect 172464 530383 172470 530395
rect 172501 530392 172513 530395
rect 172547 530392 172559 530426
rect 172501 530386 172559 530392
rect 174522 530383 174528 530435
rect 174580 530423 174586 530435
rect 174893 530426 174951 530432
rect 174893 530423 174905 530426
rect 174580 530395 174905 530423
rect 174580 530383 174586 530395
rect 174893 530392 174905 530395
rect 174939 530392 174951 530426
rect 174893 530386 174951 530392
rect 175833 530426 175891 530432
rect 175833 530392 175845 530426
rect 175879 530423 175891 530426
rect 176481 530426 176611 530432
rect 176481 530423 176493 530426
rect 175879 530395 176493 530423
rect 175879 530392 175951 530395
rect 175833 530386 175951 530392
rect 176481 530392 176493 530395
rect 176527 530392 176565 530426
rect 176599 530423 176611 530426
rect 176656 530423 176684 530463
rect 176822 530451 176828 530463
rect 176880 530451 176886 530503
rect 178754 530451 178760 530503
rect 178812 530451 178818 530503
rect 179401 530494 179459 530500
rect 179401 530491 179413 530494
rect 178864 530463 179413 530491
rect 176599 530395 176684 530423
rect 176599 530392 176611 530395
rect 176481 530386 176611 530392
rect 172869 530358 172927 530364
rect 172869 530324 172881 530358
rect 172915 530355 172927 530358
rect 174798 530355 174804 530367
rect 172915 530327 174804 530355
rect 172915 530324 172927 530327
rect 172869 530318 172927 530324
rect 174798 530315 174804 530327
rect 174856 530315 174862 530367
rect 175261 530358 175319 530364
rect 175261 530324 175273 530358
rect 175307 530355 175319 530358
rect 175442 530355 175448 530367
rect 175307 530327 175448 530355
rect 175307 530324 175319 530327
rect 175261 530318 175319 530324
rect 175442 530315 175448 530327
rect 175500 530315 175506 530367
rect 175893 530363 175951 530386
rect 176730 530383 176736 530435
rect 176788 530423 176794 530435
rect 178864 530423 178892 530463
rect 179401 530460 179413 530463
rect 179447 530460 179459 530494
rect 179401 530454 179459 530460
rect 179490 530451 179496 530503
rect 179548 530491 179554 530503
rect 180689 530494 180747 530500
rect 180689 530491 180701 530494
rect 179548 530463 180701 530491
rect 179548 530451 179554 530463
rect 180689 530460 180701 530463
rect 180735 530460 180747 530494
rect 180689 530454 180747 530460
rect 176788 530395 178892 530423
rect 180704 530423 180732 530454
rect 182986 530451 182992 530503
rect 183044 530491 183050 530503
rect 183265 530494 183323 530500
rect 183265 530491 183277 530494
rect 183044 530463 183277 530491
rect 183044 530451 183050 530463
rect 183265 530460 183277 530463
rect 183311 530460 183323 530494
rect 183265 530454 183323 530460
rect 185102 530451 185108 530503
rect 185160 530491 185166 530503
rect 185381 530494 185439 530500
rect 185381 530491 185393 530494
rect 185160 530463 185393 530491
rect 185160 530451 185166 530463
rect 185381 530460 185393 530463
rect 185427 530460 185439 530494
rect 185381 530454 185439 530460
rect 182069 530426 182127 530432
rect 182069 530423 182081 530426
rect 180704 530395 182081 530423
rect 176788 530383 176794 530395
rect 182069 530392 182081 530395
rect 182115 530392 182127 530426
rect 185289 530426 185347 530432
rect 185289 530423 185301 530426
rect 182069 530386 182127 530392
rect 182636 530395 185301 530423
rect 175893 530329 175905 530363
rect 175939 530329 175951 530363
rect 175893 530323 175951 530329
rect 176109 530358 176167 530364
rect 176109 530324 176121 530358
rect 176155 530355 176167 530358
rect 176825 530358 176883 530364
rect 176825 530355 176837 530358
rect 176155 530327 176837 530355
rect 176155 530324 176167 530327
rect 176109 530318 176167 530324
rect 176825 530324 176837 530327
rect 176871 530355 176883 530358
rect 177192 530358 177250 530364
rect 177192 530355 177204 530358
rect 176871 530327 177204 530355
rect 176871 530324 176883 530327
rect 176825 530318 176883 530324
rect 177192 530324 177204 530327
rect 177238 530324 177250 530358
rect 177192 530318 177250 530324
rect 178573 530358 178631 530364
rect 178573 530324 178585 530358
rect 178619 530355 178631 530358
rect 178938 530355 178944 530367
rect 178619 530327 178944 530355
rect 178619 530324 178631 530327
rect 178573 530318 178631 530324
rect 178938 530315 178944 530327
rect 178996 530315 179002 530367
rect 179033 530358 179091 530364
rect 179033 530324 179045 530358
rect 179079 530355 179091 530358
rect 179214 530355 179220 530367
rect 179079 530327 179220 530355
rect 179079 530324 179091 530327
rect 179033 530318 179091 530324
rect 179214 530315 179220 530327
rect 179272 530315 179278 530367
rect 179309 530358 179367 530364
rect 179309 530324 179321 530358
rect 179355 530324 179367 530358
rect 179309 530318 179367 530324
rect 180597 530358 180655 530364
rect 180597 530324 180609 530358
rect 180643 530355 180655 530358
rect 181517 530358 181575 530364
rect 180643 530327 181468 530355
rect 180643 530324 180655 530327
rect 180597 530318 180655 530324
rect 174816 530287 174844 530315
rect 175537 530290 175595 530296
rect 175537 530287 175549 530290
rect 174816 530259 175549 530287
rect 175537 530256 175549 530259
rect 175583 530256 175595 530290
rect 175537 530250 175595 530256
rect 176638 530247 176644 530299
rect 176696 530287 176702 530299
rect 177009 530290 177067 530296
rect 177009 530287 177021 530290
rect 176696 530259 177021 530287
rect 176696 530247 176702 530259
rect 177009 530256 177021 530259
rect 177055 530256 177067 530290
rect 177009 530250 177067 530256
rect 177282 530247 177288 530299
rect 177340 530247 177346 530299
rect 178202 530247 178208 530299
rect 178260 530287 178266 530299
rect 179324 530287 179352 530318
rect 178260 530259 179352 530287
rect 178260 530247 178266 530259
rect 180686 530247 180692 530299
rect 180744 530287 180750 530299
rect 181440 530296 181468 530327
rect 181517 530324 181529 530358
rect 181563 530355 181575 530358
rect 182250 530355 182256 530367
rect 181563 530327 182256 530355
rect 181563 530324 181575 530327
rect 181517 530318 181575 530324
rect 182250 530315 182256 530327
rect 182308 530355 182314 530367
rect 182636 530355 182664 530395
rect 185289 530392 185301 530395
rect 185335 530392 185347 530426
rect 185289 530386 185347 530392
rect 182308 530327 182664 530355
rect 182308 530315 182314 530327
rect 183170 530315 183176 530367
rect 183228 530315 183234 530367
rect 187126 530315 187132 530367
rect 187184 530315 187190 530367
rect 180781 530290 180839 530296
rect 180781 530287 180793 530290
rect 180744 530259 180793 530287
rect 180744 530247 180750 530259
rect 180781 530256 180793 530259
rect 180827 530287 180839 530290
rect 181241 530290 181299 530296
rect 181241 530287 181253 530290
rect 180827 530259 181253 530287
rect 180827 530256 180839 530259
rect 180781 530250 180839 530256
rect 181241 530256 181253 530259
rect 181287 530256 181299 530290
rect 181241 530250 181299 530256
rect 181425 530290 181483 530296
rect 181425 530256 181437 530290
rect 181471 530287 181483 530290
rect 182618 530287 182624 530299
rect 181471 530259 182624 530287
rect 181471 530256 181483 530259
rect 181425 530250 181483 530256
rect 182618 530247 182624 530259
rect 182676 530247 182682 530299
rect 176109 530222 176167 530228
rect 176109 530188 176121 530222
rect 176155 530219 176167 530222
rect 176733 530222 176791 530228
rect 176733 530219 176745 530222
rect 176155 530191 176745 530219
rect 176155 530188 176167 530191
rect 176109 530182 176167 530188
rect 176733 530188 176745 530191
rect 176779 530219 176791 530222
rect 177111 530222 177169 530228
rect 177111 530219 177123 530222
rect 176779 530191 177123 530219
rect 176779 530188 176791 530191
rect 176733 530182 176791 530188
rect 177111 530188 177123 530191
rect 177157 530188 177169 530222
rect 177111 530182 177169 530188
rect 181885 530222 181943 530228
rect 181885 530188 181897 530222
rect 181931 530219 181943 530222
rect 181931 530191 182756 530219
rect 181931 530188 181943 530191
rect 181885 530182 181943 530188
rect 182728 530163 182756 530191
rect 177650 530111 177656 530163
rect 177708 530111 177714 530163
rect 178294 530111 178300 530163
rect 178352 530151 178358 530163
rect 178389 530154 178447 530160
rect 178389 530151 178401 530154
rect 178352 530123 178401 530151
rect 178352 530111 178358 530123
rect 178389 530120 178401 530123
rect 178435 530120 178447 530154
rect 178389 530114 178447 530120
rect 179674 530111 179680 530163
rect 179732 530151 179738 530163
rect 180229 530154 180287 530160
rect 180229 530151 180241 530154
rect 179732 530123 180241 530151
rect 179732 530111 179738 530123
rect 180229 530120 180241 530123
rect 180275 530120 180287 530154
rect 180229 530114 180287 530120
rect 182158 530111 182164 530163
rect 182216 530111 182222 530163
rect 182710 530111 182716 530163
rect 182768 530111 182774 530163
rect 172208 530061 187480 530083
rect 172208 530052 173963 530061
rect 174015 530052 174027 530061
rect 174079 530052 174091 530061
rect 172208 530018 172237 530052
rect 172271 530018 172329 530052
rect 172363 530018 172421 530052
rect 172455 530018 172513 530052
rect 172547 530018 172605 530052
rect 172639 530018 172697 530052
rect 172731 530018 172789 530052
rect 172823 530018 172881 530052
rect 172915 530018 172973 530052
rect 173007 530018 173065 530052
rect 173099 530018 173157 530052
rect 173191 530018 173249 530052
rect 173283 530018 173341 530052
rect 173375 530018 173433 530052
rect 173467 530018 173525 530052
rect 173559 530018 173617 530052
rect 173651 530018 173709 530052
rect 173743 530018 173801 530052
rect 173835 530018 173893 530052
rect 173927 530018 173963 530052
rect 174019 530018 174027 530052
rect 172208 530009 173963 530018
rect 174015 530009 174027 530018
rect 174079 530009 174091 530018
rect 174143 530009 174155 530061
rect 174207 530009 174219 530061
rect 174271 530052 177781 530061
rect 174295 530018 174353 530052
rect 174387 530018 174445 530052
rect 174479 530018 174537 530052
rect 174571 530018 174629 530052
rect 174663 530018 174721 530052
rect 174755 530018 174813 530052
rect 174847 530018 174905 530052
rect 174939 530018 174997 530052
rect 175031 530018 175089 530052
rect 175123 530018 175181 530052
rect 175215 530018 175273 530052
rect 175307 530018 175365 530052
rect 175399 530018 175457 530052
rect 175491 530018 175549 530052
rect 175583 530018 175641 530052
rect 175675 530018 175733 530052
rect 175767 530018 175825 530052
rect 175859 530018 175917 530052
rect 175951 530018 176009 530052
rect 176043 530018 176101 530052
rect 176135 530018 176193 530052
rect 176227 530018 176285 530052
rect 176319 530018 176377 530052
rect 176411 530018 176469 530052
rect 176503 530018 176561 530052
rect 176595 530018 176653 530052
rect 176687 530018 176745 530052
rect 176779 530018 176837 530052
rect 176871 530018 176929 530052
rect 176963 530018 177021 530052
rect 177055 530018 177113 530052
rect 177147 530018 177205 530052
rect 177239 530018 177297 530052
rect 177331 530018 177389 530052
rect 177423 530018 177481 530052
rect 177515 530018 177573 530052
rect 177607 530018 177665 530052
rect 177699 530018 177757 530052
rect 174271 530009 177781 530018
rect 177833 530009 177845 530061
rect 177897 530009 177909 530061
rect 177961 530052 177973 530061
rect 178025 530052 178037 530061
rect 178089 530052 181599 530061
rect 181651 530052 181663 530061
rect 181715 530052 181727 530061
rect 178025 530018 178033 530052
rect 178089 530018 178125 530052
rect 178159 530018 178217 530052
rect 178251 530018 178309 530052
rect 178343 530018 178401 530052
rect 178435 530018 178493 530052
rect 178527 530018 178585 530052
rect 178619 530018 178677 530052
rect 178711 530018 178769 530052
rect 178803 530018 178861 530052
rect 178895 530018 178953 530052
rect 178987 530018 179045 530052
rect 179079 530018 179137 530052
rect 179171 530018 179229 530052
rect 179263 530018 179321 530052
rect 179355 530018 179413 530052
rect 179447 530018 179505 530052
rect 179539 530018 179597 530052
rect 179631 530018 179689 530052
rect 179723 530018 179781 530052
rect 179815 530018 179873 530052
rect 179907 530018 179965 530052
rect 179999 530018 180057 530052
rect 180091 530018 180149 530052
rect 180183 530018 180241 530052
rect 180275 530018 180333 530052
rect 180367 530018 180425 530052
rect 180459 530018 180517 530052
rect 180551 530018 180609 530052
rect 180643 530018 180701 530052
rect 180735 530018 180793 530052
rect 180827 530018 180885 530052
rect 180919 530018 180977 530052
rect 181011 530018 181069 530052
rect 181103 530018 181161 530052
rect 181195 530018 181253 530052
rect 181287 530018 181345 530052
rect 181379 530018 181437 530052
rect 181471 530018 181529 530052
rect 181563 530018 181599 530052
rect 181655 530018 181663 530052
rect 177961 530009 177973 530018
rect 178025 530009 178037 530018
rect 178089 530009 181599 530018
rect 181651 530009 181663 530018
rect 181715 530009 181727 530018
rect 181779 530009 181791 530061
rect 181843 530009 181855 530061
rect 181907 530052 185417 530061
rect 181931 530018 181989 530052
rect 182023 530018 182081 530052
rect 182115 530018 182173 530052
rect 182207 530018 182265 530052
rect 182299 530018 182357 530052
rect 182391 530018 182449 530052
rect 182483 530018 182541 530052
rect 182575 530018 182633 530052
rect 182667 530018 182725 530052
rect 182759 530018 182817 530052
rect 182851 530018 182909 530052
rect 182943 530018 183001 530052
rect 183035 530018 183093 530052
rect 183127 530018 183185 530052
rect 183219 530018 183277 530052
rect 183311 530018 183369 530052
rect 183403 530018 183461 530052
rect 183495 530018 183553 530052
rect 183587 530018 183645 530052
rect 183679 530018 183737 530052
rect 183771 530018 183829 530052
rect 183863 530018 183921 530052
rect 183955 530018 184013 530052
rect 184047 530018 184105 530052
rect 184139 530018 184197 530052
rect 184231 530018 184289 530052
rect 184323 530018 184381 530052
rect 184415 530018 184473 530052
rect 184507 530018 184565 530052
rect 184599 530018 184657 530052
rect 184691 530018 184749 530052
rect 184783 530018 184841 530052
rect 184875 530018 184933 530052
rect 184967 530018 185025 530052
rect 185059 530018 185117 530052
rect 185151 530018 185209 530052
rect 185243 530018 185301 530052
rect 185335 530018 185393 530052
rect 181907 530009 185417 530018
rect 185469 530009 185481 530061
rect 185533 530009 185545 530061
rect 185597 530052 185609 530061
rect 185661 530052 185673 530061
rect 185725 530052 187480 530061
rect 185661 530018 185669 530052
rect 185725 530018 185761 530052
rect 185795 530018 185853 530052
rect 185887 530018 185945 530052
rect 185979 530018 186037 530052
rect 186071 530018 186129 530052
rect 186163 530018 186221 530052
rect 186255 530018 186313 530052
rect 186347 530018 186405 530052
rect 186439 530018 186497 530052
rect 186531 530018 186589 530052
rect 186623 530018 186681 530052
rect 186715 530018 186773 530052
rect 186807 530018 186865 530052
rect 186899 530018 186957 530052
rect 186991 530018 187049 530052
rect 187083 530018 187141 530052
rect 187175 530018 187233 530052
rect 187267 530018 187325 530052
rect 187359 530018 187417 530052
rect 187451 530018 187480 530052
rect 185597 530009 185609 530018
rect 185661 530009 185673 530018
rect 185725 530009 187480 530018
rect 172208 529987 187480 530009
rect 177285 529950 177343 529956
rect 177285 529916 177297 529950
rect 177331 529947 177343 529950
rect 178202 529947 178208 529959
rect 177331 529919 178208 529947
rect 177331 529916 177343 529919
rect 177285 529910 177343 529916
rect 178202 529907 178208 529919
rect 178260 529907 178266 529959
rect 178389 529950 178447 529956
rect 178389 529916 178401 529950
rect 178435 529947 178447 529950
rect 179490 529947 179496 529959
rect 178435 529919 179496 529947
rect 178435 529916 178447 529919
rect 178389 529910 178447 529916
rect 179490 529907 179496 529919
rect 179548 529907 179554 529959
rect 180870 529907 180876 529959
rect 180928 529947 180934 529959
rect 182158 529947 182164 529959
rect 180928 529919 182164 529947
rect 180928 529907 180934 529919
rect 182158 529907 182164 529919
rect 182216 529907 182222 529959
rect 182618 529907 182624 529959
rect 182676 529907 182682 529959
rect 175711 529882 175769 529888
rect 175711 529848 175723 529882
rect 175757 529879 175769 529882
rect 176089 529882 176147 529888
rect 176089 529879 176101 529882
rect 175757 529851 176101 529879
rect 175757 529848 175769 529851
rect 175711 529842 175769 529848
rect 176089 529848 176101 529851
rect 176135 529879 176147 529882
rect 176713 529882 176771 529888
rect 176713 529879 176725 529882
rect 176135 529851 176725 529879
rect 176135 529848 176147 529851
rect 176089 529842 176147 529848
rect 176713 529848 176725 529851
rect 176759 529848 176771 529882
rect 176713 529842 176771 529848
rect 178110 529839 178116 529891
rect 178168 529879 178174 529891
rect 178297 529882 178355 529888
rect 178297 529879 178309 529882
rect 178168 529851 178309 529879
rect 178168 529839 178174 529851
rect 178297 529848 178309 529851
rect 178343 529848 178355 529882
rect 178297 529842 178355 529848
rect 178961 529882 179019 529888
rect 178961 529848 178973 529882
rect 179007 529879 179019 529882
rect 179585 529882 179643 529888
rect 179585 529879 179597 529882
rect 179007 529851 179597 529879
rect 179007 529848 179019 529851
rect 178961 529842 179019 529848
rect 179585 529848 179597 529851
rect 179631 529879 179643 529882
rect 179963 529882 180021 529888
rect 179963 529879 179975 529882
rect 179631 529851 179975 529879
rect 179631 529848 179643 529851
rect 179585 529842 179643 529848
rect 179963 529848 179975 529851
rect 180009 529848 180021 529882
rect 179963 529842 180021 529848
rect 180403 529882 180461 529888
rect 180403 529848 180415 529882
rect 180449 529879 180461 529882
rect 180781 529882 180839 529888
rect 180781 529879 180793 529882
rect 180449 529851 180793 529879
rect 180449 529848 180461 529851
rect 180403 529842 180461 529848
rect 180781 529848 180793 529851
rect 180827 529879 180839 529882
rect 181405 529882 181463 529888
rect 181405 529879 181417 529882
rect 180827 529851 181417 529879
rect 180827 529848 180839 529851
rect 180781 529842 180839 529848
rect 181405 529848 181417 529851
rect 181451 529848 181463 529882
rect 181405 529842 181463 529848
rect 174798 529771 174804 529823
rect 174856 529771 174862 529823
rect 175813 529814 175871 529820
rect 175813 529780 175825 529814
rect 175859 529811 175871 529814
rect 177653 529814 177711 529820
rect 177653 529811 177665 529814
rect 175859 529783 177420 529811
rect 175859 529780 175871 529783
rect 175813 529774 175871 529780
rect 175537 529746 175595 529752
rect 175537 529712 175549 529746
rect 175583 529712 175595 529746
rect 175537 529706 175595 529712
rect 175630 529746 175688 529752
rect 175630 529712 175642 529746
rect 175676 529743 175688 529746
rect 175997 529746 176055 529752
rect 175997 529743 176009 529746
rect 175676 529715 176009 529743
rect 175676 529712 175688 529715
rect 175630 529706 175688 529712
rect 175997 529712 176009 529715
rect 176043 529743 176055 529746
rect 176713 529746 176771 529752
rect 176713 529743 176725 529746
rect 176043 529715 176725 529743
rect 176043 529712 176055 529715
rect 175997 529706 176055 529712
rect 176713 529712 176725 529715
rect 176759 529712 176771 529746
rect 176713 529706 176771 529712
rect 175552 529675 175580 529706
rect 176822 529703 176828 529755
rect 176880 529743 176886 529755
rect 176929 529743 176987 529747
rect 176880 529741 176987 529743
rect 176880 529715 176941 529741
rect 176880 529703 176886 529715
rect 176929 529707 176941 529715
rect 176975 529707 176987 529741
rect 176929 529684 176987 529707
rect 177392 529687 177420 529783
rect 177576 529783 177665 529811
rect 177576 529687 177604 529783
rect 177653 529780 177665 529783
rect 177699 529780 177711 529814
rect 179306 529811 179312 529823
rect 177653 529774 177711 529780
rect 177944 529783 179312 529811
rect 177944 529752 177972 529783
rect 179306 529771 179312 529783
rect 179364 529771 179370 529823
rect 179858 529771 179864 529823
rect 179916 529771 179922 529823
rect 180505 529814 180563 529820
rect 180505 529780 180517 529814
rect 180551 529811 180563 529814
rect 181977 529814 182035 529820
rect 180551 529783 181836 529811
rect 180551 529780 180563 529783
rect 180505 529774 180563 529780
rect 177929 529746 177987 529752
rect 177929 529712 177941 529746
rect 177975 529712 177987 529746
rect 177929 529706 177987 529712
rect 178745 529741 178803 529747
rect 178745 529707 178757 529741
rect 178791 529707 178803 529741
rect 176269 529678 176399 529684
rect 175552 529647 176132 529675
rect 176104 529619 176132 529647
rect 176269 529644 176281 529678
rect 176315 529644 176353 529678
rect 176387 529675 176399 529678
rect 176929 529678 177047 529684
rect 176929 529675 177001 529678
rect 176387 529647 177001 529675
rect 176387 529644 176399 529647
rect 176269 529638 176399 529644
rect 175350 529567 175356 529619
rect 175408 529607 175414 529619
rect 175445 529610 175503 529616
rect 175445 529607 175457 529610
rect 175408 529579 175457 529607
rect 175408 529567 175414 529579
rect 175445 529576 175457 529579
rect 175491 529576 175503 529610
rect 175445 529570 175503 529576
rect 176086 529567 176092 529619
rect 176144 529567 176150 529619
rect 176932 529607 176960 529647
rect 176989 529644 177001 529647
rect 177035 529644 177047 529678
rect 176989 529638 177047 529644
rect 177374 529635 177380 529687
rect 177432 529635 177438 529687
rect 177558 529635 177564 529687
rect 177616 529635 177622 529687
rect 177650 529635 177656 529687
rect 177708 529675 177714 529687
rect 178745 529684 178803 529707
rect 178961 529746 179019 529752
rect 178961 529712 178973 529746
rect 179007 529743 179019 529746
rect 179677 529746 179735 529752
rect 179677 529743 179689 529746
rect 179007 529715 179689 529743
rect 179007 529712 179019 529715
rect 178961 529706 179019 529712
rect 179677 529712 179689 529715
rect 179723 529743 179735 529746
rect 180044 529746 180102 529752
rect 180044 529743 180056 529746
rect 179723 529715 180056 529743
rect 179723 529712 179735 529715
rect 179677 529706 179735 529712
rect 180044 529712 180056 529715
rect 180090 529712 180102 529746
rect 180044 529706 180102 529712
rect 180137 529746 180195 529752
rect 180137 529712 180149 529746
rect 180183 529743 180195 529746
rect 180229 529746 180287 529752
rect 180229 529743 180241 529746
rect 180183 529715 180241 529743
rect 180183 529712 180195 529715
rect 180137 529706 180195 529712
rect 180229 529712 180241 529715
rect 180275 529712 180287 529746
rect 180229 529706 180287 529712
rect 180322 529746 180380 529752
rect 180322 529712 180334 529746
rect 180368 529743 180380 529746
rect 180689 529746 180747 529752
rect 180689 529743 180701 529746
rect 180368 529715 180701 529743
rect 180368 529712 180380 529715
rect 180322 529706 180380 529712
rect 180689 529712 180701 529715
rect 180735 529743 180747 529746
rect 181405 529746 181463 529752
rect 181405 529743 181417 529746
rect 180735 529715 181417 529743
rect 180735 529712 180747 529715
rect 180689 529706 180747 529712
rect 181405 529712 181417 529715
rect 181451 529712 181463 529746
rect 181405 529706 181463 529712
rect 181621 529741 181679 529747
rect 181621 529707 181633 529741
rect 181667 529707 181679 529741
rect 177837 529678 177895 529684
rect 177837 529675 177849 529678
rect 177708 529647 177849 529675
rect 177708 529635 177714 529647
rect 177837 529644 177849 529647
rect 177883 529644 177895 529678
rect 178685 529678 178803 529684
rect 178685 529675 178697 529678
rect 177837 529638 177895 529644
rect 178404 529647 178697 529675
rect 177926 529607 177932 529619
rect 176932 529579 177932 529607
rect 177926 529567 177932 529579
rect 177984 529607 177990 529619
rect 178404 529607 178432 529647
rect 178685 529644 178697 529647
rect 178731 529675 178803 529678
rect 179333 529678 179463 529684
rect 179333 529675 179345 529678
rect 178731 529647 179345 529675
rect 178731 529644 178743 529647
rect 178685 529638 178743 529644
rect 179333 529644 179345 529647
rect 179379 529644 179417 529678
rect 179451 529644 179463 529678
rect 180244 529675 180272 529706
rect 180961 529678 181091 529684
rect 180244 529647 180548 529675
rect 179333 529638 179463 529644
rect 180520 529619 180548 529647
rect 180961 529644 180973 529678
rect 181007 529644 181045 529678
rect 181079 529675 181091 529678
rect 181514 529675 181520 529687
rect 181079 529647 181520 529675
rect 181079 529644 181091 529647
rect 180961 529638 181091 529644
rect 181514 529635 181520 529647
rect 181572 529675 181578 529687
rect 181621 529684 181679 529707
rect 181621 529678 181739 529684
rect 181621 529675 181693 529678
rect 181572 529647 181693 529675
rect 181572 529635 181578 529647
rect 181681 529644 181693 529647
rect 181727 529644 181739 529678
rect 181681 529638 181739 529644
rect 181808 529619 181836 529783
rect 181977 529780 181989 529814
rect 182023 529811 182035 529814
rect 183170 529811 183176 529823
rect 182023 529783 183176 529811
rect 182023 529780 182035 529783
rect 181977 529774 182035 529780
rect 183170 529771 183176 529783
rect 183228 529771 183234 529823
rect 177984 529579 178432 529607
rect 177984 529567 177990 529579
rect 180502 529567 180508 529619
rect 180560 529567 180566 529619
rect 181790 529567 181796 529619
rect 181848 529567 181854 529619
rect 172208 529517 187480 529539
rect 172208 529508 174623 529517
rect 172208 529474 172237 529508
rect 172271 529474 172329 529508
rect 172363 529474 172421 529508
rect 172455 529474 172513 529508
rect 172547 529474 172605 529508
rect 172639 529474 172697 529508
rect 172731 529474 172789 529508
rect 172823 529474 172881 529508
rect 172915 529474 172973 529508
rect 173007 529474 173065 529508
rect 173099 529474 173157 529508
rect 173191 529474 173249 529508
rect 173283 529474 173341 529508
rect 173375 529474 173433 529508
rect 173467 529474 173525 529508
rect 173559 529474 173617 529508
rect 173651 529474 173709 529508
rect 173743 529474 173801 529508
rect 173835 529474 173893 529508
rect 173927 529474 173985 529508
rect 174019 529474 174077 529508
rect 174111 529474 174169 529508
rect 174203 529474 174261 529508
rect 174295 529474 174353 529508
rect 174387 529474 174445 529508
rect 174479 529474 174537 529508
rect 174571 529474 174623 529508
rect 172208 529465 174623 529474
rect 174675 529465 174687 529517
rect 174739 529508 174751 529517
rect 174803 529508 174815 529517
rect 174803 529474 174813 529508
rect 174739 529465 174751 529474
rect 174803 529465 174815 529474
rect 174867 529465 174879 529517
rect 174931 529508 178441 529517
rect 174939 529474 174997 529508
rect 175031 529474 175089 529508
rect 175123 529474 175181 529508
rect 175215 529474 175273 529508
rect 175307 529474 175365 529508
rect 175399 529474 175457 529508
rect 175491 529474 175549 529508
rect 175583 529474 175641 529508
rect 175675 529474 175733 529508
rect 175767 529474 175825 529508
rect 175859 529474 175917 529508
rect 175951 529474 176009 529508
rect 176043 529474 176101 529508
rect 176135 529474 176193 529508
rect 176227 529474 176285 529508
rect 176319 529474 176377 529508
rect 176411 529474 176469 529508
rect 176503 529474 176561 529508
rect 176595 529474 176653 529508
rect 176687 529474 176745 529508
rect 176779 529474 176837 529508
rect 176871 529474 176929 529508
rect 176963 529474 177021 529508
rect 177055 529474 177113 529508
rect 177147 529474 177205 529508
rect 177239 529474 177297 529508
rect 177331 529474 177389 529508
rect 177423 529474 177481 529508
rect 177515 529474 177573 529508
rect 177607 529474 177665 529508
rect 177699 529474 177757 529508
rect 177791 529474 177849 529508
rect 177883 529474 177941 529508
rect 177975 529474 178033 529508
rect 178067 529474 178125 529508
rect 178159 529474 178217 529508
rect 178251 529474 178309 529508
rect 178343 529474 178401 529508
rect 178435 529474 178441 529508
rect 174931 529465 178441 529474
rect 178493 529508 178505 529517
rect 178493 529465 178505 529474
rect 178557 529465 178569 529517
rect 178621 529465 178633 529517
rect 178685 529508 178697 529517
rect 178749 529508 182259 529517
rect 178749 529474 178769 529508
rect 178803 529474 178861 529508
rect 178895 529474 178953 529508
rect 178987 529474 179045 529508
rect 179079 529474 179137 529508
rect 179171 529474 179229 529508
rect 179263 529474 179321 529508
rect 179355 529474 179413 529508
rect 179447 529474 179505 529508
rect 179539 529474 179597 529508
rect 179631 529474 179689 529508
rect 179723 529474 179781 529508
rect 179815 529474 179873 529508
rect 179907 529474 179965 529508
rect 179999 529474 180057 529508
rect 180091 529474 180149 529508
rect 180183 529474 180241 529508
rect 180275 529474 180333 529508
rect 180367 529474 180425 529508
rect 180459 529474 180517 529508
rect 180551 529474 180609 529508
rect 180643 529474 180701 529508
rect 180735 529474 180793 529508
rect 180827 529474 180885 529508
rect 180919 529474 180977 529508
rect 181011 529474 181069 529508
rect 181103 529474 181161 529508
rect 181195 529474 181253 529508
rect 181287 529474 181345 529508
rect 181379 529474 181437 529508
rect 181471 529474 181529 529508
rect 181563 529474 181621 529508
rect 181655 529474 181713 529508
rect 181747 529474 181805 529508
rect 181839 529474 181897 529508
rect 181931 529474 181989 529508
rect 182023 529474 182081 529508
rect 182115 529474 182173 529508
rect 182207 529474 182259 529508
rect 178685 529465 178697 529474
rect 178749 529465 182259 529474
rect 182311 529465 182323 529517
rect 182375 529508 182387 529517
rect 182439 529508 182451 529517
rect 182439 529474 182449 529508
rect 182375 529465 182387 529474
rect 182439 529465 182451 529474
rect 182503 529465 182515 529517
rect 182567 529508 186077 529517
rect 182575 529474 182633 529508
rect 182667 529474 182725 529508
rect 182759 529474 182817 529508
rect 182851 529474 182909 529508
rect 182943 529474 183001 529508
rect 183035 529474 183093 529508
rect 183127 529474 183185 529508
rect 183219 529474 183277 529508
rect 183311 529474 183369 529508
rect 183403 529474 183461 529508
rect 183495 529474 183553 529508
rect 183587 529474 183645 529508
rect 183679 529474 183737 529508
rect 183771 529474 183829 529508
rect 183863 529474 183921 529508
rect 183955 529474 184013 529508
rect 184047 529474 184105 529508
rect 184139 529474 184197 529508
rect 184231 529474 184289 529508
rect 184323 529474 184381 529508
rect 184415 529474 184473 529508
rect 184507 529474 184565 529508
rect 184599 529474 184657 529508
rect 184691 529474 184749 529508
rect 184783 529474 184841 529508
rect 184875 529474 184933 529508
rect 184967 529474 185025 529508
rect 185059 529474 185117 529508
rect 185151 529474 185209 529508
rect 185243 529474 185301 529508
rect 185335 529474 185393 529508
rect 185427 529474 185485 529508
rect 185519 529474 185577 529508
rect 185611 529474 185669 529508
rect 185703 529474 185761 529508
rect 185795 529474 185853 529508
rect 185887 529474 185945 529508
rect 185979 529474 186037 529508
rect 186071 529474 186077 529508
rect 182567 529465 186077 529474
rect 186129 529508 186141 529517
rect 186129 529465 186141 529474
rect 186193 529465 186205 529517
rect 186257 529465 186269 529517
rect 186321 529508 186333 529517
rect 186385 529508 187480 529517
rect 186385 529474 186405 529508
rect 186439 529474 186497 529508
rect 186531 529474 186589 529508
rect 186623 529474 186681 529508
rect 186715 529474 186773 529508
rect 186807 529474 186865 529508
rect 186899 529474 186957 529508
rect 186991 529474 187049 529508
rect 187083 529474 187141 529508
rect 187175 529474 187233 529508
rect 187267 529474 187325 529508
rect 187359 529474 187417 529508
rect 187451 529474 187480 529508
rect 186321 529465 186333 529474
rect 186385 529465 187480 529474
rect 172208 529443 187480 529465
rect 175350 529363 175356 529415
rect 175408 529363 175414 529415
rect 177926 529363 177932 529415
rect 177984 529403 177990 529415
rect 177984 529375 179352 529403
rect 177984 529363 177990 529375
rect 178021 529338 178079 529344
rect 178021 529304 178033 529338
rect 178067 529335 178079 529338
rect 178294 529335 178300 529347
rect 178067 529307 178300 529335
rect 178067 529304 178079 529307
rect 178021 529298 178079 529304
rect 178294 529295 178300 529307
rect 178352 529295 178358 529347
rect 178477 529338 178607 529344
rect 178477 529304 178489 529338
rect 178523 529304 178561 529338
rect 178595 529335 178607 529338
rect 179197 529338 179255 529344
rect 179197 529335 179209 529338
rect 178595 529307 179209 529335
rect 178595 529304 178607 529307
rect 178477 529298 178607 529304
rect 179137 529304 179209 529307
rect 179243 529335 179255 529338
rect 179324 529335 179352 529375
rect 179858 529363 179864 529415
rect 179916 529363 179922 529415
rect 181790 529363 181796 529415
rect 181848 529403 181854 529415
rect 182529 529406 182587 529412
rect 182529 529403 182541 529406
rect 181848 529375 182541 529403
rect 181848 529363 181854 529375
rect 182529 529372 182541 529375
rect 182575 529372 182587 529406
rect 182529 529366 182587 529372
rect 179243 529307 181560 529335
rect 179243 529304 179255 529307
rect 179137 529298 179255 529304
rect 175442 529227 175448 529279
rect 175500 529267 175506 529279
rect 176730 529267 176736 529279
rect 175500 529239 176736 529267
rect 175500 529227 175506 529239
rect 176730 529227 176736 529239
rect 176788 529227 176794 529279
rect 177650 529227 177656 529279
rect 177708 529227 177714 529279
rect 177838 529270 177896 529276
rect 177838 529236 177850 529270
rect 177884 529267 177896 529270
rect 178205 529270 178263 529276
rect 178205 529267 178217 529270
rect 177884 529239 178217 529267
rect 177884 529236 177896 529239
rect 177838 529230 177896 529236
rect 178205 529236 178217 529239
rect 178251 529267 178263 529270
rect 178921 529270 178979 529276
rect 178921 529267 178933 529270
rect 178251 529239 178933 529267
rect 178251 529236 178263 529239
rect 178205 529230 178263 529236
rect 178921 529236 178933 529239
rect 178967 529236 178979 529270
rect 178921 529230 178979 529236
rect 179137 529275 179195 529298
rect 181532 529279 181560 529307
rect 179137 529241 179149 529275
rect 179183 529241 179195 529275
rect 179137 529235 179195 529241
rect 179674 529227 179680 529279
rect 179732 529227 179738 529279
rect 180689 529270 180747 529276
rect 180689 529236 180701 529270
rect 180735 529236 180747 529270
rect 180689 529230 180747 529236
rect 173602 529159 173608 529211
rect 173660 529199 173666 529211
rect 175258 529199 175264 529211
rect 173660 529171 175264 529199
rect 173660 529159 173666 529171
rect 175258 529159 175264 529171
rect 175316 529159 175322 529211
rect 177282 529199 177288 529211
rect 176196 529171 177288 529199
rect 175813 529066 175871 529072
rect 175813 529032 175825 529066
rect 175859 529063 175871 529066
rect 175902 529063 175908 529075
rect 175859 529035 175908 529063
rect 175859 529032 175871 529035
rect 175813 529026 175871 529032
rect 175902 529023 175908 529035
rect 175960 529023 175966 529075
rect 176086 529023 176092 529075
rect 176144 529063 176150 529075
rect 176196 529072 176224 529171
rect 177282 529159 177288 529171
rect 177340 529199 177346 529211
rect 177745 529202 177803 529208
rect 177745 529199 177757 529202
rect 177340 529171 177757 529199
rect 177340 529159 177346 529171
rect 177745 529168 177757 529171
rect 177791 529168 177803 529202
rect 180704 529199 180732 529230
rect 181514 529227 181520 529279
rect 181572 529227 181578 529279
rect 182710 529227 182716 529279
rect 182768 529227 182774 529279
rect 177745 529162 177803 529168
rect 179692 529171 180732 529199
rect 177919 529134 177977 529140
rect 177919 529100 177931 529134
rect 177965 529131 177977 529134
rect 178297 529134 178355 529140
rect 178297 529131 178309 529134
rect 177965 529103 178309 529131
rect 177965 529100 177977 529103
rect 177919 529094 177977 529100
rect 178297 529100 178309 529103
rect 178343 529131 178355 529134
rect 178921 529134 178979 529140
rect 178921 529131 178933 529134
rect 178343 529103 178933 529131
rect 178343 529100 178355 529103
rect 178297 529094 178355 529100
rect 178921 529100 178933 529103
rect 178967 529100 178979 529134
rect 178921 529094 178979 529100
rect 179692 529075 179720 529171
rect 176181 529066 176239 529072
rect 176181 529063 176193 529066
rect 176144 529035 176193 529063
rect 176144 529023 176150 529035
rect 176181 529032 176193 529035
rect 176227 529032 176239 529066
rect 176181 529026 176239 529032
rect 179306 529023 179312 529075
rect 179364 529063 179370 529075
rect 179493 529066 179551 529072
rect 179493 529063 179505 529066
rect 179364 529035 179505 529063
rect 179364 529023 179370 529035
rect 179493 529032 179505 529035
rect 179539 529032 179551 529066
rect 179493 529026 179551 529032
rect 179674 529023 179680 529075
rect 179732 529023 179738 529075
rect 180502 529023 180508 529075
rect 180560 529063 180566 529075
rect 181977 529066 182035 529072
rect 181977 529063 181989 529066
rect 180560 529035 181989 529063
rect 180560 529023 180566 529035
rect 181977 529032 181989 529035
rect 182023 529032 182035 529066
rect 181977 529026 182035 529032
rect 172208 528973 187480 528995
rect 172208 528964 173963 528973
rect 174015 528964 174027 528973
rect 174079 528964 174091 528973
rect 172208 528930 172237 528964
rect 172271 528930 172329 528964
rect 172363 528930 172421 528964
rect 172455 528930 172513 528964
rect 172547 528930 172605 528964
rect 172639 528930 172697 528964
rect 172731 528930 172789 528964
rect 172823 528930 172881 528964
rect 172915 528930 172973 528964
rect 173007 528930 173065 528964
rect 173099 528930 173157 528964
rect 173191 528930 173249 528964
rect 173283 528930 173341 528964
rect 173375 528930 173433 528964
rect 173467 528930 173525 528964
rect 173559 528930 173617 528964
rect 173651 528930 173709 528964
rect 173743 528930 173801 528964
rect 173835 528930 173893 528964
rect 173927 528930 173963 528964
rect 174019 528930 174027 528964
rect 172208 528921 173963 528930
rect 174015 528921 174027 528930
rect 174079 528921 174091 528930
rect 174143 528921 174155 528973
rect 174207 528921 174219 528973
rect 174271 528964 177781 528973
rect 174295 528930 174353 528964
rect 174387 528930 174445 528964
rect 174479 528930 174537 528964
rect 174571 528930 174629 528964
rect 174663 528930 174721 528964
rect 174755 528930 174813 528964
rect 174847 528930 174905 528964
rect 174939 528930 174997 528964
rect 175031 528930 175089 528964
rect 175123 528930 175181 528964
rect 175215 528930 175273 528964
rect 175307 528930 175365 528964
rect 175399 528930 175457 528964
rect 175491 528930 175549 528964
rect 175583 528930 175641 528964
rect 175675 528930 175733 528964
rect 175767 528930 175825 528964
rect 175859 528930 175917 528964
rect 175951 528930 176009 528964
rect 176043 528930 176101 528964
rect 176135 528930 176193 528964
rect 176227 528930 176285 528964
rect 176319 528930 176377 528964
rect 176411 528930 176469 528964
rect 176503 528930 176561 528964
rect 176595 528930 176653 528964
rect 176687 528930 176745 528964
rect 176779 528930 176837 528964
rect 176871 528930 176929 528964
rect 176963 528930 177021 528964
rect 177055 528930 177113 528964
rect 177147 528930 177205 528964
rect 177239 528930 177297 528964
rect 177331 528930 177389 528964
rect 177423 528930 177481 528964
rect 177515 528930 177573 528964
rect 177607 528930 177665 528964
rect 177699 528930 177757 528964
rect 174271 528921 177781 528930
rect 177833 528921 177845 528973
rect 177897 528921 177909 528973
rect 177961 528964 177973 528973
rect 178025 528964 178037 528973
rect 178089 528964 181599 528973
rect 181651 528964 181663 528973
rect 181715 528964 181727 528973
rect 178025 528930 178033 528964
rect 178089 528930 178125 528964
rect 178159 528930 178217 528964
rect 178251 528930 178309 528964
rect 178343 528930 178401 528964
rect 178435 528930 178493 528964
rect 178527 528930 178585 528964
rect 178619 528930 178677 528964
rect 178711 528930 178769 528964
rect 178803 528930 178861 528964
rect 178895 528930 178953 528964
rect 178987 528930 179045 528964
rect 179079 528930 179137 528964
rect 179171 528930 179229 528964
rect 179263 528930 179321 528964
rect 179355 528930 179413 528964
rect 179447 528930 179505 528964
rect 179539 528930 179597 528964
rect 179631 528930 179689 528964
rect 179723 528930 179781 528964
rect 179815 528930 179873 528964
rect 179907 528930 179965 528964
rect 179999 528930 180057 528964
rect 180091 528930 180149 528964
rect 180183 528930 180241 528964
rect 180275 528930 180333 528964
rect 180367 528930 180425 528964
rect 180459 528930 180517 528964
rect 180551 528930 180609 528964
rect 180643 528930 180701 528964
rect 180735 528930 180793 528964
rect 180827 528930 180885 528964
rect 180919 528930 180977 528964
rect 181011 528930 181069 528964
rect 181103 528930 181161 528964
rect 181195 528930 181253 528964
rect 181287 528930 181345 528964
rect 181379 528930 181437 528964
rect 181471 528930 181529 528964
rect 181563 528930 181599 528964
rect 181655 528930 181663 528964
rect 177961 528921 177973 528930
rect 178025 528921 178037 528930
rect 178089 528921 181599 528930
rect 181651 528921 181663 528930
rect 181715 528921 181727 528930
rect 181779 528921 181791 528973
rect 181843 528921 181855 528973
rect 181907 528964 185417 528973
rect 181931 528930 181989 528964
rect 182023 528930 182081 528964
rect 182115 528930 182173 528964
rect 182207 528930 182265 528964
rect 182299 528930 182357 528964
rect 182391 528930 182449 528964
rect 182483 528930 182541 528964
rect 182575 528930 182633 528964
rect 182667 528930 182725 528964
rect 182759 528930 182817 528964
rect 182851 528930 182909 528964
rect 182943 528930 183001 528964
rect 183035 528930 183093 528964
rect 183127 528930 183185 528964
rect 183219 528930 183277 528964
rect 183311 528930 183369 528964
rect 183403 528930 183461 528964
rect 183495 528930 183553 528964
rect 183587 528930 183645 528964
rect 183679 528930 183737 528964
rect 183771 528930 183829 528964
rect 183863 528930 183921 528964
rect 183955 528930 184013 528964
rect 184047 528930 184105 528964
rect 184139 528930 184197 528964
rect 184231 528930 184289 528964
rect 184323 528930 184381 528964
rect 184415 528930 184473 528964
rect 184507 528930 184565 528964
rect 184599 528930 184657 528964
rect 184691 528930 184749 528964
rect 184783 528930 184841 528964
rect 184875 528930 184933 528964
rect 184967 528930 185025 528964
rect 185059 528930 185117 528964
rect 185151 528930 185209 528964
rect 185243 528930 185301 528964
rect 185335 528930 185393 528964
rect 181907 528921 185417 528930
rect 185469 528921 185481 528973
rect 185533 528921 185545 528973
rect 185597 528964 185609 528973
rect 185661 528964 185673 528973
rect 185725 528964 187480 528973
rect 185661 528930 185669 528964
rect 185725 528930 185761 528964
rect 185795 528930 185853 528964
rect 185887 528930 185945 528964
rect 185979 528930 186037 528964
rect 186071 528930 186129 528964
rect 186163 528930 186221 528964
rect 186255 528930 186313 528964
rect 186347 528930 186405 528964
rect 186439 528930 186497 528964
rect 186531 528930 186589 528964
rect 186623 528930 186681 528964
rect 186715 528930 186773 528964
rect 186807 528930 186865 528964
rect 186899 528930 186957 528964
rect 186991 528930 187049 528964
rect 187083 528930 187141 528964
rect 187175 528930 187233 528964
rect 187267 528930 187325 528964
rect 187359 528930 187417 528964
rect 187451 528930 187480 528964
rect 185597 528921 185609 528930
rect 185661 528921 185673 528930
rect 185725 528921 187480 528930
rect 172208 528899 187480 528921
rect 175258 528819 175264 528871
rect 175316 528819 175322 528871
rect 176089 528862 176147 528868
rect 176089 528828 176101 528862
rect 176135 528859 176147 528862
rect 176638 528859 176644 528871
rect 176135 528831 176644 528859
rect 176135 528828 176147 528831
rect 176089 528822 176147 528828
rect 176638 528819 176644 528831
rect 176696 528819 176702 528871
rect 177650 528819 177656 528871
rect 177708 528859 177714 528871
rect 179674 528859 179680 528871
rect 177708 528831 179680 528859
rect 177708 528819 177714 528831
rect 179674 528819 179680 528831
rect 179732 528819 179738 528871
rect 180428 528831 180640 528859
rect 175276 528723 175304 528819
rect 180428 528800 180456 528831
rect 180413 528794 180471 528800
rect 180413 528760 180425 528794
rect 180459 528760 180471 528794
rect 180413 528754 180471 528760
rect 176549 528726 176607 528732
rect 176549 528723 176561 528726
rect 175276 528695 176561 528723
rect 176549 528692 176561 528695
rect 176595 528723 176607 528726
rect 177558 528723 177564 528735
rect 176595 528695 177564 528723
rect 176595 528692 176607 528695
rect 176549 528686 176607 528692
rect 177558 528683 177564 528695
rect 177616 528723 177622 528735
rect 178018 528723 178024 528735
rect 177616 528695 178024 528723
rect 177616 528683 177622 528695
rect 178018 528683 178024 528695
rect 178076 528683 178082 528735
rect 178113 528726 178171 528732
rect 178113 528692 178125 528726
rect 178159 528723 178171 528726
rect 178202 528723 178208 528735
rect 178159 528695 178208 528723
rect 178159 528692 178171 528695
rect 178113 528686 178171 528692
rect 178202 528683 178208 528695
rect 178260 528683 178266 528735
rect 180502 528683 180508 528735
rect 180560 528683 180566 528735
rect 180612 528723 180640 528831
rect 182158 528819 182164 528871
rect 182216 528859 182222 528871
rect 182253 528862 182311 528868
rect 182253 528859 182265 528862
rect 182216 528831 182265 528859
rect 182216 528819 182222 528831
rect 182253 528828 182265 528831
rect 182299 528828 182311 528862
rect 182253 528822 182311 528828
rect 180679 528794 180737 528800
rect 180679 528760 180691 528794
rect 180725 528791 180737 528794
rect 181057 528794 181115 528800
rect 181057 528791 181069 528794
rect 180725 528763 181069 528791
rect 180725 528760 180737 528763
rect 180679 528754 180737 528760
rect 181057 528760 181069 528763
rect 181103 528791 181115 528794
rect 181681 528794 181739 528800
rect 181681 528791 181693 528794
rect 181103 528763 181693 528791
rect 181103 528760 181115 528763
rect 181057 528754 181115 528760
rect 181681 528760 181693 528763
rect 181727 528760 181739 528794
rect 181681 528754 181739 528760
rect 180781 528726 180839 528732
rect 180781 528723 180793 528726
rect 180612 528695 180793 528723
rect 180781 528692 180793 528695
rect 180827 528692 180839 528726
rect 180781 528686 180839 528692
rect 181514 528683 181520 528735
rect 181572 528723 181578 528735
rect 181572 528695 182020 528723
rect 181572 528683 181578 528695
rect 175902 528615 175908 528667
rect 175960 528615 175966 528667
rect 176181 528658 176239 528664
rect 176181 528624 176193 528658
rect 176227 528655 176239 528658
rect 176825 528658 176883 528664
rect 176227 528627 176316 528655
rect 176227 528624 176239 528627
rect 176181 528618 176239 528624
rect 176288 528531 176316 528627
rect 176825 528624 176837 528658
rect 176871 528655 176883 528658
rect 177469 528658 177527 528664
rect 177469 528655 177481 528658
rect 176871 528627 177481 528655
rect 176871 528624 176883 528627
rect 176825 528618 176883 528624
rect 177469 528624 177481 528627
rect 177515 528624 177527 528658
rect 177469 528618 177527 528624
rect 180229 528658 180287 528664
rect 180229 528624 180241 528658
rect 180275 528655 180287 528658
rect 180598 528658 180656 528664
rect 180275 528627 180548 528655
rect 180275 528624 180287 528627
rect 180229 528618 180287 528624
rect 178386 528547 178392 528599
rect 178444 528547 178450 528599
rect 180520 528587 180548 528627
rect 180598 528624 180610 528658
rect 180644 528655 180656 528658
rect 180965 528658 181023 528664
rect 180965 528655 180977 528658
rect 180644 528627 180977 528655
rect 180644 528624 180656 528627
rect 180598 528618 180656 528624
rect 180965 528624 180977 528627
rect 181011 528655 181023 528658
rect 181681 528658 181739 528664
rect 181681 528655 181693 528658
rect 181011 528627 181693 528655
rect 181011 528624 181023 528627
rect 180965 528618 181023 528624
rect 181681 528624 181693 528627
rect 181727 528624 181739 528658
rect 181681 528618 181739 528624
rect 181897 528653 181955 528659
rect 181897 528619 181909 528653
rect 181943 528619 181955 528653
rect 181897 528596 181955 528619
rect 181992 528596 182020 528695
rect 181237 528590 181367 528596
rect 180520 528559 181008 528587
rect 180980 528531 181008 528559
rect 181237 528556 181249 528590
rect 181283 528556 181321 528590
rect 181355 528587 181367 528590
rect 181897 528590 182020 528596
rect 181897 528587 181969 528590
rect 181355 528559 181969 528587
rect 181355 528556 181367 528559
rect 181237 528550 181367 528556
rect 181957 528556 181969 528559
rect 182003 528587 182020 528590
rect 186574 528587 186580 528599
rect 182003 528559 186580 528587
rect 182003 528556 182015 528559
rect 181957 528550 182015 528556
rect 186574 528547 186580 528559
rect 186632 528547 186638 528599
rect 176270 528479 176276 528531
rect 176328 528479 176334 528531
rect 176362 528479 176368 528531
rect 176420 528479 176426 528531
rect 176730 528479 176736 528531
rect 176788 528479 176794 528531
rect 177006 528479 177012 528531
rect 177064 528519 177070 528531
rect 177193 528522 177251 528528
rect 177193 528519 177205 528522
rect 177064 528491 177205 528519
rect 177064 528479 177070 528491
rect 177193 528488 177205 528491
rect 177239 528488 177251 528522
rect 177193 528482 177251 528488
rect 180962 528479 180968 528531
rect 181020 528479 181026 528531
rect 172208 528429 187480 528451
rect 172208 528420 174623 528429
rect 172208 528386 172237 528420
rect 172271 528386 172329 528420
rect 172363 528386 172421 528420
rect 172455 528386 172513 528420
rect 172547 528386 172605 528420
rect 172639 528386 172697 528420
rect 172731 528386 172789 528420
rect 172823 528386 172881 528420
rect 172915 528386 172973 528420
rect 173007 528386 173065 528420
rect 173099 528386 173157 528420
rect 173191 528386 173249 528420
rect 173283 528386 173341 528420
rect 173375 528386 173433 528420
rect 173467 528386 173525 528420
rect 173559 528386 173617 528420
rect 173651 528386 173709 528420
rect 173743 528386 173801 528420
rect 173835 528386 173893 528420
rect 173927 528386 173985 528420
rect 174019 528386 174077 528420
rect 174111 528386 174169 528420
rect 174203 528386 174261 528420
rect 174295 528386 174353 528420
rect 174387 528386 174445 528420
rect 174479 528386 174537 528420
rect 174571 528386 174623 528420
rect 172208 528377 174623 528386
rect 174675 528377 174687 528429
rect 174739 528420 174751 528429
rect 174803 528420 174815 528429
rect 174803 528386 174813 528420
rect 174739 528377 174751 528386
rect 174803 528377 174815 528386
rect 174867 528377 174879 528429
rect 174931 528420 178441 528429
rect 174939 528386 174997 528420
rect 175031 528386 175089 528420
rect 175123 528386 175181 528420
rect 175215 528386 175273 528420
rect 175307 528386 175365 528420
rect 175399 528386 175457 528420
rect 175491 528386 175549 528420
rect 175583 528386 175641 528420
rect 175675 528386 175733 528420
rect 175767 528386 175825 528420
rect 175859 528386 175917 528420
rect 175951 528386 176009 528420
rect 176043 528386 176101 528420
rect 176135 528386 176193 528420
rect 176227 528386 176285 528420
rect 176319 528386 176377 528420
rect 176411 528386 176469 528420
rect 176503 528386 176561 528420
rect 176595 528386 176653 528420
rect 176687 528386 176745 528420
rect 176779 528386 176837 528420
rect 176871 528386 176929 528420
rect 176963 528386 177021 528420
rect 177055 528386 177113 528420
rect 177147 528386 177205 528420
rect 177239 528386 177297 528420
rect 177331 528386 177389 528420
rect 177423 528386 177481 528420
rect 177515 528386 177573 528420
rect 177607 528386 177665 528420
rect 177699 528386 177757 528420
rect 177791 528386 177849 528420
rect 177883 528386 177941 528420
rect 177975 528386 178033 528420
rect 178067 528386 178125 528420
rect 178159 528386 178217 528420
rect 178251 528386 178309 528420
rect 178343 528386 178401 528420
rect 178435 528386 178441 528420
rect 174931 528377 178441 528386
rect 178493 528420 178505 528429
rect 178493 528377 178505 528386
rect 178557 528377 178569 528429
rect 178621 528377 178633 528429
rect 178685 528420 178697 528429
rect 178749 528420 182259 528429
rect 178749 528386 178769 528420
rect 178803 528386 178861 528420
rect 178895 528386 178953 528420
rect 178987 528386 179045 528420
rect 179079 528386 179137 528420
rect 179171 528386 179229 528420
rect 179263 528386 179321 528420
rect 179355 528386 179413 528420
rect 179447 528386 179505 528420
rect 179539 528386 179597 528420
rect 179631 528386 179689 528420
rect 179723 528386 179781 528420
rect 179815 528386 179873 528420
rect 179907 528386 179965 528420
rect 179999 528386 180057 528420
rect 180091 528386 180149 528420
rect 180183 528386 180241 528420
rect 180275 528386 180333 528420
rect 180367 528386 180425 528420
rect 180459 528386 180517 528420
rect 180551 528386 180609 528420
rect 180643 528386 180701 528420
rect 180735 528386 180793 528420
rect 180827 528386 180885 528420
rect 180919 528386 180977 528420
rect 181011 528386 181069 528420
rect 181103 528386 181161 528420
rect 181195 528386 181253 528420
rect 181287 528386 181345 528420
rect 181379 528386 181437 528420
rect 181471 528386 181529 528420
rect 181563 528386 181621 528420
rect 181655 528386 181713 528420
rect 181747 528386 181805 528420
rect 181839 528386 181897 528420
rect 181931 528386 181989 528420
rect 182023 528386 182081 528420
rect 182115 528386 182173 528420
rect 182207 528386 182259 528420
rect 178685 528377 178697 528386
rect 178749 528377 182259 528386
rect 182311 528377 182323 528429
rect 182375 528420 182387 528429
rect 182439 528420 182451 528429
rect 182439 528386 182449 528420
rect 182375 528377 182387 528386
rect 182439 528377 182451 528386
rect 182503 528377 182515 528429
rect 182567 528420 186077 528429
rect 182575 528386 182633 528420
rect 182667 528386 182725 528420
rect 182759 528386 182817 528420
rect 182851 528386 182909 528420
rect 182943 528386 183001 528420
rect 183035 528386 183093 528420
rect 183127 528386 183185 528420
rect 183219 528386 183277 528420
rect 183311 528386 183369 528420
rect 183403 528386 183461 528420
rect 183495 528386 183553 528420
rect 183587 528386 183645 528420
rect 183679 528386 183737 528420
rect 183771 528386 183829 528420
rect 183863 528386 183921 528420
rect 183955 528386 184013 528420
rect 184047 528386 184105 528420
rect 184139 528386 184197 528420
rect 184231 528386 184289 528420
rect 184323 528386 184381 528420
rect 184415 528386 184473 528420
rect 184507 528386 184565 528420
rect 184599 528386 184657 528420
rect 184691 528386 184749 528420
rect 184783 528386 184841 528420
rect 184875 528386 184933 528420
rect 184967 528386 185025 528420
rect 185059 528386 185117 528420
rect 185151 528386 185209 528420
rect 185243 528386 185301 528420
rect 185335 528386 185393 528420
rect 185427 528386 185485 528420
rect 185519 528386 185577 528420
rect 185611 528386 185669 528420
rect 185703 528386 185761 528420
rect 185795 528386 185853 528420
rect 185887 528386 185945 528420
rect 185979 528386 186037 528420
rect 186071 528386 186077 528420
rect 182567 528377 186077 528386
rect 186129 528420 186141 528429
rect 186129 528377 186141 528386
rect 186193 528377 186205 528429
rect 186257 528377 186269 528429
rect 186321 528420 186333 528429
rect 186385 528420 187480 528429
rect 186385 528386 186405 528420
rect 186439 528386 186497 528420
rect 186531 528386 186589 528420
rect 186623 528386 186681 528420
rect 186715 528386 186773 528420
rect 186807 528386 186865 528420
rect 186899 528386 186957 528420
rect 186991 528386 187049 528420
rect 187083 528386 187141 528420
rect 187175 528386 187233 528420
rect 187267 528386 187325 528420
rect 187359 528386 187417 528420
rect 187451 528386 187480 528420
rect 186321 528377 186333 528386
rect 186385 528377 187480 528386
rect 172208 528355 187480 528377
rect 176730 528275 176736 528327
rect 176788 528315 176794 528327
rect 177837 528318 177895 528324
rect 177837 528315 177849 528318
rect 176788 528287 177849 528315
rect 176788 528275 176794 528287
rect 177837 528284 177849 528287
rect 177883 528284 177895 528318
rect 177837 528278 177895 528284
rect 178018 528275 178024 528327
rect 178076 528275 178082 528327
rect 178938 528275 178944 528327
rect 178996 528275 179002 528327
rect 179306 528275 179312 528327
rect 179364 528315 179370 528327
rect 179401 528318 179459 528324
rect 179401 528315 179413 528318
rect 179364 528287 179413 528315
rect 179364 528275 179370 528287
rect 179401 528284 179413 528287
rect 179447 528284 179459 528318
rect 179401 528278 179459 528284
rect 180962 528275 180968 528327
rect 181020 528275 181026 528327
rect 181425 528318 181483 528324
rect 181425 528284 181437 528318
rect 181471 528315 181483 528318
rect 182158 528315 182164 528327
rect 181471 528287 182164 528315
rect 181471 528284 181483 528287
rect 181425 528278 181483 528284
rect 182158 528275 182164 528287
rect 182216 528275 182222 528327
rect 176362 528207 176368 528259
rect 176420 528207 176426 528259
rect 176822 528256 176828 528259
rect 176821 528210 176828 528256
rect 176880 528256 176886 528259
rect 176880 528250 176951 528256
rect 176880 528216 176905 528250
rect 176939 528247 176951 528250
rect 177541 528250 177599 528256
rect 177541 528247 177553 528250
rect 176939 528219 177553 528247
rect 176939 528216 176951 528219
rect 176822 528207 176828 528210
rect 176880 528210 176951 528216
rect 177481 528216 177553 528219
rect 177587 528216 177599 528250
rect 178036 528247 178064 528275
rect 178036 528219 179536 528247
rect 177481 528210 177599 528216
rect 176880 528207 176886 528210
rect 176086 528139 176092 528191
rect 176144 528139 176150 528191
rect 176182 528182 176240 528188
rect 176182 528148 176194 528182
rect 176228 528179 176240 528182
rect 176549 528182 176607 528188
rect 176549 528179 176561 528182
rect 176228 528151 176561 528179
rect 176228 528148 176240 528151
rect 176182 528142 176240 528148
rect 176549 528148 176561 528151
rect 176595 528179 176607 528182
rect 177265 528182 177323 528188
rect 177265 528179 177277 528182
rect 176595 528151 177277 528179
rect 176595 528148 176607 528151
rect 176549 528142 176607 528148
rect 177265 528148 177277 528151
rect 177311 528148 177323 528182
rect 177265 528142 177323 528148
rect 177481 528187 177539 528210
rect 177481 528153 177493 528187
rect 177527 528153 177539 528187
rect 177481 528147 177539 528153
rect 178110 528139 178116 528191
rect 178168 528139 178174 528191
rect 179309 528182 179367 528188
rect 179309 528148 179321 528182
rect 179355 528148 179367 528182
rect 179309 528142 179367 528148
rect 176263 528046 176321 528052
rect 176263 528012 176275 528046
rect 176309 528043 176321 528046
rect 176641 528046 176699 528052
rect 176641 528043 176653 528046
rect 176309 528015 176653 528043
rect 176309 528012 176321 528015
rect 176263 528006 176321 528012
rect 176641 528012 176653 528015
rect 176687 528043 176699 528046
rect 177265 528046 177323 528052
rect 177265 528043 177277 528046
rect 176687 528015 177277 528043
rect 176687 528012 176699 528015
rect 176641 528006 176699 528012
rect 177265 528012 177277 528015
rect 177311 528012 177323 528046
rect 177265 528006 177323 528012
rect 177374 528003 177380 528055
rect 177432 528043 177438 528055
rect 177929 528046 177987 528052
rect 177929 528043 177941 528046
rect 177432 528015 177941 528043
rect 177432 528003 177438 528015
rect 177929 528012 177941 528015
rect 177975 528012 177987 528046
rect 177929 528006 177987 528012
rect 178938 527935 178944 527987
rect 178996 527975 179002 527987
rect 179324 527975 179352 528142
rect 179508 528120 179536 528219
rect 181330 528139 181336 528191
rect 181388 528139 181394 528191
rect 179493 528114 179551 528120
rect 179493 528080 179505 528114
rect 179539 528111 179551 528114
rect 180686 528111 180692 528123
rect 179539 528083 180692 528111
rect 179539 528080 179551 528083
rect 179493 528074 179551 528080
rect 180686 528071 180692 528083
rect 180744 528111 180750 528123
rect 181517 528114 181575 528120
rect 181517 528111 181529 528114
rect 180744 528083 181529 528111
rect 180744 528071 180750 528083
rect 181517 528080 181529 528083
rect 181563 528080 181575 528114
rect 181517 528074 181575 528080
rect 178996 527947 179352 527975
rect 178996 527935 179002 527947
rect 172208 527885 187480 527907
rect 172208 527876 173963 527885
rect 174015 527876 174027 527885
rect 174079 527876 174091 527885
rect 172208 527842 172237 527876
rect 172271 527842 172329 527876
rect 172363 527842 172421 527876
rect 172455 527842 172513 527876
rect 172547 527842 172605 527876
rect 172639 527842 172697 527876
rect 172731 527842 172789 527876
rect 172823 527842 172881 527876
rect 172915 527842 172973 527876
rect 173007 527842 173065 527876
rect 173099 527842 173157 527876
rect 173191 527842 173249 527876
rect 173283 527842 173341 527876
rect 173375 527842 173433 527876
rect 173467 527842 173525 527876
rect 173559 527842 173617 527876
rect 173651 527842 173709 527876
rect 173743 527842 173801 527876
rect 173835 527842 173893 527876
rect 173927 527842 173963 527876
rect 174019 527842 174027 527876
rect 172208 527833 173963 527842
rect 174015 527833 174027 527842
rect 174079 527833 174091 527842
rect 174143 527833 174155 527885
rect 174207 527833 174219 527885
rect 174271 527876 177781 527885
rect 174295 527842 174353 527876
rect 174387 527842 174445 527876
rect 174479 527842 174537 527876
rect 174571 527842 174629 527876
rect 174663 527842 174721 527876
rect 174755 527842 174813 527876
rect 174847 527842 174905 527876
rect 174939 527842 174997 527876
rect 175031 527842 175089 527876
rect 175123 527842 175181 527876
rect 175215 527842 175273 527876
rect 175307 527842 175365 527876
rect 175399 527842 175457 527876
rect 175491 527842 175549 527876
rect 175583 527842 175641 527876
rect 175675 527842 175733 527876
rect 175767 527842 175825 527876
rect 175859 527842 175917 527876
rect 175951 527842 176009 527876
rect 176043 527842 176101 527876
rect 176135 527842 176193 527876
rect 176227 527842 176285 527876
rect 176319 527842 176377 527876
rect 176411 527842 176469 527876
rect 176503 527842 176561 527876
rect 176595 527842 176653 527876
rect 176687 527842 176745 527876
rect 176779 527842 176837 527876
rect 176871 527842 176929 527876
rect 176963 527842 177021 527876
rect 177055 527842 177113 527876
rect 177147 527842 177205 527876
rect 177239 527842 177297 527876
rect 177331 527842 177389 527876
rect 177423 527842 177481 527876
rect 177515 527842 177573 527876
rect 177607 527842 177665 527876
rect 177699 527842 177757 527876
rect 174271 527833 177781 527842
rect 177833 527833 177845 527885
rect 177897 527833 177909 527885
rect 177961 527876 177973 527885
rect 178025 527876 178037 527885
rect 178089 527876 181599 527885
rect 181651 527876 181663 527885
rect 181715 527876 181727 527885
rect 178025 527842 178033 527876
rect 178089 527842 178125 527876
rect 178159 527842 178217 527876
rect 178251 527842 178309 527876
rect 178343 527842 178401 527876
rect 178435 527842 178493 527876
rect 178527 527842 178585 527876
rect 178619 527842 178677 527876
rect 178711 527842 178769 527876
rect 178803 527842 178861 527876
rect 178895 527842 178953 527876
rect 178987 527842 179045 527876
rect 179079 527842 179137 527876
rect 179171 527842 179229 527876
rect 179263 527842 179321 527876
rect 179355 527842 179413 527876
rect 179447 527842 179505 527876
rect 179539 527842 179597 527876
rect 179631 527842 179689 527876
rect 179723 527842 179781 527876
rect 179815 527842 179873 527876
rect 179907 527842 179965 527876
rect 179999 527842 180057 527876
rect 180091 527842 180149 527876
rect 180183 527842 180241 527876
rect 180275 527842 180333 527876
rect 180367 527842 180425 527876
rect 180459 527842 180517 527876
rect 180551 527842 180609 527876
rect 180643 527842 180701 527876
rect 180735 527842 180793 527876
rect 180827 527842 180885 527876
rect 180919 527842 180977 527876
rect 181011 527842 181069 527876
rect 181103 527842 181161 527876
rect 181195 527842 181253 527876
rect 181287 527842 181345 527876
rect 181379 527842 181437 527876
rect 181471 527842 181529 527876
rect 181563 527842 181599 527876
rect 181655 527842 181663 527876
rect 177961 527833 177973 527842
rect 178025 527833 178037 527842
rect 178089 527833 181599 527842
rect 181651 527833 181663 527842
rect 181715 527833 181727 527842
rect 181779 527833 181791 527885
rect 181843 527833 181855 527885
rect 181907 527876 185417 527885
rect 181931 527842 181989 527876
rect 182023 527842 182081 527876
rect 182115 527842 182173 527876
rect 182207 527842 182265 527876
rect 182299 527842 182357 527876
rect 182391 527842 182449 527876
rect 182483 527842 182541 527876
rect 182575 527842 182633 527876
rect 182667 527842 182725 527876
rect 182759 527842 182817 527876
rect 182851 527842 182909 527876
rect 182943 527842 183001 527876
rect 183035 527842 183093 527876
rect 183127 527842 183185 527876
rect 183219 527842 183277 527876
rect 183311 527842 183369 527876
rect 183403 527842 183461 527876
rect 183495 527842 183553 527876
rect 183587 527842 183645 527876
rect 183679 527842 183737 527876
rect 183771 527842 183829 527876
rect 183863 527842 183921 527876
rect 183955 527842 184013 527876
rect 184047 527842 184105 527876
rect 184139 527842 184197 527876
rect 184231 527842 184289 527876
rect 184323 527842 184381 527876
rect 184415 527842 184473 527876
rect 184507 527842 184565 527876
rect 184599 527842 184657 527876
rect 184691 527842 184749 527876
rect 184783 527842 184841 527876
rect 184875 527842 184933 527876
rect 184967 527842 185025 527876
rect 185059 527842 185117 527876
rect 185151 527842 185209 527876
rect 185243 527842 185301 527876
rect 185335 527842 185393 527876
rect 181907 527833 185417 527842
rect 185469 527833 185481 527885
rect 185533 527833 185545 527885
rect 185597 527876 185609 527885
rect 185661 527876 185673 527885
rect 185725 527876 187480 527885
rect 185661 527842 185669 527876
rect 185725 527842 185761 527876
rect 185795 527842 185853 527876
rect 185887 527842 185945 527876
rect 185979 527842 186037 527876
rect 186071 527842 186129 527876
rect 186163 527842 186221 527876
rect 186255 527842 186313 527876
rect 186347 527842 186405 527876
rect 186439 527842 186497 527876
rect 186531 527842 186589 527876
rect 186623 527842 186681 527876
rect 186715 527842 186773 527876
rect 186807 527842 186865 527876
rect 186899 527842 186957 527876
rect 186991 527842 187049 527876
rect 187083 527842 187141 527876
rect 187175 527842 187233 527876
rect 187267 527842 187325 527876
rect 187359 527842 187417 527876
rect 187451 527842 187480 527876
rect 185597 527833 185609 527842
rect 185661 527833 185673 527842
rect 185725 527833 187480 527842
rect 172208 527811 187480 527833
rect 176270 527731 176276 527783
rect 176328 527771 176334 527783
rect 176365 527774 176423 527780
rect 176365 527771 176377 527774
rect 176328 527743 176377 527771
rect 176328 527731 176334 527743
rect 176365 527740 176377 527743
rect 176411 527740 176423 527774
rect 176365 527734 176423 527740
rect 178938 527731 178944 527783
rect 178996 527731 179002 527783
rect 177006 527595 177012 527647
rect 177064 527595 177070 527647
rect 179490 527595 179496 527647
rect 179548 527595 179554 527647
rect 172208 527341 187480 527363
rect 172208 527332 174623 527341
rect 172208 527298 172237 527332
rect 172271 527298 172329 527332
rect 172363 527298 172421 527332
rect 172455 527298 172513 527332
rect 172547 527298 172605 527332
rect 172639 527298 172697 527332
rect 172731 527298 172789 527332
rect 172823 527298 172881 527332
rect 172915 527298 172973 527332
rect 173007 527298 173065 527332
rect 173099 527298 173157 527332
rect 173191 527298 173249 527332
rect 173283 527298 173341 527332
rect 173375 527298 173433 527332
rect 173467 527298 173525 527332
rect 173559 527298 173617 527332
rect 173651 527298 173709 527332
rect 173743 527298 173801 527332
rect 173835 527298 173893 527332
rect 173927 527298 173985 527332
rect 174019 527298 174077 527332
rect 174111 527298 174169 527332
rect 174203 527298 174261 527332
rect 174295 527298 174353 527332
rect 174387 527298 174445 527332
rect 174479 527298 174537 527332
rect 174571 527298 174623 527332
rect 172208 527289 174623 527298
rect 174675 527289 174687 527341
rect 174739 527332 174751 527341
rect 174803 527332 174815 527341
rect 174803 527298 174813 527332
rect 174739 527289 174751 527298
rect 174803 527289 174815 527298
rect 174867 527289 174879 527341
rect 174931 527332 178441 527341
rect 174939 527298 174997 527332
rect 175031 527298 175089 527332
rect 175123 527298 175181 527332
rect 175215 527298 175273 527332
rect 175307 527298 175365 527332
rect 175399 527298 175457 527332
rect 175491 527298 175549 527332
rect 175583 527298 175641 527332
rect 175675 527298 175733 527332
rect 175767 527298 175825 527332
rect 175859 527298 175917 527332
rect 175951 527298 176009 527332
rect 176043 527298 176101 527332
rect 176135 527298 176193 527332
rect 176227 527298 176285 527332
rect 176319 527298 176377 527332
rect 176411 527298 176469 527332
rect 176503 527298 176561 527332
rect 176595 527298 176653 527332
rect 176687 527298 176745 527332
rect 176779 527298 176837 527332
rect 176871 527298 176929 527332
rect 176963 527298 177021 527332
rect 177055 527298 177113 527332
rect 177147 527298 177205 527332
rect 177239 527298 177297 527332
rect 177331 527298 177389 527332
rect 177423 527298 177481 527332
rect 177515 527298 177573 527332
rect 177607 527298 177665 527332
rect 177699 527298 177757 527332
rect 177791 527298 177849 527332
rect 177883 527298 177941 527332
rect 177975 527298 178033 527332
rect 178067 527298 178125 527332
rect 178159 527298 178217 527332
rect 178251 527298 178309 527332
rect 178343 527298 178401 527332
rect 178435 527298 178441 527332
rect 174931 527289 178441 527298
rect 178493 527332 178505 527341
rect 178493 527289 178505 527298
rect 178557 527289 178569 527341
rect 178621 527289 178633 527341
rect 178685 527332 178697 527341
rect 178749 527332 182259 527341
rect 178749 527298 178769 527332
rect 178803 527298 178861 527332
rect 178895 527298 178953 527332
rect 178987 527298 179045 527332
rect 179079 527298 179137 527332
rect 179171 527298 179229 527332
rect 179263 527298 179321 527332
rect 179355 527298 179413 527332
rect 179447 527298 179505 527332
rect 179539 527298 179597 527332
rect 179631 527298 179689 527332
rect 179723 527298 179781 527332
rect 179815 527298 179873 527332
rect 179907 527298 179965 527332
rect 179999 527298 180057 527332
rect 180091 527298 180149 527332
rect 180183 527298 180241 527332
rect 180275 527298 180333 527332
rect 180367 527298 180425 527332
rect 180459 527298 180517 527332
rect 180551 527298 180609 527332
rect 180643 527298 180701 527332
rect 180735 527298 180793 527332
rect 180827 527298 180885 527332
rect 180919 527298 180977 527332
rect 181011 527298 181069 527332
rect 181103 527298 181161 527332
rect 181195 527298 181253 527332
rect 181287 527298 181345 527332
rect 181379 527298 181437 527332
rect 181471 527298 181529 527332
rect 181563 527298 181621 527332
rect 181655 527298 181713 527332
rect 181747 527298 181805 527332
rect 181839 527298 181897 527332
rect 181931 527298 181989 527332
rect 182023 527298 182081 527332
rect 182115 527298 182173 527332
rect 182207 527298 182259 527332
rect 178685 527289 178697 527298
rect 178749 527289 182259 527298
rect 182311 527289 182323 527341
rect 182375 527332 182387 527341
rect 182439 527332 182451 527341
rect 182439 527298 182449 527332
rect 182375 527289 182387 527298
rect 182439 527289 182451 527298
rect 182503 527289 182515 527341
rect 182567 527332 186077 527341
rect 182575 527298 182633 527332
rect 182667 527298 182725 527332
rect 182759 527298 182817 527332
rect 182851 527298 182909 527332
rect 182943 527298 183001 527332
rect 183035 527298 183093 527332
rect 183127 527298 183185 527332
rect 183219 527298 183277 527332
rect 183311 527298 183369 527332
rect 183403 527298 183461 527332
rect 183495 527298 183553 527332
rect 183587 527298 183645 527332
rect 183679 527298 183737 527332
rect 183771 527298 183829 527332
rect 183863 527298 183921 527332
rect 183955 527298 184013 527332
rect 184047 527298 184105 527332
rect 184139 527298 184197 527332
rect 184231 527298 184289 527332
rect 184323 527298 184381 527332
rect 184415 527298 184473 527332
rect 184507 527298 184565 527332
rect 184599 527298 184657 527332
rect 184691 527298 184749 527332
rect 184783 527298 184841 527332
rect 184875 527298 184933 527332
rect 184967 527298 185025 527332
rect 185059 527298 185117 527332
rect 185151 527298 185209 527332
rect 185243 527298 185301 527332
rect 185335 527298 185393 527332
rect 185427 527298 185485 527332
rect 185519 527298 185577 527332
rect 185611 527298 185669 527332
rect 185703 527298 185761 527332
rect 185795 527298 185853 527332
rect 185887 527298 185945 527332
rect 185979 527298 186037 527332
rect 186071 527298 186077 527332
rect 182567 527289 186077 527298
rect 186129 527332 186141 527341
rect 186129 527289 186141 527298
rect 186193 527289 186205 527341
rect 186257 527289 186269 527341
rect 186321 527332 186333 527341
rect 186385 527332 187480 527341
rect 186385 527298 186405 527332
rect 186439 527298 186497 527332
rect 186531 527298 186589 527332
rect 186623 527298 186681 527332
rect 186715 527298 186773 527332
rect 186807 527298 186865 527332
rect 186899 527298 186957 527332
rect 186991 527298 187049 527332
rect 187083 527298 187141 527332
rect 187175 527298 187233 527332
rect 187267 527298 187325 527332
rect 187359 527298 187417 527332
rect 187451 527298 187480 527332
rect 186321 527289 186333 527298
rect 186385 527289 187480 527298
rect 172208 527267 187480 527289
rect 172208 526797 187480 526819
rect 172208 526788 173963 526797
rect 174015 526788 174027 526797
rect 174079 526788 174091 526797
rect 172208 526754 172237 526788
rect 172271 526754 172329 526788
rect 172363 526754 172421 526788
rect 172455 526754 172513 526788
rect 172547 526754 172605 526788
rect 172639 526754 172697 526788
rect 172731 526754 172789 526788
rect 172823 526754 172881 526788
rect 172915 526754 172973 526788
rect 173007 526754 173065 526788
rect 173099 526754 173157 526788
rect 173191 526754 173249 526788
rect 173283 526754 173341 526788
rect 173375 526754 173433 526788
rect 173467 526754 173525 526788
rect 173559 526754 173617 526788
rect 173651 526754 173709 526788
rect 173743 526754 173801 526788
rect 173835 526754 173893 526788
rect 173927 526754 173963 526788
rect 174019 526754 174027 526788
rect 172208 526745 173963 526754
rect 174015 526745 174027 526754
rect 174079 526745 174091 526754
rect 174143 526745 174155 526797
rect 174207 526745 174219 526797
rect 174271 526788 177781 526797
rect 174295 526754 174353 526788
rect 174387 526754 174445 526788
rect 174479 526754 174537 526788
rect 174571 526754 174629 526788
rect 174663 526754 174721 526788
rect 174755 526754 174813 526788
rect 174847 526754 174905 526788
rect 174939 526754 174997 526788
rect 175031 526754 175089 526788
rect 175123 526754 175181 526788
rect 175215 526754 175273 526788
rect 175307 526754 175365 526788
rect 175399 526754 175457 526788
rect 175491 526754 175549 526788
rect 175583 526754 175641 526788
rect 175675 526754 175733 526788
rect 175767 526754 175825 526788
rect 175859 526754 175917 526788
rect 175951 526754 176009 526788
rect 176043 526754 176101 526788
rect 176135 526754 176193 526788
rect 176227 526754 176285 526788
rect 176319 526754 176377 526788
rect 176411 526754 176469 526788
rect 176503 526754 176561 526788
rect 176595 526754 176653 526788
rect 176687 526754 176745 526788
rect 176779 526754 176837 526788
rect 176871 526754 176929 526788
rect 176963 526754 177021 526788
rect 177055 526754 177113 526788
rect 177147 526754 177205 526788
rect 177239 526754 177297 526788
rect 177331 526754 177389 526788
rect 177423 526754 177481 526788
rect 177515 526754 177573 526788
rect 177607 526754 177665 526788
rect 177699 526754 177757 526788
rect 174271 526745 177781 526754
rect 177833 526745 177845 526797
rect 177897 526745 177909 526797
rect 177961 526788 177973 526797
rect 178025 526788 178037 526797
rect 178089 526788 181599 526797
rect 181651 526788 181663 526797
rect 181715 526788 181727 526797
rect 178025 526754 178033 526788
rect 178089 526754 178125 526788
rect 178159 526754 178217 526788
rect 178251 526754 178309 526788
rect 178343 526754 178401 526788
rect 178435 526754 178493 526788
rect 178527 526754 178585 526788
rect 178619 526754 178677 526788
rect 178711 526754 178769 526788
rect 178803 526754 178861 526788
rect 178895 526754 178953 526788
rect 178987 526754 179045 526788
rect 179079 526754 179137 526788
rect 179171 526754 179229 526788
rect 179263 526754 179321 526788
rect 179355 526754 179413 526788
rect 179447 526754 179505 526788
rect 179539 526754 179597 526788
rect 179631 526754 179689 526788
rect 179723 526754 179781 526788
rect 179815 526754 179873 526788
rect 179907 526754 179965 526788
rect 179999 526754 180057 526788
rect 180091 526754 180149 526788
rect 180183 526754 180241 526788
rect 180275 526754 180333 526788
rect 180367 526754 180425 526788
rect 180459 526754 180517 526788
rect 180551 526754 180609 526788
rect 180643 526754 180701 526788
rect 180735 526754 180793 526788
rect 180827 526754 180885 526788
rect 180919 526754 180977 526788
rect 181011 526754 181069 526788
rect 181103 526754 181161 526788
rect 181195 526754 181253 526788
rect 181287 526754 181345 526788
rect 181379 526754 181437 526788
rect 181471 526754 181529 526788
rect 181563 526754 181599 526788
rect 181655 526754 181663 526788
rect 177961 526745 177973 526754
rect 178025 526745 178037 526754
rect 178089 526745 181599 526754
rect 181651 526745 181663 526754
rect 181715 526745 181727 526754
rect 181779 526745 181791 526797
rect 181843 526745 181855 526797
rect 181907 526788 185417 526797
rect 181931 526754 181989 526788
rect 182023 526754 182081 526788
rect 182115 526754 182173 526788
rect 182207 526754 182265 526788
rect 182299 526754 182357 526788
rect 182391 526754 182449 526788
rect 182483 526754 182541 526788
rect 182575 526754 182633 526788
rect 182667 526754 182725 526788
rect 182759 526754 182817 526788
rect 182851 526754 182909 526788
rect 182943 526754 183001 526788
rect 183035 526754 183093 526788
rect 183127 526754 183185 526788
rect 183219 526754 183277 526788
rect 183311 526754 183369 526788
rect 183403 526754 183461 526788
rect 183495 526754 183553 526788
rect 183587 526754 183645 526788
rect 183679 526754 183737 526788
rect 183771 526754 183829 526788
rect 183863 526754 183921 526788
rect 183955 526754 184013 526788
rect 184047 526754 184105 526788
rect 184139 526754 184197 526788
rect 184231 526754 184289 526788
rect 184323 526754 184381 526788
rect 184415 526754 184473 526788
rect 184507 526754 184565 526788
rect 184599 526754 184657 526788
rect 184691 526754 184749 526788
rect 184783 526754 184841 526788
rect 184875 526754 184933 526788
rect 184967 526754 185025 526788
rect 185059 526754 185117 526788
rect 185151 526754 185209 526788
rect 185243 526754 185301 526788
rect 185335 526754 185393 526788
rect 181907 526745 185417 526754
rect 185469 526745 185481 526797
rect 185533 526745 185545 526797
rect 185597 526788 185609 526797
rect 185661 526788 185673 526797
rect 185725 526788 187480 526797
rect 185661 526754 185669 526788
rect 185725 526754 185761 526788
rect 185795 526754 185853 526788
rect 185887 526754 185945 526788
rect 185979 526754 186037 526788
rect 186071 526754 186129 526788
rect 186163 526754 186221 526788
rect 186255 526754 186313 526788
rect 186347 526754 186405 526788
rect 186439 526754 186497 526788
rect 186531 526754 186589 526788
rect 186623 526754 186681 526788
rect 186715 526754 186773 526788
rect 186807 526754 186865 526788
rect 186899 526754 186957 526788
rect 186991 526754 187049 526788
rect 187083 526754 187141 526788
rect 187175 526754 187233 526788
rect 187267 526754 187325 526788
rect 187359 526754 187417 526788
rect 187451 526754 187480 526788
rect 185597 526745 185609 526754
rect 185661 526745 185673 526754
rect 185725 526745 187480 526754
rect 172208 526723 187480 526745
rect 172208 526253 187480 526275
rect 172208 526244 174623 526253
rect 172208 526210 172237 526244
rect 172271 526210 172329 526244
rect 172363 526210 172421 526244
rect 172455 526210 172513 526244
rect 172547 526210 172605 526244
rect 172639 526210 172697 526244
rect 172731 526210 172789 526244
rect 172823 526210 172881 526244
rect 172915 526210 172973 526244
rect 173007 526210 173065 526244
rect 173099 526210 173157 526244
rect 173191 526210 173249 526244
rect 173283 526210 173341 526244
rect 173375 526210 173433 526244
rect 173467 526210 173525 526244
rect 173559 526210 173617 526244
rect 173651 526210 173709 526244
rect 173743 526210 173801 526244
rect 173835 526210 173893 526244
rect 173927 526210 173985 526244
rect 174019 526210 174077 526244
rect 174111 526210 174169 526244
rect 174203 526210 174261 526244
rect 174295 526210 174353 526244
rect 174387 526210 174445 526244
rect 174479 526210 174537 526244
rect 174571 526210 174623 526244
rect 172208 526201 174623 526210
rect 174675 526201 174687 526253
rect 174739 526244 174751 526253
rect 174803 526244 174815 526253
rect 174803 526210 174813 526244
rect 174739 526201 174751 526210
rect 174803 526201 174815 526210
rect 174867 526201 174879 526253
rect 174931 526244 178441 526253
rect 174939 526210 174997 526244
rect 175031 526210 175089 526244
rect 175123 526210 175181 526244
rect 175215 526210 175273 526244
rect 175307 526210 175365 526244
rect 175399 526210 175457 526244
rect 175491 526210 175549 526244
rect 175583 526210 175641 526244
rect 175675 526210 175733 526244
rect 175767 526210 175825 526244
rect 175859 526210 175917 526244
rect 175951 526210 176009 526244
rect 176043 526210 176101 526244
rect 176135 526210 176193 526244
rect 176227 526210 176285 526244
rect 176319 526210 176377 526244
rect 176411 526210 176469 526244
rect 176503 526210 176561 526244
rect 176595 526210 176653 526244
rect 176687 526210 176745 526244
rect 176779 526210 176837 526244
rect 176871 526210 176929 526244
rect 176963 526210 177021 526244
rect 177055 526210 177113 526244
rect 177147 526210 177205 526244
rect 177239 526210 177297 526244
rect 177331 526210 177389 526244
rect 177423 526210 177481 526244
rect 177515 526210 177573 526244
rect 177607 526210 177665 526244
rect 177699 526210 177757 526244
rect 177791 526210 177849 526244
rect 177883 526210 177941 526244
rect 177975 526210 178033 526244
rect 178067 526210 178125 526244
rect 178159 526210 178217 526244
rect 178251 526210 178309 526244
rect 178343 526210 178401 526244
rect 178435 526210 178441 526244
rect 174931 526201 178441 526210
rect 178493 526244 178505 526253
rect 178493 526201 178505 526210
rect 178557 526201 178569 526253
rect 178621 526201 178633 526253
rect 178685 526244 178697 526253
rect 178749 526244 182259 526253
rect 178749 526210 178769 526244
rect 178803 526210 178861 526244
rect 178895 526210 178953 526244
rect 178987 526210 179045 526244
rect 179079 526210 179137 526244
rect 179171 526210 179229 526244
rect 179263 526210 179321 526244
rect 179355 526210 179413 526244
rect 179447 526210 179505 526244
rect 179539 526210 179597 526244
rect 179631 526210 179689 526244
rect 179723 526210 179781 526244
rect 179815 526210 179873 526244
rect 179907 526210 179965 526244
rect 179999 526210 180057 526244
rect 180091 526210 180149 526244
rect 180183 526210 180241 526244
rect 180275 526210 180333 526244
rect 180367 526210 180425 526244
rect 180459 526210 180517 526244
rect 180551 526210 180609 526244
rect 180643 526210 180701 526244
rect 180735 526210 180793 526244
rect 180827 526210 180885 526244
rect 180919 526210 180977 526244
rect 181011 526210 181069 526244
rect 181103 526210 181161 526244
rect 181195 526210 181253 526244
rect 181287 526210 181345 526244
rect 181379 526210 181437 526244
rect 181471 526210 181529 526244
rect 181563 526210 181621 526244
rect 181655 526210 181713 526244
rect 181747 526210 181805 526244
rect 181839 526210 181897 526244
rect 181931 526210 181989 526244
rect 182023 526210 182081 526244
rect 182115 526210 182173 526244
rect 182207 526210 182259 526244
rect 178685 526201 178697 526210
rect 178749 526201 182259 526210
rect 182311 526201 182323 526253
rect 182375 526244 182387 526253
rect 182439 526244 182451 526253
rect 182439 526210 182449 526244
rect 182375 526201 182387 526210
rect 182439 526201 182451 526210
rect 182503 526201 182515 526253
rect 182567 526244 186077 526253
rect 182575 526210 182633 526244
rect 182667 526210 182725 526244
rect 182759 526210 182817 526244
rect 182851 526210 182909 526244
rect 182943 526210 183001 526244
rect 183035 526210 183093 526244
rect 183127 526210 183185 526244
rect 183219 526210 183277 526244
rect 183311 526210 183369 526244
rect 183403 526210 183461 526244
rect 183495 526210 183553 526244
rect 183587 526210 183645 526244
rect 183679 526210 183737 526244
rect 183771 526210 183829 526244
rect 183863 526210 183921 526244
rect 183955 526210 184013 526244
rect 184047 526210 184105 526244
rect 184139 526210 184197 526244
rect 184231 526210 184289 526244
rect 184323 526210 184381 526244
rect 184415 526210 184473 526244
rect 184507 526210 184565 526244
rect 184599 526210 184657 526244
rect 184691 526210 184749 526244
rect 184783 526210 184841 526244
rect 184875 526210 184933 526244
rect 184967 526210 185025 526244
rect 185059 526210 185117 526244
rect 185151 526210 185209 526244
rect 185243 526210 185301 526244
rect 185335 526210 185393 526244
rect 185427 526210 185485 526244
rect 185519 526210 185577 526244
rect 185611 526210 185669 526244
rect 185703 526210 185761 526244
rect 185795 526210 185853 526244
rect 185887 526210 185945 526244
rect 185979 526210 186037 526244
rect 186071 526210 186077 526244
rect 182567 526201 186077 526210
rect 186129 526244 186141 526253
rect 186129 526201 186141 526210
rect 186193 526201 186205 526253
rect 186257 526201 186269 526253
rect 186321 526244 186333 526253
rect 186385 526244 187480 526253
rect 186385 526210 186405 526244
rect 186439 526210 186497 526244
rect 186531 526210 186589 526244
rect 186623 526210 186681 526244
rect 186715 526210 186773 526244
rect 186807 526210 186865 526244
rect 186899 526210 186957 526244
rect 186991 526210 187049 526244
rect 187083 526210 187141 526244
rect 187175 526210 187233 526244
rect 187267 526210 187325 526244
rect 187359 526210 187417 526244
rect 187451 526210 187480 526244
rect 186321 526201 186333 526210
rect 186385 526201 187480 526210
rect 172208 526179 187480 526201
rect 172208 525709 187480 525731
rect 172208 525700 173963 525709
rect 174015 525700 174027 525709
rect 174079 525700 174091 525709
rect 172208 525666 172237 525700
rect 172271 525666 172329 525700
rect 172363 525666 172421 525700
rect 172455 525666 172513 525700
rect 172547 525666 172605 525700
rect 172639 525666 172697 525700
rect 172731 525666 172789 525700
rect 172823 525666 172881 525700
rect 172915 525666 172973 525700
rect 173007 525666 173065 525700
rect 173099 525666 173157 525700
rect 173191 525666 173249 525700
rect 173283 525666 173341 525700
rect 173375 525666 173433 525700
rect 173467 525666 173525 525700
rect 173559 525666 173617 525700
rect 173651 525666 173709 525700
rect 173743 525666 173801 525700
rect 173835 525666 173893 525700
rect 173927 525666 173963 525700
rect 174019 525666 174027 525700
rect 172208 525657 173963 525666
rect 174015 525657 174027 525666
rect 174079 525657 174091 525666
rect 174143 525657 174155 525709
rect 174207 525657 174219 525709
rect 174271 525700 177781 525709
rect 174295 525666 174353 525700
rect 174387 525666 174445 525700
rect 174479 525666 174537 525700
rect 174571 525666 174629 525700
rect 174663 525666 174721 525700
rect 174755 525666 174813 525700
rect 174847 525666 174905 525700
rect 174939 525666 174997 525700
rect 175031 525666 175089 525700
rect 175123 525666 175181 525700
rect 175215 525666 175273 525700
rect 175307 525666 175365 525700
rect 175399 525666 175457 525700
rect 175491 525666 175549 525700
rect 175583 525666 175641 525700
rect 175675 525666 175733 525700
rect 175767 525666 175825 525700
rect 175859 525666 175917 525700
rect 175951 525666 176009 525700
rect 176043 525666 176101 525700
rect 176135 525666 176193 525700
rect 176227 525666 176285 525700
rect 176319 525666 176377 525700
rect 176411 525666 176469 525700
rect 176503 525666 176561 525700
rect 176595 525666 176653 525700
rect 176687 525666 176745 525700
rect 176779 525666 176837 525700
rect 176871 525666 176929 525700
rect 176963 525666 177021 525700
rect 177055 525666 177113 525700
rect 177147 525666 177205 525700
rect 177239 525666 177297 525700
rect 177331 525666 177389 525700
rect 177423 525666 177481 525700
rect 177515 525666 177573 525700
rect 177607 525666 177665 525700
rect 177699 525666 177757 525700
rect 174271 525657 177781 525666
rect 177833 525657 177845 525709
rect 177897 525657 177909 525709
rect 177961 525700 177973 525709
rect 178025 525700 178037 525709
rect 178089 525700 181599 525709
rect 181651 525700 181663 525709
rect 181715 525700 181727 525709
rect 178025 525666 178033 525700
rect 178089 525666 178125 525700
rect 178159 525666 178217 525700
rect 178251 525666 178309 525700
rect 178343 525666 178401 525700
rect 178435 525666 178493 525700
rect 178527 525666 178585 525700
rect 178619 525666 178677 525700
rect 178711 525666 178769 525700
rect 178803 525666 178861 525700
rect 178895 525666 178953 525700
rect 178987 525666 179045 525700
rect 179079 525666 179137 525700
rect 179171 525666 179229 525700
rect 179263 525666 179321 525700
rect 179355 525666 179413 525700
rect 179447 525666 179505 525700
rect 179539 525666 179597 525700
rect 179631 525666 179689 525700
rect 179723 525666 179781 525700
rect 179815 525666 179873 525700
rect 179907 525666 179965 525700
rect 179999 525666 180057 525700
rect 180091 525666 180149 525700
rect 180183 525666 180241 525700
rect 180275 525666 180333 525700
rect 180367 525666 180425 525700
rect 180459 525666 180517 525700
rect 180551 525666 180609 525700
rect 180643 525666 180701 525700
rect 180735 525666 180793 525700
rect 180827 525666 180885 525700
rect 180919 525666 180977 525700
rect 181011 525666 181069 525700
rect 181103 525666 181161 525700
rect 181195 525666 181253 525700
rect 181287 525666 181345 525700
rect 181379 525666 181437 525700
rect 181471 525666 181529 525700
rect 181563 525666 181599 525700
rect 181655 525666 181663 525700
rect 177961 525657 177973 525666
rect 178025 525657 178037 525666
rect 178089 525657 181599 525666
rect 181651 525657 181663 525666
rect 181715 525657 181727 525666
rect 181779 525657 181791 525709
rect 181843 525657 181855 525709
rect 181907 525700 185417 525709
rect 181931 525666 181989 525700
rect 182023 525666 182081 525700
rect 182115 525666 182173 525700
rect 182207 525666 182265 525700
rect 182299 525666 182357 525700
rect 182391 525666 182449 525700
rect 182483 525666 182541 525700
rect 182575 525666 182633 525700
rect 182667 525666 182725 525700
rect 182759 525666 182817 525700
rect 182851 525666 182909 525700
rect 182943 525666 183001 525700
rect 183035 525666 183093 525700
rect 183127 525666 183185 525700
rect 183219 525666 183277 525700
rect 183311 525666 183369 525700
rect 183403 525666 183461 525700
rect 183495 525666 183553 525700
rect 183587 525666 183645 525700
rect 183679 525666 183737 525700
rect 183771 525666 183829 525700
rect 183863 525666 183921 525700
rect 183955 525666 184013 525700
rect 184047 525666 184105 525700
rect 184139 525666 184197 525700
rect 184231 525666 184289 525700
rect 184323 525666 184381 525700
rect 184415 525666 184473 525700
rect 184507 525666 184565 525700
rect 184599 525666 184657 525700
rect 184691 525666 184749 525700
rect 184783 525666 184841 525700
rect 184875 525666 184933 525700
rect 184967 525666 185025 525700
rect 185059 525666 185117 525700
rect 185151 525666 185209 525700
rect 185243 525666 185301 525700
rect 185335 525666 185393 525700
rect 181907 525657 185417 525666
rect 185469 525657 185481 525709
rect 185533 525657 185545 525709
rect 185597 525700 185609 525709
rect 185661 525700 185673 525709
rect 185725 525700 187480 525709
rect 185661 525666 185669 525700
rect 185725 525666 185761 525700
rect 185795 525666 185853 525700
rect 185887 525666 185945 525700
rect 185979 525666 186037 525700
rect 186071 525666 186129 525700
rect 186163 525666 186221 525700
rect 186255 525666 186313 525700
rect 186347 525666 186405 525700
rect 186439 525666 186497 525700
rect 186531 525666 186589 525700
rect 186623 525666 186681 525700
rect 186715 525666 186773 525700
rect 186807 525666 186865 525700
rect 186899 525666 186957 525700
rect 186991 525666 187049 525700
rect 187083 525666 187141 525700
rect 187175 525666 187233 525700
rect 187267 525666 187325 525700
rect 187359 525666 187417 525700
rect 187451 525666 187480 525700
rect 185597 525657 185609 525666
rect 185661 525657 185673 525666
rect 185725 525657 187480 525666
rect 172208 525635 187480 525657
rect 172208 525165 187480 525187
rect 172208 525156 174623 525165
rect 172208 525122 172237 525156
rect 172271 525122 172329 525156
rect 172363 525122 172421 525156
rect 172455 525122 172513 525156
rect 172547 525122 172605 525156
rect 172639 525122 172697 525156
rect 172731 525122 172789 525156
rect 172823 525122 172881 525156
rect 172915 525122 172973 525156
rect 173007 525122 173065 525156
rect 173099 525122 173157 525156
rect 173191 525122 173249 525156
rect 173283 525122 173341 525156
rect 173375 525122 173433 525156
rect 173467 525122 173525 525156
rect 173559 525122 173617 525156
rect 173651 525122 173709 525156
rect 173743 525122 173801 525156
rect 173835 525122 173893 525156
rect 173927 525122 173985 525156
rect 174019 525122 174077 525156
rect 174111 525122 174169 525156
rect 174203 525122 174261 525156
rect 174295 525122 174353 525156
rect 174387 525122 174445 525156
rect 174479 525122 174537 525156
rect 174571 525122 174623 525156
rect 172208 525113 174623 525122
rect 174675 525113 174687 525165
rect 174739 525156 174751 525165
rect 174803 525156 174815 525165
rect 174803 525122 174813 525156
rect 174739 525113 174751 525122
rect 174803 525113 174815 525122
rect 174867 525113 174879 525165
rect 174931 525156 178441 525165
rect 174939 525122 174997 525156
rect 175031 525122 175089 525156
rect 175123 525122 175181 525156
rect 175215 525122 175273 525156
rect 175307 525122 175365 525156
rect 175399 525122 175457 525156
rect 175491 525122 175549 525156
rect 175583 525122 175641 525156
rect 175675 525122 175733 525156
rect 175767 525122 175825 525156
rect 175859 525122 175917 525156
rect 175951 525122 176009 525156
rect 176043 525122 176101 525156
rect 176135 525122 176193 525156
rect 176227 525122 176285 525156
rect 176319 525122 176377 525156
rect 176411 525122 176469 525156
rect 176503 525122 176561 525156
rect 176595 525122 176653 525156
rect 176687 525122 176745 525156
rect 176779 525122 176837 525156
rect 176871 525122 176929 525156
rect 176963 525122 177021 525156
rect 177055 525122 177113 525156
rect 177147 525122 177205 525156
rect 177239 525122 177297 525156
rect 177331 525122 177389 525156
rect 177423 525122 177481 525156
rect 177515 525122 177573 525156
rect 177607 525122 177665 525156
rect 177699 525122 177757 525156
rect 177791 525122 177849 525156
rect 177883 525122 177941 525156
rect 177975 525122 178033 525156
rect 178067 525122 178125 525156
rect 178159 525122 178217 525156
rect 178251 525122 178309 525156
rect 178343 525122 178401 525156
rect 178435 525122 178441 525156
rect 174931 525113 178441 525122
rect 178493 525156 178505 525165
rect 178493 525113 178505 525122
rect 178557 525113 178569 525165
rect 178621 525113 178633 525165
rect 178685 525156 178697 525165
rect 178749 525156 182259 525165
rect 178749 525122 178769 525156
rect 178803 525122 178861 525156
rect 178895 525122 178953 525156
rect 178987 525122 179045 525156
rect 179079 525122 179137 525156
rect 179171 525122 179229 525156
rect 179263 525122 179321 525156
rect 179355 525122 179413 525156
rect 179447 525122 179505 525156
rect 179539 525122 179597 525156
rect 179631 525122 179689 525156
rect 179723 525122 179781 525156
rect 179815 525122 179873 525156
rect 179907 525122 179965 525156
rect 179999 525122 180057 525156
rect 180091 525122 180149 525156
rect 180183 525122 180241 525156
rect 180275 525122 180333 525156
rect 180367 525122 180425 525156
rect 180459 525122 180517 525156
rect 180551 525122 180609 525156
rect 180643 525122 180701 525156
rect 180735 525122 180793 525156
rect 180827 525122 180885 525156
rect 180919 525122 180977 525156
rect 181011 525122 181069 525156
rect 181103 525122 181161 525156
rect 181195 525122 181253 525156
rect 181287 525122 181345 525156
rect 181379 525122 181437 525156
rect 181471 525122 181529 525156
rect 181563 525122 181621 525156
rect 181655 525122 181713 525156
rect 181747 525122 181805 525156
rect 181839 525122 181897 525156
rect 181931 525122 181989 525156
rect 182023 525122 182081 525156
rect 182115 525122 182173 525156
rect 182207 525122 182259 525156
rect 178685 525113 178697 525122
rect 178749 525113 182259 525122
rect 182311 525113 182323 525165
rect 182375 525156 182387 525165
rect 182439 525156 182451 525165
rect 182439 525122 182449 525156
rect 182375 525113 182387 525122
rect 182439 525113 182451 525122
rect 182503 525113 182515 525165
rect 182567 525156 186077 525165
rect 182575 525122 182633 525156
rect 182667 525122 182725 525156
rect 182759 525122 182817 525156
rect 182851 525122 182909 525156
rect 182943 525122 183001 525156
rect 183035 525122 183093 525156
rect 183127 525122 183185 525156
rect 183219 525122 183277 525156
rect 183311 525122 183369 525156
rect 183403 525122 183461 525156
rect 183495 525122 183553 525156
rect 183587 525122 183645 525156
rect 183679 525122 183737 525156
rect 183771 525122 183829 525156
rect 183863 525122 183921 525156
rect 183955 525122 184013 525156
rect 184047 525122 184105 525156
rect 184139 525122 184197 525156
rect 184231 525122 184289 525156
rect 184323 525122 184381 525156
rect 184415 525122 184473 525156
rect 184507 525122 184565 525156
rect 184599 525122 184657 525156
rect 184691 525122 184749 525156
rect 184783 525122 184841 525156
rect 184875 525122 184933 525156
rect 184967 525122 185025 525156
rect 185059 525122 185117 525156
rect 185151 525122 185209 525156
rect 185243 525122 185301 525156
rect 185335 525122 185393 525156
rect 185427 525122 185485 525156
rect 185519 525122 185577 525156
rect 185611 525122 185669 525156
rect 185703 525122 185761 525156
rect 185795 525122 185853 525156
rect 185887 525122 185945 525156
rect 185979 525122 186037 525156
rect 186071 525122 186077 525156
rect 182567 525113 186077 525122
rect 186129 525156 186141 525165
rect 186129 525113 186141 525122
rect 186193 525113 186205 525165
rect 186257 525113 186269 525165
rect 186321 525156 186333 525165
rect 186385 525156 187480 525165
rect 186385 525122 186405 525156
rect 186439 525122 186497 525156
rect 186531 525122 186589 525156
rect 186623 525122 186681 525156
rect 186715 525122 186773 525156
rect 186807 525122 186865 525156
rect 186899 525122 186957 525156
rect 186991 525122 187049 525156
rect 187083 525122 187141 525156
rect 187175 525122 187233 525156
rect 187267 525122 187325 525156
rect 187359 525122 187417 525156
rect 187451 525122 187480 525156
rect 186321 525113 186333 525122
rect 186385 525113 187480 525122
rect 172208 525091 187480 525113
rect 172208 524621 187480 524643
rect 172208 524612 173963 524621
rect 174015 524612 174027 524621
rect 174079 524612 174091 524621
rect 172208 524578 172237 524612
rect 172271 524578 172329 524612
rect 172363 524578 172421 524612
rect 172455 524578 172513 524612
rect 172547 524578 172605 524612
rect 172639 524578 172697 524612
rect 172731 524578 172789 524612
rect 172823 524578 172881 524612
rect 172915 524578 172973 524612
rect 173007 524578 173065 524612
rect 173099 524578 173157 524612
rect 173191 524578 173249 524612
rect 173283 524578 173341 524612
rect 173375 524578 173433 524612
rect 173467 524578 173525 524612
rect 173559 524578 173617 524612
rect 173651 524578 173709 524612
rect 173743 524578 173801 524612
rect 173835 524578 173893 524612
rect 173927 524578 173963 524612
rect 174019 524578 174027 524612
rect 172208 524569 173963 524578
rect 174015 524569 174027 524578
rect 174079 524569 174091 524578
rect 174143 524569 174155 524621
rect 174207 524569 174219 524621
rect 174271 524612 177781 524621
rect 174295 524578 174353 524612
rect 174387 524578 174445 524612
rect 174479 524578 174537 524612
rect 174571 524578 174629 524612
rect 174663 524578 174721 524612
rect 174755 524578 174813 524612
rect 174847 524578 174905 524612
rect 174939 524578 174997 524612
rect 175031 524578 175089 524612
rect 175123 524578 175181 524612
rect 175215 524578 175273 524612
rect 175307 524578 175365 524612
rect 175399 524578 175457 524612
rect 175491 524578 175549 524612
rect 175583 524578 175641 524612
rect 175675 524578 175733 524612
rect 175767 524578 175825 524612
rect 175859 524578 175917 524612
rect 175951 524578 176009 524612
rect 176043 524578 176101 524612
rect 176135 524578 176193 524612
rect 176227 524578 176285 524612
rect 176319 524578 176377 524612
rect 176411 524578 176469 524612
rect 176503 524578 176561 524612
rect 176595 524578 176653 524612
rect 176687 524578 176745 524612
rect 176779 524578 176837 524612
rect 176871 524578 176929 524612
rect 176963 524578 177021 524612
rect 177055 524578 177113 524612
rect 177147 524578 177205 524612
rect 177239 524578 177297 524612
rect 177331 524578 177389 524612
rect 177423 524578 177481 524612
rect 177515 524578 177573 524612
rect 177607 524578 177665 524612
rect 177699 524578 177757 524612
rect 174271 524569 177781 524578
rect 177833 524569 177845 524621
rect 177897 524569 177909 524621
rect 177961 524612 177973 524621
rect 178025 524612 178037 524621
rect 178089 524612 181599 524621
rect 181651 524612 181663 524621
rect 181715 524612 181727 524621
rect 178025 524578 178033 524612
rect 178089 524578 178125 524612
rect 178159 524578 178217 524612
rect 178251 524578 178309 524612
rect 178343 524578 178401 524612
rect 178435 524578 178493 524612
rect 178527 524578 178585 524612
rect 178619 524578 178677 524612
rect 178711 524578 178769 524612
rect 178803 524578 178861 524612
rect 178895 524578 178953 524612
rect 178987 524578 179045 524612
rect 179079 524578 179137 524612
rect 179171 524578 179229 524612
rect 179263 524578 179321 524612
rect 179355 524578 179413 524612
rect 179447 524578 179505 524612
rect 179539 524578 179597 524612
rect 179631 524578 179689 524612
rect 179723 524578 179781 524612
rect 179815 524578 179873 524612
rect 179907 524578 179965 524612
rect 179999 524578 180057 524612
rect 180091 524578 180149 524612
rect 180183 524578 180241 524612
rect 180275 524578 180333 524612
rect 180367 524578 180425 524612
rect 180459 524578 180517 524612
rect 180551 524578 180609 524612
rect 180643 524578 180701 524612
rect 180735 524578 180793 524612
rect 180827 524578 180885 524612
rect 180919 524578 180977 524612
rect 181011 524578 181069 524612
rect 181103 524578 181161 524612
rect 181195 524578 181253 524612
rect 181287 524578 181345 524612
rect 181379 524578 181437 524612
rect 181471 524578 181529 524612
rect 181563 524578 181599 524612
rect 181655 524578 181663 524612
rect 177961 524569 177973 524578
rect 178025 524569 178037 524578
rect 178089 524569 181599 524578
rect 181651 524569 181663 524578
rect 181715 524569 181727 524578
rect 181779 524569 181791 524621
rect 181843 524569 181855 524621
rect 181907 524612 185417 524621
rect 181931 524578 181989 524612
rect 182023 524578 182081 524612
rect 182115 524578 182173 524612
rect 182207 524578 182265 524612
rect 182299 524578 182357 524612
rect 182391 524578 182449 524612
rect 182483 524578 182541 524612
rect 182575 524578 182633 524612
rect 182667 524578 182725 524612
rect 182759 524578 182817 524612
rect 182851 524578 182909 524612
rect 182943 524578 183001 524612
rect 183035 524578 183093 524612
rect 183127 524578 183185 524612
rect 183219 524578 183277 524612
rect 183311 524578 183369 524612
rect 183403 524578 183461 524612
rect 183495 524578 183553 524612
rect 183587 524578 183645 524612
rect 183679 524578 183737 524612
rect 183771 524578 183829 524612
rect 183863 524578 183921 524612
rect 183955 524578 184013 524612
rect 184047 524578 184105 524612
rect 184139 524578 184197 524612
rect 184231 524578 184289 524612
rect 184323 524578 184381 524612
rect 184415 524578 184473 524612
rect 184507 524578 184565 524612
rect 184599 524578 184657 524612
rect 184691 524578 184749 524612
rect 184783 524578 184841 524612
rect 184875 524578 184933 524612
rect 184967 524578 185025 524612
rect 185059 524578 185117 524612
rect 185151 524578 185209 524612
rect 185243 524578 185301 524612
rect 185335 524578 185393 524612
rect 181907 524569 185417 524578
rect 185469 524569 185481 524621
rect 185533 524569 185545 524621
rect 185597 524612 185609 524621
rect 185661 524612 185673 524621
rect 185725 524612 187480 524621
rect 185661 524578 185669 524612
rect 185725 524578 185761 524612
rect 185795 524578 185853 524612
rect 185887 524578 185945 524612
rect 185979 524578 186037 524612
rect 186071 524578 186129 524612
rect 186163 524578 186221 524612
rect 186255 524578 186313 524612
rect 186347 524578 186405 524612
rect 186439 524578 186497 524612
rect 186531 524578 186589 524612
rect 186623 524578 186681 524612
rect 186715 524578 186773 524612
rect 186807 524578 186865 524612
rect 186899 524578 186957 524612
rect 186991 524578 187049 524612
rect 187083 524578 187141 524612
rect 187175 524578 187233 524612
rect 187267 524578 187325 524612
rect 187359 524578 187417 524612
rect 187451 524578 187480 524612
rect 185597 524569 185609 524578
rect 185661 524569 185673 524578
rect 185725 524569 187480 524578
rect 172208 524547 187480 524569
rect 172208 524077 187480 524099
rect 172208 524068 174623 524077
rect 172208 524034 172237 524068
rect 172271 524034 172329 524068
rect 172363 524034 172421 524068
rect 172455 524034 172513 524068
rect 172547 524034 172605 524068
rect 172639 524034 172697 524068
rect 172731 524034 172789 524068
rect 172823 524034 172881 524068
rect 172915 524034 172973 524068
rect 173007 524034 173065 524068
rect 173099 524034 173157 524068
rect 173191 524034 173249 524068
rect 173283 524034 173341 524068
rect 173375 524034 173433 524068
rect 173467 524034 173525 524068
rect 173559 524034 173617 524068
rect 173651 524034 173709 524068
rect 173743 524034 173801 524068
rect 173835 524034 173893 524068
rect 173927 524034 173985 524068
rect 174019 524034 174077 524068
rect 174111 524034 174169 524068
rect 174203 524034 174261 524068
rect 174295 524034 174353 524068
rect 174387 524034 174445 524068
rect 174479 524034 174537 524068
rect 174571 524034 174623 524068
rect 172208 524025 174623 524034
rect 174675 524025 174687 524077
rect 174739 524068 174751 524077
rect 174803 524068 174815 524077
rect 174803 524034 174813 524068
rect 174739 524025 174751 524034
rect 174803 524025 174815 524034
rect 174867 524025 174879 524077
rect 174931 524068 178441 524077
rect 174939 524034 174997 524068
rect 175031 524034 175089 524068
rect 175123 524034 175181 524068
rect 175215 524034 175273 524068
rect 175307 524034 175365 524068
rect 175399 524034 175457 524068
rect 175491 524034 175549 524068
rect 175583 524034 175641 524068
rect 175675 524034 175733 524068
rect 175767 524034 175825 524068
rect 175859 524034 175917 524068
rect 175951 524034 176009 524068
rect 176043 524034 176101 524068
rect 176135 524034 176193 524068
rect 176227 524034 176285 524068
rect 176319 524034 176377 524068
rect 176411 524034 176469 524068
rect 176503 524034 176561 524068
rect 176595 524034 176653 524068
rect 176687 524034 176745 524068
rect 176779 524034 176837 524068
rect 176871 524034 176929 524068
rect 176963 524034 177021 524068
rect 177055 524034 177113 524068
rect 177147 524034 177205 524068
rect 177239 524034 177297 524068
rect 177331 524034 177389 524068
rect 177423 524034 177481 524068
rect 177515 524034 177573 524068
rect 177607 524034 177665 524068
rect 177699 524034 177757 524068
rect 177791 524034 177849 524068
rect 177883 524034 177941 524068
rect 177975 524034 178033 524068
rect 178067 524034 178125 524068
rect 178159 524034 178217 524068
rect 178251 524034 178309 524068
rect 178343 524034 178401 524068
rect 178435 524034 178441 524068
rect 174931 524025 178441 524034
rect 178493 524068 178505 524077
rect 178493 524025 178505 524034
rect 178557 524025 178569 524077
rect 178621 524025 178633 524077
rect 178685 524068 178697 524077
rect 178749 524068 182259 524077
rect 178749 524034 178769 524068
rect 178803 524034 178861 524068
rect 178895 524034 178953 524068
rect 178987 524034 179045 524068
rect 179079 524034 179137 524068
rect 179171 524034 179229 524068
rect 179263 524034 179321 524068
rect 179355 524034 179413 524068
rect 179447 524034 179505 524068
rect 179539 524034 179597 524068
rect 179631 524034 179689 524068
rect 179723 524034 179781 524068
rect 179815 524034 179873 524068
rect 179907 524034 179965 524068
rect 179999 524034 180057 524068
rect 180091 524034 180149 524068
rect 180183 524034 180241 524068
rect 180275 524034 180333 524068
rect 180367 524034 180425 524068
rect 180459 524034 180517 524068
rect 180551 524034 180609 524068
rect 180643 524034 180701 524068
rect 180735 524034 180793 524068
rect 180827 524034 180885 524068
rect 180919 524034 180977 524068
rect 181011 524034 181069 524068
rect 181103 524034 181161 524068
rect 181195 524034 181253 524068
rect 181287 524034 181345 524068
rect 181379 524034 181437 524068
rect 181471 524034 181529 524068
rect 181563 524034 181621 524068
rect 181655 524034 181713 524068
rect 181747 524034 181805 524068
rect 181839 524034 181897 524068
rect 181931 524034 181989 524068
rect 182023 524034 182081 524068
rect 182115 524034 182173 524068
rect 182207 524034 182259 524068
rect 178685 524025 178697 524034
rect 178749 524025 182259 524034
rect 182311 524025 182323 524077
rect 182375 524068 182387 524077
rect 182439 524068 182451 524077
rect 182439 524034 182449 524068
rect 182375 524025 182387 524034
rect 182439 524025 182451 524034
rect 182503 524025 182515 524077
rect 182567 524068 186077 524077
rect 182575 524034 182633 524068
rect 182667 524034 182725 524068
rect 182759 524034 182817 524068
rect 182851 524034 182909 524068
rect 182943 524034 183001 524068
rect 183035 524034 183093 524068
rect 183127 524034 183185 524068
rect 183219 524034 183277 524068
rect 183311 524034 183369 524068
rect 183403 524034 183461 524068
rect 183495 524034 183553 524068
rect 183587 524034 183645 524068
rect 183679 524034 183737 524068
rect 183771 524034 183829 524068
rect 183863 524034 183921 524068
rect 183955 524034 184013 524068
rect 184047 524034 184105 524068
rect 184139 524034 184197 524068
rect 184231 524034 184289 524068
rect 184323 524034 184381 524068
rect 184415 524034 184473 524068
rect 184507 524034 184565 524068
rect 184599 524034 184657 524068
rect 184691 524034 184749 524068
rect 184783 524034 184841 524068
rect 184875 524034 184933 524068
rect 184967 524034 185025 524068
rect 185059 524034 185117 524068
rect 185151 524034 185209 524068
rect 185243 524034 185301 524068
rect 185335 524034 185393 524068
rect 185427 524034 185485 524068
rect 185519 524034 185577 524068
rect 185611 524034 185669 524068
rect 185703 524034 185761 524068
rect 185795 524034 185853 524068
rect 185887 524034 185945 524068
rect 185979 524034 186037 524068
rect 186071 524034 186077 524068
rect 182567 524025 186077 524034
rect 186129 524068 186141 524077
rect 186129 524025 186141 524034
rect 186193 524025 186205 524077
rect 186257 524025 186269 524077
rect 186321 524068 186333 524077
rect 186385 524068 187480 524077
rect 186385 524034 186405 524068
rect 186439 524034 186497 524068
rect 186531 524034 186589 524068
rect 186623 524034 186681 524068
rect 186715 524034 186773 524068
rect 186807 524034 186865 524068
rect 186899 524034 186957 524068
rect 186991 524034 187049 524068
rect 187083 524034 187141 524068
rect 187175 524034 187233 524068
rect 187267 524034 187325 524068
rect 187359 524034 187417 524068
rect 187451 524034 187480 524068
rect 186321 524025 186333 524034
rect 186385 524025 187480 524034
rect 172208 524003 187480 524025
rect 193000 524000 195000 526000
rect 192428 523570 192628 523585
rect 193000 523570 193130 524000
rect 192428 523555 193130 523570
rect 172208 523533 193130 523555
rect 172208 523524 173963 523533
rect 174015 523524 174027 523533
rect 174079 523524 174091 523533
rect 172208 523490 172237 523524
rect 172271 523490 172329 523524
rect 172363 523490 172421 523524
rect 172455 523490 172513 523524
rect 172547 523490 172605 523524
rect 172639 523490 172697 523524
rect 172731 523490 172789 523524
rect 172823 523490 172881 523524
rect 172915 523490 172973 523524
rect 173007 523490 173065 523524
rect 173099 523490 173157 523524
rect 173191 523490 173249 523524
rect 173283 523490 173341 523524
rect 173375 523490 173433 523524
rect 173467 523490 173525 523524
rect 173559 523490 173617 523524
rect 173651 523490 173709 523524
rect 173743 523490 173801 523524
rect 173835 523490 173893 523524
rect 173927 523490 173963 523524
rect 174019 523490 174027 523524
rect 172208 523481 173963 523490
rect 174015 523481 174027 523490
rect 174079 523481 174091 523490
rect 174143 523481 174155 523533
rect 174207 523481 174219 523533
rect 174271 523524 177781 523533
rect 174295 523490 174353 523524
rect 174387 523490 174445 523524
rect 174479 523490 174537 523524
rect 174571 523490 174629 523524
rect 174663 523490 174721 523524
rect 174755 523490 174813 523524
rect 174847 523490 174905 523524
rect 174939 523490 174997 523524
rect 175031 523490 175089 523524
rect 175123 523490 175181 523524
rect 175215 523490 175273 523524
rect 175307 523490 175365 523524
rect 175399 523490 175457 523524
rect 175491 523490 175549 523524
rect 175583 523490 175641 523524
rect 175675 523490 175733 523524
rect 175767 523490 175825 523524
rect 175859 523490 175917 523524
rect 175951 523490 176009 523524
rect 176043 523490 176101 523524
rect 176135 523490 176193 523524
rect 176227 523490 176285 523524
rect 176319 523490 176377 523524
rect 176411 523490 176469 523524
rect 176503 523490 176561 523524
rect 176595 523490 176653 523524
rect 176687 523490 176745 523524
rect 176779 523490 176837 523524
rect 176871 523490 176929 523524
rect 176963 523490 177021 523524
rect 177055 523490 177113 523524
rect 177147 523490 177205 523524
rect 177239 523490 177297 523524
rect 177331 523490 177389 523524
rect 177423 523490 177481 523524
rect 177515 523490 177573 523524
rect 177607 523490 177665 523524
rect 177699 523490 177757 523524
rect 174271 523481 177781 523490
rect 177833 523481 177845 523533
rect 177897 523481 177909 523533
rect 177961 523524 177973 523533
rect 178025 523524 178037 523533
rect 178089 523524 181599 523533
rect 181651 523524 181663 523533
rect 181715 523524 181727 523533
rect 178025 523490 178033 523524
rect 178089 523490 178125 523524
rect 178159 523490 178217 523524
rect 178251 523490 178309 523524
rect 178343 523490 178401 523524
rect 178435 523490 178493 523524
rect 178527 523490 178585 523524
rect 178619 523490 178677 523524
rect 178711 523490 178769 523524
rect 178803 523490 178861 523524
rect 178895 523490 178953 523524
rect 178987 523490 179045 523524
rect 179079 523490 179137 523524
rect 179171 523490 179229 523524
rect 179263 523490 179321 523524
rect 179355 523490 179413 523524
rect 179447 523490 179505 523524
rect 179539 523490 179597 523524
rect 179631 523490 179689 523524
rect 179723 523490 179781 523524
rect 179815 523490 179873 523524
rect 179907 523490 179965 523524
rect 179999 523490 180057 523524
rect 180091 523490 180149 523524
rect 180183 523490 180241 523524
rect 180275 523490 180333 523524
rect 180367 523490 180425 523524
rect 180459 523490 180517 523524
rect 180551 523490 180609 523524
rect 180643 523490 180701 523524
rect 180735 523490 180793 523524
rect 180827 523490 180885 523524
rect 180919 523490 180977 523524
rect 181011 523490 181069 523524
rect 181103 523490 181161 523524
rect 181195 523490 181253 523524
rect 181287 523490 181345 523524
rect 181379 523490 181437 523524
rect 181471 523490 181529 523524
rect 181563 523490 181599 523524
rect 181655 523490 181663 523524
rect 177961 523481 177973 523490
rect 178025 523481 178037 523490
rect 178089 523481 181599 523490
rect 181651 523481 181663 523490
rect 181715 523481 181727 523490
rect 181779 523481 181791 523533
rect 181843 523481 181855 523533
rect 181907 523524 185417 523533
rect 181931 523490 181989 523524
rect 182023 523490 182081 523524
rect 182115 523490 182173 523524
rect 182207 523490 182265 523524
rect 182299 523490 182357 523524
rect 182391 523490 182449 523524
rect 182483 523490 182541 523524
rect 182575 523490 182633 523524
rect 182667 523490 182725 523524
rect 182759 523490 182817 523524
rect 182851 523490 182909 523524
rect 182943 523490 183001 523524
rect 183035 523490 183093 523524
rect 183127 523490 183185 523524
rect 183219 523490 183277 523524
rect 183311 523490 183369 523524
rect 183403 523490 183461 523524
rect 183495 523490 183553 523524
rect 183587 523490 183645 523524
rect 183679 523490 183737 523524
rect 183771 523490 183829 523524
rect 183863 523490 183921 523524
rect 183955 523490 184013 523524
rect 184047 523490 184105 523524
rect 184139 523490 184197 523524
rect 184231 523490 184289 523524
rect 184323 523490 184381 523524
rect 184415 523490 184473 523524
rect 184507 523490 184565 523524
rect 184599 523490 184657 523524
rect 184691 523490 184749 523524
rect 184783 523490 184841 523524
rect 184875 523490 184933 523524
rect 184967 523490 185025 523524
rect 185059 523490 185117 523524
rect 185151 523490 185209 523524
rect 185243 523490 185301 523524
rect 185335 523490 185393 523524
rect 181907 523481 185417 523490
rect 185469 523481 185481 523533
rect 185533 523481 185545 523533
rect 185597 523524 185609 523533
rect 185661 523524 185673 523533
rect 185725 523524 193130 523533
rect 185661 523490 185669 523524
rect 185725 523490 185761 523524
rect 185795 523490 185853 523524
rect 185887 523490 185945 523524
rect 185979 523490 186037 523524
rect 186071 523490 186129 523524
rect 186163 523490 186221 523524
rect 186255 523490 186313 523524
rect 186347 523490 186405 523524
rect 186439 523490 186497 523524
rect 186531 523490 186589 523524
rect 186623 523490 186681 523524
rect 186715 523490 186773 523524
rect 186807 523490 186865 523524
rect 186899 523490 186957 523524
rect 186991 523490 187049 523524
rect 187083 523490 187141 523524
rect 187175 523490 187233 523524
rect 187267 523490 187325 523524
rect 187359 523490 187417 523524
rect 187451 523490 193130 523524
rect 185597 523481 185609 523490
rect 185661 523481 185673 523490
rect 185725 523481 193130 523490
rect 172208 523459 193130 523481
rect 187468 523455 193130 523459
rect 192428 523450 193130 523455
rect 192428 523395 192628 523450
rect 172208 523005 187480 523011
rect 192428 523010 192628 523065
rect 192428 523005 193020 523010
rect 172208 522989 192108 523005
rect 172208 522980 174623 522989
rect 172208 522946 172237 522980
rect 172271 522946 172329 522980
rect 172363 522946 172421 522980
rect 172455 522946 172513 522980
rect 172547 522946 172605 522980
rect 172639 522946 172697 522980
rect 172731 522946 172789 522980
rect 172823 522946 172881 522980
rect 172915 522946 172973 522980
rect 173007 522946 173065 522980
rect 173099 522946 173157 522980
rect 173191 522946 173249 522980
rect 173283 522946 173341 522980
rect 173375 522946 173433 522980
rect 173467 522946 173525 522980
rect 173559 522946 173617 522980
rect 173651 522946 173709 522980
rect 173743 522946 173801 522980
rect 173835 522946 173893 522980
rect 173927 522946 173985 522980
rect 174019 522946 174077 522980
rect 174111 522946 174169 522980
rect 174203 522946 174261 522980
rect 174295 522946 174353 522980
rect 174387 522946 174445 522980
rect 174479 522946 174537 522980
rect 174571 522946 174623 522980
rect 172208 522937 174623 522946
rect 174675 522937 174687 522989
rect 174739 522980 174751 522989
rect 174803 522980 174815 522989
rect 174803 522946 174813 522980
rect 174739 522937 174751 522946
rect 174803 522937 174815 522946
rect 174867 522937 174879 522989
rect 174931 522980 178441 522989
rect 174939 522946 174997 522980
rect 175031 522946 175089 522980
rect 175123 522946 175181 522980
rect 175215 522946 175273 522980
rect 175307 522946 175365 522980
rect 175399 522946 175457 522980
rect 175491 522946 175549 522980
rect 175583 522946 175641 522980
rect 175675 522946 175733 522980
rect 175767 522946 175825 522980
rect 175859 522946 175917 522980
rect 175951 522946 176009 522980
rect 176043 522946 176101 522980
rect 176135 522946 176193 522980
rect 176227 522946 176285 522980
rect 176319 522946 176377 522980
rect 176411 522946 176469 522980
rect 176503 522946 176561 522980
rect 176595 522946 176653 522980
rect 176687 522946 176745 522980
rect 176779 522946 176837 522980
rect 176871 522946 176929 522980
rect 176963 522946 177021 522980
rect 177055 522946 177113 522980
rect 177147 522946 177205 522980
rect 177239 522946 177297 522980
rect 177331 522946 177389 522980
rect 177423 522946 177481 522980
rect 177515 522946 177573 522980
rect 177607 522946 177665 522980
rect 177699 522946 177757 522980
rect 177791 522946 177849 522980
rect 177883 522946 177941 522980
rect 177975 522946 178033 522980
rect 178067 522946 178125 522980
rect 178159 522946 178217 522980
rect 178251 522946 178309 522980
rect 178343 522946 178401 522980
rect 178435 522946 178441 522980
rect 174931 522937 178441 522946
rect 178493 522980 178505 522989
rect 178493 522937 178505 522946
rect 178557 522937 178569 522989
rect 178621 522937 178633 522989
rect 178685 522980 178697 522989
rect 178749 522980 182259 522989
rect 178749 522946 178769 522980
rect 178803 522946 178861 522980
rect 178895 522946 178953 522980
rect 178987 522946 179045 522980
rect 179079 522946 179137 522980
rect 179171 522946 179229 522980
rect 179263 522946 179321 522980
rect 179355 522946 179413 522980
rect 179447 522946 179505 522980
rect 179539 522946 179597 522980
rect 179631 522946 179689 522980
rect 179723 522946 179781 522980
rect 179815 522946 179873 522980
rect 179907 522946 179965 522980
rect 179999 522946 180057 522980
rect 180091 522946 180149 522980
rect 180183 522946 180241 522980
rect 180275 522946 180333 522980
rect 180367 522946 180425 522980
rect 180459 522946 180517 522980
rect 180551 522946 180609 522980
rect 180643 522946 180701 522980
rect 180735 522946 180793 522980
rect 180827 522946 180885 522980
rect 180919 522946 180977 522980
rect 181011 522946 181069 522980
rect 181103 522946 181161 522980
rect 181195 522946 181253 522980
rect 181287 522946 181345 522980
rect 181379 522946 181437 522980
rect 181471 522946 181529 522980
rect 181563 522946 181621 522980
rect 181655 522946 181713 522980
rect 181747 522946 181805 522980
rect 181839 522946 181897 522980
rect 181931 522946 181989 522980
rect 182023 522946 182081 522980
rect 182115 522946 182173 522980
rect 182207 522946 182259 522980
rect 178685 522937 178697 522946
rect 178749 522937 182259 522946
rect 182311 522937 182323 522989
rect 182375 522980 182387 522989
rect 182439 522980 182451 522989
rect 182439 522946 182449 522980
rect 182375 522937 182387 522946
rect 182439 522937 182451 522946
rect 182503 522937 182515 522989
rect 182567 522980 186077 522989
rect 182575 522946 182633 522980
rect 182667 522946 182725 522980
rect 182759 522946 182817 522980
rect 182851 522946 182909 522980
rect 182943 522946 183001 522980
rect 183035 522946 183093 522980
rect 183127 522946 183185 522980
rect 183219 522946 183277 522980
rect 183311 522946 183369 522980
rect 183403 522946 183461 522980
rect 183495 522946 183553 522980
rect 183587 522946 183645 522980
rect 183679 522946 183737 522980
rect 183771 522946 183829 522980
rect 183863 522946 183921 522980
rect 183955 522946 184013 522980
rect 184047 522946 184105 522980
rect 184139 522946 184197 522980
rect 184231 522946 184289 522980
rect 184323 522946 184381 522980
rect 184415 522946 184473 522980
rect 184507 522946 184565 522980
rect 184599 522946 184657 522980
rect 184691 522946 184749 522980
rect 184783 522946 184841 522980
rect 184875 522946 184933 522980
rect 184967 522946 185025 522980
rect 185059 522946 185117 522980
rect 185151 522946 185209 522980
rect 185243 522946 185301 522980
rect 185335 522946 185393 522980
rect 185427 522946 185485 522980
rect 185519 522946 185577 522980
rect 185611 522946 185669 522980
rect 185703 522946 185761 522980
rect 185795 522946 185853 522980
rect 185887 522946 185945 522980
rect 185979 522946 186037 522980
rect 186071 522946 186077 522980
rect 182567 522937 186077 522946
rect 186129 522980 186141 522989
rect 186129 522937 186141 522946
rect 186193 522937 186205 522989
rect 186257 522937 186269 522989
rect 186321 522980 186333 522989
rect 186385 522980 192108 522989
rect 186385 522946 186405 522980
rect 186439 522946 186497 522980
rect 186531 522946 186589 522980
rect 186623 522946 186681 522980
rect 186715 522946 186773 522980
rect 186807 522946 186865 522980
rect 186899 522946 186957 522980
rect 186991 522946 187049 522980
rect 187083 522946 187141 522980
rect 187175 522946 187233 522980
rect 187267 522946 187325 522980
rect 187359 522946 187417 522980
rect 187451 522946 192108 522980
rect 186321 522937 186333 522946
rect 186385 522937 192108 522946
rect 172208 522915 192108 522937
rect 192138 523000 193020 523005
rect 192138 522915 195000 523000
rect 192428 522910 195000 522915
rect 192428 522875 192628 522910
rect 172208 522445 187480 522467
rect 172208 522436 173963 522445
rect 174015 522436 174027 522445
rect 174079 522436 174091 522445
rect 172208 522402 172237 522436
rect 172271 522402 172329 522436
rect 172363 522402 172421 522436
rect 172455 522402 172513 522436
rect 172547 522402 172605 522436
rect 172639 522402 172697 522436
rect 172731 522402 172789 522436
rect 172823 522402 172881 522436
rect 172915 522402 172973 522436
rect 173007 522402 173065 522436
rect 173099 522402 173157 522436
rect 173191 522402 173249 522436
rect 173283 522402 173341 522436
rect 173375 522402 173433 522436
rect 173467 522402 173525 522436
rect 173559 522402 173617 522436
rect 173651 522402 173709 522436
rect 173743 522402 173801 522436
rect 173835 522402 173893 522436
rect 173927 522402 173963 522436
rect 174019 522402 174027 522436
rect 172208 522393 173963 522402
rect 174015 522393 174027 522402
rect 174079 522393 174091 522402
rect 174143 522393 174155 522445
rect 174207 522393 174219 522445
rect 174271 522436 177781 522445
rect 174295 522402 174353 522436
rect 174387 522402 174445 522436
rect 174479 522402 174537 522436
rect 174571 522402 174629 522436
rect 174663 522402 174721 522436
rect 174755 522402 174813 522436
rect 174847 522402 174905 522436
rect 174939 522402 174997 522436
rect 175031 522402 175089 522436
rect 175123 522402 175181 522436
rect 175215 522402 175273 522436
rect 175307 522402 175365 522436
rect 175399 522402 175457 522436
rect 175491 522402 175549 522436
rect 175583 522402 175641 522436
rect 175675 522402 175733 522436
rect 175767 522402 175825 522436
rect 175859 522402 175917 522436
rect 175951 522402 176009 522436
rect 176043 522402 176101 522436
rect 176135 522402 176193 522436
rect 176227 522402 176285 522436
rect 176319 522402 176377 522436
rect 176411 522402 176469 522436
rect 176503 522402 176561 522436
rect 176595 522402 176653 522436
rect 176687 522402 176745 522436
rect 176779 522402 176837 522436
rect 176871 522402 176929 522436
rect 176963 522402 177021 522436
rect 177055 522402 177113 522436
rect 177147 522402 177205 522436
rect 177239 522402 177297 522436
rect 177331 522402 177389 522436
rect 177423 522402 177481 522436
rect 177515 522402 177573 522436
rect 177607 522402 177665 522436
rect 177699 522402 177757 522436
rect 174271 522393 177781 522402
rect 177833 522393 177845 522445
rect 177897 522393 177909 522445
rect 177961 522436 177973 522445
rect 178025 522436 178037 522445
rect 178089 522436 181599 522445
rect 181651 522436 181663 522445
rect 181715 522436 181727 522445
rect 178025 522402 178033 522436
rect 178089 522402 178125 522436
rect 178159 522402 178217 522436
rect 178251 522402 178309 522436
rect 178343 522402 178401 522436
rect 178435 522402 178493 522436
rect 178527 522402 178585 522436
rect 178619 522402 178677 522436
rect 178711 522402 178769 522436
rect 178803 522402 178861 522436
rect 178895 522402 178953 522436
rect 178987 522402 179045 522436
rect 179079 522402 179137 522436
rect 179171 522402 179229 522436
rect 179263 522402 179321 522436
rect 179355 522402 179413 522436
rect 179447 522402 179505 522436
rect 179539 522402 179597 522436
rect 179631 522402 179689 522436
rect 179723 522402 179781 522436
rect 179815 522402 179873 522436
rect 179907 522402 179965 522436
rect 179999 522402 180057 522436
rect 180091 522402 180149 522436
rect 180183 522402 180241 522436
rect 180275 522402 180333 522436
rect 180367 522402 180425 522436
rect 180459 522402 180517 522436
rect 180551 522402 180609 522436
rect 180643 522402 180701 522436
rect 180735 522402 180793 522436
rect 180827 522402 180885 522436
rect 180919 522402 180977 522436
rect 181011 522402 181069 522436
rect 181103 522402 181161 522436
rect 181195 522402 181253 522436
rect 181287 522402 181345 522436
rect 181379 522402 181437 522436
rect 181471 522402 181529 522436
rect 181563 522402 181599 522436
rect 181655 522402 181663 522436
rect 177961 522393 177973 522402
rect 178025 522393 178037 522402
rect 178089 522393 181599 522402
rect 181651 522393 181663 522402
rect 181715 522393 181727 522402
rect 181779 522393 181791 522445
rect 181843 522393 181855 522445
rect 181907 522436 185417 522445
rect 181931 522402 181989 522436
rect 182023 522402 182081 522436
rect 182115 522402 182173 522436
rect 182207 522402 182265 522436
rect 182299 522402 182357 522436
rect 182391 522402 182449 522436
rect 182483 522402 182541 522436
rect 182575 522402 182633 522436
rect 182667 522402 182725 522436
rect 182759 522402 182817 522436
rect 182851 522402 182909 522436
rect 182943 522402 183001 522436
rect 183035 522402 183093 522436
rect 183127 522402 183185 522436
rect 183219 522402 183277 522436
rect 183311 522402 183369 522436
rect 183403 522402 183461 522436
rect 183495 522402 183553 522436
rect 183587 522402 183645 522436
rect 183679 522402 183737 522436
rect 183771 522402 183829 522436
rect 183863 522402 183921 522436
rect 183955 522402 184013 522436
rect 184047 522402 184105 522436
rect 184139 522402 184197 522436
rect 184231 522402 184289 522436
rect 184323 522402 184381 522436
rect 184415 522402 184473 522436
rect 184507 522402 184565 522436
rect 184599 522402 184657 522436
rect 184691 522402 184749 522436
rect 184783 522402 184841 522436
rect 184875 522402 184933 522436
rect 184967 522402 185025 522436
rect 185059 522402 185117 522436
rect 185151 522402 185209 522436
rect 185243 522402 185301 522436
rect 185335 522402 185393 522436
rect 181907 522393 185417 522402
rect 185469 522393 185481 522445
rect 185533 522393 185545 522445
rect 185597 522436 185609 522445
rect 185661 522436 185673 522445
rect 185725 522436 187480 522445
rect 185661 522402 185669 522436
rect 185725 522402 185761 522436
rect 185795 522402 185853 522436
rect 185887 522402 185945 522436
rect 185979 522402 186037 522436
rect 186071 522402 186129 522436
rect 186163 522402 186221 522436
rect 186255 522402 186313 522436
rect 186347 522402 186405 522436
rect 186439 522402 186497 522436
rect 186531 522402 186589 522436
rect 186623 522402 186681 522436
rect 186715 522402 186773 522436
rect 186807 522402 186865 522436
rect 186899 522402 186957 522436
rect 186991 522402 187049 522436
rect 187083 522402 187141 522436
rect 187175 522402 187233 522436
rect 187267 522402 187325 522436
rect 187359 522402 187417 522436
rect 187451 522402 187480 522436
rect 185597 522393 185609 522402
rect 185661 522393 185673 522402
rect 185725 522393 187480 522402
rect 172208 522371 187480 522393
rect 172208 521901 187480 521923
rect 172208 521892 174623 521901
rect 172208 521858 172237 521892
rect 172271 521858 172329 521892
rect 172363 521858 172421 521892
rect 172455 521858 172513 521892
rect 172547 521858 172605 521892
rect 172639 521858 172697 521892
rect 172731 521858 172789 521892
rect 172823 521858 172881 521892
rect 172915 521858 172973 521892
rect 173007 521858 173065 521892
rect 173099 521858 173157 521892
rect 173191 521858 173249 521892
rect 173283 521858 173341 521892
rect 173375 521858 173433 521892
rect 173467 521858 173525 521892
rect 173559 521858 173617 521892
rect 173651 521858 173709 521892
rect 173743 521858 173801 521892
rect 173835 521858 173893 521892
rect 173927 521858 173985 521892
rect 174019 521858 174077 521892
rect 174111 521858 174169 521892
rect 174203 521858 174261 521892
rect 174295 521858 174353 521892
rect 174387 521858 174445 521892
rect 174479 521858 174537 521892
rect 174571 521858 174623 521892
rect 172208 521849 174623 521858
rect 174675 521849 174687 521901
rect 174739 521892 174751 521901
rect 174803 521892 174815 521901
rect 174803 521858 174813 521892
rect 174739 521849 174751 521858
rect 174803 521849 174815 521858
rect 174867 521849 174879 521901
rect 174931 521892 178441 521901
rect 174939 521858 174997 521892
rect 175031 521858 175089 521892
rect 175123 521858 175181 521892
rect 175215 521858 175273 521892
rect 175307 521858 175365 521892
rect 175399 521858 175457 521892
rect 175491 521858 175549 521892
rect 175583 521858 175641 521892
rect 175675 521858 175733 521892
rect 175767 521858 175825 521892
rect 175859 521858 175917 521892
rect 175951 521858 176009 521892
rect 176043 521858 176101 521892
rect 176135 521858 176193 521892
rect 176227 521858 176285 521892
rect 176319 521858 176377 521892
rect 176411 521858 176469 521892
rect 176503 521858 176561 521892
rect 176595 521858 176653 521892
rect 176687 521858 176745 521892
rect 176779 521858 176837 521892
rect 176871 521858 176929 521892
rect 176963 521858 177021 521892
rect 177055 521858 177113 521892
rect 177147 521858 177205 521892
rect 177239 521858 177297 521892
rect 177331 521858 177389 521892
rect 177423 521858 177481 521892
rect 177515 521858 177573 521892
rect 177607 521858 177665 521892
rect 177699 521858 177757 521892
rect 177791 521858 177849 521892
rect 177883 521858 177941 521892
rect 177975 521858 178033 521892
rect 178067 521858 178125 521892
rect 178159 521858 178217 521892
rect 178251 521858 178309 521892
rect 178343 521858 178401 521892
rect 178435 521858 178441 521892
rect 174931 521849 178441 521858
rect 178493 521892 178505 521901
rect 178493 521849 178505 521858
rect 178557 521849 178569 521901
rect 178621 521849 178633 521901
rect 178685 521892 178697 521901
rect 178749 521892 182259 521901
rect 178749 521858 178769 521892
rect 178803 521858 178861 521892
rect 178895 521858 178953 521892
rect 178987 521858 179045 521892
rect 179079 521858 179137 521892
rect 179171 521858 179229 521892
rect 179263 521858 179321 521892
rect 179355 521858 179413 521892
rect 179447 521858 179505 521892
rect 179539 521858 179597 521892
rect 179631 521858 179689 521892
rect 179723 521858 179781 521892
rect 179815 521858 179873 521892
rect 179907 521858 179965 521892
rect 179999 521858 180057 521892
rect 180091 521858 180149 521892
rect 180183 521858 180241 521892
rect 180275 521858 180333 521892
rect 180367 521858 180425 521892
rect 180459 521858 180517 521892
rect 180551 521858 180609 521892
rect 180643 521858 180701 521892
rect 180735 521858 180793 521892
rect 180827 521858 180885 521892
rect 180919 521858 180977 521892
rect 181011 521858 181069 521892
rect 181103 521858 181161 521892
rect 181195 521858 181253 521892
rect 181287 521858 181345 521892
rect 181379 521858 181437 521892
rect 181471 521858 181529 521892
rect 181563 521858 181621 521892
rect 181655 521858 181713 521892
rect 181747 521858 181805 521892
rect 181839 521858 181897 521892
rect 181931 521858 181989 521892
rect 182023 521858 182081 521892
rect 182115 521858 182173 521892
rect 182207 521858 182259 521892
rect 178685 521849 178697 521858
rect 178749 521849 182259 521858
rect 182311 521849 182323 521901
rect 182375 521892 182387 521901
rect 182439 521892 182451 521901
rect 182439 521858 182449 521892
rect 182375 521849 182387 521858
rect 182439 521849 182451 521858
rect 182503 521849 182515 521901
rect 182567 521892 186077 521901
rect 182575 521858 182633 521892
rect 182667 521858 182725 521892
rect 182759 521858 182817 521892
rect 182851 521858 182909 521892
rect 182943 521858 183001 521892
rect 183035 521858 183093 521892
rect 183127 521858 183185 521892
rect 183219 521858 183277 521892
rect 183311 521858 183369 521892
rect 183403 521858 183461 521892
rect 183495 521858 183553 521892
rect 183587 521858 183645 521892
rect 183679 521858 183737 521892
rect 183771 521858 183829 521892
rect 183863 521858 183921 521892
rect 183955 521858 184013 521892
rect 184047 521858 184105 521892
rect 184139 521858 184197 521892
rect 184231 521858 184289 521892
rect 184323 521858 184381 521892
rect 184415 521858 184473 521892
rect 184507 521858 184565 521892
rect 184599 521858 184657 521892
rect 184691 521858 184749 521892
rect 184783 521858 184841 521892
rect 184875 521858 184933 521892
rect 184967 521858 185025 521892
rect 185059 521858 185117 521892
rect 185151 521858 185209 521892
rect 185243 521858 185301 521892
rect 185335 521858 185393 521892
rect 185427 521858 185485 521892
rect 185519 521858 185577 521892
rect 185611 521858 185669 521892
rect 185703 521858 185761 521892
rect 185795 521858 185853 521892
rect 185887 521858 185945 521892
rect 185979 521858 186037 521892
rect 186071 521858 186077 521892
rect 182567 521849 186077 521858
rect 186129 521892 186141 521901
rect 186129 521849 186141 521858
rect 186193 521849 186205 521901
rect 186257 521849 186269 521901
rect 186321 521892 186333 521901
rect 186385 521892 187480 521901
rect 186385 521858 186405 521892
rect 186439 521858 186497 521892
rect 186531 521858 186589 521892
rect 186623 521858 186681 521892
rect 186715 521858 186773 521892
rect 186807 521858 186865 521892
rect 186899 521858 186957 521892
rect 186991 521858 187049 521892
rect 187083 521858 187141 521892
rect 187175 521858 187233 521892
rect 187267 521858 187325 521892
rect 187359 521858 187417 521892
rect 187451 521858 187480 521892
rect 186321 521849 186333 521858
rect 186385 521849 187480 521858
rect 172208 521827 187480 521849
rect 172208 521357 187480 521379
rect 172208 521348 173963 521357
rect 174015 521348 174027 521357
rect 174079 521348 174091 521357
rect 172208 521314 172237 521348
rect 172271 521314 172329 521348
rect 172363 521314 172421 521348
rect 172455 521314 172513 521348
rect 172547 521314 172605 521348
rect 172639 521314 172697 521348
rect 172731 521314 172789 521348
rect 172823 521314 172881 521348
rect 172915 521314 172973 521348
rect 173007 521314 173065 521348
rect 173099 521314 173157 521348
rect 173191 521314 173249 521348
rect 173283 521314 173341 521348
rect 173375 521314 173433 521348
rect 173467 521314 173525 521348
rect 173559 521314 173617 521348
rect 173651 521314 173709 521348
rect 173743 521314 173801 521348
rect 173835 521314 173893 521348
rect 173927 521314 173963 521348
rect 174019 521314 174027 521348
rect 172208 521305 173963 521314
rect 174015 521305 174027 521314
rect 174079 521305 174091 521314
rect 174143 521305 174155 521357
rect 174207 521305 174219 521357
rect 174271 521348 177781 521357
rect 174295 521314 174353 521348
rect 174387 521314 174445 521348
rect 174479 521314 174537 521348
rect 174571 521314 174629 521348
rect 174663 521314 174721 521348
rect 174755 521314 174813 521348
rect 174847 521314 174905 521348
rect 174939 521314 174997 521348
rect 175031 521314 175089 521348
rect 175123 521314 175181 521348
rect 175215 521314 175273 521348
rect 175307 521314 175365 521348
rect 175399 521314 175457 521348
rect 175491 521314 175549 521348
rect 175583 521314 175641 521348
rect 175675 521314 175733 521348
rect 175767 521314 175825 521348
rect 175859 521314 175917 521348
rect 175951 521314 176009 521348
rect 176043 521314 176101 521348
rect 176135 521314 176193 521348
rect 176227 521314 176285 521348
rect 176319 521314 176377 521348
rect 176411 521314 176469 521348
rect 176503 521314 176561 521348
rect 176595 521314 176653 521348
rect 176687 521314 176745 521348
rect 176779 521314 176837 521348
rect 176871 521314 176929 521348
rect 176963 521314 177021 521348
rect 177055 521314 177113 521348
rect 177147 521314 177205 521348
rect 177239 521314 177297 521348
rect 177331 521314 177389 521348
rect 177423 521314 177481 521348
rect 177515 521314 177573 521348
rect 177607 521314 177665 521348
rect 177699 521314 177757 521348
rect 174271 521305 177781 521314
rect 177833 521305 177845 521357
rect 177897 521305 177909 521357
rect 177961 521348 177973 521357
rect 178025 521348 178037 521357
rect 178089 521348 181599 521357
rect 181651 521348 181663 521357
rect 181715 521348 181727 521357
rect 178025 521314 178033 521348
rect 178089 521314 178125 521348
rect 178159 521314 178217 521348
rect 178251 521314 178309 521348
rect 178343 521314 178401 521348
rect 178435 521314 178493 521348
rect 178527 521314 178585 521348
rect 178619 521314 178677 521348
rect 178711 521314 178769 521348
rect 178803 521314 178861 521348
rect 178895 521314 178953 521348
rect 178987 521314 179045 521348
rect 179079 521314 179137 521348
rect 179171 521314 179229 521348
rect 179263 521314 179321 521348
rect 179355 521314 179413 521348
rect 179447 521314 179505 521348
rect 179539 521314 179597 521348
rect 179631 521314 179689 521348
rect 179723 521314 179781 521348
rect 179815 521314 179873 521348
rect 179907 521314 179965 521348
rect 179999 521314 180057 521348
rect 180091 521314 180149 521348
rect 180183 521314 180241 521348
rect 180275 521314 180333 521348
rect 180367 521314 180425 521348
rect 180459 521314 180517 521348
rect 180551 521314 180609 521348
rect 180643 521314 180701 521348
rect 180735 521314 180793 521348
rect 180827 521314 180885 521348
rect 180919 521314 180977 521348
rect 181011 521314 181069 521348
rect 181103 521314 181161 521348
rect 181195 521314 181253 521348
rect 181287 521314 181345 521348
rect 181379 521314 181437 521348
rect 181471 521314 181529 521348
rect 181563 521314 181599 521348
rect 181655 521314 181663 521348
rect 177961 521305 177973 521314
rect 178025 521305 178037 521314
rect 178089 521305 181599 521314
rect 181651 521305 181663 521314
rect 181715 521305 181727 521314
rect 181779 521305 181791 521357
rect 181843 521305 181855 521357
rect 181907 521348 185417 521357
rect 181931 521314 181989 521348
rect 182023 521314 182081 521348
rect 182115 521314 182173 521348
rect 182207 521314 182265 521348
rect 182299 521314 182357 521348
rect 182391 521314 182449 521348
rect 182483 521314 182541 521348
rect 182575 521314 182633 521348
rect 182667 521314 182725 521348
rect 182759 521314 182817 521348
rect 182851 521314 182909 521348
rect 182943 521314 183001 521348
rect 183035 521314 183093 521348
rect 183127 521314 183185 521348
rect 183219 521314 183277 521348
rect 183311 521314 183369 521348
rect 183403 521314 183461 521348
rect 183495 521314 183553 521348
rect 183587 521314 183645 521348
rect 183679 521314 183737 521348
rect 183771 521314 183829 521348
rect 183863 521314 183921 521348
rect 183955 521314 184013 521348
rect 184047 521314 184105 521348
rect 184139 521314 184197 521348
rect 184231 521314 184289 521348
rect 184323 521314 184381 521348
rect 184415 521314 184473 521348
rect 184507 521314 184565 521348
rect 184599 521314 184657 521348
rect 184691 521314 184749 521348
rect 184783 521314 184841 521348
rect 184875 521314 184933 521348
rect 184967 521314 185025 521348
rect 185059 521314 185117 521348
rect 185151 521314 185209 521348
rect 185243 521314 185301 521348
rect 185335 521314 185393 521348
rect 181907 521305 185417 521314
rect 185469 521305 185481 521357
rect 185533 521305 185545 521357
rect 185597 521348 185609 521357
rect 185661 521348 185673 521357
rect 185725 521348 187480 521357
rect 185661 521314 185669 521348
rect 185725 521314 185761 521348
rect 185795 521314 185853 521348
rect 185887 521314 185945 521348
rect 185979 521314 186037 521348
rect 186071 521314 186129 521348
rect 186163 521314 186221 521348
rect 186255 521314 186313 521348
rect 186347 521314 186405 521348
rect 186439 521314 186497 521348
rect 186531 521314 186589 521348
rect 186623 521314 186681 521348
rect 186715 521314 186773 521348
rect 186807 521314 186865 521348
rect 186899 521314 186957 521348
rect 186991 521314 187049 521348
rect 187083 521314 187141 521348
rect 187175 521314 187233 521348
rect 187267 521314 187325 521348
rect 187359 521314 187417 521348
rect 187451 521314 187480 521348
rect 185597 521305 185609 521314
rect 185661 521305 185673 521314
rect 185725 521305 187480 521314
rect 172208 521283 187480 521305
rect 193000 521000 195000 522910
rect 172208 520813 187480 520835
rect 172208 520804 174623 520813
rect 172208 520770 172237 520804
rect 172271 520770 172329 520804
rect 172363 520770 172421 520804
rect 172455 520770 172513 520804
rect 172547 520770 172605 520804
rect 172639 520770 172697 520804
rect 172731 520770 172789 520804
rect 172823 520770 172881 520804
rect 172915 520770 172973 520804
rect 173007 520770 173065 520804
rect 173099 520770 173157 520804
rect 173191 520770 173249 520804
rect 173283 520770 173341 520804
rect 173375 520770 173433 520804
rect 173467 520770 173525 520804
rect 173559 520770 173617 520804
rect 173651 520770 173709 520804
rect 173743 520770 173801 520804
rect 173835 520770 173893 520804
rect 173927 520770 173985 520804
rect 174019 520770 174077 520804
rect 174111 520770 174169 520804
rect 174203 520770 174261 520804
rect 174295 520770 174353 520804
rect 174387 520770 174445 520804
rect 174479 520770 174537 520804
rect 174571 520770 174623 520804
rect 172208 520761 174623 520770
rect 174675 520761 174687 520813
rect 174739 520804 174751 520813
rect 174803 520804 174815 520813
rect 174803 520770 174813 520804
rect 174739 520761 174751 520770
rect 174803 520761 174815 520770
rect 174867 520761 174879 520813
rect 174931 520804 178441 520813
rect 174939 520770 174997 520804
rect 175031 520770 175089 520804
rect 175123 520770 175181 520804
rect 175215 520770 175273 520804
rect 175307 520770 175365 520804
rect 175399 520770 175457 520804
rect 175491 520770 175549 520804
rect 175583 520770 175641 520804
rect 175675 520770 175733 520804
rect 175767 520770 175825 520804
rect 175859 520770 175917 520804
rect 175951 520770 176009 520804
rect 176043 520770 176101 520804
rect 176135 520770 176193 520804
rect 176227 520770 176285 520804
rect 176319 520770 176377 520804
rect 176411 520770 176469 520804
rect 176503 520770 176561 520804
rect 176595 520770 176653 520804
rect 176687 520770 176745 520804
rect 176779 520770 176837 520804
rect 176871 520770 176929 520804
rect 176963 520770 177021 520804
rect 177055 520770 177113 520804
rect 177147 520770 177205 520804
rect 177239 520770 177297 520804
rect 177331 520770 177389 520804
rect 177423 520770 177481 520804
rect 177515 520770 177573 520804
rect 177607 520770 177665 520804
rect 177699 520770 177757 520804
rect 177791 520770 177849 520804
rect 177883 520770 177941 520804
rect 177975 520770 178033 520804
rect 178067 520770 178125 520804
rect 178159 520770 178217 520804
rect 178251 520770 178309 520804
rect 178343 520770 178401 520804
rect 178435 520770 178441 520804
rect 174931 520761 178441 520770
rect 178493 520804 178505 520813
rect 178493 520761 178505 520770
rect 178557 520761 178569 520813
rect 178621 520761 178633 520813
rect 178685 520804 178697 520813
rect 178749 520804 182259 520813
rect 178749 520770 178769 520804
rect 178803 520770 178861 520804
rect 178895 520770 178953 520804
rect 178987 520770 179045 520804
rect 179079 520770 179137 520804
rect 179171 520770 179229 520804
rect 179263 520770 179321 520804
rect 179355 520770 179413 520804
rect 179447 520770 179505 520804
rect 179539 520770 179597 520804
rect 179631 520770 179689 520804
rect 179723 520770 179781 520804
rect 179815 520770 179873 520804
rect 179907 520770 179965 520804
rect 179999 520770 180057 520804
rect 180091 520770 180149 520804
rect 180183 520770 180241 520804
rect 180275 520770 180333 520804
rect 180367 520770 180425 520804
rect 180459 520770 180517 520804
rect 180551 520770 180609 520804
rect 180643 520770 180701 520804
rect 180735 520770 180793 520804
rect 180827 520770 180885 520804
rect 180919 520770 180977 520804
rect 181011 520770 181069 520804
rect 181103 520770 181161 520804
rect 181195 520770 181253 520804
rect 181287 520770 181345 520804
rect 181379 520770 181437 520804
rect 181471 520770 181529 520804
rect 181563 520770 181621 520804
rect 181655 520770 181713 520804
rect 181747 520770 181805 520804
rect 181839 520770 181897 520804
rect 181931 520770 181989 520804
rect 182023 520770 182081 520804
rect 182115 520770 182173 520804
rect 182207 520770 182259 520804
rect 178685 520761 178697 520770
rect 178749 520761 182259 520770
rect 182311 520761 182323 520813
rect 182375 520804 182387 520813
rect 182439 520804 182451 520813
rect 182439 520770 182449 520804
rect 182375 520761 182387 520770
rect 182439 520761 182451 520770
rect 182503 520761 182515 520813
rect 182567 520804 186077 520813
rect 182575 520770 182633 520804
rect 182667 520770 182725 520804
rect 182759 520770 182817 520804
rect 182851 520770 182909 520804
rect 182943 520770 183001 520804
rect 183035 520770 183093 520804
rect 183127 520770 183185 520804
rect 183219 520770 183277 520804
rect 183311 520770 183369 520804
rect 183403 520770 183461 520804
rect 183495 520770 183553 520804
rect 183587 520770 183645 520804
rect 183679 520770 183737 520804
rect 183771 520770 183829 520804
rect 183863 520770 183921 520804
rect 183955 520770 184013 520804
rect 184047 520770 184105 520804
rect 184139 520770 184197 520804
rect 184231 520770 184289 520804
rect 184323 520770 184381 520804
rect 184415 520770 184473 520804
rect 184507 520770 184565 520804
rect 184599 520770 184657 520804
rect 184691 520770 184749 520804
rect 184783 520770 184841 520804
rect 184875 520770 184933 520804
rect 184967 520770 185025 520804
rect 185059 520770 185117 520804
rect 185151 520770 185209 520804
rect 185243 520770 185301 520804
rect 185335 520770 185393 520804
rect 185427 520770 185485 520804
rect 185519 520770 185577 520804
rect 185611 520770 185669 520804
rect 185703 520770 185761 520804
rect 185795 520770 185853 520804
rect 185887 520770 185945 520804
rect 185979 520770 186037 520804
rect 186071 520770 186077 520804
rect 182567 520761 186077 520770
rect 186129 520804 186141 520813
rect 186129 520761 186141 520770
rect 186193 520761 186205 520813
rect 186257 520761 186269 520813
rect 186321 520804 186333 520813
rect 186385 520804 187480 520813
rect 186385 520770 186405 520804
rect 186439 520770 186497 520804
rect 186531 520770 186589 520804
rect 186623 520770 186681 520804
rect 186715 520770 186773 520804
rect 186807 520770 186865 520804
rect 186899 520770 186957 520804
rect 186991 520770 187049 520804
rect 187083 520770 187141 520804
rect 187175 520770 187233 520804
rect 187267 520770 187325 520804
rect 187359 520770 187417 520804
rect 187451 520770 187480 520804
rect 186321 520761 186333 520770
rect 186385 520761 187480 520770
rect 172208 520739 187480 520761
rect 172208 520269 187480 520291
rect 172208 520260 173963 520269
rect 174015 520260 174027 520269
rect 174079 520260 174091 520269
rect 172208 520226 172237 520260
rect 172271 520226 172329 520260
rect 172363 520226 172421 520260
rect 172455 520226 172513 520260
rect 172547 520226 172605 520260
rect 172639 520226 172697 520260
rect 172731 520226 172789 520260
rect 172823 520226 172881 520260
rect 172915 520226 172973 520260
rect 173007 520226 173065 520260
rect 173099 520226 173157 520260
rect 173191 520226 173249 520260
rect 173283 520226 173341 520260
rect 173375 520226 173433 520260
rect 173467 520226 173525 520260
rect 173559 520226 173617 520260
rect 173651 520226 173709 520260
rect 173743 520226 173801 520260
rect 173835 520226 173893 520260
rect 173927 520226 173963 520260
rect 174019 520226 174027 520260
rect 172208 520217 173963 520226
rect 174015 520217 174027 520226
rect 174079 520217 174091 520226
rect 174143 520217 174155 520269
rect 174207 520217 174219 520269
rect 174271 520260 177781 520269
rect 174295 520226 174353 520260
rect 174387 520226 174445 520260
rect 174479 520226 174537 520260
rect 174571 520226 174629 520260
rect 174663 520226 174721 520260
rect 174755 520226 174813 520260
rect 174847 520226 174905 520260
rect 174939 520226 174997 520260
rect 175031 520226 175089 520260
rect 175123 520226 175181 520260
rect 175215 520226 175273 520260
rect 175307 520226 175365 520260
rect 175399 520226 175457 520260
rect 175491 520226 175549 520260
rect 175583 520226 175641 520260
rect 175675 520226 175733 520260
rect 175767 520226 175825 520260
rect 175859 520226 175917 520260
rect 175951 520226 176009 520260
rect 176043 520226 176101 520260
rect 176135 520226 176193 520260
rect 176227 520226 176285 520260
rect 176319 520226 176377 520260
rect 176411 520226 176469 520260
rect 176503 520226 176561 520260
rect 176595 520226 176653 520260
rect 176687 520226 176745 520260
rect 176779 520226 176837 520260
rect 176871 520226 176929 520260
rect 176963 520226 177021 520260
rect 177055 520226 177113 520260
rect 177147 520226 177205 520260
rect 177239 520226 177297 520260
rect 177331 520226 177389 520260
rect 177423 520226 177481 520260
rect 177515 520226 177573 520260
rect 177607 520226 177665 520260
rect 177699 520226 177757 520260
rect 174271 520217 177781 520226
rect 177833 520217 177845 520269
rect 177897 520217 177909 520269
rect 177961 520260 177973 520269
rect 178025 520260 178037 520269
rect 178089 520260 181599 520269
rect 181651 520260 181663 520269
rect 181715 520260 181727 520269
rect 178025 520226 178033 520260
rect 178089 520226 178125 520260
rect 178159 520226 178217 520260
rect 178251 520226 178309 520260
rect 178343 520226 178401 520260
rect 178435 520226 178493 520260
rect 178527 520226 178585 520260
rect 178619 520226 178677 520260
rect 178711 520226 178769 520260
rect 178803 520226 178861 520260
rect 178895 520226 178953 520260
rect 178987 520226 179045 520260
rect 179079 520226 179137 520260
rect 179171 520226 179229 520260
rect 179263 520226 179321 520260
rect 179355 520226 179413 520260
rect 179447 520226 179505 520260
rect 179539 520226 179597 520260
rect 179631 520226 179689 520260
rect 179723 520226 179781 520260
rect 179815 520226 179873 520260
rect 179907 520226 179965 520260
rect 179999 520226 180057 520260
rect 180091 520226 180149 520260
rect 180183 520226 180241 520260
rect 180275 520226 180333 520260
rect 180367 520226 180425 520260
rect 180459 520226 180517 520260
rect 180551 520226 180609 520260
rect 180643 520226 180701 520260
rect 180735 520226 180793 520260
rect 180827 520226 180885 520260
rect 180919 520226 180977 520260
rect 181011 520226 181069 520260
rect 181103 520226 181161 520260
rect 181195 520226 181253 520260
rect 181287 520226 181345 520260
rect 181379 520226 181437 520260
rect 181471 520226 181529 520260
rect 181563 520226 181599 520260
rect 181655 520226 181663 520260
rect 177961 520217 177973 520226
rect 178025 520217 178037 520226
rect 178089 520217 181599 520226
rect 181651 520217 181663 520226
rect 181715 520217 181727 520226
rect 181779 520217 181791 520269
rect 181843 520217 181855 520269
rect 181907 520260 185417 520269
rect 181931 520226 181989 520260
rect 182023 520226 182081 520260
rect 182115 520226 182173 520260
rect 182207 520226 182265 520260
rect 182299 520226 182357 520260
rect 182391 520226 182449 520260
rect 182483 520226 182541 520260
rect 182575 520226 182633 520260
rect 182667 520226 182725 520260
rect 182759 520226 182817 520260
rect 182851 520226 182909 520260
rect 182943 520226 183001 520260
rect 183035 520226 183093 520260
rect 183127 520226 183185 520260
rect 183219 520226 183277 520260
rect 183311 520226 183369 520260
rect 183403 520226 183461 520260
rect 183495 520226 183553 520260
rect 183587 520226 183645 520260
rect 183679 520226 183737 520260
rect 183771 520226 183829 520260
rect 183863 520226 183921 520260
rect 183955 520226 184013 520260
rect 184047 520226 184105 520260
rect 184139 520226 184197 520260
rect 184231 520226 184289 520260
rect 184323 520226 184381 520260
rect 184415 520226 184473 520260
rect 184507 520226 184565 520260
rect 184599 520226 184657 520260
rect 184691 520226 184749 520260
rect 184783 520226 184841 520260
rect 184875 520226 184933 520260
rect 184967 520226 185025 520260
rect 185059 520226 185117 520260
rect 185151 520226 185209 520260
rect 185243 520226 185301 520260
rect 185335 520226 185393 520260
rect 181907 520217 185417 520226
rect 185469 520217 185481 520269
rect 185533 520217 185545 520269
rect 185597 520260 185609 520269
rect 185661 520260 185673 520269
rect 185725 520260 187480 520269
rect 185661 520226 185669 520260
rect 185725 520226 185761 520260
rect 185795 520226 185853 520260
rect 185887 520226 185945 520260
rect 185979 520226 186037 520260
rect 186071 520226 186129 520260
rect 186163 520226 186221 520260
rect 186255 520226 186313 520260
rect 186347 520226 186405 520260
rect 186439 520226 186497 520260
rect 186531 520226 186589 520260
rect 186623 520226 186681 520260
rect 186715 520226 186773 520260
rect 186807 520226 186865 520260
rect 186899 520226 186957 520260
rect 186991 520226 187049 520260
rect 187083 520226 187141 520260
rect 187175 520226 187233 520260
rect 187267 520226 187325 520260
rect 187359 520226 187417 520260
rect 187451 520226 187480 520260
rect 185597 520217 185609 520226
rect 185661 520217 185673 520226
rect 185725 520217 187480 520226
rect 172208 520195 187480 520217
rect 172208 519725 187480 519747
rect 172208 519716 174623 519725
rect 172208 519682 172237 519716
rect 172271 519682 172329 519716
rect 172363 519682 172421 519716
rect 172455 519682 172513 519716
rect 172547 519682 172605 519716
rect 172639 519682 172697 519716
rect 172731 519682 172789 519716
rect 172823 519682 172881 519716
rect 172915 519682 172973 519716
rect 173007 519682 173065 519716
rect 173099 519682 173157 519716
rect 173191 519682 173249 519716
rect 173283 519682 173341 519716
rect 173375 519682 173433 519716
rect 173467 519682 173525 519716
rect 173559 519682 173617 519716
rect 173651 519682 173709 519716
rect 173743 519682 173801 519716
rect 173835 519682 173893 519716
rect 173927 519682 173985 519716
rect 174019 519682 174077 519716
rect 174111 519682 174169 519716
rect 174203 519682 174261 519716
rect 174295 519682 174353 519716
rect 174387 519682 174445 519716
rect 174479 519682 174537 519716
rect 174571 519682 174623 519716
rect 172208 519673 174623 519682
rect 174675 519673 174687 519725
rect 174739 519716 174751 519725
rect 174803 519716 174815 519725
rect 174803 519682 174813 519716
rect 174739 519673 174751 519682
rect 174803 519673 174815 519682
rect 174867 519673 174879 519725
rect 174931 519716 178441 519725
rect 174939 519682 174997 519716
rect 175031 519682 175089 519716
rect 175123 519682 175181 519716
rect 175215 519682 175273 519716
rect 175307 519682 175365 519716
rect 175399 519682 175457 519716
rect 175491 519682 175549 519716
rect 175583 519682 175641 519716
rect 175675 519682 175733 519716
rect 175767 519682 175825 519716
rect 175859 519682 175917 519716
rect 175951 519682 176009 519716
rect 176043 519682 176101 519716
rect 176135 519682 176193 519716
rect 176227 519682 176285 519716
rect 176319 519682 176377 519716
rect 176411 519682 176469 519716
rect 176503 519682 176561 519716
rect 176595 519682 176653 519716
rect 176687 519682 176745 519716
rect 176779 519682 176837 519716
rect 176871 519682 176929 519716
rect 176963 519682 177021 519716
rect 177055 519682 177113 519716
rect 177147 519682 177205 519716
rect 177239 519682 177297 519716
rect 177331 519682 177389 519716
rect 177423 519682 177481 519716
rect 177515 519682 177573 519716
rect 177607 519682 177665 519716
rect 177699 519682 177757 519716
rect 177791 519682 177849 519716
rect 177883 519682 177941 519716
rect 177975 519682 178033 519716
rect 178067 519682 178125 519716
rect 178159 519682 178217 519716
rect 178251 519682 178309 519716
rect 178343 519682 178401 519716
rect 178435 519682 178441 519716
rect 174931 519673 178441 519682
rect 178493 519716 178505 519725
rect 178493 519673 178505 519682
rect 178557 519673 178569 519725
rect 178621 519673 178633 519725
rect 178685 519716 178697 519725
rect 178749 519716 182259 519725
rect 178749 519682 178769 519716
rect 178803 519682 178861 519716
rect 178895 519682 178953 519716
rect 178987 519682 179045 519716
rect 179079 519682 179137 519716
rect 179171 519682 179229 519716
rect 179263 519682 179321 519716
rect 179355 519682 179413 519716
rect 179447 519682 179505 519716
rect 179539 519682 179597 519716
rect 179631 519682 179689 519716
rect 179723 519682 179781 519716
rect 179815 519682 179873 519716
rect 179907 519682 179965 519716
rect 179999 519682 180057 519716
rect 180091 519682 180149 519716
rect 180183 519682 180241 519716
rect 180275 519682 180333 519716
rect 180367 519682 180425 519716
rect 180459 519682 180517 519716
rect 180551 519682 180609 519716
rect 180643 519682 180701 519716
rect 180735 519682 180793 519716
rect 180827 519682 180885 519716
rect 180919 519682 180977 519716
rect 181011 519682 181069 519716
rect 181103 519682 181161 519716
rect 181195 519682 181253 519716
rect 181287 519682 181345 519716
rect 181379 519682 181437 519716
rect 181471 519682 181529 519716
rect 181563 519682 181621 519716
rect 181655 519682 181713 519716
rect 181747 519682 181805 519716
rect 181839 519682 181897 519716
rect 181931 519682 181989 519716
rect 182023 519682 182081 519716
rect 182115 519682 182173 519716
rect 182207 519682 182259 519716
rect 178685 519673 178697 519682
rect 178749 519673 182259 519682
rect 182311 519673 182323 519725
rect 182375 519716 182387 519725
rect 182439 519716 182451 519725
rect 182439 519682 182449 519716
rect 182375 519673 182387 519682
rect 182439 519673 182451 519682
rect 182503 519673 182515 519725
rect 182567 519716 186077 519725
rect 182575 519682 182633 519716
rect 182667 519682 182725 519716
rect 182759 519682 182817 519716
rect 182851 519682 182909 519716
rect 182943 519682 183001 519716
rect 183035 519682 183093 519716
rect 183127 519682 183185 519716
rect 183219 519682 183277 519716
rect 183311 519682 183369 519716
rect 183403 519682 183461 519716
rect 183495 519682 183553 519716
rect 183587 519682 183645 519716
rect 183679 519682 183737 519716
rect 183771 519682 183829 519716
rect 183863 519682 183921 519716
rect 183955 519682 184013 519716
rect 184047 519682 184105 519716
rect 184139 519682 184197 519716
rect 184231 519682 184289 519716
rect 184323 519682 184381 519716
rect 184415 519682 184473 519716
rect 184507 519682 184565 519716
rect 184599 519682 184657 519716
rect 184691 519682 184749 519716
rect 184783 519682 184841 519716
rect 184875 519682 184933 519716
rect 184967 519682 185025 519716
rect 185059 519682 185117 519716
rect 185151 519682 185209 519716
rect 185243 519682 185301 519716
rect 185335 519682 185393 519716
rect 185427 519682 185485 519716
rect 185519 519682 185577 519716
rect 185611 519682 185669 519716
rect 185703 519682 185761 519716
rect 185795 519682 185853 519716
rect 185887 519682 185945 519716
rect 185979 519682 186037 519716
rect 186071 519682 186077 519716
rect 182567 519673 186077 519682
rect 186129 519716 186141 519725
rect 186129 519673 186141 519682
rect 186193 519673 186205 519725
rect 186257 519673 186269 519725
rect 186321 519716 186333 519725
rect 186385 519716 187480 519725
rect 186385 519682 186405 519716
rect 186439 519682 186497 519716
rect 186531 519682 186589 519716
rect 186623 519682 186681 519716
rect 186715 519682 186773 519716
rect 186807 519682 186865 519716
rect 186899 519682 186957 519716
rect 186991 519682 187049 519716
rect 187083 519682 187141 519716
rect 187175 519682 187233 519716
rect 187267 519682 187325 519716
rect 187359 519682 187417 519716
rect 187451 519682 187480 519716
rect 186321 519673 186333 519682
rect 186385 519673 187480 519682
rect 172208 519651 187480 519673
rect 172208 519181 187480 519203
rect 172208 519172 173963 519181
rect 174015 519172 174027 519181
rect 174079 519172 174091 519181
rect 172208 519138 172237 519172
rect 172271 519138 172329 519172
rect 172363 519138 172421 519172
rect 172455 519138 172513 519172
rect 172547 519138 172605 519172
rect 172639 519138 172697 519172
rect 172731 519138 172789 519172
rect 172823 519138 172881 519172
rect 172915 519138 172973 519172
rect 173007 519138 173065 519172
rect 173099 519138 173157 519172
rect 173191 519138 173249 519172
rect 173283 519138 173341 519172
rect 173375 519138 173433 519172
rect 173467 519138 173525 519172
rect 173559 519138 173617 519172
rect 173651 519138 173709 519172
rect 173743 519138 173801 519172
rect 173835 519138 173893 519172
rect 173927 519138 173963 519172
rect 174019 519138 174027 519172
rect 172208 519129 173963 519138
rect 174015 519129 174027 519138
rect 174079 519129 174091 519138
rect 174143 519129 174155 519181
rect 174207 519129 174219 519181
rect 174271 519172 177781 519181
rect 174295 519138 174353 519172
rect 174387 519138 174445 519172
rect 174479 519138 174537 519172
rect 174571 519138 174629 519172
rect 174663 519138 174721 519172
rect 174755 519138 174813 519172
rect 174847 519138 174905 519172
rect 174939 519138 174997 519172
rect 175031 519138 175089 519172
rect 175123 519138 175181 519172
rect 175215 519138 175273 519172
rect 175307 519138 175365 519172
rect 175399 519138 175457 519172
rect 175491 519138 175549 519172
rect 175583 519138 175641 519172
rect 175675 519138 175733 519172
rect 175767 519138 175825 519172
rect 175859 519138 175917 519172
rect 175951 519138 176009 519172
rect 176043 519138 176101 519172
rect 176135 519138 176193 519172
rect 176227 519138 176285 519172
rect 176319 519138 176377 519172
rect 176411 519138 176469 519172
rect 176503 519138 176561 519172
rect 176595 519138 176653 519172
rect 176687 519138 176745 519172
rect 176779 519138 176837 519172
rect 176871 519138 176929 519172
rect 176963 519138 177021 519172
rect 177055 519138 177113 519172
rect 177147 519138 177205 519172
rect 177239 519138 177297 519172
rect 177331 519138 177389 519172
rect 177423 519138 177481 519172
rect 177515 519138 177573 519172
rect 177607 519138 177665 519172
rect 177699 519138 177757 519172
rect 174271 519129 177781 519138
rect 177833 519129 177845 519181
rect 177897 519129 177909 519181
rect 177961 519172 177973 519181
rect 178025 519172 178037 519181
rect 178089 519172 181599 519181
rect 181651 519172 181663 519181
rect 181715 519172 181727 519181
rect 178025 519138 178033 519172
rect 178089 519138 178125 519172
rect 178159 519138 178217 519172
rect 178251 519138 178309 519172
rect 178343 519138 178401 519172
rect 178435 519138 178493 519172
rect 178527 519138 178585 519172
rect 178619 519138 178677 519172
rect 178711 519138 178769 519172
rect 178803 519138 178861 519172
rect 178895 519138 178953 519172
rect 178987 519138 179045 519172
rect 179079 519138 179137 519172
rect 179171 519138 179229 519172
rect 179263 519138 179321 519172
rect 179355 519138 179413 519172
rect 179447 519138 179505 519172
rect 179539 519138 179597 519172
rect 179631 519138 179689 519172
rect 179723 519138 179781 519172
rect 179815 519138 179873 519172
rect 179907 519138 179965 519172
rect 179999 519138 180057 519172
rect 180091 519138 180149 519172
rect 180183 519138 180241 519172
rect 180275 519138 180333 519172
rect 180367 519138 180425 519172
rect 180459 519138 180517 519172
rect 180551 519138 180609 519172
rect 180643 519138 180701 519172
rect 180735 519138 180793 519172
rect 180827 519138 180885 519172
rect 180919 519138 180977 519172
rect 181011 519138 181069 519172
rect 181103 519138 181161 519172
rect 181195 519138 181253 519172
rect 181287 519138 181345 519172
rect 181379 519138 181437 519172
rect 181471 519138 181529 519172
rect 181563 519138 181599 519172
rect 181655 519138 181663 519172
rect 177961 519129 177973 519138
rect 178025 519129 178037 519138
rect 178089 519129 181599 519138
rect 181651 519129 181663 519138
rect 181715 519129 181727 519138
rect 181779 519129 181791 519181
rect 181843 519129 181855 519181
rect 181907 519172 185417 519181
rect 181931 519138 181989 519172
rect 182023 519138 182081 519172
rect 182115 519138 182173 519172
rect 182207 519138 182265 519172
rect 182299 519138 182357 519172
rect 182391 519138 182449 519172
rect 182483 519138 182541 519172
rect 182575 519138 182633 519172
rect 182667 519138 182725 519172
rect 182759 519138 182817 519172
rect 182851 519138 182909 519172
rect 182943 519138 183001 519172
rect 183035 519138 183093 519172
rect 183127 519138 183185 519172
rect 183219 519138 183277 519172
rect 183311 519138 183369 519172
rect 183403 519138 183461 519172
rect 183495 519138 183553 519172
rect 183587 519138 183645 519172
rect 183679 519138 183737 519172
rect 183771 519138 183829 519172
rect 183863 519138 183921 519172
rect 183955 519138 184013 519172
rect 184047 519138 184105 519172
rect 184139 519138 184197 519172
rect 184231 519138 184289 519172
rect 184323 519138 184381 519172
rect 184415 519138 184473 519172
rect 184507 519138 184565 519172
rect 184599 519138 184657 519172
rect 184691 519138 184749 519172
rect 184783 519138 184841 519172
rect 184875 519138 184933 519172
rect 184967 519138 185025 519172
rect 185059 519138 185117 519172
rect 185151 519138 185209 519172
rect 185243 519138 185301 519172
rect 185335 519138 185393 519172
rect 181907 519129 185417 519138
rect 185469 519129 185481 519181
rect 185533 519129 185545 519181
rect 185597 519172 185609 519181
rect 185661 519172 185673 519181
rect 185725 519172 187480 519181
rect 185661 519138 185669 519172
rect 185725 519138 185761 519172
rect 185795 519138 185853 519172
rect 185887 519138 185945 519172
rect 185979 519138 186037 519172
rect 186071 519138 186129 519172
rect 186163 519138 186221 519172
rect 186255 519138 186313 519172
rect 186347 519138 186405 519172
rect 186439 519138 186497 519172
rect 186531 519138 186589 519172
rect 186623 519138 186681 519172
rect 186715 519138 186773 519172
rect 186807 519138 186865 519172
rect 186899 519138 186957 519172
rect 186991 519138 187049 519172
rect 187083 519138 187141 519172
rect 187175 519138 187233 519172
rect 187267 519138 187325 519172
rect 187359 519138 187417 519172
rect 187451 519138 187480 519172
rect 185597 519129 185609 519138
rect 185661 519129 185673 519138
rect 185725 519129 187480 519138
rect 172208 519107 187480 519129
rect 172208 518637 187480 518659
rect 172208 518628 174623 518637
rect 172208 518594 172237 518628
rect 172271 518594 172329 518628
rect 172363 518594 172421 518628
rect 172455 518594 172513 518628
rect 172547 518594 172605 518628
rect 172639 518594 172697 518628
rect 172731 518594 172789 518628
rect 172823 518594 172881 518628
rect 172915 518594 172973 518628
rect 173007 518594 173065 518628
rect 173099 518594 173157 518628
rect 173191 518594 173249 518628
rect 173283 518594 173341 518628
rect 173375 518594 173433 518628
rect 173467 518594 173525 518628
rect 173559 518594 173617 518628
rect 173651 518594 173709 518628
rect 173743 518594 173801 518628
rect 173835 518594 173893 518628
rect 173927 518594 173985 518628
rect 174019 518594 174077 518628
rect 174111 518594 174169 518628
rect 174203 518594 174261 518628
rect 174295 518594 174353 518628
rect 174387 518594 174445 518628
rect 174479 518594 174537 518628
rect 174571 518594 174623 518628
rect 172208 518585 174623 518594
rect 174675 518585 174687 518637
rect 174739 518628 174751 518637
rect 174803 518628 174815 518637
rect 174803 518594 174813 518628
rect 174739 518585 174751 518594
rect 174803 518585 174815 518594
rect 174867 518585 174879 518637
rect 174931 518628 178441 518637
rect 174939 518594 174997 518628
rect 175031 518594 175089 518628
rect 175123 518594 175181 518628
rect 175215 518594 175273 518628
rect 175307 518594 175365 518628
rect 175399 518594 175457 518628
rect 175491 518594 175549 518628
rect 175583 518594 175641 518628
rect 175675 518594 175733 518628
rect 175767 518594 175825 518628
rect 175859 518594 175917 518628
rect 175951 518594 176009 518628
rect 176043 518594 176101 518628
rect 176135 518594 176193 518628
rect 176227 518594 176285 518628
rect 176319 518594 176377 518628
rect 176411 518594 176469 518628
rect 176503 518594 176561 518628
rect 176595 518594 176653 518628
rect 176687 518594 176745 518628
rect 176779 518594 176837 518628
rect 176871 518594 176929 518628
rect 176963 518594 177021 518628
rect 177055 518594 177113 518628
rect 177147 518594 177205 518628
rect 177239 518594 177297 518628
rect 177331 518594 177389 518628
rect 177423 518594 177481 518628
rect 177515 518594 177573 518628
rect 177607 518594 177665 518628
rect 177699 518594 177757 518628
rect 177791 518594 177849 518628
rect 177883 518594 177941 518628
rect 177975 518594 178033 518628
rect 178067 518594 178125 518628
rect 178159 518594 178217 518628
rect 178251 518594 178309 518628
rect 178343 518594 178401 518628
rect 178435 518594 178441 518628
rect 174931 518585 178441 518594
rect 178493 518628 178505 518637
rect 178493 518585 178505 518594
rect 178557 518585 178569 518637
rect 178621 518585 178633 518637
rect 178685 518628 178697 518637
rect 178749 518628 182259 518637
rect 178749 518594 178769 518628
rect 178803 518594 178861 518628
rect 178895 518594 178953 518628
rect 178987 518594 179045 518628
rect 179079 518594 179137 518628
rect 179171 518594 179229 518628
rect 179263 518594 179321 518628
rect 179355 518594 179413 518628
rect 179447 518594 179505 518628
rect 179539 518594 179597 518628
rect 179631 518594 179689 518628
rect 179723 518594 179781 518628
rect 179815 518594 179873 518628
rect 179907 518594 179965 518628
rect 179999 518594 180057 518628
rect 180091 518594 180149 518628
rect 180183 518594 180241 518628
rect 180275 518594 180333 518628
rect 180367 518594 180425 518628
rect 180459 518594 180517 518628
rect 180551 518594 180609 518628
rect 180643 518594 180701 518628
rect 180735 518594 180793 518628
rect 180827 518594 180885 518628
rect 180919 518594 180977 518628
rect 181011 518594 181069 518628
rect 181103 518594 181161 518628
rect 181195 518594 181253 518628
rect 181287 518594 181345 518628
rect 181379 518594 181437 518628
rect 181471 518594 181529 518628
rect 181563 518594 181621 518628
rect 181655 518594 181713 518628
rect 181747 518594 181805 518628
rect 181839 518594 181897 518628
rect 181931 518594 181989 518628
rect 182023 518594 182081 518628
rect 182115 518594 182173 518628
rect 182207 518594 182259 518628
rect 178685 518585 178697 518594
rect 178749 518585 182259 518594
rect 182311 518585 182323 518637
rect 182375 518628 182387 518637
rect 182439 518628 182451 518637
rect 182439 518594 182449 518628
rect 182375 518585 182387 518594
rect 182439 518585 182451 518594
rect 182503 518585 182515 518637
rect 182567 518628 186077 518637
rect 182575 518594 182633 518628
rect 182667 518594 182725 518628
rect 182759 518594 182817 518628
rect 182851 518594 182909 518628
rect 182943 518594 183001 518628
rect 183035 518594 183093 518628
rect 183127 518594 183185 518628
rect 183219 518594 183277 518628
rect 183311 518594 183369 518628
rect 183403 518594 183461 518628
rect 183495 518594 183553 518628
rect 183587 518594 183645 518628
rect 183679 518594 183737 518628
rect 183771 518594 183829 518628
rect 183863 518594 183921 518628
rect 183955 518594 184013 518628
rect 184047 518594 184105 518628
rect 184139 518594 184197 518628
rect 184231 518594 184289 518628
rect 184323 518594 184381 518628
rect 184415 518594 184473 518628
rect 184507 518594 184565 518628
rect 184599 518594 184657 518628
rect 184691 518594 184749 518628
rect 184783 518594 184841 518628
rect 184875 518594 184933 518628
rect 184967 518594 185025 518628
rect 185059 518594 185117 518628
rect 185151 518594 185209 518628
rect 185243 518594 185301 518628
rect 185335 518594 185393 518628
rect 185427 518594 185485 518628
rect 185519 518594 185577 518628
rect 185611 518594 185669 518628
rect 185703 518594 185761 518628
rect 185795 518594 185853 518628
rect 185887 518594 185945 518628
rect 185979 518594 186037 518628
rect 186071 518594 186077 518628
rect 182567 518585 186077 518594
rect 186129 518628 186141 518637
rect 186129 518585 186141 518594
rect 186193 518585 186205 518637
rect 186257 518585 186269 518637
rect 186321 518628 186333 518637
rect 186385 518628 187480 518637
rect 186385 518594 186405 518628
rect 186439 518594 186497 518628
rect 186531 518594 186589 518628
rect 186623 518594 186681 518628
rect 186715 518594 186773 518628
rect 186807 518594 186865 518628
rect 186899 518594 186957 518628
rect 186991 518594 187049 518628
rect 187083 518594 187141 518628
rect 187175 518594 187233 518628
rect 187267 518594 187325 518628
rect 187359 518594 187417 518628
rect 187451 518594 187480 518628
rect 186321 518585 186333 518594
rect 186385 518585 187480 518594
rect 172208 518563 187480 518585
rect 172208 518093 187480 518115
rect 172208 518084 173963 518093
rect 174015 518084 174027 518093
rect 174079 518084 174091 518093
rect 172208 518050 172237 518084
rect 172271 518050 172329 518084
rect 172363 518050 172421 518084
rect 172455 518050 172513 518084
rect 172547 518050 172605 518084
rect 172639 518050 172697 518084
rect 172731 518050 172789 518084
rect 172823 518050 172881 518084
rect 172915 518050 172973 518084
rect 173007 518050 173065 518084
rect 173099 518050 173157 518084
rect 173191 518050 173249 518084
rect 173283 518050 173341 518084
rect 173375 518050 173433 518084
rect 173467 518050 173525 518084
rect 173559 518050 173617 518084
rect 173651 518050 173709 518084
rect 173743 518050 173801 518084
rect 173835 518050 173893 518084
rect 173927 518050 173963 518084
rect 174019 518050 174027 518084
rect 172208 518041 173963 518050
rect 174015 518041 174027 518050
rect 174079 518041 174091 518050
rect 174143 518041 174155 518093
rect 174207 518041 174219 518093
rect 174271 518084 177781 518093
rect 174295 518050 174353 518084
rect 174387 518050 174445 518084
rect 174479 518050 174537 518084
rect 174571 518050 174629 518084
rect 174663 518050 174721 518084
rect 174755 518050 174813 518084
rect 174847 518050 174905 518084
rect 174939 518050 174997 518084
rect 175031 518050 175089 518084
rect 175123 518050 175181 518084
rect 175215 518050 175273 518084
rect 175307 518050 175365 518084
rect 175399 518050 175457 518084
rect 175491 518050 175549 518084
rect 175583 518050 175641 518084
rect 175675 518050 175733 518084
rect 175767 518050 175825 518084
rect 175859 518050 175917 518084
rect 175951 518050 176009 518084
rect 176043 518050 176101 518084
rect 176135 518050 176193 518084
rect 176227 518050 176285 518084
rect 176319 518050 176377 518084
rect 176411 518050 176469 518084
rect 176503 518050 176561 518084
rect 176595 518050 176653 518084
rect 176687 518050 176745 518084
rect 176779 518050 176837 518084
rect 176871 518050 176929 518084
rect 176963 518050 177021 518084
rect 177055 518050 177113 518084
rect 177147 518050 177205 518084
rect 177239 518050 177297 518084
rect 177331 518050 177389 518084
rect 177423 518050 177481 518084
rect 177515 518050 177573 518084
rect 177607 518050 177665 518084
rect 177699 518050 177757 518084
rect 174271 518041 177781 518050
rect 177833 518041 177845 518093
rect 177897 518041 177909 518093
rect 177961 518084 177973 518093
rect 178025 518084 178037 518093
rect 178089 518084 181599 518093
rect 181651 518084 181663 518093
rect 181715 518084 181727 518093
rect 178025 518050 178033 518084
rect 178089 518050 178125 518084
rect 178159 518050 178217 518084
rect 178251 518050 178309 518084
rect 178343 518050 178401 518084
rect 178435 518050 178493 518084
rect 178527 518050 178585 518084
rect 178619 518050 178677 518084
rect 178711 518050 178769 518084
rect 178803 518050 178861 518084
rect 178895 518050 178953 518084
rect 178987 518050 179045 518084
rect 179079 518050 179137 518084
rect 179171 518050 179229 518084
rect 179263 518050 179321 518084
rect 179355 518050 179413 518084
rect 179447 518050 179505 518084
rect 179539 518050 179597 518084
rect 179631 518050 179689 518084
rect 179723 518050 179781 518084
rect 179815 518050 179873 518084
rect 179907 518050 179965 518084
rect 179999 518050 180057 518084
rect 180091 518050 180149 518084
rect 180183 518050 180241 518084
rect 180275 518050 180333 518084
rect 180367 518050 180425 518084
rect 180459 518050 180517 518084
rect 180551 518050 180609 518084
rect 180643 518050 180701 518084
rect 180735 518050 180793 518084
rect 180827 518050 180885 518084
rect 180919 518050 180977 518084
rect 181011 518050 181069 518084
rect 181103 518050 181161 518084
rect 181195 518050 181253 518084
rect 181287 518050 181345 518084
rect 181379 518050 181437 518084
rect 181471 518050 181529 518084
rect 181563 518050 181599 518084
rect 181655 518050 181663 518084
rect 177961 518041 177973 518050
rect 178025 518041 178037 518050
rect 178089 518041 181599 518050
rect 181651 518041 181663 518050
rect 181715 518041 181727 518050
rect 181779 518041 181791 518093
rect 181843 518041 181855 518093
rect 181907 518084 185417 518093
rect 181931 518050 181989 518084
rect 182023 518050 182081 518084
rect 182115 518050 182173 518084
rect 182207 518050 182265 518084
rect 182299 518050 182357 518084
rect 182391 518050 182449 518084
rect 182483 518050 182541 518084
rect 182575 518050 182633 518084
rect 182667 518050 182725 518084
rect 182759 518050 182817 518084
rect 182851 518050 182909 518084
rect 182943 518050 183001 518084
rect 183035 518050 183093 518084
rect 183127 518050 183185 518084
rect 183219 518050 183277 518084
rect 183311 518050 183369 518084
rect 183403 518050 183461 518084
rect 183495 518050 183553 518084
rect 183587 518050 183645 518084
rect 183679 518050 183737 518084
rect 183771 518050 183829 518084
rect 183863 518050 183921 518084
rect 183955 518050 184013 518084
rect 184047 518050 184105 518084
rect 184139 518050 184197 518084
rect 184231 518050 184289 518084
rect 184323 518050 184381 518084
rect 184415 518050 184473 518084
rect 184507 518050 184565 518084
rect 184599 518050 184657 518084
rect 184691 518050 184749 518084
rect 184783 518050 184841 518084
rect 184875 518050 184933 518084
rect 184967 518050 185025 518084
rect 185059 518050 185117 518084
rect 185151 518050 185209 518084
rect 185243 518050 185301 518084
rect 185335 518050 185393 518084
rect 181907 518041 185417 518050
rect 185469 518041 185481 518093
rect 185533 518041 185545 518093
rect 185597 518084 185609 518093
rect 185661 518084 185673 518093
rect 185725 518084 187480 518093
rect 185661 518050 185669 518084
rect 185725 518050 185761 518084
rect 185795 518050 185853 518084
rect 185887 518050 185945 518084
rect 185979 518050 186037 518084
rect 186071 518050 186129 518084
rect 186163 518050 186221 518084
rect 186255 518050 186313 518084
rect 186347 518050 186405 518084
rect 186439 518050 186497 518084
rect 186531 518050 186589 518084
rect 186623 518050 186681 518084
rect 186715 518050 186773 518084
rect 186807 518050 186865 518084
rect 186899 518050 186957 518084
rect 186991 518050 187049 518084
rect 187083 518050 187141 518084
rect 187175 518050 187233 518084
rect 187267 518050 187325 518084
rect 187359 518050 187417 518084
rect 187451 518050 187480 518084
rect 185597 518041 185609 518050
rect 185661 518041 185673 518050
rect 185725 518041 187480 518050
rect 172208 518019 187480 518041
rect 172208 517549 187480 517571
rect 172208 517540 174623 517549
rect 172208 517506 172237 517540
rect 172271 517506 172329 517540
rect 172363 517506 172421 517540
rect 172455 517506 172513 517540
rect 172547 517506 172605 517540
rect 172639 517506 172697 517540
rect 172731 517506 172789 517540
rect 172823 517506 172881 517540
rect 172915 517506 172973 517540
rect 173007 517506 173065 517540
rect 173099 517506 173157 517540
rect 173191 517506 173249 517540
rect 173283 517506 173341 517540
rect 173375 517506 173433 517540
rect 173467 517506 173525 517540
rect 173559 517506 173617 517540
rect 173651 517506 173709 517540
rect 173743 517506 173801 517540
rect 173835 517506 173893 517540
rect 173927 517506 173985 517540
rect 174019 517506 174077 517540
rect 174111 517506 174169 517540
rect 174203 517506 174261 517540
rect 174295 517506 174353 517540
rect 174387 517506 174445 517540
rect 174479 517506 174537 517540
rect 174571 517506 174623 517540
rect 172208 517497 174623 517506
rect 174675 517497 174687 517549
rect 174739 517540 174751 517549
rect 174803 517540 174815 517549
rect 174803 517506 174813 517540
rect 174739 517497 174751 517506
rect 174803 517497 174815 517506
rect 174867 517497 174879 517549
rect 174931 517540 178441 517549
rect 174939 517506 174997 517540
rect 175031 517506 175089 517540
rect 175123 517506 175181 517540
rect 175215 517506 175273 517540
rect 175307 517506 175365 517540
rect 175399 517506 175457 517540
rect 175491 517506 175549 517540
rect 175583 517506 175641 517540
rect 175675 517506 175733 517540
rect 175767 517506 175825 517540
rect 175859 517506 175917 517540
rect 175951 517506 176009 517540
rect 176043 517506 176101 517540
rect 176135 517506 176193 517540
rect 176227 517506 176285 517540
rect 176319 517506 176377 517540
rect 176411 517506 176469 517540
rect 176503 517506 176561 517540
rect 176595 517506 176653 517540
rect 176687 517506 176745 517540
rect 176779 517506 176837 517540
rect 176871 517506 176929 517540
rect 176963 517506 177021 517540
rect 177055 517506 177113 517540
rect 177147 517506 177205 517540
rect 177239 517506 177297 517540
rect 177331 517506 177389 517540
rect 177423 517506 177481 517540
rect 177515 517506 177573 517540
rect 177607 517506 177665 517540
rect 177699 517506 177757 517540
rect 177791 517506 177849 517540
rect 177883 517506 177941 517540
rect 177975 517506 178033 517540
rect 178067 517506 178125 517540
rect 178159 517506 178217 517540
rect 178251 517506 178309 517540
rect 178343 517506 178401 517540
rect 178435 517506 178441 517540
rect 174931 517497 178441 517506
rect 178493 517540 178505 517549
rect 178493 517497 178505 517506
rect 178557 517497 178569 517549
rect 178621 517497 178633 517549
rect 178685 517540 178697 517549
rect 178749 517540 182259 517549
rect 178749 517506 178769 517540
rect 178803 517506 178861 517540
rect 178895 517506 178953 517540
rect 178987 517506 179045 517540
rect 179079 517506 179137 517540
rect 179171 517506 179229 517540
rect 179263 517506 179321 517540
rect 179355 517506 179413 517540
rect 179447 517506 179505 517540
rect 179539 517506 179597 517540
rect 179631 517506 179689 517540
rect 179723 517506 179781 517540
rect 179815 517506 179873 517540
rect 179907 517506 179965 517540
rect 179999 517506 180057 517540
rect 180091 517506 180149 517540
rect 180183 517506 180241 517540
rect 180275 517506 180333 517540
rect 180367 517506 180425 517540
rect 180459 517506 180517 517540
rect 180551 517506 180609 517540
rect 180643 517506 180701 517540
rect 180735 517506 180793 517540
rect 180827 517506 180885 517540
rect 180919 517506 180977 517540
rect 181011 517506 181069 517540
rect 181103 517506 181161 517540
rect 181195 517506 181253 517540
rect 181287 517506 181345 517540
rect 181379 517506 181437 517540
rect 181471 517506 181529 517540
rect 181563 517506 181621 517540
rect 181655 517506 181713 517540
rect 181747 517506 181805 517540
rect 181839 517506 181897 517540
rect 181931 517506 181989 517540
rect 182023 517506 182081 517540
rect 182115 517506 182173 517540
rect 182207 517506 182259 517540
rect 178685 517497 178697 517506
rect 178749 517497 182259 517506
rect 182311 517497 182323 517549
rect 182375 517540 182387 517549
rect 182439 517540 182451 517549
rect 182439 517506 182449 517540
rect 182375 517497 182387 517506
rect 182439 517497 182451 517506
rect 182503 517497 182515 517549
rect 182567 517540 186077 517549
rect 182575 517506 182633 517540
rect 182667 517506 182725 517540
rect 182759 517506 182817 517540
rect 182851 517506 182909 517540
rect 182943 517506 183001 517540
rect 183035 517506 183093 517540
rect 183127 517506 183185 517540
rect 183219 517506 183277 517540
rect 183311 517506 183369 517540
rect 183403 517506 183461 517540
rect 183495 517506 183553 517540
rect 183587 517506 183645 517540
rect 183679 517506 183737 517540
rect 183771 517506 183829 517540
rect 183863 517506 183921 517540
rect 183955 517506 184013 517540
rect 184047 517506 184105 517540
rect 184139 517506 184197 517540
rect 184231 517506 184289 517540
rect 184323 517506 184381 517540
rect 184415 517506 184473 517540
rect 184507 517506 184565 517540
rect 184599 517506 184657 517540
rect 184691 517506 184749 517540
rect 184783 517506 184841 517540
rect 184875 517506 184933 517540
rect 184967 517506 185025 517540
rect 185059 517506 185117 517540
rect 185151 517506 185209 517540
rect 185243 517506 185301 517540
rect 185335 517506 185393 517540
rect 185427 517506 185485 517540
rect 185519 517506 185577 517540
rect 185611 517506 185669 517540
rect 185703 517506 185761 517540
rect 185795 517506 185853 517540
rect 185887 517506 185945 517540
rect 185979 517506 186037 517540
rect 186071 517506 186077 517540
rect 182567 517497 186077 517506
rect 186129 517540 186141 517549
rect 186129 517497 186141 517506
rect 186193 517497 186205 517549
rect 186257 517497 186269 517549
rect 186321 517540 186333 517549
rect 186385 517540 187480 517549
rect 186385 517506 186405 517540
rect 186439 517506 186497 517540
rect 186531 517506 186589 517540
rect 186623 517506 186681 517540
rect 186715 517506 186773 517540
rect 186807 517506 186865 517540
rect 186899 517506 186957 517540
rect 186991 517506 187049 517540
rect 187083 517506 187141 517540
rect 187175 517506 187233 517540
rect 187267 517506 187325 517540
rect 187359 517506 187417 517540
rect 187451 517506 187480 517540
rect 186321 517497 186333 517506
rect 186385 517497 187480 517506
rect 172208 517475 187480 517497
rect 177650 517395 177656 517447
rect 177708 517435 177714 517447
rect 178294 517435 178300 517447
rect 177708 517407 178300 517435
rect 177708 517395 177714 517407
rect 178294 517395 178300 517407
rect 178352 517395 178358 517447
rect 172208 517005 187480 517027
rect 172208 516996 173963 517005
rect 174015 516996 174027 517005
rect 174079 516996 174091 517005
rect 172208 516962 172237 516996
rect 172271 516962 172329 516996
rect 172363 516962 172421 516996
rect 172455 516962 172513 516996
rect 172547 516962 172605 516996
rect 172639 516962 172697 516996
rect 172731 516962 172789 516996
rect 172823 516962 172881 516996
rect 172915 516962 172973 516996
rect 173007 516962 173065 516996
rect 173099 516962 173157 516996
rect 173191 516962 173249 516996
rect 173283 516962 173341 516996
rect 173375 516962 173433 516996
rect 173467 516962 173525 516996
rect 173559 516962 173617 516996
rect 173651 516962 173709 516996
rect 173743 516962 173801 516996
rect 173835 516962 173893 516996
rect 173927 516962 173963 516996
rect 174019 516962 174027 516996
rect 172208 516953 173963 516962
rect 174015 516953 174027 516962
rect 174079 516953 174091 516962
rect 174143 516953 174155 517005
rect 174207 516953 174219 517005
rect 174271 516996 177781 517005
rect 174295 516962 174353 516996
rect 174387 516962 174445 516996
rect 174479 516962 174537 516996
rect 174571 516962 174629 516996
rect 174663 516962 174721 516996
rect 174755 516962 174813 516996
rect 174847 516962 174905 516996
rect 174939 516962 174997 516996
rect 175031 516962 175089 516996
rect 175123 516962 175181 516996
rect 175215 516962 175273 516996
rect 175307 516962 175365 516996
rect 175399 516962 175457 516996
rect 175491 516962 175549 516996
rect 175583 516962 175641 516996
rect 175675 516962 175733 516996
rect 175767 516962 175825 516996
rect 175859 516962 175917 516996
rect 175951 516962 176009 516996
rect 176043 516962 176101 516996
rect 176135 516962 176193 516996
rect 176227 516962 176285 516996
rect 176319 516962 176377 516996
rect 176411 516962 176469 516996
rect 176503 516962 176561 516996
rect 176595 516962 176653 516996
rect 176687 516962 176745 516996
rect 176779 516962 176837 516996
rect 176871 516962 176929 516996
rect 176963 516962 177021 516996
rect 177055 516962 177113 516996
rect 177147 516962 177205 516996
rect 177239 516962 177297 516996
rect 177331 516962 177389 516996
rect 177423 516962 177481 516996
rect 177515 516962 177573 516996
rect 177607 516962 177665 516996
rect 177699 516962 177757 516996
rect 174271 516953 177781 516962
rect 177833 516953 177845 517005
rect 177897 516953 177909 517005
rect 177961 516996 177973 517005
rect 178025 516996 178037 517005
rect 178089 516996 181599 517005
rect 181651 516996 181663 517005
rect 181715 516996 181727 517005
rect 178025 516962 178033 516996
rect 178089 516962 178125 516996
rect 178159 516962 178217 516996
rect 178251 516962 178309 516996
rect 178343 516962 178401 516996
rect 178435 516962 178493 516996
rect 178527 516962 178585 516996
rect 178619 516962 178677 516996
rect 178711 516962 178769 516996
rect 178803 516962 178861 516996
rect 178895 516962 178953 516996
rect 178987 516962 179045 516996
rect 179079 516962 179137 516996
rect 179171 516962 179229 516996
rect 179263 516962 179321 516996
rect 179355 516962 179413 516996
rect 179447 516962 179505 516996
rect 179539 516962 179597 516996
rect 179631 516962 179689 516996
rect 179723 516962 179781 516996
rect 179815 516962 179873 516996
rect 179907 516962 179965 516996
rect 179999 516962 180057 516996
rect 180091 516962 180149 516996
rect 180183 516962 180241 516996
rect 180275 516962 180333 516996
rect 180367 516962 180425 516996
rect 180459 516962 180517 516996
rect 180551 516962 180609 516996
rect 180643 516962 180701 516996
rect 180735 516962 180793 516996
rect 180827 516962 180885 516996
rect 180919 516962 180977 516996
rect 181011 516962 181069 516996
rect 181103 516962 181161 516996
rect 181195 516962 181253 516996
rect 181287 516962 181345 516996
rect 181379 516962 181437 516996
rect 181471 516962 181529 516996
rect 181563 516962 181599 516996
rect 181655 516962 181663 516996
rect 177961 516953 177973 516962
rect 178025 516953 178037 516962
rect 178089 516953 181599 516962
rect 181651 516953 181663 516962
rect 181715 516953 181727 516962
rect 181779 516953 181791 517005
rect 181843 516953 181855 517005
rect 181907 516996 185417 517005
rect 181931 516962 181989 516996
rect 182023 516962 182081 516996
rect 182115 516962 182173 516996
rect 182207 516962 182265 516996
rect 182299 516962 182357 516996
rect 182391 516962 182449 516996
rect 182483 516962 182541 516996
rect 182575 516962 182633 516996
rect 182667 516962 182725 516996
rect 182759 516962 182817 516996
rect 182851 516962 182909 516996
rect 182943 516962 183001 516996
rect 183035 516962 183093 516996
rect 183127 516962 183185 516996
rect 183219 516962 183277 516996
rect 183311 516962 183369 516996
rect 183403 516962 183461 516996
rect 183495 516962 183553 516996
rect 183587 516962 183645 516996
rect 183679 516962 183737 516996
rect 183771 516962 183829 516996
rect 183863 516962 183921 516996
rect 183955 516962 184013 516996
rect 184047 516962 184105 516996
rect 184139 516962 184197 516996
rect 184231 516962 184289 516996
rect 184323 516962 184381 516996
rect 184415 516962 184473 516996
rect 184507 516962 184565 516996
rect 184599 516962 184657 516996
rect 184691 516962 184749 516996
rect 184783 516962 184841 516996
rect 184875 516962 184933 516996
rect 184967 516962 185025 516996
rect 185059 516962 185117 516996
rect 185151 516962 185209 516996
rect 185243 516962 185301 516996
rect 185335 516962 185393 516996
rect 181907 516953 185417 516962
rect 185469 516953 185481 517005
rect 185533 516953 185545 517005
rect 185597 516996 185609 517005
rect 185661 516996 185673 517005
rect 185725 516996 187480 517005
rect 185661 516962 185669 516996
rect 185725 516962 185761 516996
rect 185795 516962 185853 516996
rect 185887 516962 185945 516996
rect 185979 516962 186037 516996
rect 186071 516962 186129 516996
rect 186163 516962 186221 516996
rect 186255 516962 186313 516996
rect 186347 516962 186405 516996
rect 186439 516962 186497 516996
rect 186531 516962 186589 516996
rect 186623 516962 186681 516996
rect 186715 516962 186773 516996
rect 186807 516962 186865 516996
rect 186899 516962 186957 516996
rect 186991 516962 187049 516996
rect 187083 516962 187141 516996
rect 187175 516962 187233 516996
rect 187267 516962 187325 516996
rect 187359 516962 187417 516996
rect 187451 516962 187480 516996
rect 185597 516953 185609 516962
rect 185661 516953 185673 516962
rect 185725 516953 187480 516962
rect 172208 516931 187480 516953
rect 172208 516461 187480 516483
rect 172208 516452 174623 516461
rect 172208 516418 172237 516452
rect 172271 516418 172329 516452
rect 172363 516418 172421 516452
rect 172455 516418 172513 516452
rect 172547 516418 172605 516452
rect 172639 516418 172697 516452
rect 172731 516418 172789 516452
rect 172823 516418 172881 516452
rect 172915 516418 172973 516452
rect 173007 516418 173065 516452
rect 173099 516418 173157 516452
rect 173191 516418 173249 516452
rect 173283 516418 173341 516452
rect 173375 516418 173433 516452
rect 173467 516418 173525 516452
rect 173559 516418 173617 516452
rect 173651 516418 173709 516452
rect 173743 516418 173801 516452
rect 173835 516418 173893 516452
rect 173927 516418 173985 516452
rect 174019 516418 174077 516452
rect 174111 516418 174169 516452
rect 174203 516418 174261 516452
rect 174295 516418 174353 516452
rect 174387 516418 174445 516452
rect 174479 516418 174537 516452
rect 174571 516418 174623 516452
rect 172208 516409 174623 516418
rect 174675 516409 174687 516461
rect 174739 516452 174751 516461
rect 174803 516452 174815 516461
rect 174803 516418 174813 516452
rect 174739 516409 174751 516418
rect 174803 516409 174815 516418
rect 174867 516409 174879 516461
rect 174931 516452 178441 516461
rect 174939 516418 174997 516452
rect 175031 516418 175089 516452
rect 175123 516418 175181 516452
rect 175215 516418 175273 516452
rect 175307 516418 175365 516452
rect 175399 516418 175457 516452
rect 175491 516418 175549 516452
rect 175583 516418 175641 516452
rect 175675 516418 175733 516452
rect 175767 516418 175825 516452
rect 175859 516418 175917 516452
rect 175951 516418 176009 516452
rect 176043 516418 176101 516452
rect 176135 516418 176193 516452
rect 176227 516418 176285 516452
rect 176319 516418 176377 516452
rect 176411 516418 176469 516452
rect 176503 516418 176561 516452
rect 176595 516418 176653 516452
rect 176687 516418 176745 516452
rect 176779 516418 176837 516452
rect 176871 516418 176929 516452
rect 176963 516418 177021 516452
rect 177055 516418 177113 516452
rect 177147 516418 177205 516452
rect 177239 516418 177297 516452
rect 177331 516418 177389 516452
rect 177423 516418 177481 516452
rect 177515 516418 177573 516452
rect 177607 516418 177665 516452
rect 177699 516418 177757 516452
rect 177791 516418 177849 516452
rect 177883 516418 177941 516452
rect 177975 516418 178033 516452
rect 178067 516418 178125 516452
rect 178159 516418 178217 516452
rect 178251 516418 178309 516452
rect 178343 516418 178401 516452
rect 178435 516418 178441 516452
rect 174931 516409 178441 516418
rect 178493 516452 178505 516461
rect 178493 516409 178505 516418
rect 178557 516409 178569 516461
rect 178621 516409 178633 516461
rect 178685 516452 178697 516461
rect 178749 516452 182259 516461
rect 178749 516418 178769 516452
rect 178803 516418 178861 516452
rect 178895 516418 178953 516452
rect 178987 516418 179045 516452
rect 179079 516418 179137 516452
rect 179171 516418 179229 516452
rect 179263 516418 179321 516452
rect 179355 516418 179413 516452
rect 179447 516418 179505 516452
rect 179539 516418 179597 516452
rect 179631 516418 179689 516452
rect 179723 516418 179781 516452
rect 179815 516418 179873 516452
rect 179907 516418 179965 516452
rect 179999 516418 180057 516452
rect 180091 516418 180149 516452
rect 180183 516418 180241 516452
rect 180275 516418 180333 516452
rect 180367 516418 180425 516452
rect 180459 516418 180517 516452
rect 180551 516418 180609 516452
rect 180643 516418 180701 516452
rect 180735 516418 180793 516452
rect 180827 516418 180885 516452
rect 180919 516418 180977 516452
rect 181011 516418 181069 516452
rect 181103 516418 181161 516452
rect 181195 516418 181253 516452
rect 181287 516418 181345 516452
rect 181379 516418 181437 516452
rect 181471 516418 181529 516452
rect 181563 516418 181621 516452
rect 181655 516418 181713 516452
rect 181747 516418 181805 516452
rect 181839 516418 181897 516452
rect 181931 516418 181989 516452
rect 182023 516418 182081 516452
rect 182115 516418 182173 516452
rect 182207 516418 182259 516452
rect 178685 516409 178697 516418
rect 178749 516409 182259 516418
rect 182311 516409 182323 516461
rect 182375 516452 182387 516461
rect 182439 516452 182451 516461
rect 182439 516418 182449 516452
rect 182375 516409 182387 516418
rect 182439 516409 182451 516418
rect 182503 516409 182515 516461
rect 182567 516452 186077 516461
rect 182575 516418 182633 516452
rect 182667 516418 182725 516452
rect 182759 516418 182817 516452
rect 182851 516418 182909 516452
rect 182943 516418 183001 516452
rect 183035 516418 183093 516452
rect 183127 516418 183185 516452
rect 183219 516418 183277 516452
rect 183311 516418 183369 516452
rect 183403 516418 183461 516452
rect 183495 516418 183553 516452
rect 183587 516418 183645 516452
rect 183679 516418 183737 516452
rect 183771 516418 183829 516452
rect 183863 516418 183921 516452
rect 183955 516418 184013 516452
rect 184047 516418 184105 516452
rect 184139 516418 184197 516452
rect 184231 516418 184289 516452
rect 184323 516418 184381 516452
rect 184415 516418 184473 516452
rect 184507 516418 184565 516452
rect 184599 516418 184657 516452
rect 184691 516418 184749 516452
rect 184783 516418 184841 516452
rect 184875 516418 184933 516452
rect 184967 516418 185025 516452
rect 185059 516418 185117 516452
rect 185151 516418 185209 516452
rect 185243 516418 185301 516452
rect 185335 516418 185393 516452
rect 185427 516418 185485 516452
rect 185519 516418 185577 516452
rect 185611 516418 185669 516452
rect 185703 516418 185761 516452
rect 185795 516418 185853 516452
rect 185887 516418 185945 516452
rect 185979 516418 186037 516452
rect 186071 516418 186077 516452
rect 182567 516409 186077 516418
rect 186129 516452 186141 516461
rect 186129 516409 186141 516418
rect 186193 516409 186205 516461
rect 186257 516409 186269 516461
rect 186321 516452 186333 516461
rect 186385 516452 187480 516461
rect 186385 516418 186405 516452
rect 186439 516418 186497 516452
rect 186531 516418 186589 516452
rect 186623 516418 186681 516452
rect 186715 516418 186773 516452
rect 186807 516418 186865 516452
rect 186899 516418 186957 516452
rect 186991 516418 187049 516452
rect 187083 516418 187141 516452
rect 187175 516418 187233 516452
rect 187267 516418 187325 516452
rect 187359 516418 187417 516452
rect 187451 516418 187480 516452
rect 186321 516409 186333 516418
rect 186385 516409 187480 516418
rect 172208 516387 187480 516409
rect 172208 515917 187480 515939
rect 172208 515908 173963 515917
rect 174015 515908 174027 515917
rect 174079 515908 174091 515917
rect 172208 515874 172237 515908
rect 172271 515874 172329 515908
rect 172363 515874 172421 515908
rect 172455 515874 172513 515908
rect 172547 515874 172605 515908
rect 172639 515874 172697 515908
rect 172731 515874 172789 515908
rect 172823 515874 172881 515908
rect 172915 515874 172973 515908
rect 173007 515874 173065 515908
rect 173099 515874 173157 515908
rect 173191 515874 173249 515908
rect 173283 515874 173341 515908
rect 173375 515874 173433 515908
rect 173467 515874 173525 515908
rect 173559 515874 173617 515908
rect 173651 515874 173709 515908
rect 173743 515874 173801 515908
rect 173835 515874 173893 515908
rect 173927 515874 173963 515908
rect 174019 515874 174027 515908
rect 172208 515865 173963 515874
rect 174015 515865 174027 515874
rect 174079 515865 174091 515874
rect 174143 515865 174155 515917
rect 174207 515865 174219 515917
rect 174271 515908 177781 515917
rect 174295 515874 174353 515908
rect 174387 515874 174445 515908
rect 174479 515874 174537 515908
rect 174571 515874 174629 515908
rect 174663 515874 174721 515908
rect 174755 515874 174813 515908
rect 174847 515874 174905 515908
rect 174939 515874 174997 515908
rect 175031 515874 175089 515908
rect 175123 515874 175181 515908
rect 175215 515874 175273 515908
rect 175307 515874 175365 515908
rect 175399 515874 175457 515908
rect 175491 515874 175549 515908
rect 175583 515874 175641 515908
rect 175675 515874 175733 515908
rect 175767 515874 175825 515908
rect 175859 515874 175917 515908
rect 175951 515874 176009 515908
rect 176043 515874 176101 515908
rect 176135 515874 176193 515908
rect 176227 515874 176285 515908
rect 176319 515874 176377 515908
rect 176411 515874 176469 515908
rect 176503 515874 176561 515908
rect 176595 515874 176653 515908
rect 176687 515874 176745 515908
rect 176779 515874 176837 515908
rect 176871 515874 176929 515908
rect 176963 515874 177021 515908
rect 177055 515874 177113 515908
rect 177147 515874 177205 515908
rect 177239 515874 177297 515908
rect 177331 515874 177389 515908
rect 177423 515874 177481 515908
rect 177515 515874 177573 515908
rect 177607 515874 177665 515908
rect 177699 515874 177757 515908
rect 174271 515865 177781 515874
rect 177833 515865 177845 515917
rect 177897 515865 177909 515917
rect 177961 515908 177973 515917
rect 178025 515908 178037 515917
rect 178089 515908 181599 515917
rect 181651 515908 181663 515917
rect 181715 515908 181727 515917
rect 178025 515874 178033 515908
rect 178089 515874 178125 515908
rect 178159 515874 178217 515908
rect 178251 515874 178309 515908
rect 178343 515874 178401 515908
rect 178435 515874 178493 515908
rect 178527 515874 178585 515908
rect 178619 515874 178677 515908
rect 178711 515874 178769 515908
rect 178803 515874 178861 515908
rect 178895 515874 178953 515908
rect 178987 515874 179045 515908
rect 179079 515874 179137 515908
rect 179171 515874 179229 515908
rect 179263 515874 179321 515908
rect 179355 515874 179413 515908
rect 179447 515874 179505 515908
rect 179539 515874 179597 515908
rect 179631 515874 179689 515908
rect 179723 515874 179781 515908
rect 179815 515874 179873 515908
rect 179907 515874 179965 515908
rect 179999 515874 180057 515908
rect 180091 515874 180149 515908
rect 180183 515874 180241 515908
rect 180275 515874 180333 515908
rect 180367 515874 180425 515908
rect 180459 515874 180517 515908
rect 180551 515874 180609 515908
rect 180643 515874 180701 515908
rect 180735 515874 180793 515908
rect 180827 515874 180885 515908
rect 180919 515874 180977 515908
rect 181011 515874 181069 515908
rect 181103 515874 181161 515908
rect 181195 515874 181253 515908
rect 181287 515874 181345 515908
rect 181379 515874 181437 515908
rect 181471 515874 181529 515908
rect 181563 515874 181599 515908
rect 181655 515874 181663 515908
rect 177961 515865 177973 515874
rect 178025 515865 178037 515874
rect 178089 515865 181599 515874
rect 181651 515865 181663 515874
rect 181715 515865 181727 515874
rect 181779 515865 181791 515917
rect 181843 515865 181855 515917
rect 181907 515908 185417 515917
rect 181931 515874 181989 515908
rect 182023 515874 182081 515908
rect 182115 515874 182173 515908
rect 182207 515874 182265 515908
rect 182299 515874 182357 515908
rect 182391 515874 182449 515908
rect 182483 515874 182541 515908
rect 182575 515874 182633 515908
rect 182667 515874 182725 515908
rect 182759 515874 182817 515908
rect 182851 515874 182909 515908
rect 182943 515874 183001 515908
rect 183035 515874 183093 515908
rect 183127 515874 183185 515908
rect 183219 515874 183277 515908
rect 183311 515874 183369 515908
rect 183403 515874 183461 515908
rect 183495 515874 183553 515908
rect 183587 515874 183645 515908
rect 183679 515874 183737 515908
rect 183771 515874 183829 515908
rect 183863 515874 183921 515908
rect 183955 515874 184013 515908
rect 184047 515874 184105 515908
rect 184139 515874 184197 515908
rect 184231 515874 184289 515908
rect 184323 515874 184381 515908
rect 184415 515874 184473 515908
rect 184507 515874 184565 515908
rect 184599 515874 184657 515908
rect 184691 515874 184749 515908
rect 184783 515874 184841 515908
rect 184875 515874 184933 515908
rect 184967 515874 185025 515908
rect 185059 515874 185117 515908
rect 185151 515874 185209 515908
rect 185243 515874 185301 515908
rect 185335 515874 185393 515908
rect 181907 515865 185417 515874
rect 185469 515865 185481 515917
rect 185533 515865 185545 515917
rect 185597 515908 185609 515917
rect 185661 515908 185673 515917
rect 185725 515908 187480 515917
rect 185661 515874 185669 515908
rect 185725 515874 185761 515908
rect 185795 515874 185853 515908
rect 185887 515874 185945 515908
rect 185979 515874 186037 515908
rect 186071 515874 186129 515908
rect 186163 515874 186221 515908
rect 186255 515874 186313 515908
rect 186347 515874 186405 515908
rect 186439 515874 186497 515908
rect 186531 515874 186589 515908
rect 186623 515874 186681 515908
rect 186715 515874 186773 515908
rect 186807 515874 186865 515908
rect 186899 515874 186957 515908
rect 186991 515874 187049 515908
rect 187083 515874 187141 515908
rect 187175 515874 187233 515908
rect 187267 515874 187325 515908
rect 187359 515874 187417 515908
rect 187451 515874 187480 515908
rect 185597 515865 185609 515874
rect 185661 515865 185673 515874
rect 185725 515865 187480 515874
rect 172208 515843 187480 515865
rect 173602 515763 173608 515815
rect 173660 515763 173666 515815
rect 181330 515763 181336 515815
rect 181388 515803 181394 515815
rect 182069 515806 182127 515812
rect 182069 515803 182081 515806
rect 181388 515775 182081 515803
rect 181388 515763 181394 515775
rect 182069 515772 182081 515775
rect 182115 515772 182127 515806
rect 182069 515766 182127 515772
rect 186574 515763 186580 515815
rect 186632 515763 186638 515815
rect 182253 515602 182311 515608
rect 182253 515599 182265 515602
rect 182176 515571 182265 515599
rect 173326 515491 173332 515543
rect 173384 515531 173390 515543
rect 173513 515534 173571 515540
rect 173513 515531 173525 515534
rect 173384 515503 173525 515531
rect 173384 515491 173390 515503
rect 173513 515500 173525 515503
rect 173559 515500 173571 515534
rect 173513 515494 173571 515500
rect 182176 515475 182204 515571
rect 182253 515568 182265 515571
rect 182299 515568 182311 515602
rect 182253 515562 182311 515568
rect 186482 515491 186488 515543
rect 186540 515491 186546 515543
rect 182158 515423 182164 515475
rect 182216 515423 182222 515475
rect 172208 515373 187480 515395
rect 172208 515364 174623 515373
rect 172208 515330 172237 515364
rect 172271 515330 172329 515364
rect 172363 515330 172421 515364
rect 172455 515330 172513 515364
rect 172547 515330 172605 515364
rect 172639 515330 172697 515364
rect 172731 515330 172789 515364
rect 172823 515330 172881 515364
rect 172915 515330 172973 515364
rect 173007 515330 173065 515364
rect 173099 515330 173157 515364
rect 173191 515330 173249 515364
rect 173283 515330 173341 515364
rect 173375 515330 173433 515364
rect 173467 515330 173525 515364
rect 173559 515330 173617 515364
rect 173651 515330 173709 515364
rect 173743 515330 173801 515364
rect 173835 515330 173893 515364
rect 173927 515330 173985 515364
rect 174019 515330 174077 515364
rect 174111 515330 174169 515364
rect 174203 515330 174261 515364
rect 174295 515330 174353 515364
rect 174387 515330 174445 515364
rect 174479 515330 174537 515364
rect 174571 515330 174623 515364
rect 172208 515321 174623 515330
rect 174675 515321 174687 515373
rect 174739 515364 174751 515373
rect 174803 515364 174815 515373
rect 174803 515330 174813 515364
rect 174739 515321 174751 515330
rect 174803 515321 174815 515330
rect 174867 515321 174879 515373
rect 174931 515364 178441 515373
rect 174939 515330 174997 515364
rect 175031 515330 175089 515364
rect 175123 515330 175181 515364
rect 175215 515330 175273 515364
rect 175307 515330 175365 515364
rect 175399 515330 175457 515364
rect 175491 515330 175549 515364
rect 175583 515330 175641 515364
rect 175675 515330 175733 515364
rect 175767 515330 175825 515364
rect 175859 515330 175917 515364
rect 175951 515330 176009 515364
rect 176043 515330 176101 515364
rect 176135 515330 176193 515364
rect 176227 515330 176285 515364
rect 176319 515330 176377 515364
rect 176411 515330 176469 515364
rect 176503 515330 176561 515364
rect 176595 515330 176653 515364
rect 176687 515330 176745 515364
rect 176779 515330 176837 515364
rect 176871 515330 176929 515364
rect 176963 515330 177021 515364
rect 177055 515330 177113 515364
rect 177147 515330 177205 515364
rect 177239 515330 177297 515364
rect 177331 515330 177389 515364
rect 177423 515330 177481 515364
rect 177515 515330 177573 515364
rect 177607 515330 177665 515364
rect 177699 515330 177757 515364
rect 177791 515330 177849 515364
rect 177883 515330 177941 515364
rect 177975 515330 178033 515364
rect 178067 515330 178125 515364
rect 178159 515330 178217 515364
rect 178251 515330 178309 515364
rect 178343 515330 178401 515364
rect 178435 515330 178441 515364
rect 174931 515321 178441 515330
rect 178493 515364 178505 515373
rect 178493 515321 178505 515330
rect 178557 515321 178569 515373
rect 178621 515321 178633 515373
rect 178685 515364 178697 515373
rect 178749 515364 182259 515373
rect 178749 515330 178769 515364
rect 178803 515330 178861 515364
rect 178895 515330 178953 515364
rect 178987 515330 179045 515364
rect 179079 515330 179137 515364
rect 179171 515330 179229 515364
rect 179263 515330 179321 515364
rect 179355 515330 179413 515364
rect 179447 515330 179505 515364
rect 179539 515330 179597 515364
rect 179631 515330 179689 515364
rect 179723 515330 179781 515364
rect 179815 515330 179873 515364
rect 179907 515330 179965 515364
rect 179999 515330 180057 515364
rect 180091 515330 180149 515364
rect 180183 515330 180241 515364
rect 180275 515330 180333 515364
rect 180367 515330 180425 515364
rect 180459 515330 180517 515364
rect 180551 515330 180609 515364
rect 180643 515330 180701 515364
rect 180735 515330 180793 515364
rect 180827 515330 180885 515364
rect 180919 515330 180977 515364
rect 181011 515330 181069 515364
rect 181103 515330 181161 515364
rect 181195 515330 181253 515364
rect 181287 515330 181345 515364
rect 181379 515330 181437 515364
rect 181471 515330 181529 515364
rect 181563 515330 181621 515364
rect 181655 515330 181713 515364
rect 181747 515330 181805 515364
rect 181839 515330 181897 515364
rect 181931 515330 181989 515364
rect 182023 515330 182081 515364
rect 182115 515330 182173 515364
rect 182207 515330 182259 515364
rect 178685 515321 178697 515330
rect 178749 515321 182259 515330
rect 182311 515321 182323 515373
rect 182375 515364 182387 515373
rect 182439 515364 182451 515373
rect 182439 515330 182449 515364
rect 182375 515321 182387 515330
rect 182439 515321 182451 515330
rect 182503 515321 182515 515373
rect 182567 515364 186077 515373
rect 182575 515330 182633 515364
rect 182667 515330 182725 515364
rect 182759 515330 182817 515364
rect 182851 515330 182909 515364
rect 182943 515330 183001 515364
rect 183035 515330 183093 515364
rect 183127 515330 183185 515364
rect 183219 515330 183277 515364
rect 183311 515330 183369 515364
rect 183403 515330 183461 515364
rect 183495 515330 183553 515364
rect 183587 515330 183645 515364
rect 183679 515330 183737 515364
rect 183771 515330 183829 515364
rect 183863 515330 183921 515364
rect 183955 515330 184013 515364
rect 184047 515330 184105 515364
rect 184139 515330 184197 515364
rect 184231 515330 184289 515364
rect 184323 515330 184381 515364
rect 184415 515330 184473 515364
rect 184507 515330 184565 515364
rect 184599 515330 184657 515364
rect 184691 515330 184749 515364
rect 184783 515330 184841 515364
rect 184875 515330 184933 515364
rect 184967 515330 185025 515364
rect 185059 515330 185117 515364
rect 185151 515330 185209 515364
rect 185243 515330 185301 515364
rect 185335 515330 185393 515364
rect 185427 515330 185485 515364
rect 185519 515330 185577 515364
rect 185611 515330 185669 515364
rect 185703 515330 185761 515364
rect 185795 515330 185853 515364
rect 185887 515330 185945 515364
rect 185979 515330 186037 515364
rect 186071 515330 186077 515364
rect 182567 515321 186077 515330
rect 186129 515364 186141 515373
rect 186129 515321 186141 515330
rect 186193 515321 186205 515373
rect 186257 515321 186269 515373
rect 186321 515364 186333 515373
rect 186385 515364 187480 515373
rect 186385 515330 186405 515364
rect 186439 515330 186497 515364
rect 186531 515330 186589 515364
rect 186623 515330 186681 515364
rect 186715 515330 186773 515364
rect 186807 515330 186865 515364
rect 186899 515330 186957 515364
rect 186991 515330 187049 515364
rect 187083 515330 187141 515364
rect 187175 515330 187233 515364
rect 187267 515330 187325 515364
rect 187359 515330 187417 515364
rect 187451 515330 187480 515364
rect 186321 515321 186333 515330
rect 186385 515321 187480 515330
rect 172208 515299 187480 515321
rect 173000 512810 173250 513000
rect 173450 512810 175000 513000
rect 173000 509000 175000 512810
rect 1990 507000 2000 509000
rect 4000 507000 175000 509000
rect 177000 512810 177580 513000
rect 177780 512810 179000 513000
rect 177000 506000 179000 512810
rect 5000 504000 179000 506000
rect 181000 512810 181910 513000
rect 182110 512810 183000 513000
rect 5000 466000 7000 504000
rect 181000 503000 183000 512810
rect 1990 464000 2000 466000
rect 4000 464000 7000 466000
rect 8000 501000 183000 503000
rect 185000 512810 186230 513000
rect 186430 512810 187000 513000
rect 8000 423000 10000 501000
rect 185000 500000 187000 512810
rect 1990 421000 2000 423000
rect 4000 421000 10000 423000
rect 11000 498000 187000 500000
rect 11000 380000 13000 498000
rect 1990 378000 2000 380000
rect 4000 378000 13000 380000
<< rmetal1 >>
rect 192108 522915 192138 523005
<< via1 >>
rect 18000 699000 20000 701000
rect 70000 699000 72000 701000
rect 122000 699000 124000 701000
rect 3000 682000 5000 684000
rect 146000 626000 148000 628000
rect 154000 551000 156000 553000
rect 146000 544000 148000 546000
rect 154000 538000 156000 540000
rect 161388 538545 161508 538665
rect 163028 538665 163328 538865
rect 159398 538215 159478 538295
rect 165888 540895 165943 540995
rect 165943 540895 165977 540995
rect 165977 540895 165998 540995
rect 165888 540775 165943 540875
rect 165943 540775 165977 540875
rect 165977 540775 165998 540875
rect 165888 540655 165943 540755
rect 165943 540655 165977 540755
rect 165977 540655 165998 540755
rect 166688 540065 166868 540245
rect 161688 537706 161748 537735
rect 161688 537675 161698 537706
rect 161698 537675 161732 537706
rect 161732 537675 161748 537706
rect 162878 537885 162938 537945
rect 165898 538705 166038 538805
rect 166688 539125 166868 539305
rect 157418 536845 157508 536925
rect 161788 536825 161848 536905
rect 158478 536395 158578 536555
rect 161088 536465 161168 536545
rect 160198 535435 160348 535575
rect 163838 535905 164048 536235
rect 166928 536045 167258 536265
rect 166718 535425 166848 535555
rect 166898 535415 167028 535545
rect 167078 535395 167208 535525
rect 166698 535235 166828 535365
rect 166888 535225 167018 535355
rect 167088 535215 167218 535345
rect 169688 540895 169743 540995
rect 169743 540895 169777 540995
rect 169777 540895 169798 540995
rect 169688 540775 169743 540875
rect 169743 540775 169777 540875
rect 169777 540775 169798 540875
rect 169688 540655 169743 540755
rect 169743 540655 169777 540755
rect 169777 540655 169798 540755
rect 170488 540065 170668 540245
rect 169698 538705 169838 538805
rect 170488 539125 170668 539305
rect 169568 535975 169868 536255
rect 173388 540895 173443 540995
rect 173443 540895 173477 540995
rect 173477 540895 173498 540995
rect 173388 540775 173443 540875
rect 173443 540775 173477 540875
rect 173477 540775 173498 540875
rect 173388 540655 173443 540755
rect 173443 540655 173477 540755
rect 173477 540655 173498 540755
rect 174188 540075 174368 540255
rect 173398 538705 173538 538805
rect 174188 539125 174368 539305
rect 172608 535975 172938 536265
rect 176888 540895 176943 540995
rect 176943 540895 176977 540995
rect 176977 540895 176998 540995
rect 176888 540775 176943 540875
rect 176943 540775 176977 540875
rect 176977 540775 176998 540875
rect 176888 540655 176943 540755
rect 176943 540655 176977 540755
rect 176977 540655 176998 540755
rect 177698 540065 177878 540245
rect 176898 538705 177038 538805
rect 177688 539125 177868 539305
rect 175278 536019 175358 536255
rect 175358 536019 175396 536255
rect 175396 536019 175498 536255
rect 175278 535945 175498 536019
rect 172358 532565 172488 532735
rect 174488 532575 174618 532745
rect 176578 532565 176708 532735
rect 180488 540895 180543 540995
rect 180543 540895 180577 540995
rect 180577 540895 180598 540995
rect 180488 540775 180543 540875
rect 180543 540775 180577 540875
rect 180577 540775 180598 540875
rect 180488 540655 180543 540755
rect 180543 540655 180577 540755
rect 180577 540655 180598 540755
rect 181288 540065 181468 540245
rect 180498 538705 180638 538805
rect 181288 539125 181468 539305
rect 178868 535965 179068 536275
rect 183788 540895 183843 540995
rect 183843 540895 183877 540995
rect 183877 540895 183898 540995
rect 183788 540775 183843 540875
rect 183843 540775 183877 540875
rect 183877 540775 183898 540875
rect 183788 540655 183843 540755
rect 183843 540655 183877 540755
rect 183877 540655 183898 540755
rect 184588 540065 184768 540245
rect 183798 538705 183938 538805
rect 184588 539125 184768 539305
rect 182188 536025 182388 536285
rect 187088 540895 187143 540995
rect 187143 540895 187177 540995
rect 187177 540895 187198 540995
rect 187088 540775 187143 540875
rect 187143 540775 187177 540875
rect 187177 540775 187198 540875
rect 187088 540655 187143 540755
rect 187143 540655 187177 540755
rect 187177 540655 187198 540755
rect 187898 540065 188078 540245
rect 187098 538705 187238 538805
rect 187888 539125 188068 539305
rect 185488 536145 185698 536265
rect 178698 532565 178828 532735
rect 180868 532565 180998 532735
rect 190388 540895 190443 540995
rect 190443 540895 190477 540995
rect 190477 540895 190498 540995
rect 190388 540775 190443 540875
rect 190443 540775 190477 540875
rect 190477 540775 190498 540875
rect 190388 540655 190443 540755
rect 190443 540655 190477 540755
rect 190477 540655 190498 540755
rect 191188 540065 191368 540245
rect 190398 538705 190538 538805
rect 191198 539135 191378 539315
rect 188778 536035 188998 536275
rect 182958 532565 183088 532735
rect 185058 532605 185188 532775
rect 191808 540065 191988 540245
rect 191818 539125 191998 539305
rect 187168 532595 187268 532735
rect 174623 530596 174675 530605
rect 174623 530562 174629 530596
rect 174629 530562 174663 530596
rect 174663 530562 174675 530596
rect 174623 530553 174675 530562
rect 174687 530596 174739 530605
rect 174751 530596 174803 530605
rect 174815 530596 174867 530605
rect 174687 530562 174721 530596
rect 174721 530562 174739 530596
rect 174751 530562 174755 530596
rect 174755 530562 174803 530596
rect 174815 530562 174847 530596
rect 174847 530562 174867 530596
rect 174687 530553 174739 530562
rect 174751 530553 174803 530562
rect 174815 530553 174867 530562
rect 174879 530596 174931 530605
rect 174879 530562 174905 530596
rect 174905 530562 174931 530596
rect 174879 530553 174931 530562
rect 178441 530553 178493 530605
rect 178505 530596 178557 530605
rect 178505 530562 178527 530596
rect 178527 530562 178557 530596
rect 178505 530553 178557 530562
rect 178569 530596 178621 530605
rect 178569 530562 178585 530596
rect 178585 530562 178619 530596
rect 178619 530562 178621 530596
rect 178569 530553 178621 530562
rect 178633 530596 178685 530605
rect 178697 530596 178749 530605
rect 182259 530596 182311 530605
rect 178633 530562 178677 530596
rect 178677 530562 178685 530596
rect 178697 530562 178711 530596
rect 178711 530562 178749 530596
rect 182259 530562 182265 530596
rect 182265 530562 182299 530596
rect 182299 530562 182311 530596
rect 178633 530553 178685 530562
rect 178697 530553 178749 530562
rect 182259 530553 182311 530562
rect 182323 530596 182375 530605
rect 182387 530596 182439 530605
rect 182451 530596 182503 530605
rect 182323 530562 182357 530596
rect 182357 530562 182375 530596
rect 182387 530562 182391 530596
rect 182391 530562 182439 530596
rect 182451 530562 182483 530596
rect 182483 530562 182503 530596
rect 182323 530553 182375 530562
rect 182387 530553 182439 530562
rect 182451 530553 182503 530562
rect 182515 530596 182567 530605
rect 182515 530562 182541 530596
rect 182541 530562 182567 530596
rect 182515 530553 182567 530562
rect 186077 530553 186129 530605
rect 186141 530596 186193 530605
rect 186141 530562 186163 530596
rect 186163 530562 186193 530596
rect 186141 530553 186193 530562
rect 186205 530596 186257 530605
rect 186205 530562 186221 530596
rect 186221 530562 186255 530596
rect 186255 530562 186257 530596
rect 186205 530553 186257 530562
rect 186269 530596 186321 530605
rect 186333 530596 186385 530605
rect 186269 530562 186313 530596
rect 186313 530562 186321 530596
rect 186333 530562 186347 530596
rect 186347 530562 186385 530596
rect 186269 530553 186321 530562
rect 186333 530553 186385 530562
rect 172412 530383 172464 530435
rect 174528 530383 174580 530435
rect 176828 530451 176880 530503
rect 178760 530494 178812 530503
rect 178760 530460 178769 530494
rect 178769 530460 178803 530494
rect 178803 530460 178812 530494
rect 178760 530451 178812 530460
rect 174804 530315 174856 530367
rect 175448 530315 175500 530367
rect 176736 530383 176788 530435
rect 179496 530451 179548 530503
rect 182992 530451 183044 530503
rect 185108 530451 185160 530503
rect 178944 530315 178996 530367
rect 179220 530315 179272 530367
rect 176644 530247 176696 530299
rect 177288 530290 177340 530299
rect 177288 530256 177297 530290
rect 177297 530256 177331 530290
rect 177331 530256 177340 530290
rect 177288 530247 177340 530256
rect 178208 530290 178260 530299
rect 178208 530256 178217 530290
rect 178217 530256 178251 530290
rect 178251 530256 178260 530290
rect 178208 530247 178260 530256
rect 180692 530247 180744 530299
rect 182256 530315 182308 530367
rect 183176 530358 183228 530367
rect 183176 530324 183185 530358
rect 183185 530324 183219 530358
rect 183219 530324 183228 530358
rect 183176 530315 183228 530324
rect 187132 530358 187184 530367
rect 187132 530324 187141 530358
rect 187141 530324 187175 530358
rect 187175 530324 187184 530358
rect 187132 530315 187184 530324
rect 182624 530247 182676 530299
rect 177656 530154 177708 530163
rect 177656 530120 177665 530154
rect 177665 530120 177699 530154
rect 177699 530120 177708 530154
rect 177656 530111 177708 530120
rect 178300 530111 178352 530163
rect 179680 530111 179732 530163
rect 182164 530154 182216 530163
rect 182164 530120 182173 530154
rect 182173 530120 182207 530154
rect 182207 530120 182216 530154
rect 182164 530111 182216 530120
rect 182716 530111 182768 530163
rect 173963 530052 174015 530061
rect 174027 530052 174079 530061
rect 174091 530052 174143 530061
rect 173963 530018 173985 530052
rect 173985 530018 174015 530052
rect 174027 530018 174077 530052
rect 174077 530018 174079 530052
rect 174091 530018 174111 530052
rect 174111 530018 174143 530052
rect 173963 530009 174015 530018
rect 174027 530009 174079 530018
rect 174091 530009 174143 530018
rect 174155 530052 174207 530061
rect 174155 530018 174169 530052
rect 174169 530018 174203 530052
rect 174203 530018 174207 530052
rect 174155 530009 174207 530018
rect 174219 530052 174271 530061
rect 177781 530052 177833 530061
rect 174219 530018 174261 530052
rect 174261 530018 174271 530052
rect 177781 530018 177791 530052
rect 177791 530018 177833 530052
rect 174219 530009 174271 530018
rect 177781 530009 177833 530018
rect 177845 530052 177897 530061
rect 177845 530018 177849 530052
rect 177849 530018 177883 530052
rect 177883 530018 177897 530052
rect 177845 530009 177897 530018
rect 177909 530052 177961 530061
rect 177973 530052 178025 530061
rect 178037 530052 178089 530061
rect 181599 530052 181651 530061
rect 181663 530052 181715 530061
rect 181727 530052 181779 530061
rect 177909 530018 177941 530052
rect 177941 530018 177961 530052
rect 177973 530018 177975 530052
rect 177975 530018 178025 530052
rect 178037 530018 178067 530052
rect 178067 530018 178089 530052
rect 181599 530018 181621 530052
rect 181621 530018 181651 530052
rect 181663 530018 181713 530052
rect 181713 530018 181715 530052
rect 181727 530018 181747 530052
rect 181747 530018 181779 530052
rect 177909 530009 177961 530018
rect 177973 530009 178025 530018
rect 178037 530009 178089 530018
rect 181599 530009 181651 530018
rect 181663 530009 181715 530018
rect 181727 530009 181779 530018
rect 181791 530052 181843 530061
rect 181791 530018 181805 530052
rect 181805 530018 181839 530052
rect 181839 530018 181843 530052
rect 181791 530009 181843 530018
rect 181855 530052 181907 530061
rect 185417 530052 185469 530061
rect 181855 530018 181897 530052
rect 181897 530018 181907 530052
rect 185417 530018 185427 530052
rect 185427 530018 185469 530052
rect 181855 530009 181907 530018
rect 185417 530009 185469 530018
rect 185481 530052 185533 530061
rect 185481 530018 185485 530052
rect 185485 530018 185519 530052
rect 185519 530018 185533 530052
rect 185481 530009 185533 530018
rect 185545 530052 185597 530061
rect 185609 530052 185661 530061
rect 185673 530052 185725 530061
rect 185545 530018 185577 530052
rect 185577 530018 185597 530052
rect 185609 530018 185611 530052
rect 185611 530018 185661 530052
rect 185673 530018 185703 530052
rect 185703 530018 185725 530052
rect 185545 530009 185597 530018
rect 185609 530009 185661 530018
rect 185673 530009 185725 530018
rect 178208 529907 178260 529959
rect 179496 529907 179548 529959
rect 180876 529907 180928 529959
rect 182164 529907 182216 529959
rect 182624 529950 182676 529959
rect 182624 529916 182633 529950
rect 182633 529916 182667 529950
rect 182667 529916 182676 529950
rect 182624 529907 182676 529916
rect 178116 529839 178168 529891
rect 174804 529814 174856 529823
rect 174804 529780 174813 529814
rect 174813 529780 174847 529814
rect 174847 529780 174856 529814
rect 174804 529771 174856 529780
rect 176828 529703 176880 529755
rect 179312 529771 179364 529823
rect 179864 529814 179916 529823
rect 179864 529780 179873 529814
rect 179873 529780 179907 529814
rect 179907 529780 179916 529814
rect 179864 529771 179916 529780
rect 175356 529567 175408 529619
rect 176092 529567 176144 529619
rect 177380 529635 177432 529687
rect 177564 529635 177616 529687
rect 177656 529635 177708 529687
rect 177932 529567 177984 529619
rect 181520 529635 181572 529687
rect 183176 529814 183228 529823
rect 183176 529780 183185 529814
rect 183185 529780 183219 529814
rect 183219 529780 183228 529814
rect 183176 529771 183228 529780
rect 180508 529567 180560 529619
rect 181796 529567 181848 529619
rect 174623 529508 174675 529517
rect 174623 529474 174629 529508
rect 174629 529474 174663 529508
rect 174663 529474 174675 529508
rect 174623 529465 174675 529474
rect 174687 529508 174739 529517
rect 174751 529508 174803 529517
rect 174815 529508 174867 529517
rect 174687 529474 174721 529508
rect 174721 529474 174739 529508
rect 174751 529474 174755 529508
rect 174755 529474 174803 529508
rect 174815 529474 174847 529508
rect 174847 529474 174867 529508
rect 174687 529465 174739 529474
rect 174751 529465 174803 529474
rect 174815 529465 174867 529474
rect 174879 529508 174931 529517
rect 174879 529474 174905 529508
rect 174905 529474 174931 529508
rect 174879 529465 174931 529474
rect 178441 529465 178493 529517
rect 178505 529508 178557 529517
rect 178505 529474 178527 529508
rect 178527 529474 178557 529508
rect 178505 529465 178557 529474
rect 178569 529508 178621 529517
rect 178569 529474 178585 529508
rect 178585 529474 178619 529508
rect 178619 529474 178621 529508
rect 178569 529465 178621 529474
rect 178633 529508 178685 529517
rect 178697 529508 178749 529517
rect 182259 529508 182311 529517
rect 178633 529474 178677 529508
rect 178677 529474 178685 529508
rect 178697 529474 178711 529508
rect 178711 529474 178749 529508
rect 182259 529474 182265 529508
rect 182265 529474 182299 529508
rect 182299 529474 182311 529508
rect 178633 529465 178685 529474
rect 178697 529465 178749 529474
rect 182259 529465 182311 529474
rect 182323 529508 182375 529517
rect 182387 529508 182439 529517
rect 182451 529508 182503 529517
rect 182323 529474 182357 529508
rect 182357 529474 182375 529508
rect 182387 529474 182391 529508
rect 182391 529474 182439 529508
rect 182451 529474 182483 529508
rect 182483 529474 182503 529508
rect 182323 529465 182375 529474
rect 182387 529465 182439 529474
rect 182451 529465 182503 529474
rect 182515 529508 182567 529517
rect 182515 529474 182541 529508
rect 182541 529474 182567 529508
rect 182515 529465 182567 529474
rect 186077 529465 186129 529517
rect 186141 529508 186193 529517
rect 186141 529474 186163 529508
rect 186163 529474 186193 529508
rect 186141 529465 186193 529474
rect 186205 529508 186257 529517
rect 186205 529474 186221 529508
rect 186221 529474 186255 529508
rect 186255 529474 186257 529508
rect 186205 529465 186257 529474
rect 186269 529508 186321 529517
rect 186333 529508 186385 529517
rect 186269 529474 186313 529508
rect 186313 529474 186321 529508
rect 186333 529474 186347 529508
rect 186347 529474 186385 529508
rect 186269 529465 186321 529474
rect 186333 529465 186385 529474
rect 175356 529406 175408 529415
rect 175356 529372 175365 529406
rect 175365 529372 175399 529406
rect 175399 529372 175408 529406
rect 175356 529363 175408 529372
rect 177932 529363 177984 529415
rect 178300 529295 178352 529347
rect 179864 529406 179916 529415
rect 179864 529372 179873 529406
rect 179873 529372 179907 529406
rect 179907 529372 179916 529406
rect 179864 529363 179916 529372
rect 181796 529363 181848 529415
rect 175448 529270 175500 529279
rect 175448 529236 175457 529270
rect 175457 529236 175491 529270
rect 175491 529236 175500 529270
rect 175448 529227 175500 529236
rect 176736 529227 176788 529279
rect 177656 529270 177708 529279
rect 177656 529236 177665 529270
rect 177665 529236 177699 529270
rect 177699 529236 177708 529270
rect 177656 529227 177708 529236
rect 179680 529270 179732 529279
rect 179680 529236 179689 529270
rect 179689 529236 179723 529270
rect 179723 529236 179732 529270
rect 179680 529227 179732 529236
rect 173608 529159 173660 529211
rect 175264 529202 175316 529211
rect 175264 529168 175273 529202
rect 175273 529168 175307 529202
rect 175307 529168 175316 529202
rect 175264 529159 175316 529168
rect 175908 529023 175960 529075
rect 176092 529023 176144 529075
rect 177288 529159 177340 529211
rect 181520 529227 181572 529279
rect 182716 529270 182768 529279
rect 182716 529236 182725 529270
rect 182725 529236 182759 529270
rect 182759 529236 182768 529270
rect 182716 529227 182768 529236
rect 179312 529023 179364 529075
rect 179680 529023 179732 529075
rect 180508 529023 180560 529075
rect 173963 528964 174015 528973
rect 174027 528964 174079 528973
rect 174091 528964 174143 528973
rect 173963 528930 173985 528964
rect 173985 528930 174015 528964
rect 174027 528930 174077 528964
rect 174077 528930 174079 528964
rect 174091 528930 174111 528964
rect 174111 528930 174143 528964
rect 173963 528921 174015 528930
rect 174027 528921 174079 528930
rect 174091 528921 174143 528930
rect 174155 528964 174207 528973
rect 174155 528930 174169 528964
rect 174169 528930 174203 528964
rect 174203 528930 174207 528964
rect 174155 528921 174207 528930
rect 174219 528964 174271 528973
rect 177781 528964 177833 528973
rect 174219 528930 174261 528964
rect 174261 528930 174271 528964
rect 177781 528930 177791 528964
rect 177791 528930 177833 528964
rect 174219 528921 174271 528930
rect 177781 528921 177833 528930
rect 177845 528964 177897 528973
rect 177845 528930 177849 528964
rect 177849 528930 177883 528964
rect 177883 528930 177897 528964
rect 177845 528921 177897 528930
rect 177909 528964 177961 528973
rect 177973 528964 178025 528973
rect 178037 528964 178089 528973
rect 181599 528964 181651 528973
rect 181663 528964 181715 528973
rect 181727 528964 181779 528973
rect 177909 528930 177941 528964
rect 177941 528930 177961 528964
rect 177973 528930 177975 528964
rect 177975 528930 178025 528964
rect 178037 528930 178067 528964
rect 178067 528930 178089 528964
rect 181599 528930 181621 528964
rect 181621 528930 181651 528964
rect 181663 528930 181713 528964
rect 181713 528930 181715 528964
rect 181727 528930 181747 528964
rect 181747 528930 181779 528964
rect 177909 528921 177961 528930
rect 177973 528921 178025 528930
rect 178037 528921 178089 528930
rect 181599 528921 181651 528930
rect 181663 528921 181715 528930
rect 181727 528921 181779 528930
rect 181791 528964 181843 528973
rect 181791 528930 181805 528964
rect 181805 528930 181839 528964
rect 181839 528930 181843 528964
rect 181791 528921 181843 528930
rect 181855 528964 181907 528973
rect 185417 528964 185469 528973
rect 181855 528930 181897 528964
rect 181897 528930 181907 528964
rect 185417 528930 185427 528964
rect 185427 528930 185469 528964
rect 181855 528921 181907 528930
rect 185417 528921 185469 528930
rect 185481 528964 185533 528973
rect 185481 528930 185485 528964
rect 185485 528930 185519 528964
rect 185519 528930 185533 528964
rect 185481 528921 185533 528930
rect 185545 528964 185597 528973
rect 185609 528964 185661 528973
rect 185673 528964 185725 528973
rect 185545 528930 185577 528964
rect 185577 528930 185597 528964
rect 185609 528930 185611 528964
rect 185611 528930 185661 528964
rect 185673 528930 185703 528964
rect 185703 528930 185725 528964
rect 185545 528921 185597 528930
rect 185609 528921 185661 528930
rect 185673 528921 185725 528930
rect 175264 528819 175316 528871
rect 176644 528819 176696 528871
rect 177656 528819 177708 528871
rect 179680 528862 179732 528871
rect 179680 528828 179689 528862
rect 179689 528828 179723 528862
rect 179723 528828 179732 528862
rect 179680 528819 179732 528828
rect 177564 528683 177616 528735
rect 178024 528683 178076 528735
rect 178208 528683 178260 528735
rect 180508 528726 180560 528735
rect 180508 528692 180517 528726
rect 180517 528692 180551 528726
rect 180551 528692 180560 528726
rect 180508 528683 180560 528692
rect 182164 528819 182216 528871
rect 181520 528683 181572 528735
rect 175908 528658 175960 528667
rect 175908 528624 175917 528658
rect 175917 528624 175951 528658
rect 175951 528624 175960 528658
rect 175908 528615 175960 528624
rect 178392 528590 178444 528599
rect 178392 528556 178401 528590
rect 178401 528556 178435 528590
rect 178435 528556 178444 528590
rect 178392 528547 178444 528556
rect 186580 528547 186632 528599
rect 176276 528479 176328 528531
rect 176368 528522 176420 528531
rect 176368 528488 176377 528522
rect 176377 528488 176411 528522
rect 176411 528488 176420 528522
rect 176368 528479 176420 528488
rect 176736 528522 176788 528531
rect 176736 528488 176745 528522
rect 176745 528488 176779 528522
rect 176779 528488 176788 528522
rect 176736 528479 176788 528488
rect 177012 528479 177064 528531
rect 180968 528479 181020 528531
rect 174623 528420 174675 528429
rect 174623 528386 174629 528420
rect 174629 528386 174663 528420
rect 174663 528386 174675 528420
rect 174623 528377 174675 528386
rect 174687 528420 174739 528429
rect 174751 528420 174803 528429
rect 174815 528420 174867 528429
rect 174687 528386 174721 528420
rect 174721 528386 174739 528420
rect 174751 528386 174755 528420
rect 174755 528386 174803 528420
rect 174815 528386 174847 528420
rect 174847 528386 174867 528420
rect 174687 528377 174739 528386
rect 174751 528377 174803 528386
rect 174815 528377 174867 528386
rect 174879 528420 174931 528429
rect 174879 528386 174905 528420
rect 174905 528386 174931 528420
rect 174879 528377 174931 528386
rect 178441 528377 178493 528429
rect 178505 528420 178557 528429
rect 178505 528386 178527 528420
rect 178527 528386 178557 528420
rect 178505 528377 178557 528386
rect 178569 528420 178621 528429
rect 178569 528386 178585 528420
rect 178585 528386 178619 528420
rect 178619 528386 178621 528420
rect 178569 528377 178621 528386
rect 178633 528420 178685 528429
rect 178697 528420 178749 528429
rect 182259 528420 182311 528429
rect 178633 528386 178677 528420
rect 178677 528386 178685 528420
rect 178697 528386 178711 528420
rect 178711 528386 178749 528420
rect 182259 528386 182265 528420
rect 182265 528386 182299 528420
rect 182299 528386 182311 528420
rect 178633 528377 178685 528386
rect 178697 528377 178749 528386
rect 182259 528377 182311 528386
rect 182323 528420 182375 528429
rect 182387 528420 182439 528429
rect 182451 528420 182503 528429
rect 182323 528386 182357 528420
rect 182357 528386 182375 528420
rect 182387 528386 182391 528420
rect 182391 528386 182439 528420
rect 182451 528386 182483 528420
rect 182483 528386 182503 528420
rect 182323 528377 182375 528386
rect 182387 528377 182439 528386
rect 182451 528377 182503 528386
rect 182515 528420 182567 528429
rect 182515 528386 182541 528420
rect 182541 528386 182567 528420
rect 182515 528377 182567 528386
rect 186077 528377 186129 528429
rect 186141 528420 186193 528429
rect 186141 528386 186163 528420
rect 186163 528386 186193 528420
rect 186141 528377 186193 528386
rect 186205 528420 186257 528429
rect 186205 528386 186221 528420
rect 186221 528386 186255 528420
rect 186255 528386 186257 528420
rect 186205 528377 186257 528386
rect 186269 528420 186321 528429
rect 186333 528420 186385 528429
rect 186269 528386 186313 528420
rect 186313 528386 186321 528420
rect 186333 528386 186347 528420
rect 186347 528386 186385 528420
rect 186269 528377 186321 528386
rect 186333 528377 186385 528386
rect 176736 528275 176788 528327
rect 178024 528275 178076 528327
rect 178944 528318 178996 528327
rect 178944 528284 178953 528318
rect 178953 528284 178987 528318
rect 178987 528284 178996 528318
rect 178944 528275 178996 528284
rect 179312 528275 179364 528327
rect 180968 528318 181020 528327
rect 180968 528284 180977 528318
rect 180977 528284 181011 528318
rect 181011 528284 181020 528318
rect 180968 528275 181020 528284
rect 182164 528275 182216 528327
rect 176368 528250 176420 528259
rect 176368 528216 176377 528250
rect 176377 528216 176411 528250
rect 176411 528216 176420 528250
rect 176368 528207 176420 528216
rect 176828 528250 176880 528259
rect 176828 528216 176833 528250
rect 176833 528216 176867 528250
rect 176867 528216 176880 528250
rect 176828 528207 176880 528216
rect 176092 528182 176144 528191
rect 176092 528148 176101 528182
rect 176101 528148 176135 528182
rect 176135 528148 176144 528182
rect 176092 528139 176144 528148
rect 178116 528182 178168 528191
rect 178116 528148 178125 528182
rect 178125 528148 178159 528182
rect 178159 528148 178168 528182
rect 178116 528139 178168 528148
rect 177380 528003 177432 528055
rect 178944 527935 178996 527987
rect 181336 528182 181388 528191
rect 181336 528148 181345 528182
rect 181345 528148 181379 528182
rect 181379 528148 181388 528182
rect 181336 528139 181388 528148
rect 180692 528071 180744 528123
rect 173963 527876 174015 527885
rect 174027 527876 174079 527885
rect 174091 527876 174143 527885
rect 173963 527842 173985 527876
rect 173985 527842 174015 527876
rect 174027 527842 174077 527876
rect 174077 527842 174079 527876
rect 174091 527842 174111 527876
rect 174111 527842 174143 527876
rect 173963 527833 174015 527842
rect 174027 527833 174079 527842
rect 174091 527833 174143 527842
rect 174155 527876 174207 527885
rect 174155 527842 174169 527876
rect 174169 527842 174203 527876
rect 174203 527842 174207 527876
rect 174155 527833 174207 527842
rect 174219 527876 174271 527885
rect 177781 527876 177833 527885
rect 174219 527842 174261 527876
rect 174261 527842 174271 527876
rect 177781 527842 177791 527876
rect 177791 527842 177833 527876
rect 174219 527833 174271 527842
rect 177781 527833 177833 527842
rect 177845 527876 177897 527885
rect 177845 527842 177849 527876
rect 177849 527842 177883 527876
rect 177883 527842 177897 527876
rect 177845 527833 177897 527842
rect 177909 527876 177961 527885
rect 177973 527876 178025 527885
rect 178037 527876 178089 527885
rect 181599 527876 181651 527885
rect 181663 527876 181715 527885
rect 181727 527876 181779 527885
rect 177909 527842 177941 527876
rect 177941 527842 177961 527876
rect 177973 527842 177975 527876
rect 177975 527842 178025 527876
rect 178037 527842 178067 527876
rect 178067 527842 178089 527876
rect 181599 527842 181621 527876
rect 181621 527842 181651 527876
rect 181663 527842 181713 527876
rect 181713 527842 181715 527876
rect 181727 527842 181747 527876
rect 181747 527842 181779 527876
rect 177909 527833 177961 527842
rect 177973 527833 178025 527842
rect 178037 527833 178089 527842
rect 181599 527833 181651 527842
rect 181663 527833 181715 527842
rect 181727 527833 181779 527842
rect 181791 527876 181843 527885
rect 181791 527842 181805 527876
rect 181805 527842 181839 527876
rect 181839 527842 181843 527876
rect 181791 527833 181843 527842
rect 181855 527876 181907 527885
rect 185417 527876 185469 527885
rect 181855 527842 181897 527876
rect 181897 527842 181907 527876
rect 185417 527842 185427 527876
rect 185427 527842 185469 527876
rect 181855 527833 181907 527842
rect 185417 527833 185469 527842
rect 185481 527876 185533 527885
rect 185481 527842 185485 527876
rect 185485 527842 185519 527876
rect 185519 527842 185533 527876
rect 185481 527833 185533 527842
rect 185545 527876 185597 527885
rect 185609 527876 185661 527885
rect 185673 527876 185725 527885
rect 185545 527842 185577 527876
rect 185577 527842 185597 527876
rect 185609 527842 185611 527876
rect 185611 527842 185661 527876
rect 185673 527842 185703 527876
rect 185703 527842 185725 527876
rect 185545 527833 185597 527842
rect 185609 527833 185661 527842
rect 185673 527833 185725 527842
rect 176276 527731 176328 527783
rect 178944 527774 178996 527783
rect 178944 527740 178953 527774
rect 178953 527740 178987 527774
rect 178987 527740 178996 527774
rect 178944 527731 178996 527740
rect 177012 527638 177064 527647
rect 177012 527604 177021 527638
rect 177021 527604 177055 527638
rect 177055 527604 177064 527638
rect 177012 527595 177064 527604
rect 179496 527638 179548 527647
rect 179496 527604 179505 527638
rect 179505 527604 179539 527638
rect 179539 527604 179548 527638
rect 179496 527595 179548 527604
rect 174623 527332 174675 527341
rect 174623 527298 174629 527332
rect 174629 527298 174663 527332
rect 174663 527298 174675 527332
rect 174623 527289 174675 527298
rect 174687 527332 174739 527341
rect 174751 527332 174803 527341
rect 174815 527332 174867 527341
rect 174687 527298 174721 527332
rect 174721 527298 174739 527332
rect 174751 527298 174755 527332
rect 174755 527298 174803 527332
rect 174815 527298 174847 527332
rect 174847 527298 174867 527332
rect 174687 527289 174739 527298
rect 174751 527289 174803 527298
rect 174815 527289 174867 527298
rect 174879 527332 174931 527341
rect 174879 527298 174905 527332
rect 174905 527298 174931 527332
rect 174879 527289 174931 527298
rect 178441 527289 178493 527341
rect 178505 527332 178557 527341
rect 178505 527298 178527 527332
rect 178527 527298 178557 527332
rect 178505 527289 178557 527298
rect 178569 527332 178621 527341
rect 178569 527298 178585 527332
rect 178585 527298 178619 527332
rect 178619 527298 178621 527332
rect 178569 527289 178621 527298
rect 178633 527332 178685 527341
rect 178697 527332 178749 527341
rect 182259 527332 182311 527341
rect 178633 527298 178677 527332
rect 178677 527298 178685 527332
rect 178697 527298 178711 527332
rect 178711 527298 178749 527332
rect 182259 527298 182265 527332
rect 182265 527298 182299 527332
rect 182299 527298 182311 527332
rect 178633 527289 178685 527298
rect 178697 527289 178749 527298
rect 182259 527289 182311 527298
rect 182323 527332 182375 527341
rect 182387 527332 182439 527341
rect 182451 527332 182503 527341
rect 182323 527298 182357 527332
rect 182357 527298 182375 527332
rect 182387 527298 182391 527332
rect 182391 527298 182439 527332
rect 182451 527298 182483 527332
rect 182483 527298 182503 527332
rect 182323 527289 182375 527298
rect 182387 527289 182439 527298
rect 182451 527289 182503 527298
rect 182515 527332 182567 527341
rect 182515 527298 182541 527332
rect 182541 527298 182567 527332
rect 182515 527289 182567 527298
rect 186077 527289 186129 527341
rect 186141 527332 186193 527341
rect 186141 527298 186163 527332
rect 186163 527298 186193 527332
rect 186141 527289 186193 527298
rect 186205 527332 186257 527341
rect 186205 527298 186221 527332
rect 186221 527298 186255 527332
rect 186255 527298 186257 527332
rect 186205 527289 186257 527298
rect 186269 527332 186321 527341
rect 186333 527332 186385 527341
rect 186269 527298 186313 527332
rect 186313 527298 186321 527332
rect 186333 527298 186347 527332
rect 186347 527298 186385 527332
rect 186269 527289 186321 527298
rect 186333 527289 186385 527298
rect 173963 526788 174015 526797
rect 174027 526788 174079 526797
rect 174091 526788 174143 526797
rect 173963 526754 173985 526788
rect 173985 526754 174015 526788
rect 174027 526754 174077 526788
rect 174077 526754 174079 526788
rect 174091 526754 174111 526788
rect 174111 526754 174143 526788
rect 173963 526745 174015 526754
rect 174027 526745 174079 526754
rect 174091 526745 174143 526754
rect 174155 526788 174207 526797
rect 174155 526754 174169 526788
rect 174169 526754 174203 526788
rect 174203 526754 174207 526788
rect 174155 526745 174207 526754
rect 174219 526788 174271 526797
rect 177781 526788 177833 526797
rect 174219 526754 174261 526788
rect 174261 526754 174271 526788
rect 177781 526754 177791 526788
rect 177791 526754 177833 526788
rect 174219 526745 174271 526754
rect 177781 526745 177833 526754
rect 177845 526788 177897 526797
rect 177845 526754 177849 526788
rect 177849 526754 177883 526788
rect 177883 526754 177897 526788
rect 177845 526745 177897 526754
rect 177909 526788 177961 526797
rect 177973 526788 178025 526797
rect 178037 526788 178089 526797
rect 181599 526788 181651 526797
rect 181663 526788 181715 526797
rect 181727 526788 181779 526797
rect 177909 526754 177941 526788
rect 177941 526754 177961 526788
rect 177973 526754 177975 526788
rect 177975 526754 178025 526788
rect 178037 526754 178067 526788
rect 178067 526754 178089 526788
rect 181599 526754 181621 526788
rect 181621 526754 181651 526788
rect 181663 526754 181713 526788
rect 181713 526754 181715 526788
rect 181727 526754 181747 526788
rect 181747 526754 181779 526788
rect 177909 526745 177961 526754
rect 177973 526745 178025 526754
rect 178037 526745 178089 526754
rect 181599 526745 181651 526754
rect 181663 526745 181715 526754
rect 181727 526745 181779 526754
rect 181791 526788 181843 526797
rect 181791 526754 181805 526788
rect 181805 526754 181839 526788
rect 181839 526754 181843 526788
rect 181791 526745 181843 526754
rect 181855 526788 181907 526797
rect 185417 526788 185469 526797
rect 181855 526754 181897 526788
rect 181897 526754 181907 526788
rect 185417 526754 185427 526788
rect 185427 526754 185469 526788
rect 181855 526745 181907 526754
rect 185417 526745 185469 526754
rect 185481 526788 185533 526797
rect 185481 526754 185485 526788
rect 185485 526754 185519 526788
rect 185519 526754 185533 526788
rect 185481 526745 185533 526754
rect 185545 526788 185597 526797
rect 185609 526788 185661 526797
rect 185673 526788 185725 526797
rect 185545 526754 185577 526788
rect 185577 526754 185597 526788
rect 185609 526754 185611 526788
rect 185611 526754 185661 526788
rect 185673 526754 185703 526788
rect 185703 526754 185725 526788
rect 185545 526745 185597 526754
rect 185609 526745 185661 526754
rect 185673 526745 185725 526754
rect 174623 526244 174675 526253
rect 174623 526210 174629 526244
rect 174629 526210 174663 526244
rect 174663 526210 174675 526244
rect 174623 526201 174675 526210
rect 174687 526244 174739 526253
rect 174751 526244 174803 526253
rect 174815 526244 174867 526253
rect 174687 526210 174721 526244
rect 174721 526210 174739 526244
rect 174751 526210 174755 526244
rect 174755 526210 174803 526244
rect 174815 526210 174847 526244
rect 174847 526210 174867 526244
rect 174687 526201 174739 526210
rect 174751 526201 174803 526210
rect 174815 526201 174867 526210
rect 174879 526244 174931 526253
rect 174879 526210 174905 526244
rect 174905 526210 174931 526244
rect 174879 526201 174931 526210
rect 178441 526201 178493 526253
rect 178505 526244 178557 526253
rect 178505 526210 178527 526244
rect 178527 526210 178557 526244
rect 178505 526201 178557 526210
rect 178569 526244 178621 526253
rect 178569 526210 178585 526244
rect 178585 526210 178619 526244
rect 178619 526210 178621 526244
rect 178569 526201 178621 526210
rect 178633 526244 178685 526253
rect 178697 526244 178749 526253
rect 182259 526244 182311 526253
rect 178633 526210 178677 526244
rect 178677 526210 178685 526244
rect 178697 526210 178711 526244
rect 178711 526210 178749 526244
rect 182259 526210 182265 526244
rect 182265 526210 182299 526244
rect 182299 526210 182311 526244
rect 178633 526201 178685 526210
rect 178697 526201 178749 526210
rect 182259 526201 182311 526210
rect 182323 526244 182375 526253
rect 182387 526244 182439 526253
rect 182451 526244 182503 526253
rect 182323 526210 182357 526244
rect 182357 526210 182375 526244
rect 182387 526210 182391 526244
rect 182391 526210 182439 526244
rect 182451 526210 182483 526244
rect 182483 526210 182503 526244
rect 182323 526201 182375 526210
rect 182387 526201 182439 526210
rect 182451 526201 182503 526210
rect 182515 526244 182567 526253
rect 182515 526210 182541 526244
rect 182541 526210 182567 526244
rect 182515 526201 182567 526210
rect 186077 526201 186129 526253
rect 186141 526244 186193 526253
rect 186141 526210 186163 526244
rect 186163 526210 186193 526244
rect 186141 526201 186193 526210
rect 186205 526244 186257 526253
rect 186205 526210 186221 526244
rect 186221 526210 186255 526244
rect 186255 526210 186257 526244
rect 186205 526201 186257 526210
rect 186269 526244 186321 526253
rect 186333 526244 186385 526253
rect 186269 526210 186313 526244
rect 186313 526210 186321 526244
rect 186333 526210 186347 526244
rect 186347 526210 186385 526244
rect 186269 526201 186321 526210
rect 186333 526201 186385 526210
rect 173963 525700 174015 525709
rect 174027 525700 174079 525709
rect 174091 525700 174143 525709
rect 173963 525666 173985 525700
rect 173985 525666 174015 525700
rect 174027 525666 174077 525700
rect 174077 525666 174079 525700
rect 174091 525666 174111 525700
rect 174111 525666 174143 525700
rect 173963 525657 174015 525666
rect 174027 525657 174079 525666
rect 174091 525657 174143 525666
rect 174155 525700 174207 525709
rect 174155 525666 174169 525700
rect 174169 525666 174203 525700
rect 174203 525666 174207 525700
rect 174155 525657 174207 525666
rect 174219 525700 174271 525709
rect 177781 525700 177833 525709
rect 174219 525666 174261 525700
rect 174261 525666 174271 525700
rect 177781 525666 177791 525700
rect 177791 525666 177833 525700
rect 174219 525657 174271 525666
rect 177781 525657 177833 525666
rect 177845 525700 177897 525709
rect 177845 525666 177849 525700
rect 177849 525666 177883 525700
rect 177883 525666 177897 525700
rect 177845 525657 177897 525666
rect 177909 525700 177961 525709
rect 177973 525700 178025 525709
rect 178037 525700 178089 525709
rect 181599 525700 181651 525709
rect 181663 525700 181715 525709
rect 181727 525700 181779 525709
rect 177909 525666 177941 525700
rect 177941 525666 177961 525700
rect 177973 525666 177975 525700
rect 177975 525666 178025 525700
rect 178037 525666 178067 525700
rect 178067 525666 178089 525700
rect 181599 525666 181621 525700
rect 181621 525666 181651 525700
rect 181663 525666 181713 525700
rect 181713 525666 181715 525700
rect 181727 525666 181747 525700
rect 181747 525666 181779 525700
rect 177909 525657 177961 525666
rect 177973 525657 178025 525666
rect 178037 525657 178089 525666
rect 181599 525657 181651 525666
rect 181663 525657 181715 525666
rect 181727 525657 181779 525666
rect 181791 525700 181843 525709
rect 181791 525666 181805 525700
rect 181805 525666 181839 525700
rect 181839 525666 181843 525700
rect 181791 525657 181843 525666
rect 181855 525700 181907 525709
rect 185417 525700 185469 525709
rect 181855 525666 181897 525700
rect 181897 525666 181907 525700
rect 185417 525666 185427 525700
rect 185427 525666 185469 525700
rect 181855 525657 181907 525666
rect 185417 525657 185469 525666
rect 185481 525700 185533 525709
rect 185481 525666 185485 525700
rect 185485 525666 185519 525700
rect 185519 525666 185533 525700
rect 185481 525657 185533 525666
rect 185545 525700 185597 525709
rect 185609 525700 185661 525709
rect 185673 525700 185725 525709
rect 185545 525666 185577 525700
rect 185577 525666 185597 525700
rect 185609 525666 185611 525700
rect 185611 525666 185661 525700
rect 185673 525666 185703 525700
rect 185703 525666 185725 525700
rect 185545 525657 185597 525666
rect 185609 525657 185661 525666
rect 185673 525657 185725 525666
rect 174623 525156 174675 525165
rect 174623 525122 174629 525156
rect 174629 525122 174663 525156
rect 174663 525122 174675 525156
rect 174623 525113 174675 525122
rect 174687 525156 174739 525165
rect 174751 525156 174803 525165
rect 174815 525156 174867 525165
rect 174687 525122 174721 525156
rect 174721 525122 174739 525156
rect 174751 525122 174755 525156
rect 174755 525122 174803 525156
rect 174815 525122 174847 525156
rect 174847 525122 174867 525156
rect 174687 525113 174739 525122
rect 174751 525113 174803 525122
rect 174815 525113 174867 525122
rect 174879 525156 174931 525165
rect 174879 525122 174905 525156
rect 174905 525122 174931 525156
rect 174879 525113 174931 525122
rect 178441 525113 178493 525165
rect 178505 525156 178557 525165
rect 178505 525122 178527 525156
rect 178527 525122 178557 525156
rect 178505 525113 178557 525122
rect 178569 525156 178621 525165
rect 178569 525122 178585 525156
rect 178585 525122 178619 525156
rect 178619 525122 178621 525156
rect 178569 525113 178621 525122
rect 178633 525156 178685 525165
rect 178697 525156 178749 525165
rect 182259 525156 182311 525165
rect 178633 525122 178677 525156
rect 178677 525122 178685 525156
rect 178697 525122 178711 525156
rect 178711 525122 178749 525156
rect 182259 525122 182265 525156
rect 182265 525122 182299 525156
rect 182299 525122 182311 525156
rect 178633 525113 178685 525122
rect 178697 525113 178749 525122
rect 182259 525113 182311 525122
rect 182323 525156 182375 525165
rect 182387 525156 182439 525165
rect 182451 525156 182503 525165
rect 182323 525122 182357 525156
rect 182357 525122 182375 525156
rect 182387 525122 182391 525156
rect 182391 525122 182439 525156
rect 182451 525122 182483 525156
rect 182483 525122 182503 525156
rect 182323 525113 182375 525122
rect 182387 525113 182439 525122
rect 182451 525113 182503 525122
rect 182515 525156 182567 525165
rect 182515 525122 182541 525156
rect 182541 525122 182567 525156
rect 182515 525113 182567 525122
rect 186077 525113 186129 525165
rect 186141 525156 186193 525165
rect 186141 525122 186163 525156
rect 186163 525122 186193 525156
rect 186141 525113 186193 525122
rect 186205 525156 186257 525165
rect 186205 525122 186221 525156
rect 186221 525122 186255 525156
rect 186255 525122 186257 525156
rect 186205 525113 186257 525122
rect 186269 525156 186321 525165
rect 186333 525156 186385 525165
rect 186269 525122 186313 525156
rect 186313 525122 186321 525156
rect 186333 525122 186347 525156
rect 186347 525122 186385 525156
rect 186269 525113 186321 525122
rect 186333 525113 186385 525122
rect 173963 524612 174015 524621
rect 174027 524612 174079 524621
rect 174091 524612 174143 524621
rect 173963 524578 173985 524612
rect 173985 524578 174015 524612
rect 174027 524578 174077 524612
rect 174077 524578 174079 524612
rect 174091 524578 174111 524612
rect 174111 524578 174143 524612
rect 173963 524569 174015 524578
rect 174027 524569 174079 524578
rect 174091 524569 174143 524578
rect 174155 524612 174207 524621
rect 174155 524578 174169 524612
rect 174169 524578 174203 524612
rect 174203 524578 174207 524612
rect 174155 524569 174207 524578
rect 174219 524612 174271 524621
rect 177781 524612 177833 524621
rect 174219 524578 174261 524612
rect 174261 524578 174271 524612
rect 177781 524578 177791 524612
rect 177791 524578 177833 524612
rect 174219 524569 174271 524578
rect 177781 524569 177833 524578
rect 177845 524612 177897 524621
rect 177845 524578 177849 524612
rect 177849 524578 177883 524612
rect 177883 524578 177897 524612
rect 177845 524569 177897 524578
rect 177909 524612 177961 524621
rect 177973 524612 178025 524621
rect 178037 524612 178089 524621
rect 181599 524612 181651 524621
rect 181663 524612 181715 524621
rect 181727 524612 181779 524621
rect 177909 524578 177941 524612
rect 177941 524578 177961 524612
rect 177973 524578 177975 524612
rect 177975 524578 178025 524612
rect 178037 524578 178067 524612
rect 178067 524578 178089 524612
rect 181599 524578 181621 524612
rect 181621 524578 181651 524612
rect 181663 524578 181713 524612
rect 181713 524578 181715 524612
rect 181727 524578 181747 524612
rect 181747 524578 181779 524612
rect 177909 524569 177961 524578
rect 177973 524569 178025 524578
rect 178037 524569 178089 524578
rect 181599 524569 181651 524578
rect 181663 524569 181715 524578
rect 181727 524569 181779 524578
rect 181791 524612 181843 524621
rect 181791 524578 181805 524612
rect 181805 524578 181839 524612
rect 181839 524578 181843 524612
rect 181791 524569 181843 524578
rect 181855 524612 181907 524621
rect 185417 524612 185469 524621
rect 181855 524578 181897 524612
rect 181897 524578 181907 524612
rect 185417 524578 185427 524612
rect 185427 524578 185469 524612
rect 181855 524569 181907 524578
rect 185417 524569 185469 524578
rect 185481 524612 185533 524621
rect 185481 524578 185485 524612
rect 185485 524578 185519 524612
rect 185519 524578 185533 524612
rect 185481 524569 185533 524578
rect 185545 524612 185597 524621
rect 185609 524612 185661 524621
rect 185673 524612 185725 524621
rect 185545 524578 185577 524612
rect 185577 524578 185597 524612
rect 185609 524578 185611 524612
rect 185611 524578 185661 524612
rect 185673 524578 185703 524612
rect 185703 524578 185725 524612
rect 185545 524569 185597 524578
rect 185609 524569 185661 524578
rect 185673 524569 185725 524578
rect 174623 524068 174675 524077
rect 174623 524034 174629 524068
rect 174629 524034 174663 524068
rect 174663 524034 174675 524068
rect 174623 524025 174675 524034
rect 174687 524068 174739 524077
rect 174751 524068 174803 524077
rect 174815 524068 174867 524077
rect 174687 524034 174721 524068
rect 174721 524034 174739 524068
rect 174751 524034 174755 524068
rect 174755 524034 174803 524068
rect 174815 524034 174847 524068
rect 174847 524034 174867 524068
rect 174687 524025 174739 524034
rect 174751 524025 174803 524034
rect 174815 524025 174867 524034
rect 174879 524068 174931 524077
rect 174879 524034 174905 524068
rect 174905 524034 174931 524068
rect 174879 524025 174931 524034
rect 178441 524025 178493 524077
rect 178505 524068 178557 524077
rect 178505 524034 178527 524068
rect 178527 524034 178557 524068
rect 178505 524025 178557 524034
rect 178569 524068 178621 524077
rect 178569 524034 178585 524068
rect 178585 524034 178619 524068
rect 178619 524034 178621 524068
rect 178569 524025 178621 524034
rect 178633 524068 178685 524077
rect 178697 524068 178749 524077
rect 182259 524068 182311 524077
rect 178633 524034 178677 524068
rect 178677 524034 178685 524068
rect 178697 524034 178711 524068
rect 178711 524034 178749 524068
rect 182259 524034 182265 524068
rect 182265 524034 182299 524068
rect 182299 524034 182311 524068
rect 178633 524025 178685 524034
rect 178697 524025 178749 524034
rect 182259 524025 182311 524034
rect 182323 524068 182375 524077
rect 182387 524068 182439 524077
rect 182451 524068 182503 524077
rect 182323 524034 182357 524068
rect 182357 524034 182375 524068
rect 182387 524034 182391 524068
rect 182391 524034 182439 524068
rect 182451 524034 182483 524068
rect 182483 524034 182503 524068
rect 182323 524025 182375 524034
rect 182387 524025 182439 524034
rect 182451 524025 182503 524034
rect 182515 524068 182567 524077
rect 182515 524034 182541 524068
rect 182541 524034 182567 524068
rect 182515 524025 182567 524034
rect 186077 524025 186129 524077
rect 186141 524068 186193 524077
rect 186141 524034 186163 524068
rect 186163 524034 186193 524068
rect 186141 524025 186193 524034
rect 186205 524068 186257 524077
rect 186205 524034 186221 524068
rect 186221 524034 186255 524068
rect 186255 524034 186257 524068
rect 186205 524025 186257 524034
rect 186269 524068 186321 524077
rect 186333 524068 186385 524077
rect 186269 524034 186313 524068
rect 186313 524034 186321 524068
rect 186333 524034 186347 524068
rect 186347 524034 186385 524068
rect 186269 524025 186321 524034
rect 186333 524025 186385 524034
rect 173963 523524 174015 523533
rect 174027 523524 174079 523533
rect 174091 523524 174143 523533
rect 173963 523490 173985 523524
rect 173985 523490 174015 523524
rect 174027 523490 174077 523524
rect 174077 523490 174079 523524
rect 174091 523490 174111 523524
rect 174111 523490 174143 523524
rect 173963 523481 174015 523490
rect 174027 523481 174079 523490
rect 174091 523481 174143 523490
rect 174155 523524 174207 523533
rect 174155 523490 174169 523524
rect 174169 523490 174203 523524
rect 174203 523490 174207 523524
rect 174155 523481 174207 523490
rect 174219 523524 174271 523533
rect 177781 523524 177833 523533
rect 174219 523490 174261 523524
rect 174261 523490 174271 523524
rect 177781 523490 177791 523524
rect 177791 523490 177833 523524
rect 174219 523481 174271 523490
rect 177781 523481 177833 523490
rect 177845 523524 177897 523533
rect 177845 523490 177849 523524
rect 177849 523490 177883 523524
rect 177883 523490 177897 523524
rect 177845 523481 177897 523490
rect 177909 523524 177961 523533
rect 177973 523524 178025 523533
rect 178037 523524 178089 523533
rect 181599 523524 181651 523533
rect 181663 523524 181715 523533
rect 181727 523524 181779 523533
rect 177909 523490 177941 523524
rect 177941 523490 177961 523524
rect 177973 523490 177975 523524
rect 177975 523490 178025 523524
rect 178037 523490 178067 523524
rect 178067 523490 178089 523524
rect 181599 523490 181621 523524
rect 181621 523490 181651 523524
rect 181663 523490 181713 523524
rect 181713 523490 181715 523524
rect 181727 523490 181747 523524
rect 181747 523490 181779 523524
rect 177909 523481 177961 523490
rect 177973 523481 178025 523490
rect 178037 523481 178089 523490
rect 181599 523481 181651 523490
rect 181663 523481 181715 523490
rect 181727 523481 181779 523490
rect 181791 523524 181843 523533
rect 181791 523490 181805 523524
rect 181805 523490 181839 523524
rect 181839 523490 181843 523524
rect 181791 523481 181843 523490
rect 181855 523524 181907 523533
rect 185417 523524 185469 523533
rect 181855 523490 181897 523524
rect 181897 523490 181907 523524
rect 185417 523490 185427 523524
rect 185427 523490 185469 523524
rect 181855 523481 181907 523490
rect 185417 523481 185469 523490
rect 185481 523524 185533 523533
rect 185481 523490 185485 523524
rect 185485 523490 185519 523524
rect 185519 523490 185533 523524
rect 185481 523481 185533 523490
rect 185545 523524 185597 523533
rect 185609 523524 185661 523533
rect 185673 523524 185725 523533
rect 185545 523490 185577 523524
rect 185577 523490 185597 523524
rect 185609 523490 185611 523524
rect 185611 523490 185661 523524
rect 185673 523490 185703 523524
rect 185703 523490 185725 523524
rect 185545 523481 185597 523490
rect 185609 523481 185661 523490
rect 185673 523481 185725 523490
rect 174623 522980 174675 522989
rect 174623 522946 174629 522980
rect 174629 522946 174663 522980
rect 174663 522946 174675 522980
rect 174623 522937 174675 522946
rect 174687 522980 174739 522989
rect 174751 522980 174803 522989
rect 174815 522980 174867 522989
rect 174687 522946 174721 522980
rect 174721 522946 174739 522980
rect 174751 522946 174755 522980
rect 174755 522946 174803 522980
rect 174815 522946 174847 522980
rect 174847 522946 174867 522980
rect 174687 522937 174739 522946
rect 174751 522937 174803 522946
rect 174815 522937 174867 522946
rect 174879 522980 174931 522989
rect 174879 522946 174905 522980
rect 174905 522946 174931 522980
rect 174879 522937 174931 522946
rect 178441 522937 178493 522989
rect 178505 522980 178557 522989
rect 178505 522946 178527 522980
rect 178527 522946 178557 522980
rect 178505 522937 178557 522946
rect 178569 522980 178621 522989
rect 178569 522946 178585 522980
rect 178585 522946 178619 522980
rect 178619 522946 178621 522980
rect 178569 522937 178621 522946
rect 178633 522980 178685 522989
rect 178697 522980 178749 522989
rect 182259 522980 182311 522989
rect 178633 522946 178677 522980
rect 178677 522946 178685 522980
rect 178697 522946 178711 522980
rect 178711 522946 178749 522980
rect 182259 522946 182265 522980
rect 182265 522946 182299 522980
rect 182299 522946 182311 522980
rect 178633 522937 178685 522946
rect 178697 522937 178749 522946
rect 182259 522937 182311 522946
rect 182323 522980 182375 522989
rect 182387 522980 182439 522989
rect 182451 522980 182503 522989
rect 182323 522946 182357 522980
rect 182357 522946 182375 522980
rect 182387 522946 182391 522980
rect 182391 522946 182439 522980
rect 182451 522946 182483 522980
rect 182483 522946 182503 522980
rect 182323 522937 182375 522946
rect 182387 522937 182439 522946
rect 182451 522937 182503 522946
rect 182515 522980 182567 522989
rect 182515 522946 182541 522980
rect 182541 522946 182567 522980
rect 182515 522937 182567 522946
rect 186077 522937 186129 522989
rect 186141 522980 186193 522989
rect 186141 522946 186163 522980
rect 186163 522946 186193 522980
rect 186141 522937 186193 522946
rect 186205 522980 186257 522989
rect 186205 522946 186221 522980
rect 186221 522946 186255 522980
rect 186255 522946 186257 522980
rect 186205 522937 186257 522946
rect 186269 522980 186321 522989
rect 186333 522980 186385 522989
rect 186269 522946 186313 522980
rect 186313 522946 186321 522980
rect 186333 522946 186347 522980
rect 186347 522946 186385 522980
rect 186269 522937 186321 522946
rect 186333 522937 186385 522946
rect 173963 522436 174015 522445
rect 174027 522436 174079 522445
rect 174091 522436 174143 522445
rect 173963 522402 173985 522436
rect 173985 522402 174015 522436
rect 174027 522402 174077 522436
rect 174077 522402 174079 522436
rect 174091 522402 174111 522436
rect 174111 522402 174143 522436
rect 173963 522393 174015 522402
rect 174027 522393 174079 522402
rect 174091 522393 174143 522402
rect 174155 522436 174207 522445
rect 174155 522402 174169 522436
rect 174169 522402 174203 522436
rect 174203 522402 174207 522436
rect 174155 522393 174207 522402
rect 174219 522436 174271 522445
rect 177781 522436 177833 522445
rect 174219 522402 174261 522436
rect 174261 522402 174271 522436
rect 177781 522402 177791 522436
rect 177791 522402 177833 522436
rect 174219 522393 174271 522402
rect 177781 522393 177833 522402
rect 177845 522436 177897 522445
rect 177845 522402 177849 522436
rect 177849 522402 177883 522436
rect 177883 522402 177897 522436
rect 177845 522393 177897 522402
rect 177909 522436 177961 522445
rect 177973 522436 178025 522445
rect 178037 522436 178089 522445
rect 181599 522436 181651 522445
rect 181663 522436 181715 522445
rect 181727 522436 181779 522445
rect 177909 522402 177941 522436
rect 177941 522402 177961 522436
rect 177973 522402 177975 522436
rect 177975 522402 178025 522436
rect 178037 522402 178067 522436
rect 178067 522402 178089 522436
rect 181599 522402 181621 522436
rect 181621 522402 181651 522436
rect 181663 522402 181713 522436
rect 181713 522402 181715 522436
rect 181727 522402 181747 522436
rect 181747 522402 181779 522436
rect 177909 522393 177961 522402
rect 177973 522393 178025 522402
rect 178037 522393 178089 522402
rect 181599 522393 181651 522402
rect 181663 522393 181715 522402
rect 181727 522393 181779 522402
rect 181791 522436 181843 522445
rect 181791 522402 181805 522436
rect 181805 522402 181839 522436
rect 181839 522402 181843 522436
rect 181791 522393 181843 522402
rect 181855 522436 181907 522445
rect 185417 522436 185469 522445
rect 181855 522402 181897 522436
rect 181897 522402 181907 522436
rect 185417 522402 185427 522436
rect 185427 522402 185469 522436
rect 181855 522393 181907 522402
rect 185417 522393 185469 522402
rect 185481 522436 185533 522445
rect 185481 522402 185485 522436
rect 185485 522402 185519 522436
rect 185519 522402 185533 522436
rect 185481 522393 185533 522402
rect 185545 522436 185597 522445
rect 185609 522436 185661 522445
rect 185673 522436 185725 522445
rect 185545 522402 185577 522436
rect 185577 522402 185597 522436
rect 185609 522402 185611 522436
rect 185611 522402 185661 522436
rect 185673 522402 185703 522436
rect 185703 522402 185725 522436
rect 185545 522393 185597 522402
rect 185609 522393 185661 522402
rect 185673 522393 185725 522402
rect 174623 521892 174675 521901
rect 174623 521858 174629 521892
rect 174629 521858 174663 521892
rect 174663 521858 174675 521892
rect 174623 521849 174675 521858
rect 174687 521892 174739 521901
rect 174751 521892 174803 521901
rect 174815 521892 174867 521901
rect 174687 521858 174721 521892
rect 174721 521858 174739 521892
rect 174751 521858 174755 521892
rect 174755 521858 174803 521892
rect 174815 521858 174847 521892
rect 174847 521858 174867 521892
rect 174687 521849 174739 521858
rect 174751 521849 174803 521858
rect 174815 521849 174867 521858
rect 174879 521892 174931 521901
rect 174879 521858 174905 521892
rect 174905 521858 174931 521892
rect 174879 521849 174931 521858
rect 178441 521849 178493 521901
rect 178505 521892 178557 521901
rect 178505 521858 178527 521892
rect 178527 521858 178557 521892
rect 178505 521849 178557 521858
rect 178569 521892 178621 521901
rect 178569 521858 178585 521892
rect 178585 521858 178619 521892
rect 178619 521858 178621 521892
rect 178569 521849 178621 521858
rect 178633 521892 178685 521901
rect 178697 521892 178749 521901
rect 182259 521892 182311 521901
rect 178633 521858 178677 521892
rect 178677 521858 178685 521892
rect 178697 521858 178711 521892
rect 178711 521858 178749 521892
rect 182259 521858 182265 521892
rect 182265 521858 182299 521892
rect 182299 521858 182311 521892
rect 178633 521849 178685 521858
rect 178697 521849 178749 521858
rect 182259 521849 182311 521858
rect 182323 521892 182375 521901
rect 182387 521892 182439 521901
rect 182451 521892 182503 521901
rect 182323 521858 182357 521892
rect 182357 521858 182375 521892
rect 182387 521858 182391 521892
rect 182391 521858 182439 521892
rect 182451 521858 182483 521892
rect 182483 521858 182503 521892
rect 182323 521849 182375 521858
rect 182387 521849 182439 521858
rect 182451 521849 182503 521858
rect 182515 521892 182567 521901
rect 182515 521858 182541 521892
rect 182541 521858 182567 521892
rect 182515 521849 182567 521858
rect 186077 521849 186129 521901
rect 186141 521892 186193 521901
rect 186141 521858 186163 521892
rect 186163 521858 186193 521892
rect 186141 521849 186193 521858
rect 186205 521892 186257 521901
rect 186205 521858 186221 521892
rect 186221 521858 186255 521892
rect 186255 521858 186257 521892
rect 186205 521849 186257 521858
rect 186269 521892 186321 521901
rect 186333 521892 186385 521901
rect 186269 521858 186313 521892
rect 186313 521858 186321 521892
rect 186333 521858 186347 521892
rect 186347 521858 186385 521892
rect 186269 521849 186321 521858
rect 186333 521849 186385 521858
rect 173963 521348 174015 521357
rect 174027 521348 174079 521357
rect 174091 521348 174143 521357
rect 173963 521314 173985 521348
rect 173985 521314 174015 521348
rect 174027 521314 174077 521348
rect 174077 521314 174079 521348
rect 174091 521314 174111 521348
rect 174111 521314 174143 521348
rect 173963 521305 174015 521314
rect 174027 521305 174079 521314
rect 174091 521305 174143 521314
rect 174155 521348 174207 521357
rect 174155 521314 174169 521348
rect 174169 521314 174203 521348
rect 174203 521314 174207 521348
rect 174155 521305 174207 521314
rect 174219 521348 174271 521357
rect 177781 521348 177833 521357
rect 174219 521314 174261 521348
rect 174261 521314 174271 521348
rect 177781 521314 177791 521348
rect 177791 521314 177833 521348
rect 174219 521305 174271 521314
rect 177781 521305 177833 521314
rect 177845 521348 177897 521357
rect 177845 521314 177849 521348
rect 177849 521314 177883 521348
rect 177883 521314 177897 521348
rect 177845 521305 177897 521314
rect 177909 521348 177961 521357
rect 177973 521348 178025 521357
rect 178037 521348 178089 521357
rect 181599 521348 181651 521357
rect 181663 521348 181715 521357
rect 181727 521348 181779 521357
rect 177909 521314 177941 521348
rect 177941 521314 177961 521348
rect 177973 521314 177975 521348
rect 177975 521314 178025 521348
rect 178037 521314 178067 521348
rect 178067 521314 178089 521348
rect 181599 521314 181621 521348
rect 181621 521314 181651 521348
rect 181663 521314 181713 521348
rect 181713 521314 181715 521348
rect 181727 521314 181747 521348
rect 181747 521314 181779 521348
rect 177909 521305 177961 521314
rect 177973 521305 178025 521314
rect 178037 521305 178089 521314
rect 181599 521305 181651 521314
rect 181663 521305 181715 521314
rect 181727 521305 181779 521314
rect 181791 521348 181843 521357
rect 181791 521314 181805 521348
rect 181805 521314 181839 521348
rect 181839 521314 181843 521348
rect 181791 521305 181843 521314
rect 181855 521348 181907 521357
rect 185417 521348 185469 521357
rect 181855 521314 181897 521348
rect 181897 521314 181907 521348
rect 185417 521314 185427 521348
rect 185427 521314 185469 521348
rect 181855 521305 181907 521314
rect 185417 521305 185469 521314
rect 185481 521348 185533 521357
rect 185481 521314 185485 521348
rect 185485 521314 185519 521348
rect 185519 521314 185533 521348
rect 185481 521305 185533 521314
rect 185545 521348 185597 521357
rect 185609 521348 185661 521357
rect 185673 521348 185725 521357
rect 185545 521314 185577 521348
rect 185577 521314 185597 521348
rect 185609 521314 185611 521348
rect 185611 521314 185661 521348
rect 185673 521314 185703 521348
rect 185703 521314 185725 521348
rect 185545 521305 185597 521314
rect 185609 521305 185661 521314
rect 185673 521305 185725 521314
rect 174623 520804 174675 520813
rect 174623 520770 174629 520804
rect 174629 520770 174663 520804
rect 174663 520770 174675 520804
rect 174623 520761 174675 520770
rect 174687 520804 174739 520813
rect 174751 520804 174803 520813
rect 174815 520804 174867 520813
rect 174687 520770 174721 520804
rect 174721 520770 174739 520804
rect 174751 520770 174755 520804
rect 174755 520770 174803 520804
rect 174815 520770 174847 520804
rect 174847 520770 174867 520804
rect 174687 520761 174739 520770
rect 174751 520761 174803 520770
rect 174815 520761 174867 520770
rect 174879 520804 174931 520813
rect 174879 520770 174905 520804
rect 174905 520770 174931 520804
rect 174879 520761 174931 520770
rect 178441 520761 178493 520813
rect 178505 520804 178557 520813
rect 178505 520770 178527 520804
rect 178527 520770 178557 520804
rect 178505 520761 178557 520770
rect 178569 520804 178621 520813
rect 178569 520770 178585 520804
rect 178585 520770 178619 520804
rect 178619 520770 178621 520804
rect 178569 520761 178621 520770
rect 178633 520804 178685 520813
rect 178697 520804 178749 520813
rect 182259 520804 182311 520813
rect 178633 520770 178677 520804
rect 178677 520770 178685 520804
rect 178697 520770 178711 520804
rect 178711 520770 178749 520804
rect 182259 520770 182265 520804
rect 182265 520770 182299 520804
rect 182299 520770 182311 520804
rect 178633 520761 178685 520770
rect 178697 520761 178749 520770
rect 182259 520761 182311 520770
rect 182323 520804 182375 520813
rect 182387 520804 182439 520813
rect 182451 520804 182503 520813
rect 182323 520770 182357 520804
rect 182357 520770 182375 520804
rect 182387 520770 182391 520804
rect 182391 520770 182439 520804
rect 182451 520770 182483 520804
rect 182483 520770 182503 520804
rect 182323 520761 182375 520770
rect 182387 520761 182439 520770
rect 182451 520761 182503 520770
rect 182515 520804 182567 520813
rect 182515 520770 182541 520804
rect 182541 520770 182567 520804
rect 182515 520761 182567 520770
rect 186077 520761 186129 520813
rect 186141 520804 186193 520813
rect 186141 520770 186163 520804
rect 186163 520770 186193 520804
rect 186141 520761 186193 520770
rect 186205 520804 186257 520813
rect 186205 520770 186221 520804
rect 186221 520770 186255 520804
rect 186255 520770 186257 520804
rect 186205 520761 186257 520770
rect 186269 520804 186321 520813
rect 186333 520804 186385 520813
rect 186269 520770 186313 520804
rect 186313 520770 186321 520804
rect 186333 520770 186347 520804
rect 186347 520770 186385 520804
rect 186269 520761 186321 520770
rect 186333 520761 186385 520770
rect 173963 520260 174015 520269
rect 174027 520260 174079 520269
rect 174091 520260 174143 520269
rect 173963 520226 173985 520260
rect 173985 520226 174015 520260
rect 174027 520226 174077 520260
rect 174077 520226 174079 520260
rect 174091 520226 174111 520260
rect 174111 520226 174143 520260
rect 173963 520217 174015 520226
rect 174027 520217 174079 520226
rect 174091 520217 174143 520226
rect 174155 520260 174207 520269
rect 174155 520226 174169 520260
rect 174169 520226 174203 520260
rect 174203 520226 174207 520260
rect 174155 520217 174207 520226
rect 174219 520260 174271 520269
rect 177781 520260 177833 520269
rect 174219 520226 174261 520260
rect 174261 520226 174271 520260
rect 177781 520226 177791 520260
rect 177791 520226 177833 520260
rect 174219 520217 174271 520226
rect 177781 520217 177833 520226
rect 177845 520260 177897 520269
rect 177845 520226 177849 520260
rect 177849 520226 177883 520260
rect 177883 520226 177897 520260
rect 177845 520217 177897 520226
rect 177909 520260 177961 520269
rect 177973 520260 178025 520269
rect 178037 520260 178089 520269
rect 181599 520260 181651 520269
rect 181663 520260 181715 520269
rect 181727 520260 181779 520269
rect 177909 520226 177941 520260
rect 177941 520226 177961 520260
rect 177973 520226 177975 520260
rect 177975 520226 178025 520260
rect 178037 520226 178067 520260
rect 178067 520226 178089 520260
rect 181599 520226 181621 520260
rect 181621 520226 181651 520260
rect 181663 520226 181713 520260
rect 181713 520226 181715 520260
rect 181727 520226 181747 520260
rect 181747 520226 181779 520260
rect 177909 520217 177961 520226
rect 177973 520217 178025 520226
rect 178037 520217 178089 520226
rect 181599 520217 181651 520226
rect 181663 520217 181715 520226
rect 181727 520217 181779 520226
rect 181791 520260 181843 520269
rect 181791 520226 181805 520260
rect 181805 520226 181839 520260
rect 181839 520226 181843 520260
rect 181791 520217 181843 520226
rect 181855 520260 181907 520269
rect 185417 520260 185469 520269
rect 181855 520226 181897 520260
rect 181897 520226 181907 520260
rect 185417 520226 185427 520260
rect 185427 520226 185469 520260
rect 181855 520217 181907 520226
rect 185417 520217 185469 520226
rect 185481 520260 185533 520269
rect 185481 520226 185485 520260
rect 185485 520226 185519 520260
rect 185519 520226 185533 520260
rect 185481 520217 185533 520226
rect 185545 520260 185597 520269
rect 185609 520260 185661 520269
rect 185673 520260 185725 520269
rect 185545 520226 185577 520260
rect 185577 520226 185597 520260
rect 185609 520226 185611 520260
rect 185611 520226 185661 520260
rect 185673 520226 185703 520260
rect 185703 520226 185725 520260
rect 185545 520217 185597 520226
rect 185609 520217 185661 520226
rect 185673 520217 185725 520226
rect 174623 519716 174675 519725
rect 174623 519682 174629 519716
rect 174629 519682 174663 519716
rect 174663 519682 174675 519716
rect 174623 519673 174675 519682
rect 174687 519716 174739 519725
rect 174751 519716 174803 519725
rect 174815 519716 174867 519725
rect 174687 519682 174721 519716
rect 174721 519682 174739 519716
rect 174751 519682 174755 519716
rect 174755 519682 174803 519716
rect 174815 519682 174847 519716
rect 174847 519682 174867 519716
rect 174687 519673 174739 519682
rect 174751 519673 174803 519682
rect 174815 519673 174867 519682
rect 174879 519716 174931 519725
rect 174879 519682 174905 519716
rect 174905 519682 174931 519716
rect 174879 519673 174931 519682
rect 178441 519673 178493 519725
rect 178505 519716 178557 519725
rect 178505 519682 178527 519716
rect 178527 519682 178557 519716
rect 178505 519673 178557 519682
rect 178569 519716 178621 519725
rect 178569 519682 178585 519716
rect 178585 519682 178619 519716
rect 178619 519682 178621 519716
rect 178569 519673 178621 519682
rect 178633 519716 178685 519725
rect 178697 519716 178749 519725
rect 182259 519716 182311 519725
rect 178633 519682 178677 519716
rect 178677 519682 178685 519716
rect 178697 519682 178711 519716
rect 178711 519682 178749 519716
rect 182259 519682 182265 519716
rect 182265 519682 182299 519716
rect 182299 519682 182311 519716
rect 178633 519673 178685 519682
rect 178697 519673 178749 519682
rect 182259 519673 182311 519682
rect 182323 519716 182375 519725
rect 182387 519716 182439 519725
rect 182451 519716 182503 519725
rect 182323 519682 182357 519716
rect 182357 519682 182375 519716
rect 182387 519682 182391 519716
rect 182391 519682 182439 519716
rect 182451 519682 182483 519716
rect 182483 519682 182503 519716
rect 182323 519673 182375 519682
rect 182387 519673 182439 519682
rect 182451 519673 182503 519682
rect 182515 519716 182567 519725
rect 182515 519682 182541 519716
rect 182541 519682 182567 519716
rect 182515 519673 182567 519682
rect 186077 519673 186129 519725
rect 186141 519716 186193 519725
rect 186141 519682 186163 519716
rect 186163 519682 186193 519716
rect 186141 519673 186193 519682
rect 186205 519716 186257 519725
rect 186205 519682 186221 519716
rect 186221 519682 186255 519716
rect 186255 519682 186257 519716
rect 186205 519673 186257 519682
rect 186269 519716 186321 519725
rect 186333 519716 186385 519725
rect 186269 519682 186313 519716
rect 186313 519682 186321 519716
rect 186333 519682 186347 519716
rect 186347 519682 186385 519716
rect 186269 519673 186321 519682
rect 186333 519673 186385 519682
rect 173963 519172 174015 519181
rect 174027 519172 174079 519181
rect 174091 519172 174143 519181
rect 173963 519138 173985 519172
rect 173985 519138 174015 519172
rect 174027 519138 174077 519172
rect 174077 519138 174079 519172
rect 174091 519138 174111 519172
rect 174111 519138 174143 519172
rect 173963 519129 174015 519138
rect 174027 519129 174079 519138
rect 174091 519129 174143 519138
rect 174155 519172 174207 519181
rect 174155 519138 174169 519172
rect 174169 519138 174203 519172
rect 174203 519138 174207 519172
rect 174155 519129 174207 519138
rect 174219 519172 174271 519181
rect 177781 519172 177833 519181
rect 174219 519138 174261 519172
rect 174261 519138 174271 519172
rect 177781 519138 177791 519172
rect 177791 519138 177833 519172
rect 174219 519129 174271 519138
rect 177781 519129 177833 519138
rect 177845 519172 177897 519181
rect 177845 519138 177849 519172
rect 177849 519138 177883 519172
rect 177883 519138 177897 519172
rect 177845 519129 177897 519138
rect 177909 519172 177961 519181
rect 177973 519172 178025 519181
rect 178037 519172 178089 519181
rect 181599 519172 181651 519181
rect 181663 519172 181715 519181
rect 181727 519172 181779 519181
rect 177909 519138 177941 519172
rect 177941 519138 177961 519172
rect 177973 519138 177975 519172
rect 177975 519138 178025 519172
rect 178037 519138 178067 519172
rect 178067 519138 178089 519172
rect 181599 519138 181621 519172
rect 181621 519138 181651 519172
rect 181663 519138 181713 519172
rect 181713 519138 181715 519172
rect 181727 519138 181747 519172
rect 181747 519138 181779 519172
rect 177909 519129 177961 519138
rect 177973 519129 178025 519138
rect 178037 519129 178089 519138
rect 181599 519129 181651 519138
rect 181663 519129 181715 519138
rect 181727 519129 181779 519138
rect 181791 519172 181843 519181
rect 181791 519138 181805 519172
rect 181805 519138 181839 519172
rect 181839 519138 181843 519172
rect 181791 519129 181843 519138
rect 181855 519172 181907 519181
rect 185417 519172 185469 519181
rect 181855 519138 181897 519172
rect 181897 519138 181907 519172
rect 185417 519138 185427 519172
rect 185427 519138 185469 519172
rect 181855 519129 181907 519138
rect 185417 519129 185469 519138
rect 185481 519172 185533 519181
rect 185481 519138 185485 519172
rect 185485 519138 185519 519172
rect 185519 519138 185533 519172
rect 185481 519129 185533 519138
rect 185545 519172 185597 519181
rect 185609 519172 185661 519181
rect 185673 519172 185725 519181
rect 185545 519138 185577 519172
rect 185577 519138 185597 519172
rect 185609 519138 185611 519172
rect 185611 519138 185661 519172
rect 185673 519138 185703 519172
rect 185703 519138 185725 519172
rect 185545 519129 185597 519138
rect 185609 519129 185661 519138
rect 185673 519129 185725 519138
rect 174623 518628 174675 518637
rect 174623 518594 174629 518628
rect 174629 518594 174663 518628
rect 174663 518594 174675 518628
rect 174623 518585 174675 518594
rect 174687 518628 174739 518637
rect 174751 518628 174803 518637
rect 174815 518628 174867 518637
rect 174687 518594 174721 518628
rect 174721 518594 174739 518628
rect 174751 518594 174755 518628
rect 174755 518594 174803 518628
rect 174815 518594 174847 518628
rect 174847 518594 174867 518628
rect 174687 518585 174739 518594
rect 174751 518585 174803 518594
rect 174815 518585 174867 518594
rect 174879 518628 174931 518637
rect 174879 518594 174905 518628
rect 174905 518594 174931 518628
rect 174879 518585 174931 518594
rect 178441 518585 178493 518637
rect 178505 518628 178557 518637
rect 178505 518594 178527 518628
rect 178527 518594 178557 518628
rect 178505 518585 178557 518594
rect 178569 518628 178621 518637
rect 178569 518594 178585 518628
rect 178585 518594 178619 518628
rect 178619 518594 178621 518628
rect 178569 518585 178621 518594
rect 178633 518628 178685 518637
rect 178697 518628 178749 518637
rect 182259 518628 182311 518637
rect 178633 518594 178677 518628
rect 178677 518594 178685 518628
rect 178697 518594 178711 518628
rect 178711 518594 178749 518628
rect 182259 518594 182265 518628
rect 182265 518594 182299 518628
rect 182299 518594 182311 518628
rect 178633 518585 178685 518594
rect 178697 518585 178749 518594
rect 182259 518585 182311 518594
rect 182323 518628 182375 518637
rect 182387 518628 182439 518637
rect 182451 518628 182503 518637
rect 182323 518594 182357 518628
rect 182357 518594 182375 518628
rect 182387 518594 182391 518628
rect 182391 518594 182439 518628
rect 182451 518594 182483 518628
rect 182483 518594 182503 518628
rect 182323 518585 182375 518594
rect 182387 518585 182439 518594
rect 182451 518585 182503 518594
rect 182515 518628 182567 518637
rect 182515 518594 182541 518628
rect 182541 518594 182567 518628
rect 182515 518585 182567 518594
rect 186077 518585 186129 518637
rect 186141 518628 186193 518637
rect 186141 518594 186163 518628
rect 186163 518594 186193 518628
rect 186141 518585 186193 518594
rect 186205 518628 186257 518637
rect 186205 518594 186221 518628
rect 186221 518594 186255 518628
rect 186255 518594 186257 518628
rect 186205 518585 186257 518594
rect 186269 518628 186321 518637
rect 186333 518628 186385 518637
rect 186269 518594 186313 518628
rect 186313 518594 186321 518628
rect 186333 518594 186347 518628
rect 186347 518594 186385 518628
rect 186269 518585 186321 518594
rect 186333 518585 186385 518594
rect 173963 518084 174015 518093
rect 174027 518084 174079 518093
rect 174091 518084 174143 518093
rect 173963 518050 173985 518084
rect 173985 518050 174015 518084
rect 174027 518050 174077 518084
rect 174077 518050 174079 518084
rect 174091 518050 174111 518084
rect 174111 518050 174143 518084
rect 173963 518041 174015 518050
rect 174027 518041 174079 518050
rect 174091 518041 174143 518050
rect 174155 518084 174207 518093
rect 174155 518050 174169 518084
rect 174169 518050 174203 518084
rect 174203 518050 174207 518084
rect 174155 518041 174207 518050
rect 174219 518084 174271 518093
rect 177781 518084 177833 518093
rect 174219 518050 174261 518084
rect 174261 518050 174271 518084
rect 177781 518050 177791 518084
rect 177791 518050 177833 518084
rect 174219 518041 174271 518050
rect 177781 518041 177833 518050
rect 177845 518084 177897 518093
rect 177845 518050 177849 518084
rect 177849 518050 177883 518084
rect 177883 518050 177897 518084
rect 177845 518041 177897 518050
rect 177909 518084 177961 518093
rect 177973 518084 178025 518093
rect 178037 518084 178089 518093
rect 181599 518084 181651 518093
rect 181663 518084 181715 518093
rect 181727 518084 181779 518093
rect 177909 518050 177941 518084
rect 177941 518050 177961 518084
rect 177973 518050 177975 518084
rect 177975 518050 178025 518084
rect 178037 518050 178067 518084
rect 178067 518050 178089 518084
rect 181599 518050 181621 518084
rect 181621 518050 181651 518084
rect 181663 518050 181713 518084
rect 181713 518050 181715 518084
rect 181727 518050 181747 518084
rect 181747 518050 181779 518084
rect 177909 518041 177961 518050
rect 177973 518041 178025 518050
rect 178037 518041 178089 518050
rect 181599 518041 181651 518050
rect 181663 518041 181715 518050
rect 181727 518041 181779 518050
rect 181791 518084 181843 518093
rect 181791 518050 181805 518084
rect 181805 518050 181839 518084
rect 181839 518050 181843 518084
rect 181791 518041 181843 518050
rect 181855 518084 181907 518093
rect 185417 518084 185469 518093
rect 181855 518050 181897 518084
rect 181897 518050 181907 518084
rect 185417 518050 185427 518084
rect 185427 518050 185469 518084
rect 181855 518041 181907 518050
rect 185417 518041 185469 518050
rect 185481 518084 185533 518093
rect 185481 518050 185485 518084
rect 185485 518050 185519 518084
rect 185519 518050 185533 518084
rect 185481 518041 185533 518050
rect 185545 518084 185597 518093
rect 185609 518084 185661 518093
rect 185673 518084 185725 518093
rect 185545 518050 185577 518084
rect 185577 518050 185597 518084
rect 185609 518050 185611 518084
rect 185611 518050 185661 518084
rect 185673 518050 185703 518084
rect 185703 518050 185725 518084
rect 185545 518041 185597 518050
rect 185609 518041 185661 518050
rect 185673 518041 185725 518050
rect 174623 517540 174675 517549
rect 174623 517506 174629 517540
rect 174629 517506 174663 517540
rect 174663 517506 174675 517540
rect 174623 517497 174675 517506
rect 174687 517540 174739 517549
rect 174751 517540 174803 517549
rect 174815 517540 174867 517549
rect 174687 517506 174721 517540
rect 174721 517506 174739 517540
rect 174751 517506 174755 517540
rect 174755 517506 174803 517540
rect 174815 517506 174847 517540
rect 174847 517506 174867 517540
rect 174687 517497 174739 517506
rect 174751 517497 174803 517506
rect 174815 517497 174867 517506
rect 174879 517540 174931 517549
rect 174879 517506 174905 517540
rect 174905 517506 174931 517540
rect 174879 517497 174931 517506
rect 178441 517497 178493 517549
rect 178505 517540 178557 517549
rect 178505 517506 178527 517540
rect 178527 517506 178557 517540
rect 178505 517497 178557 517506
rect 178569 517540 178621 517549
rect 178569 517506 178585 517540
rect 178585 517506 178619 517540
rect 178619 517506 178621 517540
rect 178569 517497 178621 517506
rect 178633 517540 178685 517549
rect 178697 517540 178749 517549
rect 182259 517540 182311 517549
rect 178633 517506 178677 517540
rect 178677 517506 178685 517540
rect 178697 517506 178711 517540
rect 178711 517506 178749 517540
rect 182259 517506 182265 517540
rect 182265 517506 182299 517540
rect 182299 517506 182311 517540
rect 178633 517497 178685 517506
rect 178697 517497 178749 517506
rect 182259 517497 182311 517506
rect 182323 517540 182375 517549
rect 182387 517540 182439 517549
rect 182451 517540 182503 517549
rect 182323 517506 182357 517540
rect 182357 517506 182375 517540
rect 182387 517506 182391 517540
rect 182391 517506 182439 517540
rect 182451 517506 182483 517540
rect 182483 517506 182503 517540
rect 182323 517497 182375 517506
rect 182387 517497 182439 517506
rect 182451 517497 182503 517506
rect 182515 517540 182567 517549
rect 182515 517506 182541 517540
rect 182541 517506 182567 517540
rect 182515 517497 182567 517506
rect 186077 517497 186129 517549
rect 186141 517540 186193 517549
rect 186141 517506 186163 517540
rect 186163 517506 186193 517540
rect 186141 517497 186193 517506
rect 186205 517540 186257 517549
rect 186205 517506 186221 517540
rect 186221 517506 186255 517540
rect 186255 517506 186257 517540
rect 186205 517497 186257 517506
rect 186269 517540 186321 517549
rect 186333 517540 186385 517549
rect 186269 517506 186313 517540
rect 186313 517506 186321 517540
rect 186333 517506 186347 517540
rect 186347 517506 186385 517540
rect 186269 517497 186321 517506
rect 186333 517497 186385 517506
rect 177656 517395 177708 517447
rect 178300 517395 178352 517447
rect 173963 516996 174015 517005
rect 174027 516996 174079 517005
rect 174091 516996 174143 517005
rect 173963 516962 173985 516996
rect 173985 516962 174015 516996
rect 174027 516962 174077 516996
rect 174077 516962 174079 516996
rect 174091 516962 174111 516996
rect 174111 516962 174143 516996
rect 173963 516953 174015 516962
rect 174027 516953 174079 516962
rect 174091 516953 174143 516962
rect 174155 516996 174207 517005
rect 174155 516962 174169 516996
rect 174169 516962 174203 516996
rect 174203 516962 174207 516996
rect 174155 516953 174207 516962
rect 174219 516996 174271 517005
rect 177781 516996 177833 517005
rect 174219 516962 174261 516996
rect 174261 516962 174271 516996
rect 177781 516962 177791 516996
rect 177791 516962 177833 516996
rect 174219 516953 174271 516962
rect 177781 516953 177833 516962
rect 177845 516996 177897 517005
rect 177845 516962 177849 516996
rect 177849 516962 177883 516996
rect 177883 516962 177897 516996
rect 177845 516953 177897 516962
rect 177909 516996 177961 517005
rect 177973 516996 178025 517005
rect 178037 516996 178089 517005
rect 181599 516996 181651 517005
rect 181663 516996 181715 517005
rect 181727 516996 181779 517005
rect 177909 516962 177941 516996
rect 177941 516962 177961 516996
rect 177973 516962 177975 516996
rect 177975 516962 178025 516996
rect 178037 516962 178067 516996
rect 178067 516962 178089 516996
rect 181599 516962 181621 516996
rect 181621 516962 181651 516996
rect 181663 516962 181713 516996
rect 181713 516962 181715 516996
rect 181727 516962 181747 516996
rect 181747 516962 181779 516996
rect 177909 516953 177961 516962
rect 177973 516953 178025 516962
rect 178037 516953 178089 516962
rect 181599 516953 181651 516962
rect 181663 516953 181715 516962
rect 181727 516953 181779 516962
rect 181791 516996 181843 517005
rect 181791 516962 181805 516996
rect 181805 516962 181839 516996
rect 181839 516962 181843 516996
rect 181791 516953 181843 516962
rect 181855 516996 181907 517005
rect 185417 516996 185469 517005
rect 181855 516962 181897 516996
rect 181897 516962 181907 516996
rect 185417 516962 185427 516996
rect 185427 516962 185469 516996
rect 181855 516953 181907 516962
rect 185417 516953 185469 516962
rect 185481 516996 185533 517005
rect 185481 516962 185485 516996
rect 185485 516962 185519 516996
rect 185519 516962 185533 516996
rect 185481 516953 185533 516962
rect 185545 516996 185597 517005
rect 185609 516996 185661 517005
rect 185673 516996 185725 517005
rect 185545 516962 185577 516996
rect 185577 516962 185597 516996
rect 185609 516962 185611 516996
rect 185611 516962 185661 516996
rect 185673 516962 185703 516996
rect 185703 516962 185725 516996
rect 185545 516953 185597 516962
rect 185609 516953 185661 516962
rect 185673 516953 185725 516962
rect 174623 516452 174675 516461
rect 174623 516418 174629 516452
rect 174629 516418 174663 516452
rect 174663 516418 174675 516452
rect 174623 516409 174675 516418
rect 174687 516452 174739 516461
rect 174751 516452 174803 516461
rect 174815 516452 174867 516461
rect 174687 516418 174721 516452
rect 174721 516418 174739 516452
rect 174751 516418 174755 516452
rect 174755 516418 174803 516452
rect 174815 516418 174847 516452
rect 174847 516418 174867 516452
rect 174687 516409 174739 516418
rect 174751 516409 174803 516418
rect 174815 516409 174867 516418
rect 174879 516452 174931 516461
rect 174879 516418 174905 516452
rect 174905 516418 174931 516452
rect 174879 516409 174931 516418
rect 178441 516409 178493 516461
rect 178505 516452 178557 516461
rect 178505 516418 178527 516452
rect 178527 516418 178557 516452
rect 178505 516409 178557 516418
rect 178569 516452 178621 516461
rect 178569 516418 178585 516452
rect 178585 516418 178619 516452
rect 178619 516418 178621 516452
rect 178569 516409 178621 516418
rect 178633 516452 178685 516461
rect 178697 516452 178749 516461
rect 182259 516452 182311 516461
rect 178633 516418 178677 516452
rect 178677 516418 178685 516452
rect 178697 516418 178711 516452
rect 178711 516418 178749 516452
rect 182259 516418 182265 516452
rect 182265 516418 182299 516452
rect 182299 516418 182311 516452
rect 178633 516409 178685 516418
rect 178697 516409 178749 516418
rect 182259 516409 182311 516418
rect 182323 516452 182375 516461
rect 182387 516452 182439 516461
rect 182451 516452 182503 516461
rect 182323 516418 182357 516452
rect 182357 516418 182375 516452
rect 182387 516418 182391 516452
rect 182391 516418 182439 516452
rect 182451 516418 182483 516452
rect 182483 516418 182503 516452
rect 182323 516409 182375 516418
rect 182387 516409 182439 516418
rect 182451 516409 182503 516418
rect 182515 516452 182567 516461
rect 182515 516418 182541 516452
rect 182541 516418 182567 516452
rect 182515 516409 182567 516418
rect 186077 516409 186129 516461
rect 186141 516452 186193 516461
rect 186141 516418 186163 516452
rect 186163 516418 186193 516452
rect 186141 516409 186193 516418
rect 186205 516452 186257 516461
rect 186205 516418 186221 516452
rect 186221 516418 186255 516452
rect 186255 516418 186257 516452
rect 186205 516409 186257 516418
rect 186269 516452 186321 516461
rect 186333 516452 186385 516461
rect 186269 516418 186313 516452
rect 186313 516418 186321 516452
rect 186333 516418 186347 516452
rect 186347 516418 186385 516452
rect 186269 516409 186321 516418
rect 186333 516409 186385 516418
rect 173963 515908 174015 515917
rect 174027 515908 174079 515917
rect 174091 515908 174143 515917
rect 173963 515874 173985 515908
rect 173985 515874 174015 515908
rect 174027 515874 174077 515908
rect 174077 515874 174079 515908
rect 174091 515874 174111 515908
rect 174111 515874 174143 515908
rect 173963 515865 174015 515874
rect 174027 515865 174079 515874
rect 174091 515865 174143 515874
rect 174155 515908 174207 515917
rect 174155 515874 174169 515908
rect 174169 515874 174203 515908
rect 174203 515874 174207 515908
rect 174155 515865 174207 515874
rect 174219 515908 174271 515917
rect 177781 515908 177833 515917
rect 174219 515874 174261 515908
rect 174261 515874 174271 515908
rect 177781 515874 177791 515908
rect 177791 515874 177833 515908
rect 174219 515865 174271 515874
rect 177781 515865 177833 515874
rect 177845 515908 177897 515917
rect 177845 515874 177849 515908
rect 177849 515874 177883 515908
rect 177883 515874 177897 515908
rect 177845 515865 177897 515874
rect 177909 515908 177961 515917
rect 177973 515908 178025 515917
rect 178037 515908 178089 515917
rect 181599 515908 181651 515917
rect 181663 515908 181715 515917
rect 181727 515908 181779 515917
rect 177909 515874 177941 515908
rect 177941 515874 177961 515908
rect 177973 515874 177975 515908
rect 177975 515874 178025 515908
rect 178037 515874 178067 515908
rect 178067 515874 178089 515908
rect 181599 515874 181621 515908
rect 181621 515874 181651 515908
rect 181663 515874 181713 515908
rect 181713 515874 181715 515908
rect 181727 515874 181747 515908
rect 181747 515874 181779 515908
rect 177909 515865 177961 515874
rect 177973 515865 178025 515874
rect 178037 515865 178089 515874
rect 181599 515865 181651 515874
rect 181663 515865 181715 515874
rect 181727 515865 181779 515874
rect 181791 515908 181843 515917
rect 181791 515874 181805 515908
rect 181805 515874 181839 515908
rect 181839 515874 181843 515908
rect 181791 515865 181843 515874
rect 181855 515908 181907 515917
rect 185417 515908 185469 515917
rect 181855 515874 181897 515908
rect 181897 515874 181907 515908
rect 185417 515874 185427 515908
rect 185427 515874 185469 515908
rect 181855 515865 181907 515874
rect 185417 515865 185469 515874
rect 185481 515908 185533 515917
rect 185481 515874 185485 515908
rect 185485 515874 185519 515908
rect 185519 515874 185533 515908
rect 185481 515865 185533 515874
rect 185545 515908 185597 515917
rect 185609 515908 185661 515917
rect 185673 515908 185725 515917
rect 185545 515874 185577 515908
rect 185577 515874 185597 515908
rect 185609 515874 185611 515908
rect 185611 515874 185661 515908
rect 185673 515874 185703 515908
rect 185703 515874 185725 515908
rect 185545 515865 185597 515874
rect 185609 515865 185661 515874
rect 185673 515865 185725 515874
rect 173608 515806 173660 515815
rect 173608 515772 173617 515806
rect 173617 515772 173651 515806
rect 173651 515772 173660 515806
rect 173608 515763 173660 515772
rect 181336 515763 181388 515815
rect 186580 515806 186632 515815
rect 186580 515772 186589 515806
rect 186589 515772 186623 515806
rect 186623 515772 186632 515806
rect 186580 515763 186632 515772
rect 173332 515491 173384 515543
rect 186488 515534 186540 515543
rect 186488 515500 186497 515534
rect 186497 515500 186531 515534
rect 186531 515500 186540 515534
rect 186488 515491 186540 515500
rect 182164 515423 182216 515475
rect 174623 515364 174675 515373
rect 174623 515330 174629 515364
rect 174629 515330 174663 515364
rect 174663 515330 174675 515364
rect 174623 515321 174675 515330
rect 174687 515364 174739 515373
rect 174751 515364 174803 515373
rect 174815 515364 174867 515373
rect 174687 515330 174721 515364
rect 174721 515330 174739 515364
rect 174751 515330 174755 515364
rect 174755 515330 174803 515364
rect 174815 515330 174847 515364
rect 174847 515330 174867 515364
rect 174687 515321 174739 515330
rect 174751 515321 174803 515330
rect 174815 515321 174867 515330
rect 174879 515364 174931 515373
rect 174879 515330 174905 515364
rect 174905 515330 174931 515364
rect 174879 515321 174931 515330
rect 178441 515321 178493 515373
rect 178505 515364 178557 515373
rect 178505 515330 178527 515364
rect 178527 515330 178557 515364
rect 178505 515321 178557 515330
rect 178569 515364 178621 515373
rect 178569 515330 178585 515364
rect 178585 515330 178619 515364
rect 178619 515330 178621 515364
rect 178569 515321 178621 515330
rect 178633 515364 178685 515373
rect 178697 515364 178749 515373
rect 182259 515364 182311 515373
rect 178633 515330 178677 515364
rect 178677 515330 178685 515364
rect 178697 515330 178711 515364
rect 178711 515330 178749 515364
rect 182259 515330 182265 515364
rect 182265 515330 182299 515364
rect 182299 515330 182311 515364
rect 178633 515321 178685 515330
rect 178697 515321 178749 515330
rect 182259 515321 182311 515330
rect 182323 515364 182375 515373
rect 182387 515364 182439 515373
rect 182451 515364 182503 515373
rect 182323 515330 182357 515364
rect 182357 515330 182375 515364
rect 182387 515330 182391 515364
rect 182391 515330 182439 515364
rect 182451 515330 182483 515364
rect 182483 515330 182503 515364
rect 182323 515321 182375 515330
rect 182387 515321 182439 515330
rect 182451 515321 182503 515330
rect 182515 515364 182567 515373
rect 182515 515330 182541 515364
rect 182541 515330 182567 515364
rect 182515 515321 182567 515330
rect 186077 515321 186129 515373
rect 186141 515364 186193 515373
rect 186141 515330 186163 515364
rect 186163 515330 186193 515364
rect 186141 515321 186193 515330
rect 186205 515364 186257 515373
rect 186205 515330 186221 515364
rect 186221 515330 186255 515364
rect 186255 515330 186257 515364
rect 186205 515321 186257 515330
rect 186269 515364 186321 515373
rect 186333 515364 186385 515373
rect 186269 515330 186313 515364
rect 186313 515330 186321 515364
rect 186333 515330 186347 515364
rect 186347 515330 186385 515364
rect 186269 515321 186321 515330
rect 186333 515321 186385 515330
rect 173250 512810 173450 513000
rect 2000 507000 4000 509000
rect 177580 512810 177780 513000
rect 181910 512810 182110 513000
rect 2000 464000 4000 466000
rect 186230 512810 186430 513000
rect 2000 421000 4000 423000
rect 2000 378000 4000 380000
<< metal2 >>
rect 18000 701000 20000 701010
rect 18000 698990 20000 699000
rect 70000 701000 72000 701010
rect 70000 698990 72000 699000
rect 122000 701000 124000 701010
rect 122000 698990 124000 699000
rect 3000 684000 5000 684010
rect 3000 681990 5000 682000
rect 146000 628000 148000 628010
rect 146000 546000 148000 626000
rect 146000 543990 148000 544000
rect 154000 553000 156000 553010
rect 154000 540000 156000 551000
rect 165878 540995 166008 541025
rect 165878 540895 165888 540995
rect 165998 540895 166008 540995
rect 165878 540875 166008 540895
rect 165878 540775 165888 540875
rect 165998 540775 166008 540875
rect 165878 540755 166008 540775
rect 165878 540655 165888 540755
rect 165998 540655 166008 540755
rect 165878 540635 166008 540655
rect 169678 540995 169808 541025
rect 169678 540895 169688 540995
rect 169798 540895 169808 540995
rect 169678 540875 169808 540895
rect 169678 540775 169688 540875
rect 169798 540775 169808 540875
rect 169678 540755 169808 540775
rect 169678 540655 169688 540755
rect 169798 540655 169808 540755
rect 169678 540635 169808 540655
rect 173378 540995 173508 541025
rect 173378 540895 173388 540995
rect 173498 540895 173508 540995
rect 173378 540875 173508 540895
rect 173378 540775 173388 540875
rect 173498 540775 173508 540875
rect 173378 540755 173508 540775
rect 173378 540655 173388 540755
rect 173498 540655 173508 540755
rect 173378 540635 173508 540655
rect 176878 540995 177008 541025
rect 176878 540895 176888 540995
rect 176998 540895 177008 540995
rect 176878 540875 177008 540895
rect 176878 540775 176888 540875
rect 176998 540775 177008 540875
rect 176878 540755 177008 540775
rect 176878 540655 176888 540755
rect 176998 540655 177008 540755
rect 176878 540635 177008 540655
rect 180478 540995 180608 541025
rect 180478 540895 180488 540995
rect 180598 540895 180608 540995
rect 180478 540875 180608 540895
rect 180478 540775 180488 540875
rect 180598 540775 180608 540875
rect 180478 540755 180608 540775
rect 180478 540655 180488 540755
rect 180598 540655 180608 540755
rect 180478 540635 180608 540655
rect 183778 540995 183908 541025
rect 183778 540895 183788 540995
rect 183898 540895 183908 540995
rect 183778 540875 183908 540895
rect 183778 540775 183788 540875
rect 183898 540775 183908 540875
rect 183778 540755 183908 540775
rect 183778 540655 183788 540755
rect 183898 540655 183908 540755
rect 183778 540635 183908 540655
rect 187078 540995 187208 541025
rect 187078 540895 187088 540995
rect 187198 540895 187208 540995
rect 187078 540875 187208 540895
rect 187078 540775 187088 540875
rect 187198 540775 187208 540875
rect 187078 540755 187208 540775
rect 187078 540655 187088 540755
rect 187198 540655 187208 540755
rect 187078 540635 187208 540655
rect 190378 540995 190508 541025
rect 190378 540895 190388 540995
rect 190498 540895 190508 540995
rect 190378 540875 190508 540895
rect 190378 540775 190388 540875
rect 190498 540775 190508 540875
rect 190378 540755 190508 540775
rect 190378 540655 190388 540755
rect 190498 540655 190508 540755
rect 190378 540635 190508 540655
rect 163028 538865 163328 538875
rect 161378 538665 161528 538675
rect 159388 538655 159488 538665
rect 159388 538555 159398 538655
rect 159478 538555 159488 538655
rect 159388 538340 159488 538555
rect 161378 538545 161388 538665
rect 161508 538545 161528 538665
rect 165928 538815 166008 540635
rect 166678 540245 166878 540255
rect 166678 540065 166688 540245
rect 166868 540065 166878 540245
rect 166678 540055 166878 540065
rect 166678 539305 166878 539315
rect 166678 539125 166688 539305
rect 166868 539125 166878 539305
rect 166678 539115 166878 539125
rect 169728 538815 169808 540635
rect 170478 540245 170678 540255
rect 170478 540065 170488 540245
rect 170668 540065 170678 540245
rect 170478 540055 170678 540065
rect 170478 539305 170678 539315
rect 170478 539125 170488 539305
rect 170668 539125 170678 539305
rect 170478 539115 170678 539125
rect 173428 538815 173508 540635
rect 174178 540255 174378 540265
rect 174178 540075 174188 540255
rect 174368 540075 174378 540255
rect 174178 540065 174378 540075
rect 174178 539305 174378 539315
rect 174178 539125 174188 539305
rect 174368 539125 174378 539305
rect 174178 539115 174378 539125
rect 176928 538815 177008 540635
rect 177688 540245 177888 540255
rect 177688 540065 177698 540245
rect 177878 540065 177888 540245
rect 177688 540055 177888 540065
rect 177678 539305 177878 539315
rect 177678 539125 177688 539305
rect 177868 539125 177878 539305
rect 177678 539115 177878 539125
rect 180528 538815 180608 540635
rect 181278 540245 181478 540255
rect 181278 540065 181288 540245
rect 181468 540065 181478 540245
rect 181278 540055 181478 540065
rect 181278 539305 181478 539315
rect 181278 539125 181288 539305
rect 181468 539125 181478 539305
rect 181278 539115 181478 539125
rect 183828 538815 183908 540635
rect 184578 540245 184778 540255
rect 184578 540065 184588 540245
rect 184768 540065 184778 540245
rect 184578 540055 184778 540065
rect 184578 539305 184778 539315
rect 184578 539125 184588 539305
rect 184768 539125 184778 539305
rect 184578 539115 184778 539125
rect 187128 538815 187208 540635
rect 187888 540245 188088 540255
rect 187888 540065 187898 540245
rect 188078 540065 188088 540245
rect 187888 540055 188088 540065
rect 187878 539305 188078 539315
rect 187878 539125 187888 539305
rect 188068 539125 188078 539305
rect 187878 539115 188078 539125
rect 190428 538815 190508 540635
rect 191178 540245 191378 540255
rect 191178 540065 191188 540245
rect 191368 540065 191378 540245
rect 191178 540055 191378 540065
rect 191778 540245 191998 540255
rect 191778 540065 191808 540245
rect 191988 540065 191998 540245
rect 191778 540055 191998 540065
rect 191188 539315 191388 539325
rect 191188 539135 191198 539315
rect 191378 539135 191388 539315
rect 191188 539125 191388 539135
rect 191808 539305 192008 539315
rect 191808 539125 191818 539305
rect 191998 539125 192008 539305
rect 191808 539115 192008 539125
rect 165878 538805 166058 538815
rect 165878 538705 165898 538805
rect 166038 538705 166058 538805
rect 165878 538695 166058 538705
rect 169678 538805 169858 538815
rect 169678 538705 169698 538805
rect 169838 538705 169858 538805
rect 169678 538695 169858 538705
rect 173378 538805 173558 538815
rect 173378 538705 173398 538805
rect 173538 538705 173558 538805
rect 173378 538695 173558 538705
rect 176878 538805 177058 538815
rect 176878 538705 176898 538805
rect 177038 538705 177058 538805
rect 176878 538695 177058 538705
rect 180478 538805 180658 538815
rect 180478 538705 180498 538805
rect 180638 538705 180658 538805
rect 180478 538695 180658 538705
rect 183778 538805 183958 538815
rect 183778 538705 183798 538805
rect 183938 538705 183958 538805
rect 183778 538695 183958 538705
rect 187078 538805 187258 538815
rect 187078 538705 187098 538805
rect 187238 538705 187258 538805
rect 187078 538695 187258 538705
rect 190378 538805 190558 538815
rect 190378 538705 190398 538805
rect 190538 538705 190558 538805
rect 190378 538695 190558 538705
rect 163028 538655 163328 538665
rect 161378 538535 161528 538545
rect 154000 537990 156000 538000
rect 159383 538295 159493 538340
rect 159383 538215 159398 538295
rect 159478 538215 159493 538295
rect 159383 536935 159493 538215
rect 162868 537945 162948 537955
rect 162868 537935 162878 537945
rect 161688 537885 162878 537935
rect 162938 537885 162948 537945
rect 161688 537745 161738 537885
rect 162868 537875 162948 537885
rect 161678 537735 161758 537745
rect 161678 537675 161688 537735
rect 161748 537675 161758 537735
rect 161678 537665 161758 537675
rect 157413 536925 159493 536935
rect 157413 536845 157418 536925
rect 157508 536845 159493 536925
rect 161768 536905 161868 536925
rect 161768 536885 161788 536905
rect 157413 536825 159493 536845
rect 161088 536825 161788 536885
rect 161848 536825 161868 536905
rect 157418 534975 157498 536825
rect 158478 536565 158588 536825
rect 161088 536805 161868 536825
rect 161088 536565 161168 536805
rect 158468 536555 158598 536565
rect 158468 536395 158478 536555
rect 158578 536395 158598 536555
rect 161068 536545 161188 536565
rect 161068 536465 161088 536545
rect 161168 536465 161188 536545
rect 161068 536445 161188 536465
rect 158468 536375 158598 536395
rect 163818 536285 189028 536295
rect 163818 536275 182188 536285
rect 163818 536265 178868 536275
rect 163818 536235 166928 536265
rect 163818 535905 163838 536235
rect 164048 536045 166928 536235
rect 167258 536255 172608 536265
rect 167258 536045 169568 536255
rect 164048 535975 169568 536045
rect 169868 535975 172608 536255
rect 172938 536255 178868 536265
rect 172938 535975 175278 536255
rect 164048 535945 175278 535975
rect 175498 535965 178868 536255
rect 179068 536025 182188 536275
rect 182388 536275 189028 536285
rect 182388 536265 188778 536275
rect 182388 536145 185488 536265
rect 185698 536145 188778 536265
rect 182388 536035 188778 536145
rect 188998 536035 189028 536275
rect 182388 536025 189028 536035
rect 179068 535965 189028 536025
rect 175498 535945 189028 535965
rect 164048 535905 189028 535945
rect 163818 535875 189028 535905
rect 160168 535575 160368 535605
rect 163528 535575 167238 535605
rect 160168 535435 160198 535575
rect 160348 535565 160368 535575
rect 160168 535425 160208 535435
rect 160358 535425 160368 535565
rect 160168 535415 160368 535425
rect 163478 535555 167238 535575
rect 163478 535425 166718 535555
rect 166848 535545 167238 535555
rect 166848 535425 166898 535545
rect 163478 535415 166898 535425
rect 167028 535525 167238 535545
rect 167028 535415 167078 535525
rect 163478 535395 167078 535415
rect 167208 535395 167238 535525
rect 163478 535365 167238 535395
rect 163478 535235 166698 535365
rect 166828 535355 167238 535365
rect 166828 535235 166888 535355
rect 163478 535225 166888 535235
rect 167018 535345 167238 535355
rect 167018 535225 167088 535345
rect 163478 535215 167088 535225
rect 167218 535215 167238 535345
rect 163478 535185 167238 535215
rect 163478 534975 163898 535185
rect 157418 534555 163898 534975
rect 185058 532775 185188 532785
rect 172410 532745 172466 532755
rect 174488 532745 174618 532755
rect 176642 532745 176698 532755
rect 178758 532745 178814 532755
rect 180874 532745 180930 532755
rect 182990 532745 183046 532755
rect 172358 532735 172488 532745
rect 174488 532565 174618 532575
rect 176578 532735 176708 532745
rect 172358 532555 172488 532565
rect 172410 531955 172466 532555
rect 174526 531955 174582 532565
rect 176578 532555 176708 532565
rect 178698 532735 178828 532745
rect 178698 532555 178828 532565
rect 180868 532735 180998 532745
rect 180868 532555 180998 532565
rect 182958 532735 183088 532745
rect 187222 532745 187278 532755
rect 185058 532595 185188 532605
rect 187168 532735 187288 532745
rect 187268 532595 187288 532735
rect 182958 532555 183088 532565
rect 176642 531955 176698 532555
rect 178758 531955 178814 532555
rect 180874 531955 180930 532555
rect 182990 531955 183046 532555
rect 185106 531955 185162 532595
rect 187168 532575 187288 532595
rect 187222 531955 187278 532575
rect 172424 530441 172452 531955
rect 174540 530441 174568 531955
rect 176656 531613 176684 531955
rect 178772 531613 178800 531955
rect 176656 531585 176776 531613
rect 178772 531585 178892 531613
rect 174623 530607 174931 530616
rect 174623 530605 174629 530607
rect 174685 530605 174709 530607
rect 174765 530605 174789 530607
rect 174845 530605 174869 530607
rect 174925 530605 174931 530607
rect 174685 530553 174687 530605
rect 174867 530553 174869 530605
rect 174623 530551 174629 530553
rect 174685 530551 174709 530553
rect 174765 530551 174789 530553
rect 174845 530551 174869 530553
rect 174925 530551 174931 530553
rect 174623 530542 174931 530551
rect 176748 530441 176776 531585
rect 178441 530607 178749 530616
rect 178441 530605 178447 530607
rect 178503 530605 178527 530607
rect 178583 530605 178607 530607
rect 178663 530605 178687 530607
rect 178743 530605 178749 530607
rect 178503 530553 178505 530605
rect 178685 530553 178687 530605
rect 178441 530551 178447 530553
rect 178503 530551 178527 530553
rect 178583 530551 178607 530553
rect 178663 530551 178687 530553
rect 178743 530551 178749 530553
rect 178441 530542 178749 530551
rect 178864 530525 178892 531585
rect 178772 530509 178892 530525
rect 176828 530503 176880 530509
rect 176828 530445 176880 530451
rect 178760 530503 178892 530509
rect 178812 530497 178892 530503
rect 179496 530503 179548 530509
rect 178760 530445 178812 530451
rect 179496 530445 179548 530451
rect 172412 530435 172464 530441
rect 172412 530377 172464 530383
rect 174528 530435 174580 530441
rect 174528 530377 174580 530383
rect 176736 530435 176788 530441
rect 176736 530377 176788 530383
rect 174804 530367 174856 530373
rect 174804 530309 174856 530315
rect 175448 530367 175500 530373
rect 175448 530309 175500 530315
rect 173963 530063 174271 530072
rect 173963 530061 173969 530063
rect 174025 530061 174049 530063
rect 174105 530061 174129 530063
rect 174185 530061 174209 530063
rect 174265 530061 174271 530063
rect 174025 530009 174027 530061
rect 174207 530009 174209 530061
rect 173963 530007 173969 530009
rect 174025 530007 174049 530009
rect 174105 530007 174129 530009
rect 174185 530007 174209 530009
rect 174265 530007 174271 530009
rect 173963 529998 174271 530007
rect 174816 529829 174844 530309
rect 174804 529823 174856 529829
rect 174804 529765 174856 529771
rect 175356 529619 175408 529625
rect 175356 529561 175408 529567
rect 174623 529519 174931 529528
rect 174623 529517 174629 529519
rect 174685 529517 174709 529519
rect 174765 529517 174789 529519
rect 174845 529517 174869 529519
rect 174925 529517 174931 529519
rect 174685 529465 174687 529517
rect 174867 529465 174869 529517
rect 174623 529463 174629 529465
rect 174685 529463 174709 529465
rect 174765 529463 174789 529465
rect 174845 529463 174869 529465
rect 174925 529463 174931 529465
rect 174623 529454 174931 529463
rect 175368 529421 175396 529561
rect 175356 529415 175408 529421
rect 175356 529357 175408 529363
rect 175460 529285 175488 530309
rect 176644 530299 176696 530305
rect 176644 530241 176696 530247
rect 176092 529619 176144 529625
rect 176092 529561 176144 529567
rect 175448 529279 175500 529285
rect 175448 529221 175500 529227
rect 173608 529211 173660 529217
rect 173608 529153 173660 529159
rect 175264 529211 175316 529217
rect 175264 529153 175316 529159
rect 173620 515821 173648 529153
rect 173963 528975 174271 528984
rect 173963 528973 173969 528975
rect 174025 528973 174049 528975
rect 174105 528973 174129 528975
rect 174185 528973 174209 528975
rect 174265 528973 174271 528975
rect 174025 528921 174027 528973
rect 174207 528921 174209 528973
rect 173963 528919 173969 528921
rect 174025 528919 174049 528921
rect 174105 528919 174129 528921
rect 174185 528919 174209 528921
rect 174265 528919 174271 528921
rect 173963 528910 174271 528919
rect 175276 528877 175304 529153
rect 176104 529081 176132 529561
rect 175908 529075 175960 529081
rect 175908 529017 175960 529023
rect 176092 529075 176144 529081
rect 176092 529017 176144 529023
rect 175264 528871 175316 528877
rect 175264 528813 175316 528819
rect 175920 528673 175948 529017
rect 175908 528667 175960 528673
rect 175908 528609 175960 528615
rect 174623 528431 174931 528440
rect 174623 528429 174629 528431
rect 174685 528429 174709 528431
rect 174765 528429 174789 528431
rect 174845 528429 174869 528431
rect 174925 528429 174931 528431
rect 174685 528377 174687 528429
rect 174867 528377 174869 528429
rect 174623 528375 174629 528377
rect 174685 528375 174709 528377
rect 174765 528375 174789 528377
rect 174845 528375 174869 528377
rect 174925 528375 174931 528377
rect 174623 528366 174931 528375
rect 176104 528197 176132 529017
rect 176656 528877 176684 530241
rect 176840 529761 176868 530445
rect 178944 530367 178996 530373
rect 178944 530309 178996 530315
rect 179220 530367 179272 530373
rect 179220 530309 179272 530315
rect 177288 530299 177340 530305
rect 177288 530241 177340 530247
rect 178208 530299 178260 530305
rect 178208 530241 178260 530247
rect 176828 529755 176880 529761
rect 176828 529697 176880 529703
rect 176736 529279 176788 529285
rect 176736 529221 176788 529227
rect 176644 528871 176696 528877
rect 176644 528813 176696 528819
rect 176748 528537 176776 529221
rect 176276 528531 176328 528537
rect 176276 528473 176328 528479
rect 176368 528531 176420 528537
rect 176368 528473 176420 528479
rect 176736 528531 176788 528537
rect 176736 528473 176788 528479
rect 176092 528191 176144 528197
rect 176092 528133 176144 528139
rect 173963 527887 174271 527896
rect 173963 527885 173969 527887
rect 174025 527885 174049 527887
rect 174105 527885 174129 527887
rect 174185 527885 174209 527887
rect 174265 527885 174271 527887
rect 174025 527833 174027 527885
rect 174207 527833 174209 527885
rect 173963 527831 173969 527833
rect 174025 527831 174049 527833
rect 174105 527831 174129 527833
rect 174185 527831 174209 527833
rect 174265 527831 174271 527833
rect 173963 527822 174271 527831
rect 176288 527789 176316 528473
rect 176380 528265 176408 528473
rect 176748 528333 176776 528473
rect 176736 528327 176788 528333
rect 176736 528269 176788 528275
rect 176840 528265 176868 529697
rect 177300 529217 177328 530241
rect 177656 530163 177708 530169
rect 177656 530105 177708 530111
rect 177668 529693 177696 530105
rect 177781 530063 178089 530072
rect 177781 530061 177787 530063
rect 177843 530061 177867 530063
rect 177923 530061 177947 530063
rect 178003 530061 178027 530063
rect 178083 530061 178089 530063
rect 177843 530009 177845 530061
rect 178025 530009 178027 530061
rect 177781 530007 177787 530009
rect 177843 530007 177867 530009
rect 177923 530007 177947 530009
rect 178003 530007 178027 530009
rect 178083 530007 178089 530009
rect 177781 529998 178089 530007
rect 178220 529965 178248 530241
rect 178300 530163 178352 530169
rect 178300 530105 178352 530111
rect 178208 529959 178260 529965
rect 178208 529901 178260 529907
rect 178116 529891 178168 529897
rect 178116 529833 178168 529839
rect 177380 529687 177432 529693
rect 177380 529629 177432 529635
rect 177564 529687 177616 529693
rect 177564 529629 177616 529635
rect 177656 529687 177708 529693
rect 177656 529629 177708 529635
rect 177288 529211 177340 529217
rect 177288 529153 177340 529159
rect 177012 528531 177064 528537
rect 177012 528473 177064 528479
rect 176368 528259 176420 528265
rect 176368 528201 176420 528207
rect 176828 528259 176880 528265
rect 176828 528201 176880 528207
rect 176276 527783 176328 527789
rect 176276 527725 176328 527731
rect 177024 527653 177052 528473
rect 177392 528061 177420 529629
rect 177576 528741 177604 529629
rect 177932 529619 177984 529625
rect 177932 529561 177984 529567
rect 177944 529421 177972 529561
rect 177932 529415 177984 529421
rect 177932 529357 177984 529363
rect 177656 529279 177708 529285
rect 177656 529221 177708 529227
rect 177668 528877 177696 529221
rect 177781 528975 178089 528984
rect 177781 528973 177787 528975
rect 177843 528973 177867 528975
rect 177923 528973 177947 528975
rect 178003 528973 178027 528975
rect 178083 528973 178089 528975
rect 177843 528921 177845 528973
rect 178025 528921 178027 528973
rect 177781 528919 177787 528921
rect 177843 528919 177867 528921
rect 177923 528919 177947 528921
rect 178003 528919 178027 528921
rect 178083 528919 178089 528921
rect 177781 528910 178089 528919
rect 177656 528871 177708 528877
rect 177656 528813 177708 528819
rect 177564 528735 177616 528741
rect 177564 528677 177616 528683
rect 178024 528735 178076 528741
rect 178024 528677 178076 528683
rect 178036 528333 178064 528677
rect 178024 528327 178076 528333
rect 178024 528269 178076 528275
rect 178128 528197 178156 529833
rect 178220 528741 178248 529901
rect 178312 529353 178340 530105
rect 178441 529519 178749 529528
rect 178441 529517 178447 529519
rect 178503 529517 178527 529519
rect 178583 529517 178607 529519
rect 178663 529517 178687 529519
rect 178743 529517 178749 529519
rect 178503 529465 178505 529517
rect 178685 529465 178687 529517
rect 178441 529463 178447 529465
rect 178503 529463 178527 529465
rect 178583 529463 178607 529465
rect 178663 529463 178687 529465
rect 178743 529463 178749 529465
rect 178441 529454 178749 529463
rect 178300 529347 178352 529353
rect 178300 529289 178352 529295
rect 178208 528735 178260 528741
rect 178208 528677 178260 528683
rect 178312 528605 178432 528621
rect 178312 528599 178444 528605
rect 178312 528593 178392 528599
rect 178116 528191 178168 528197
rect 178116 528133 178168 528139
rect 177380 528055 177432 528061
rect 177380 527997 177432 528003
rect 177781 527887 178089 527896
rect 177781 527885 177787 527887
rect 177843 527885 177867 527887
rect 177923 527885 177947 527887
rect 178003 527885 178027 527887
rect 178083 527885 178089 527887
rect 177843 527833 177845 527885
rect 178025 527833 178027 527885
rect 177781 527831 177787 527833
rect 177843 527831 177867 527833
rect 177923 527831 177947 527833
rect 178003 527831 178027 527833
rect 178083 527831 178089 527833
rect 177781 527822 178089 527831
rect 177012 527647 177064 527653
rect 177012 527589 177064 527595
rect 174623 527343 174931 527352
rect 174623 527341 174629 527343
rect 174685 527341 174709 527343
rect 174765 527341 174789 527343
rect 174845 527341 174869 527343
rect 174925 527341 174931 527343
rect 174685 527289 174687 527341
rect 174867 527289 174869 527341
rect 174623 527287 174629 527289
rect 174685 527287 174709 527289
rect 174765 527287 174789 527289
rect 174845 527287 174869 527289
rect 174925 527287 174931 527289
rect 174623 527278 174931 527287
rect 173963 526799 174271 526808
rect 173963 526797 173969 526799
rect 174025 526797 174049 526799
rect 174105 526797 174129 526799
rect 174185 526797 174209 526799
rect 174265 526797 174271 526799
rect 174025 526745 174027 526797
rect 174207 526745 174209 526797
rect 173963 526743 173969 526745
rect 174025 526743 174049 526745
rect 174105 526743 174129 526745
rect 174185 526743 174209 526745
rect 174265 526743 174271 526745
rect 173963 526734 174271 526743
rect 177781 526799 178089 526808
rect 177781 526797 177787 526799
rect 177843 526797 177867 526799
rect 177923 526797 177947 526799
rect 178003 526797 178027 526799
rect 178083 526797 178089 526799
rect 177843 526745 177845 526797
rect 178025 526745 178027 526797
rect 177781 526743 177787 526745
rect 177843 526743 177867 526745
rect 177923 526743 177947 526745
rect 178003 526743 178027 526745
rect 178083 526743 178089 526745
rect 177781 526734 178089 526743
rect 174623 526255 174931 526264
rect 174623 526253 174629 526255
rect 174685 526253 174709 526255
rect 174765 526253 174789 526255
rect 174845 526253 174869 526255
rect 174925 526253 174931 526255
rect 174685 526201 174687 526253
rect 174867 526201 174869 526253
rect 174623 526199 174629 526201
rect 174685 526199 174709 526201
rect 174765 526199 174789 526201
rect 174845 526199 174869 526201
rect 174925 526199 174931 526201
rect 174623 526190 174931 526199
rect 173963 525711 174271 525720
rect 173963 525709 173969 525711
rect 174025 525709 174049 525711
rect 174105 525709 174129 525711
rect 174185 525709 174209 525711
rect 174265 525709 174271 525711
rect 174025 525657 174027 525709
rect 174207 525657 174209 525709
rect 173963 525655 173969 525657
rect 174025 525655 174049 525657
rect 174105 525655 174129 525657
rect 174185 525655 174209 525657
rect 174265 525655 174271 525657
rect 173963 525646 174271 525655
rect 177781 525711 178089 525720
rect 177781 525709 177787 525711
rect 177843 525709 177867 525711
rect 177923 525709 177947 525711
rect 178003 525709 178027 525711
rect 178083 525709 178089 525711
rect 177843 525657 177845 525709
rect 178025 525657 178027 525709
rect 177781 525655 177787 525657
rect 177843 525655 177867 525657
rect 177923 525655 177947 525657
rect 178003 525655 178027 525657
rect 178083 525655 178089 525657
rect 177781 525646 178089 525655
rect 174623 525167 174931 525176
rect 174623 525165 174629 525167
rect 174685 525165 174709 525167
rect 174765 525165 174789 525167
rect 174845 525165 174869 525167
rect 174925 525165 174931 525167
rect 174685 525113 174687 525165
rect 174867 525113 174869 525165
rect 174623 525111 174629 525113
rect 174685 525111 174709 525113
rect 174765 525111 174789 525113
rect 174845 525111 174869 525113
rect 174925 525111 174931 525113
rect 174623 525102 174931 525111
rect 173963 524623 174271 524632
rect 173963 524621 173969 524623
rect 174025 524621 174049 524623
rect 174105 524621 174129 524623
rect 174185 524621 174209 524623
rect 174265 524621 174271 524623
rect 174025 524569 174027 524621
rect 174207 524569 174209 524621
rect 173963 524567 173969 524569
rect 174025 524567 174049 524569
rect 174105 524567 174129 524569
rect 174185 524567 174209 524569
rect 174265 524567 174271 524569
rect 173963 524558 174271 524567
rect 177781 524623 178089 524632
rect 177781 524621 177787 524623
rect 177843 524621 177867 524623
rect 177923 524621 177947 524623
rect 178003 524621 178027 524623
rect 178083 524621 178089 524623
rect 177843 524569 177845 524621
rect 178025 524569 178027 524621
rect 177781 524567 177787 524569
rect 177843 524567 177867 524569
rect 177923 524567 177947 524569
rect 178003 524567 178027 524569
rect 178083 524567 178089 524569
rect 177781 524558 178089 524567
rect 174623 524079 174931 524088
rect 174623 524077 174629 524079
rect 174685 524077 174709 524079
rect 174765 524077 174789 524079
rect 174845 524077 174869 524079
rect 174925 524077 174931 524079
rect 174685 524025 174687 524077
rect 174867 524025 174869 524077
rect 174623 524023 174629 524025
rect 174685 524023 174709 524025
rect 174765 524023 174789 524025
rect 174845 524023 174869 524025
rect 174925 524023 174931 524025
rect 174623 524014 174931 524023
rect 173963 523535 174271 523544
rect 173963 523533 173969 523535
rect 174025 523533 174049 523535
rect 174105 523533 174129 523535
rect 174185 523533 174209 523535
rect 174265 523533 174271 523535
rect 174025 523481 174027 523533
rect 174207 523481 174209 523533
rect 173963 523479 173969 523481
rect 174025 523479 174049 523481
rect 174105 523479 174129 523481
rect 174185 523479 174209 523481
rect 174265 523479 174271 523481
rect 173963 523470 174271 523479
rect 177781 523535 178089 523544
rect 177781 523533 177787 523535
rect 177843 523533 177867 523535
rect 177923 523533 177947 523535
rect 178003 523533 178027 523535
rect 178083 523533 178089 523535
rect 177843 523481 177845 523533
rect 178025 523481 178027 523533
rect 177781 523479 177787 523481
rect 177843 523479 177867 523481
rect 177923 523479 177947 523481
rect 178003 523479 178027 523481
rect 178083 523479 178089 523481
rect 177781 523470 178089 523479
rect 174623 522991 174931 523000
rect 174623 522989 174629 522991
rect 174685 522989 174709 522991
rect 174765 522989 174789 522991
rect 174845 522989 174869 522991
rect 174925 522989 174931 522991
rect 174685 522937 174687 522989
rect 174867 522937 174869 522989
rect 174623 522935 174629 522937
rect 174685 522935 174709 522937
rect 174765 522935 174789 522937
rect 174845 522935 174869 522937
rect 174925 522935 174931 522937
rect 174623 522926 174931 522935
rect 173963 522447 174271 522456
rect 173963 522445 173969 522447
rect 174025 522445 174049 522447
rect 174105 522445 174129 522447
rect 174185 522445 174209 522447
rect 174265 522445 174271 522447
rect 174025 522393 174027 522445
rect 174207 522393 174209 522445
rect 173963 522391 173969 522393
rect 174025 522391 174049 522393
rect 174105 522391 174129 522393
rect 174185 522391 174209 522393
rect 174265 522391 174271 522393
rect 173963 522382 174271 522391
rect 177781 522447 178089 522456
rect 177781 522445 177787 522447
rect 177843 522445 177867 522447
rect 177923 522445 177947 522447
rect 178003 522445 178027 522447
rect 178083 522445 178089 522447
rect 177843 522393 177845 522445
rect 178025 522393 178027 522445
rect 177781 522391 177787 522393
rect 177843 522391 177867 522393
rect 177923 522391 177947 522393
rect 178003 522391 178027 522393
rect 178083 522391 178089 522393
rect 177781 522382 178089 522391
rect 174623 521903 174931 521912
rect 174623 521901 174629 521903
rect 174685 521901 174709 521903
rect 174765 521901 174789 521903
rect 174845 521901 174869 521903
rect 174925 521901 174931 521903
rect 174685 521849 174687 521901
rect 174867 521849 174869 521901
rect 174623 521847 174629 521849
rect 174685 521847 174709 521849
rect 174765 521847 174789 521849
rect 174845 521847 174869 521849
rect 174925 521847 174931 521849
rect 174623 521838 174931 521847
rect 173963 521359 174271 521368
rect 173963 521357 173969 521359
rect 174025 521357 174049 521359
rect 174105 521357 174129 521359
rect 174185 521357 174209 521359
rect 174265 521357 174271 521359
rect 174025 521305 174027 521357
rect 174207 521305 174209 521357
rect 173963 521303 173969 521305
rect 174025 521303 174049 521305
rect 174105 521303 174129 521305
rect 174185 521303 174209 521305
rect 174265 521303 174271 521305
rect 173963 521294 174271 521303
rect 177781 521359 178089 521368
rect 177781 521357 177787 521359
rect 177843 521357 177867 521359
rect 177923 521357 177947 521359
rect 178003 521357 178027 521359
rect 178083 521357 178089 521359
rect 177843 521305 177845 521357
rect 178025 521305 178027 521357
rect 177781 521303 177787 521305
rect 177843 521303 177867 521305
rect 177923 521303 177947 521305
rect 178003 521303 178027 521305
rect 178083 521303 178089 521305
rect 177781 521294 178089 521303
rect 174623 520815 174931 520824
rect 174623 520813 174629 520815
rect 174685 520813 174709 520815
rect 174765 520813 174789 520815
rect 174845 520813 174869 520815
rect 174925 520813 174931 520815
rect 174685 520761 174687 520813
rect 174867 520761 174869 520813
rect 174623 520759 174629 520761
rect 174685 520759 174709 520761
rect 174765 520759 174789 520761
rect 174845 520759 174869 520761
rect 174925 520759 174931 520761
rect 174623 520750 174931 520759
rect 173963 520271 174271 520280
rect 173963 520269 173969 520271
rect 174025 520269 174049 520271
rect 174105 520269 174129 520271
rect 174185 520269 174209 520271
rect 174265 520269 174271 520271
rect 174025 520217 174027 520269
rect 174207 520217 174209 520269
rect 173963 520215 173969 520217
rect 174025 520215 174049 520217
rect 174105 520215 174129 520217
rect 174185 520215 174209 520217
rect 174265 520215 174271 520217
rect 173963 520206 174271 520215
rect 177781 520271 178089 520280
rect 177781 520269 177787 520271
rect 177843 520269 177867 520271
rect 177923 520269 177947 520271
rect 178003 520269 178027 520271
rect 178083 520269 178089 520271
rect 177843 520217 177845 520269
rect 178025 520217 178027 520269
rect 177781 520215 177787 520217
rect 177843 520215 177867 520217
rect 177923 520215 177947 520217
rect 178003 520215 178027 520217
rect 178083 520215 178089 520217
rect 177781 520206 178089 520215
rect 174623 519727 174931 519736
rect 174623 519725 174629 519727
rect 174685 519725 174709 519727
rect 174765 519725 174789 519727
rect 174845 519725 174869 519727
rect 174925 519725 174931 519727
rect 174685 519673 174687 519725
rect 174867 519673 174869 519725
rect 174623 519671 174629 519673
rect 174685 519671 174709 519673
rect 174765 519671 174789 519673
rect 174845 519671 174869 519673
rect 174925 519671 174931 519673
rect 174623 519662 174931 519671
rect 173963 519183 174271 519192
rect 173963 519181 173969 519183
rect 174025 519181 174049 519183
rect 174105 519181 174129 519183
rect 174185 519181 174209 519183
rect 174265 519181 174271 519183
rect 174025 519129 174027 519181
rect 174207 519129 174209 519181
rect 173963 519127 173969 519129
rect 174025 519127 174049 519129
rect 174105 519127 174129 519129
rect 174185 519127 174209 519129
rect 174265 519127 174271 519129
rect 173963 519118 174271 519127
rect 177781 519183 178089 519192
rect 177781 519181 177787 519183
rect 177843 519181 177867 519183
rect 177923 519181 177947 519183
rect 178003 519181 178027 519183
rect 178083 519181 178089 519183
rect 177843 519129 177845 519181
rect 178025 519129 178027 519181
rect 177781 519127 177787 519129
rect 177843 519127 177867 519129
rect 177923 519127 177947 519129
rect 178003 519127 178027 519129
rect 178083 519127 178089 519129
rect 177781 519118 178089 519127
rect 174623 518639 174931 518648
rect 174623 518637 174629 518639
rect 174685 518637 174709 518639
rect 174765 518637 174789 518639
rect 174845 518637 174869 518639
rect 174925 518637 174931 518639
rect 174685 518585 174687 518637
rect 174867 518585 174869 518637
rect 174623 518583 174629 518585
rect 174685 518583 174709 518585
rect 174765 518583 174789 518585
rect 174845 518583 174869 518585
rect 174925 518583 174931 518585
rect 174623 518574 174931 518583
rect 173963 518095 174271 518104
rect 173963 518093 173969 518095
rect 174025 518093 174049 518095
rect 174105 518093 174129 518095
rect 174185 518093 174209 518095
rect 174265 518093 174271 518095
rect 174025 518041 174027 518093
rect 174207 518041 174209 518093
rect 173963 518039 173969 518041
rect 174025 518039 174049 518041
rect 174105 518039 174129 518041
rect 174185 518039 174209 518041
rect 174265 518039 174271 518041
rect 173963 518030 174271 518039
rect 177781 518095 178089 518104
rect 177781 518093 177787 518095
rect 177843 518093 177867 518095
rect 177923 518093 177947 518095
rect 178003 518093 178027 518095
rect 178083 518093 178089 518095
rect 177843 518041 177845 518093
rect 178025 518041 178027 518093
rect 177781 518039 177787 518041
rect 177843 518039 177867 518041
rect 177923 518039 177947 518041
rect 178003 518039 178027 518041
rect 178083 518039 178089 518041
rect 177781 518030 178089 518039
rect 174623 517551 174931 517560
rect 174623 517549 174629 517551
rect 174685 517549 174709 517551
rect 174765 517549 174789 517551
rect 174845 517549 174869 517551
rect 174925 517549 174931 517551
rect 174685 517497 174687 517549
rect 174867 517497 174869 517549
rect 174623 517495 174629 517497
rect 174685 517495 174709 517497
rect 174765 517495 174789 517497
rect 174845 517495 174869 517497
rect 174925 517495 174931 517497
rect 174623 517486 174931 517495
rect 178312 517453 178340 528593
rect 178392 528541 178444 528547
rect 178441 528431 178749 528440
rect 178441 528429 178447 528431
rect 178503 528429 178527 528431
rect 178583 528429 178607 528431
rect 178663 528429 178687 528431
rect 178743 528429 178749 528431
rect 178503 528377 178505 528429
rect 178685 528377 178687 528429
rect 178441 528375 178447 528377
rect 178503 528375 178527 528377
rect 178583 528375 178607 528377
rect 178663 528375 178687 528377
rect 178743 528375 178749 528377
rect 178441 528366 178749 528375
rect 178956 528333 178984 530309
rect 179232 530253 179260 530309
rect 179232 530225 179352 530253
rect 179324 529829 179352 530225
rect 179508 529965 179536 530445
rect 180692 530299 180744 530305
rect 180692 530241 180744 530247
rect 179680 530163 179732 530169
rect 179680 530105 179732 530111
rect 179496 529959 179548 529965
rect 179496 529901 179548 529907
rect 179312 529823 179364 529829
rect 179312 529765 179364 529771
rect 179324 529081 179352 529765
rect 179312 529075 179364 529081
rect 179312 529017 179364 529023
rect 179324 528333 179352 529017
rect 178944 528327 178996 528333
rect 178944 528269 178996 528275
rect 179312 528327 179364 528333
rect 179312 528269 179364 528275
rect 178944 527987 178996 527993
rect 178944 527929 178996 527935
rect 178956 527789 178984 527929
rect 178944 527783 178996 527789
rect 178944 527725 178996 527731
rect 179508 527653 179536 529901
rect 179692 529285 179720 530105
rect 179864 529823 179916 529829
rect 179864 529765 179916 529771
rect 179876 529421 179904 529765
rect 180508 529619 180560 529625
rect 180508 529561 180560 529567
rect 179864 529415 179916 529421
rect 179864 529357 179916 529363
rect 179680 529279 179732 529285
rect 179680 529221 179732 529227
rect 180520 529081 180548 529561
rect 179680 529075 179732 529081
rect 179680 529017 179732 529023
rect 180508 529075 180560 529081
rect 180508 529017 180560 529023
rect 179692 528877 179720 529017
rect 179680 528871 179732 528877
rect 179680 528813 179732 528819
rect 180520 528741 180548 529017
rect 180508 528735 180560 528741
rect 180508 528677 180560 528683
rect 180704 528129 180732 530241
rect 180888 529965 180916 531955
rect 182259 530607 182567 530616
rect 182259 530605 182265 530607
rect 182321 530605 182345 530607
rect 182401 530605 182425 530607
rect 182481 530605 182505 530607
rect 182561 530605 182567 530607
rect 182321 530553 182323 530605
rect 182503 530553 182505 530605
rect 182259 530551 182265 530553
rect 182321 530551 182345 530553
rect 182401 530551 182425 530553
rect 182481 530551 182505 530553
rect 182561 530551 182567 530553
rect 182259 530542 182567 530551
rect 183004 530509 183032 531955
rect 185120 530509 185148 531955
rect 187236 531477 187264 531955
rect 187144 531449 187264 531477
rect 186077 530607 186385 530616
rect 186077 530605 186083 530607
rect 186139 530605 186163 530607
rect 186219 530605 186243 530607
rect 186299 530605 186323 530607
rect 186379 530605 186385 530607
rect 186139 530553 186141 530605
rect 186321 530553 186323 530605
rect 186077 530551 186083 530553
rect 186139 530551 186163 530553
rect 186219 530551 186243 530553
rect 186299 530551 186323 530553
rect 186379 530551 186385 530553
rect 186077 530542 186385 530551
rect 182992 530503 183044 530509
rect 182992 530445 183044 530451
rect 185108 530503 185160 530509
rect 185108 530445 185160 530451
rect 187144 530373 187172 531449
rect 182256 530367 182308 530373
rect 182256 530309 182308 530315
rect 183176 530367 183228 530373
rect 183176 530309 183228 530315
rect 187132 530367 187184 530373
rect 187132 530309 187184 530315
rect 182164 530163 182216 530169
rect 182164 530105 182216 530111
rect 181599 530063 181907 530072
rect 181599 530061 181605 530063
rect 181661 530061 181685 530063
rect 181741 530061 181765 530063
rect 181821 530061 181845 530063
rect 181901 530061 181907 530063
rect 181661 530009 181663 530061
rect 181843 530009 181845 530061
rect 181599 530007 181605 530009
rect 181661 530007 181685 530009
rect 181741 530007 181765 530009
rect 181821 530007 181845 530009
rect 181901 530007 181907 530009
rect 181599 529998 181907 530007
rect 182176 529965 182204 530105
rect 180876 529959 180928 529965
rect 180876 529901 180928 529907
rect 182164 529959 182216 529965
rect 182164 529901 182216 529907
rect 181520 529687 181572 529693
rect 181520 529629 181572 529635
rect 181532 529285 181560 529629
rect 181796 529619 181848 529625
rect 182268 529607 182296 530309
rect 182624 530299 182676 530305
rect 182624 530241 182676 530247
rect 182636 529965 182664 530241
rect 182716 530163 182768 530169
rect 182716 530105 182768 530111
rect 182624 529959 182676 529965
rect 182624 529901 182676 529907
rect 181796 529561 181848 529567
rect 182176 529579 182296 529607
rect 181808 529421 181836 529561
rect 181796 529415 181848 529421
rect 181796 529357 181848 529363
rect 181520 529279 181572 529285
rect 181520 529221 181572 529227
rect 181532 528741 181560 529221
rect 181599 528975 181907 528984
rect 181599 528973 181605 528975
rect 181661 528973 181685 528975
rect 181741 528973 181765 528975
rect 181821 528973 181845 528975
rect 181901 528973 181907 528975
rect 181661 528921 181663 528973
rect 181843 528921 181845 528973
rect 181599 528919 181605 528921
rect 181661 528919 181685 528921
rect 181741 528919 181765 528921
rect 181821 528919 181845 528921
rect 181901 528919 181907 528921
rect 181599 528910 181907 528919
rect 182176 528877 182204 529579
rect 182259 529519 182567 529528
rect 182259 529517 182265 529519
rect 182321 529517 182345 529519
rect 182401 529517 182425 529519
rect 182481 529517 182505 529519
rect 182561 529517 182567 529519
rect 182321 529465 182323 529517
rect 182503 529465 182505 529517
rect 182259 529463 182265 529465
rect 182321 529463 182345 529465
rect 182401 529463 182425 529465
rect 182481 529463 182505 529465
rect 182561 529463 182567 529465
rect 182259 529454 182567 529463
rect 182728 529285 182756 530105
rect 183188 529829 183216 530309
rect 185417 530063 185725 530072
rect 185417 530061 185423 530063
rect 185479 530061 185503 530063
rect 185559 530061 185583 530063
rect 185639 530061 185663 530063
rect 185719 530061 185725 530063
rect 185479 530009 185481 530061
rect 185661 530009 185663 530061
rect 185417 530007 185423 530009
rect 185479 530007 185503 530009
rect 185559 530007 185583 530009
rect 185639 530007 185663 530009
rect 185719 530007 185725 530009
rect 185417 529998 185725 530007
rect 183176 529823 183228 529829
rect 183176 529765 183228 529771
rect 186077 529519 186385 529528
rect 186077 529517 186083 529519
rect 186139 529517 186163 529519
rect 186219 529517 186243 529519
rect 186299 529517 186323 529519
rect 186379 529517 186385 529519
rect 186139 529465 186141 529517
rect 186321 529465 186323 529517
rect 186077 529463 186083 529465
rect 186139 529463 186163 529465
rect 186219 529463 186243 529465
rect 186299 529463 186323 529465
rect 186379 529463 186385 529465
rect 186077 529454 186385 529463
rect 182716 529279 182768 529285
rect 182716 529221 182768 529227
rect 185417 528975 185725 528984
rect 185417 528973 185423 528975
rect 185479 528973 185503 528975
rect 185559 528973 185583 528975
rect 185639 528973 185663 528975
rect 185719 528973 185725 528975
rect 185479 528921 185481 528973
rect 185661 528921 185663 528973
rect 185417 528919 185423 528921
rect 185479 528919 185503 528921
rect 185559 528919 185583 528921
rect 185639 528919 185663 528921
rect 185719 528919 185725 528921
rect 185417 528910 185725 528919
rect 182164 528871 182216 528877
rect 182164 528813 182216 528819
rect 181520 528735 181572 528741
rect 181520 528677 181572 528683
rect 180968 528531 181020 528537
rect 180968 528473 181020 528479
rect 180980 528333 181008 528473
rect 182176 528333 182204 528813
rect 186580 528599 186632 528605
rect 186580 528541 186632 528547
rect 182259 528431 182567 528440
rect 182259 528429 182265 528431
rect 182321 528429 182345 528431
rect 182401 528429 182425 528431
rect 182481 528429 182505 528431
rect 182561 528429 182567 528431
rect 182321 528377 182323 528429
rect 182503 528377 182505 528429
rect 182259 528375 182265 528377
rect 182321 528375 182345 528377
rect 182401 528375 182425 528377
rect 182481 528375 182505 528377
rect 182561 528375 182567 528377
rect 182259 528366 182567 528375
rect 186077 528431 186385 528440
rect 186077 528429 186083 528431
rect 186139 528429 186163 528431
rect 186219 528429 186243 528431
rect 186299 528429 186323 528431
rect 186379 528429 186385 528431
rect 186139 528377 186141 528429
rect 186321 528377 186323 528429
rect 186077 528375 186083 528377
rect 186139 528375 186163 528377
rect 186219 528375 186243 528377
rect 186299 528375 186323 528377
rect 186379 528375 186385 528377
rect 186077 528366 186385 528375
rect 180968 528327 181020 528333
rect 180968 528269 181020 528275
rect 182164 528327 182216 528333
rect 182164 528269 182216 528275
rect 181336 528191 181388 528197
rect 181336 528133 181388 528139
rect 180692 528123 180744 528129
rect 180692 528065 180744 528071
rect 179496 527647 179548 527653
rect 179496 527589 179548 527595
rect 178441 527343 178749 527352
rect 178441 527341 178447 527343
rect 178503 527341 178527 527343
rect 178583 527341 178607 527343
rect 178663 527341 178687 527343
rect 178743 527341 178749 527343
rect 178503 527289 178505 527341
rect 178685 527289 178687 527341
rect 178441 527287 178447 527289
rect 178503 527287 178527 527289
rect 178583 527287 178607 527289
rect 178663 527287 178687 527289
rect 178743 527287 178749 527289
rect 178441 527278 178749 527287
rect 178441 526255 178749 526264
rect 178441 526253 178447 526255
rect 178503 526253 178527 526255
rect 178583 526253 178607 526255
rect 178663 526253 178687 526255
rect 178743 526253 178749 526255
rect 178503 526201 178505 526253
rect 178685 526201 178687 526253
rect 178441 526199 178447 526201
rect 178503 526199 178527 526201
rect 178583 526199 178607 526201
rect 178663 526199 178687 526201
rect 178743 526199 178749 526201
rect 178441 526190 178749 526199
rect 178441 525167 178749 525176
rect 178441 525165 178447 525167
rect 178503 525165 178527 525167
rect 178583 525165 178607 525167
rect 178663 525165 178687 525167
rect 178743 525165 178749 525167
rect 178503 525113 178505 525165
rect 178685 525113 178687 525165
rect 178441 525111 178447 525113
rect 178503 525111 178527 525113
rect 178583 525111 178607 525113
rect 178663 525111 178687 525113
rect 178743 525111 178749 525113
rect 178441 525102 178749 525111
rect 178441 524079 178749 524088
rect 178441 524077 178447 524079
rect 178503 524077 178527 524079
rect 178583 524077 178607 524079
rect 178663 524077 178687 524079
rect 178743 524077 178749 524079
rect 178503 524025 178505 524077
rect 178685 524025 178687 524077
rect 178441 524023 178447 524025
rect 178503 524023 178527 524025
rect 178583 524023 178607 524025
rect 178663 524023 178687 524025
rect 178743 524023 178749 524025
rect 178441 524014 178749 524023
rect 178441 522991 178749 523000
rect 178441 522989 178447 522991
rect 178503 522989 178527 522991
rect 178583 522989 178607 522991
rect 178663 522989 178687 522991
rect 178743 522989 178749 522991
rect 178503 522937 178505 522989
rect 178685 522937 178687 522989
rect 178441 522935 178447 522937
rect 178503 522935 178527 522937
rect 178583 522935 178607 522937
rect 178663 522935 178687 522937
rect 178743 522935 178749 522937
rect 178441 522926 178749 522935
rect 178441 521903 178749 521912
rect 178441 521901 178447 521903
rect 178503 521901 178527 521903
rect 178583 521901 178607 521903
rect 178663 521901 178687 521903
rect 178743 521901 178749 521903
rect 178503 521849 178505 521901
rect 178685 521849 178687 521901
rect 178441 521847 178447 521849
rect 178503 521847 178527 521849
rect 178583 521847 178607 521849
rect 178663 521847 178687 521849
rect 178743 521847 178749 521849
rect 178441 521838 178749 521847
rect 178441 520815 178749 520824
rect 178441 520813 178447 520815
rect 178503 520813 178527 520815
rect 178583 520813 178607 520815
rect 178663 520813 178687 520815
rect 178743 520813 178749 520815
rect 178503 520761 178505 520813
rect 178685 520761 178687 520813
rect 178441 520759 178447 520761
rect 178503 520759 178527 520761
rect 178583 520759 178607 520761
rect 178663 520759 178687 520761
rect 178743 520759 178749 520761
rect 178441 520750 178749 520759
rect 178441 519727 178749 519736
rect 178441 519725 178447 519727
rect 178503 519725 178527 519727
rect 178583 519725 178607 519727
rect 178663 519725 178687 519727
rect 178743 519725 178749 519727
rect 178503 519673 178505 519725
rect 178685 519673 178687 519725
rect 178441 519671 178447 519673
rect 178503 519671 178527 519673
rect 178583 519671 178607 519673
rect 178663 519671 178687 519673
rect 178743 519671 178749 519673
rect 178441 519662 178749 519671
rect 178441 518639 178749 518648
rect 178441 518637 178447 518639
rect 178503 518637 178527 518639
rect 178583 518637 178607 518639
rect 178663 518637 178687 518639
rect 178743 518637 178749 518639
rect 178503 518585 178505 518637
rect 178685 518585 178687 518637
rect 178441 518583 178447 518585
rect 178503 518583 178527 518585
rect 178583 518583 178607 518585
rect 178663 518583 178687 518585
rect 178743 518583 178749 518585
rect 178441 518574 178749 518583
rect 178441 517551 178749 517560
rect 178441 517549 178447 517551
rect 178503 517549 178527 517551
rect 178583 517549 178607 517551
rect 178663 517549 178687 517551
rect 178743 517549 178749 517551
rect 178503 517497 178505 517549
rect 178685 517497 178687 517549
rect 178441 517495 178447 517497
rect 178503 517495 178527 517497
rect 178583 517495 178607 517497
rect 178663 517495 178687 517497
rect 178743 517495 178749 517497
rect 178441 517486 178749 517495
rect 177656 517447 177708 517453
rect 177656 517389 177708 517395
rect 178300 517447 178352 517453
rect 178300 517389 178352 517395
rect 173963 517007 174271 517016
rect 173963 517005 173969 517007
rect 174025 517005 174049 517007
rect 174105 517005 174129 517007
rect 174185 517005 174209 517007
rect 174265 517005 174271 517007
rect 174025 516953 174027 517005
rect 174207 516953 174209 517005
rect 173963 516951 173969 516953
rect 174025 516951 174049 516953
rect 174105 516951 174129 516953
rect 174185 516951 174209 516953
rect 174265 516951 174271 516953
rect 173963 516942 174271 516951
rect 174623 516463 174931 516472
rect 174623 516461 174629 516463
rect 174685 516461 174709 516463
rect 174765 516461 174789 516463
rect 174845 516461 174869 516463
rect 174925 516461 174931 516463
rect 174685 516409 174687 516461
rect 174867 516409 174869 516461
rect 174623 516407 174629 516409
rect 174685 516407 174709 516409
rect 174765 516407 174789 516409
rect 174845 516407 174869 516409
rect 174925 516407 174931 516409
rect 174623 516398 174931 516407
rect 173963 515919 174271 515928
rect 173963 515917 173969 515919
rect 174025 515917 174049 515919
rect 174105 515917 174129 515919
rect 174185 515917 174209 515919
rect 174265 515917 174271 515919
rect 174025 515865 174027 515917
rect 174207 515865 174209 515917
rect 173963 515863 173969 515865
rect 174025 515863 174049 515865
rect 174105 515863 174129 515865
rect 174185 515863 174209 515865
rect 174265 515863 174271 515865
rect 173963 515854 174271 515863
rect 173608 515815 173660 515821
rect 173608 515757 173660 515763
rect 173332 515543 173384 515549
rect 173332 515485 173384 515491
rect 173344 513899 173372 515485
rect 174623 515375 174931 515384
rect 174623 515373 174629 515375
rect 174685 515373 174709 515375
rect 174765 515373 174789 515375
rect 174845 515373 174869 515375
rect 174925 515373 174931 515375
rect 174685 515321 174687 515373
rect 174867 515321 174869 515373
rect 174623 515319 174629 515321
rect 174685 515319 174709 515321
rect 174765 515319 174789 515321
rect 174845 515319 174869 515321
rect 174925 515319 174931 515321
rect 174623 515310 174931 515319
rect 177668 513899 177696 517389
rect 177781 517007 178089 517016
rect 177781 517005 177787 517007
rect 177843 517005 177867 517007
rect 177923 517005 177947 517007
rect 178003 517005 178027 517007
rect 178083 517005 178089 517007
rect 177843 516953 177845 517005
rect 178025 516953 178027 517005
rect 177781 516951 177787 516953
rect 177843 516951 177867 516953
rect 177923 516951 177947 516953
rect 178003 516951 178027 516953
rect 178083 516951 178089 516953
rect 177781 516942 178089 516951
rect 178441 516463 178749 516472
rect 178441 516461 178447 516463
rect 178503 516461 178527 516463
rect 178583 516461 178607 516463
rect 178663 516461 178687 516463
rect 178743 516461 178749 516463
rect 178503 516409 178505 516461
rect 178685 516409 178687 516461
rect 178441 516407 178447 516409
rect 178503 516407 178527 516409
rect 178583 516407 178607 516409
rect 178663 516407 178687 516409
rect 178743 516407 178749 516409
rect 178441 516398 178749 516407
rect 177781 515919 178089 515928
rect 177781 515917 177787 515919
rect 177843 515917 177867 515919
rect 177923 515917 177947 515919
rect 178003 515917 178027 515919
rect 178083 515917 178089 515919
rect 177843 515865 177845 515917
rect 178025 515865 178027 515917
rect 177781 515863 177787 515865
rect 177843 515863 177867 515865
rect 177923 515863 177947 515865
rect 178003 515863 178027 515865
rect 178083 515863 178089 515865
rect 177781 515854 178089 515863
rect 181348 515821 181376 528133
rect 181599 527887 181907 527896
rect 181599 527885 181605 527887
rect 181661 527885 181685 527887
rect 181741 527885 181765 527887
rect 181821 527885 181845 527887
rect 181901 527885 181907 527887
rect 181661 527833 181663 527885
rect 181843 527833 181845 527885
rect 181599 527831 181605 527833
rect 181661 527831 181685 527833
rect 181741 527831 181765 527833
rect 181821 527831 181845 527833
rect 181901 527831 181907 527833
rect 181599 527822 181907 527831
rect 185417 527887 185725 527896
rect 185417 527885 185423 527887
rect 185479 527885 185503 527887
rect 185559 527885 185583 527887
rect 185639 527885 185663 527887
rect 185719 527885 185725 527887
rect 185479 527833 185481 527885
rect 185661 527833 185663 527885
rect 185417 527831 185423 527833
rect 185479 527831 185503 527833
rect 185559 527831 185583 527833
rect 185639 527831 185663 527833
rect 185719 527831 185725 527833
rect 185417 527822 185725 527831
rect 182259 527343 182567 527352
rect 182259 527341 182265 527343
rect 182321 527341 182345 527343
rect 182401 527341 182425 527343
rect 182481 527341 182505 527343
rect 182561 527341 182567 527343
rect 182321 527289 182323 527341
rect 182503 527289 182505 527341
rect 182259 527287 182265 527289
rect 182321 527287 182345 527289
rect 182401 527287 182425 527289
rect 182481 527287 182505 527289
rect 182561 527287 182567 527289
rect 182259 527278 182567 527287
rect 186077 527343 186385 527352
rect 186077 527341 186083 527343
rect 186139 527341 186163 527343
rect 186219 527341 186243 527343
rect 186299 527341 186323 527343
rect 186379 527341 186385 527343
rect 186139 527289 186141 527341
rect 186321 527289 186323 527341
rect 186077 527287 186083 527289
rect 186139 527287 186163 527289
rect 186219 527287 186243 527289
rect 186299 527287 186323 527289
rect 186379 527287 186385 527289
rect 186077 527278 186385 527287
rect 181599 526799 181907 526808
rect 181599 526797 181605 526799
rect 181661 526797 181685 526799
rect 181741 526797 181765 526799
rect 181821 526797 181845 526799
rect 181901 526797 181907 526799
rect 181661 526745 181663 526797
rect 181843 526745 181845 526797
rect 181599 526743 181605 526745
rect 181661 526743 181685 526745
rect 181741 526743 181765 526745
rect 181821 526743 181845 526745
rect 181901 526743 181907 526745
rect 181599 526734 181907 526743
rect 185417 526799 185725 526808
rect 185417 526797 185423 526799
rect 185479 526797 185503 526799
rect 185559 526797 185583 526799
rect 185639 526797 185663 526799
rect 185719 526797 185725 526799
rect 185479 526745 185481 526797
rect 185661 526745 185663 526797
rect 185417 526743 185423 526745
rect 185479 526743 185503 526745
rect 185559 526743 185583 526745
rect 185639 526743 185663 526745
rect 185719 526743 185725 526745
rect 185417 526734 185725 526743
rect 182259 526255 182567 526264
rect 182259 526253 182265 526255
rect 182321 526253 182345 526255
rect 182401 526253 182425 526255
rect 182481 526253 182505 526255
rect 182561 526253 182567 526255
rect 182321 526201 182323 526253
rect 182503 526201 182505 526253
rect 182259 526199 182265 526201
rect 182321 526199 182345 526201
rect 182401 526199 182425 526201
rect 182481 526199 182505 526201
rect 182561 526199 182567 526201
rect 182259 526190 182567 526199
rect 186077 526255 186385 526264
rect 186077 526253 186083 526255
rect 186139 526253 186163 526255
rect 186219 526253 186243 526255
rect 186299 526253 186323 526255
rect 186379 526253 186385 526255
rect 186139 526201 186141 526253
rect 186321 526201 186323 526253
rect 186077 526199 186083 526201
rect 186139 526199 186163 526201
rect 186219 526199 186243 526201
rect 186299 526199 186323 526201
rect 186379 526199 186385 526201
rect 186077 526190 186385 526199
rect 181599 525711 181907 525720
rect 181599 525709 181605 525711
rect 181661 525709 181685 525711
rect 181741 525709 181765 525711
rect 181821 525709 181845 525711
rect 181901 525709 181907 525711
rect 181661 525657 181663 525709
rect 181843 525657 181845 525709
rect 181599 525655 181605 525657
rect 181661 525655 181685 525657
rect 181741 525655 181765 525657
rect 181821 525655 181845 525657
rect 181901 525655 181907 525657
rect 181599 525646 181907 525655
rect 185417 525711 185725 525720
rect 185417 525709 185423 525711
rect 185479 525709 185503 525711
rect 185559 525709 185583 525711
rect 185639 525709 185663 525711
rect 185719 525709 185725 525711
rect 185479 525657 185481 525709
rect 185661 525657 185663 525709
rect 185417 525655 185423 525657
rect 185479 525655 185503 525657
rect 185559 525655 185583 525657
rect 185639 525655 185663 525657
rect 185719 525655 185725 525657
rect 185417 525646 185725 525655
rect 182259 525167 182567 525176
rect 182259 525165 182265 525167
rect 182321 525165 182345 525167
rect 182401 525165 182425 525167
rect 182481 525165 182505 525167
rect 182561 525165 182567 525167
rect 182321 525113 182323 525165
rect 182503 525113 182505 525165
rect 182259 525111 182265 525113
rect 182321 525111 182345 525113
rect 182401 525111 182425 525113
rect 182481 525111 182505 525113
rect 182561 525111 182567 525113
rect 182259 525102 182567 525111
rect 186077 525167 186385 525176
rect 186077 525165 186083 525167
rect 186139 525165 186163 525167
rect 186219 525165 186243 525167
rect 186299 525165 186323 525167
rect 186379 525165 186385 525167
rect 186139 525113 186141 525165
rect 186321 525113 186323 525165
rect 186077 525111 186083 525113
rect 186139 525111 186163 525113
rect 186219 525111 186243 525113
rect 186299 525111 186323 525113
rect 186379 525111 186385 525113
rect 186077 525102 186385 525111
rect 181599 524623 181907 524632
rect 181599 524621 181605 524623
rect 181661 524621 181685 524623
rect 181741 524621 181765 524623
rect 181821 524621 181845 524623
rect 181901 524621 181907 524623
rect 181661 524569 181663 524621
rect 181843 524569 181845 524621
rect 181599 524567 181605 524569
rect 181661 524567 181685 524569
rect 181741 524567 181765 524569
rect 181821 524567 181845 524569
rect 181901 524567 181907 524569
rect 181599 524558 181907 524567
rect 185417 524623 185725 524632
rect 185417 524621 185423 524623
rect 185479 524621 185503 524623
rect 185559 524621 185583 524623
rect 185639 524621 185663 524623
rect 185719 524621 185725 524623
rect 185479 524569 185481 524621
rect 185661 524569 185663 524621
rect 185417 524567 185423 524569
rect 185479 524567 185503 524569
rect 185559 524567 185583 524569
rect 185639 524567 185663 524569
rect 185719 524567 185725 524569
rect 185417 524558 185725 524567
rect 182259 524079 182567 524088
rect 182259 524077 182265 524079
rect 182321 524077 182345 524079
rect 182401 524077 182425 524079
rect 182481 524077 182505 524079
rect 182561 524077 182567 524079
rect 182321 524025 182323 524077
rect 182503 524025 182505 524077
rect 182259 524023 182265 524025
rect 182321 524023 182345 524025
rect 182401 524023 182425 524025
rect 182481 524023 182505 524025
rect 182561 524023 182567 524025
rect 182259 524014 182567 524023
rect 186077 524079 186385 524088
rect 186077 524077 186083 524079
rect 186139 524077 186163 524079
rect 186219 524077 186243 524079
rect 186299 524077 186323 524079
rect 186379 524077 186385 524079
rect 186139 524025 186141 524077
rect 186321 524025 186323 524077
rect 186077 524023 186083 524025
rect 186139 524023 186163 524025
rect 186219 524023 186243 524025
rect 186299 524023 186323 524025
rect 186379 524023 186385 524025
rect 186077 524014 186385 524023
rect 181599 523535 181907 523544
rect 181599 523533 181605 523535
rect 181661 523533 181685 523535
rect 181741 523533 181765 523535
rect 181821 523533 181845 523535
rect 181901 523533 181907 523535
rect 181661 523481 181663 523533
rect 181843 523481 181845 523533
rect 181599 523479 181605 523481
rect 181661 523479 181685 523481
rect 181741 523479 181765 523481
rect 181821 523479 181845 523481
rect 181901 523479 181907 523481
rect 181599 523470 181907 523479
rect 185417 523535 185725 523544
rect 185417 523533 185423 523535
rect 185479 523533 185503 523535
rect 185559 523533 185583 523535
rect 185639 523533 185663 523535
rect 185719 523533 185725 523535
rect 185479 523481 185481 523533
rect 185661 523481 185663 523533
rect 185417 523479 185423 523481
rect 185479 523479 185503 523481
rect 185559 523479 185583 523481
rect 185639 523479 185663 523481
rect 185719 523479 185725 523481
rect 185417 523470 185725 523479
rect 182259 522991 182567 523000
rect 182259 522989 182265 522991
rect 182321 522989 182345 522991
rect 182401 522989 182425 522991
rect 182481 522989 182505 522991
rect 182561 522989 182567 522991
rect 182321 522937 182323 522989
rect 182503 522937 182505 522989
rect 182259 522935 182265 522937
rect 182321 522935 182345 522937
rect 182401 522935 182425 522937
rect 182481 522935 182505 522937
rect 182561 522935 182567 522937
rect 182259 522926 182567 522935
rect 186077 522991 186385 523000
rect 186077 522989 186083 522991
rect 186139 522989 186163 522991
rect 186219 522989 186243 522991
rect 186299 522989 186323 522991
rect 186379 522989 186385 522991
rect 186139 522937 186141 522989
rect 186321 522937 186323 522989
rect 186077 522935 186083 522937
rect 186139 522935 186163 522937
rect 186219 522935 186243 522937
rect 186299 522935 186323 522937
rect 186379 522935 186385 522937
rect 186077 522926 186385 522935
rect 181599 522447 181907 522456
rect 181599 522445 181605 522447
rect 181661 522445 181685 522447
rect 181741 522445 181765 522447
rect 181821 522445 181845 522447
rect 181901 522445 181907 522447
rect 181661 522393 181663 522445
rect 181843 522393 181845 522445
rect 181599 522391 181605 522393
rect 181661 522391 181685 522393
rect 181741 522391 181765 522393
rect 181821 522391 181845 522393
rect 181901 522391 181907 522393
rect 181599 522382 181907 522391
rect 185417 522447 185725 522456
rect 185417 522445 185423 522447
rect 185479 522445 185503 522447
rect 185559 522445 185583 522447
rect 185639 522445 185663 522447
rect 185719 522445 185725 522447
rect 185479 522393 185481 522445
rect 185661 522393 185663 522445
rect 185417 522391 185423 522393
rect 185479 522391 185503 522393
rect 185559 522391 185583 522393
rect 185639 522391 185663 522393
rect 185719 522391 185725 522393
rect 185417 522382 185725 522391
rect 182259 521903 182567 521912
rect 182259 521901 182265 521903
rect 182321 521901 182345 521903
rect 182401 521901 182425 521903
rect 182481 521901 182505 521903
rect 182561 521901 182567 521903
rect 182321 521849 182323 521901
rect 182503 521849 182505 521901
rect 182259 521847 182265 521849
rect 182321 521847 182345 521849
rect 182401 521847 182425 521849
rect 182481 521847 182505 521849
rect 182561 521847 182567 521849
rect 182259 521838 182567 521847
rect 186077 521903 186385 521912
rect 186077 521901 186083 521903
rect 186139 521901 186163 521903
rect 186219 521901 186243 521903
rect 186299 521901 186323 521903
rect 186379 521901 186385 521903
rect 186139 521849 186141 521901
rect 186321 521849 186323 521901
rect 186077 521847 186083 521849
rect 186139 521847 186163 521849
rect 186219 521847 186243 521849
rect 186299 521847 186323 521849
rect 186379 521847 186385 521849
rect 186077 521838 186385 521847
rect 181599 521359 181907 521368
rect 181599 521357 181605 521359
rect 181661 521357 181685 521359
rect 181741 521357 181765 521359
rect 181821 521357 181845 521359
rect 181901 521357 181907 521359
rect 181661 521305 181663 521357
rect 181843 521305 181845 521357
rect 181599 521303 181605 521305
rect 181661 521303 181685 521305
rect 181741 521303 181765 521305
rect 181821 521303 181845 521305
rect 181901 521303 181907 521305
rect 181599 521294 181907 521303
rect 185417 521359 185725 521368
rect 185417 521357 185423 521359
rect 185479 521357 185503 521359
rect 185559 521357 185583 521359
rect 185639 521357 185663 521359
rect 185719 521357 185725 521359
rect 185479 521305 185481 521357
rect 185661 521305 185663 521357
rect 185417 521303 185423 521305
rect 185479 521303 185503 521305
rect 185559 521303 185583 521305
rect 185639 521303 185663 521305
rect 185719 521303 185725 521305
rect 185417 521294 185725 521303
rect 182259 520815 182567 520824
rect 182259 520813 182265 520815
rect 182321 520813 182345 520815
rect 182401 520813 182425 520815
rect 182481 520813 182505 520815
rect 182561 520813 182567 520815
rect 182321 520761 182323 520813
rect 182503 520761 182505 520813
rect 182259 520759 182265 520761
rect 182321 520759 182345 520761
rect 182401 520759 182425 520761
rect 182481 520759 182505 520761
rect 182561 520759 182567 520761
rect 182259 520750 182567 520759
rect 186077 520815 186385 520824
rect 186077 520813 186083 520815
rect 186139 520813 186163 520815
rect 186219 520813 186243 520815
rect 186299 520813 186323 520815
rect 186379 520813 186385 520815
rect 186139 520761 186141 520813
rect 186321 520761 186323 520813
rect 186077 520759 186083 520761
rect 186139 520759 186163 520761
rect 186219 520759 186243 520761
rect 186299 520759 186323 520761
rect 186379 520759 186385 520761
rect 186077 520750 186385 520759
rect 181599 520271 181907 520280
rect 181599 520269 181605 520271
rect 181661 520269 181685 520271
rect 181741 520269 181765 520271
rect 181821 520269 181845 520271
rect 181901 520269 181907 520271
rect 181661 520217 181663 520269
rect 181843 520217 181845 520269
rect 181599 520215 181605 520217
rect 181661 520215 181685 520217
rect 181741 520215 181765 520217
rect 181821 520215 181845 520217
rect 181901 520215 181907 520217
rect 181599 520206 181907 520215
rect 185417 520271 185725 520280
rect 185417 520269 185423 520271
rect 185479 520269 185503 520271
rect 185559 520269 185583 520271
rect 185639 520269 185663 520271
rect 185719 520269 185725 520271
rect 185479 520217 185481 520269
rect 185661 520217 185663 520269
rect 185417 520215 185423 520217
rect 185479 520215 185503 520217
rect 185559 520215 185583 520217
rect 185639 520215 185663 520217
rect 185719 520215 185725 520217
rect 185417 520206 185725 520215
rect 182259 519727 182567 519736
rect 182259 519725 182265 519727
rect 182321 519725 182345 519727
rect 182401 519725 182425 519727
rect 182481 519725 182505 519727
rect 182561 519725 182567 519727
rect 182321 519673 182323 519725
rect 182503 519673 182505 519725
rect 182259 519671 182265 519673
rect 182321 519671 182345 519673
rect 182401 519671 182425 519673
rect 182481 519671 182505 519673
rect 182561 519671 182567 519673
rect 182259 519662 182567 519671
rect 186077 519727 186385 519736
rect 186077 519725 186083 519727
rect 186139 519725 186163 519727
rect 186219 519725 186243 519727
rect 186299 519725 186323 519727
rect 186379 519725 186385 519727
rect 186139 519673 186141 519725
rect 186321 519673 186323 519725
rect 186077 519671 186083 519673
rect 186139 519671 186163 519673
rect 186219 519671 186243 519673
rect 186299 519671 186323 519673
rect 186379 519671 186385 519673
rect 186077 519662 186385 519671
rect 181599 519183 181907 519192
rect 181599 519181 181605 519183
rect 181661 519181 181685 519183
rect 181741 519181 181765 519183
rect 181821 519181 181845 519183
rect 181901 519181 181907 519183
rect 181661 519129 181663 519181
rect 181843 519129 181845 519181
rect 181599 519127 181605 519129
rect 181661 519127 181685 519129
rect 181741 519127 181765 519129
rect 181821 519127 181845 519129
rect 181901 519127 181907 519129
rect 181599 519118 181907 519127
rect 185417 519183 185725 519192
rect 185417 519181 185423 519183
rect 185479 519181 185503 519183
rect 185559 519181 185583 519183
rect 185639 519181 185663 519183
rect 185719 519181 185725 519183
rect 185479 519129 185481 519181
rect 185661 519129 185663 519181
rect 185417 519127 185423 519129
rect 185479 519127 185503 519129
rect 185559 519127 185583 519129
rect 185639 519127 185663 519129
rect 185719 519127 185725 519129
rect 185417 519118 185725 519127
rect 182259 518639 182567 518648
rect 182259 518637 182265 518639
rect 182321 518637 182345 518639
rect 182401 518637 182425 518639
rect 182481 518637 182505 518639
rect 182561 518637 182567 518639
rect 182321 518585 182323 518637
rect 182503 518585 182505 518637
rect 182259 518583 182265 518585
rect 182321 518583 182345 518585
rect 182401 518583 182425 518585
rect 182481 518583 182505 518585
rect 182561 518583 182567 518585
rect 182259 518574 182567 518583
rect 186077 518639 186385 518648
rect 186077 518637 186083 518639
rect 186139 518637 186163 518639
rect 186219 518637 186243 518639
rect 186299 518637 186323 518639
rect 186379 518637 186385 518639
rect 186139 518585 186141 518637
rect 186321 518585 186323 518637
rect 186077 518583 186083 518585
rect 186139 518583 186163 518585
rect 186219 518583 186243 518585
rect 186299 518583 186323 518585
rect 186379 518583 186385 518585
rect 186077 518574 186385 518583
rect 181599 518095 181907 518104
rect 181599 518093 181605 518095
rect 181661 518093 181685 518095
rect 181741 518093 181765 518095
rect 181821 518093 181845 518095
rect 181901 518093 181907 518095
rect 181661 518041 181663 518093
rect 181843 518041 181845 518093
rect 181599 518039 181605 518041
rect 181661 518039 181685 518041
rect 181741 518039 181765 518041
rect 181821 518039 181845 518041
rect 181901 518039 181907 518041
rect 181599 518030 181907 518039
rect 185417 518095 185725 518104
rect 185417 518093 185423 518095
rect 185479 518093 185503 518095
rect 185559 518093 185583 518095
rect 185639 518093 185663 518095
rect 185719 518093 185725 518095
rect 185479 518041 185481 518093
rect 185661 518041 185663 518093
rect 185417 518039 185423 518041
rect 185479 518039 185503 518041
rect 185559 518039 185583 518041
rect 185639 518039 185663 518041
rect 185719 518039 185725 518041
rect 185417 518030 185725 518039
rect 182259 517551 182567 517560
rect 182259 517549 182265 517551
rect 182321 517549 182345 517551
rect 182401 517549 182425 517551
rect 182481 517549 182505 517551
rect 182561 517549 182567 517551
rect 182321 517497 182323 517549
rect 182503 517497 182505 517549
rect 182259 517495 182265 517497
rect 182321 517495 182345 517497
rect 182401 517495 182425 517497
rect 182481 517495 182505 517497
rect 182561 517495 182567 517497
rect 182259 517486 182567 517495
rect 186077 517551 186385 517560
rect 186077 517549 186083 517551
rect 186139 517549 186163 517551
rect 186219 517549 186243 517551
rect 186299 517549 186323 517551
rect 186379 517549 186385 517551
rect 186139 517497 186141 517549
rect 186321 517497 186323 517549
rect 186077 517495 186083 517497
rect 186139 517495 186163 517497
rect 186219 517495 186243 517497
rect 186299 517495 186323 517497
rect 186379 517495 186385 517497
rect 186077 517486 186385 517495
rect 181599 517007 181907 517016
rect 181599 517005 181605 517007
rect 181661 517005 181685 517007
rect 181741 517005 181765 517007
rect 181821 517005 181845 517007
rect 181901 517005 181907 517007
rect 181661 516953 181663 517005
rect 181843 516953 181845 517005
rect 181599 516951 181605 516953
rect 181661 516951 181685 516953
rect 181741 516951 181765 516953
rect 181821 516951 181845 516953
rect 181901 516951 181907 516953
rect 181599 516942 181907 516951
rect 185417 517007 185725 517016
rect 185417 517005 185423 517007
rect 185479 517005 185503 517007
rect 185559 517005 185583 517007
rect 185639 517005 185663 517007
rect 185719 517005 185725 517007
rect 185479 516953 185481 517005
rect 185661 516953 185663 517005
rect 185417 516951 185423 516953
rect 185479 516951 185503 516953
rect 185559 516951 185583 516953
rect 185639 516951 185663 516953
rect 185719 516951 185725 516953
rect 185417 516942 185725 516951
rect 182259 516463 182567 516472
rect 182259 516461 182265 516463
rect 182321 516461 182345 516463
rect 182401 516461 182425 516463
rect 182481 516461 182505 516463
rect 182561 516461 182567 516463
rect 182321 516409 182323 516461
rect 182503 516409 182505 516461
rect 182259 516407 182265 516409
rect 182321 516407 182345 516409
rect 182401 516407 182425 516409
rect 182481 516407 182505 516409
rect 182561 516407 182567 516409
rect 182259 516398 182567 516407
rect 186077 516463 186385 516472
rect 186077 516461 186083 516463
rect 186139 516461 186163 516463
rect 186219 516461 186243 516463
rect 186299 516461 186323 516463
rect 186379 516461 186385 516463
rect 186139 516409 186141 516461
rect 186321 516409 186323 516461
rect 186077 516407 186083 516409
rect 186139 516407 186163 516409
rect 186219 516407 186243 516409
rect 186299 516407 186323 516409
rect 186379 516407 186385 516409
rect 186077 516398 186385 516407
rect 181599 515919 181907 515928
rect 181599 515917 181605 515919
rect 181661 515917 181685 515919
rect 181741 515917 181765 515919
rect 181821 515917 181845 515919
rect 181901 515917 181907 515919
rect 181661 515865 181663 515917
rect 181843 515865 181845 515917
rect 181599 515863 181605 515865
rect 181661 515863 181685 515865
rect 181741 515863 181765 515865
rect 181821 515863 181845 515865
rect 181901 515863 181907 515865
rect 181599 515854 181907 515863
rect 185417 515919 185725 515928
rect 185417 515917 185423 515919
rect 185479 515917 185503 515919
rect 185559 515917 185583 515919
rect 185639 515917 185663 515919
rect 185719 515917 185725 515919
rect 185479 515865 185481 515917
rect 185661 515865 185663 515917
rect 185417 515863 185423 515865
rect 185479 515863 185503 515865
rect 185559 515863 185583 515865
rect 185639 515863 185663 515865
rect 185719 515863 185725 515865
rect 185417 515854 185725 515863
rect 186592 515821 186620 528541
rect 181336 515815 181388 515821
rect 181336 515757 181388 515763
rect 186580 515815 186632 515821
rect 186580 515757 186632 515763
rect 186488 515543 186540 515549
rect 186488 515485 186540 515491
rect 182164 515475 182216 515481
rect 182084 515423 182164 515429
rect 182084 515417 182216 515423
rect 182084 515401 182204 515417
rect 178441 515375 178749 515384
rect 178441 515373 178447 515375
rect 178503 515373 178527 515375
rect 178583 515373 178607 515375
rect 178663 515373 178687 515375
rect 178743 515373 178749 515375
rect 178503 515321 178505 515373
rect 178685 515321 178687 515373
rect 178441 515319 178447 515321
rect 178503 515319 178527 515321
rect 178583 515319 178607 515321
rect 178663 515319 178687 515321
rect 178743 515319 178749 515321
rect 178441 515310 178749 515319
rect 173330 513285 173386 513899
rect 177654 513285 177710 513899
rect 181978 513797 182034 513899
rect 182084 513797 182112 515401
rect 182259 515375 182567 515384
rect 182259 515373 182265 515375
rect 182321 515373 182345 515375
rect 182401 515373 182425 515375
rect 182481 515373 182505 515375
rect 182561 515373 182567 515375
rect 182321 515321 182323 515373
rect 182503 515321 182505 515373
rect 182259 515319 182265 515321
rect 182321 515319 182345 515321
rect 182401 515319 182425 515321
rect 182481 515319 182505 515321
rect 182561 515319 182567 515321
rect 182259 515310 182567 515319
rect 186077 515375 186385 515384
rect 186077 515373 186083 515375
rect 186139 515373 186163 515375
rect 186219 515373 186243 515375
rect 186299 515373 186323 515375
rect 186379 515373 186385 515375
rect 186139 515321 186141 515373
rect 186321 515321 186323 515373
rect 186077 515319 186083 515321
rect 186139 515319 186163 515321
rect 186219 515319 186243 515321
rect 186299 515319 186323 515321
rect 186379 515319 186385 515321
rect 186077 515310 186385 515319
rect 181978 513769 182112 513797
rect 186302 513797 186358 513899
rect 186500 513797 186528 515485
rect 186302 513769 186528 513797
rect 181978 513285 182034 513769
rect 173248 513120 173448 513285
rect 177578 513280 177778 513285
rect 181908 513280 182108 513285
rect 173248 513095 173450 513120
rect 177578 513095 177780 513280
rect 181908 513095 182110 513280
rect 186302 513245 186358 513769
rect 173250 513000 173450 513095
rect 173250 512800 173450 512810
rect 177580 513000 177780 513095
rect 177580 512800 177780 512810
rect 181910 513000 182110 513095
rect 186228 513240 186428 513245
rect 186228 513055 186430 513240
rect 181910 512800 182110 512810
rect 186230 513000 186430 513055
rect 186230 512800 186430 512810
rect 2000 509000 4000 509010
rect 2000 506990 4000 507000
rect 2000 466000 4000 466010
rect 2000 463990 4000 464000
rect 2000 423000 4000 423010
rect 2000 420990 4000 421000
rect 2000 380000 4000 380010
rect 2000 377990 4000 378000
<< via2 >>
rect 18000 699000 20000 701000
rect 70000 699000 72000 701000
rect 122000 699000 124000 701000
rect 3000 682000 5000 684000
rect 159398 538555 159478 538655
rect 161388 538545 161508 538665
rect 163028 538665 163328 538865
rect 166688 540065 166868 540245
rect 166688 539125 166868 539305
rect 170488 540065 170668 540245
rect 170488 539125 170668 539305
rect 174188 540075 174368 540255
rect 174188 539125 174368 539305
rect 177698 540065 177878 540245
rect 177688 539125 177868 539305
rect 181288 540065 181468 540245
rect 181288 539125 181468 539305
rect 184588 540065 184768 540245
rect 184588 539125 184768 539305
rect 187898 540065 188078 540245
rect 187888 539125 188068 539305
rect 191188 540065 191368 540245
rect 191808 540065 191988 540245
rect 191198 539135 191378 539315
rect 191818 539125 191998 539305
rect 160208 535435 160348 535565
rect 160348 535435 160358 535565
rect 160208 535425 160358 535435
rect 174629 530605 174685 530607
rect 174709 530605 174765 530607
rect 174789 530605 174845 530607
rect 174869 530605 174925 530607
rect 174629 530553 174675 530605
rect 174675 530553 174685 530605
rect 174709 530553 174739 530605
rect 174739 530553 174751 530605
rect 174751 530553 174765 530605
rect 174789 530553 174803 530605
rect 174803 530553 174815 530605
rect 174815 530553 174845 530605
rect 174869 530553 174879 530605
rect 174879 530553 174925 530605
rect 174629 530551 174685 530553
rect 174709 530551 174765 530553
rect 174789 530551 174845 530553
rect 174869 530551 174925 530553
rect 178447 530605 178503 530607
rect 178527 530605 178583 530607
rect 178607 530605 178663 530607
rect 178687 530605 178743 530607
rect 178447 530553 178493 530605
rect 178493 530553 178503 530605
rect 178527 530553 178557 530605
rect 178557 530553 178569 530605
rect 178569 530553 178583 530605
rect 178607 530553 178621 530605
rect 178621 530553 178633 530605
rect 178633 530553 178663 530605
rect 178687 530553 178697 530605
rect 178697 530553 178743 530605
rect 178447 530551 178503 530553
rect 178527 530551 178583 530553
rect 178607 530551 178663 530553
rect 178687 530551 178743 530553
rect 173969 530061 174025 530063
rect 174049 530061 174105 530063
rect 174129 530061 174185 530063
rect 174209 530061 174265 530063
rect 173969 530009 174015 530061
rect 174015 530009 174025 530061
rect 174049 530009 174079 530061
rect 174079 530009 174091 530061
rect 174091 530009 174105 530061
rect 174129 530009 174143 530061
rect 174143 530009 174155 530061
rect 174155 530009 174185 530061
rect 174209 530009 174219 530061
rect 174219 530009 174265 530061
rect 173969 530007 174025 530009
rect 174049 530007 174105 530009
rect 174129 530007 174185 530009
rect 174209 530007 174265 530009
rect 174629 529517 174685 529519
rect 174709 529517 174765 529519
rect 174789 529517 174845 529519
rect 174869 529517 174925 529519
rect 174629 529465 174675 529517
rect 174675 529465 174685 529517
rect 174709 529465 174739 529517
rect 174739 529465 174751 529517
rect 174751 529465 174765 529517
rect 174789 529465 174803 529517
rect 174803 529465 174815 529517
rect 174815 529465 174845 529517
rect 174869 529465 174879 529517
rect 174879 529465 174925 529517
rect 174629 529463 174685 529465
rect 174709 529463 174765 529465
rect 174789 529463 174845 529465
rect 174869 529463 174925 529465
rect 173969 528973 174025 528975
rect 174049 528973 174105 528975
rect 174129 528973 174185 528975
rect 174209 528973 174265 528975
rect 173969 528921 174015 528973
rect 174015 528921 174025 528973
rect 174049 528921 174079 528973
rect 174079 528921 174091 528973
rect 174091 528921 174105 528973
rect 174129 528921 174143 528973
rect 174143 528921 174155 528973
rect 174155 528921 174185 528973
rect 174209 528921 174219 528973
rect 174219 528921 174265 528973
rect 173969 528919 174025 528921
rect 174049 528919 174105 528921
rect 174129 528919 174185 528921
rect 174209 528919 174265 528921
rect 174629 528429 174685 528431
rect 174709 528429 174765 528431
rect 174789 528429 174845 528431
rect 174869 528429 174925 528431
rect 174629 528377 174675 528429
rect 174675 528377 174685 528429
rect 174709 528377 174739 528429
rect 174739 528377 174751 528429
rect 174751 528377 174765 528429
rect 174789 528377 174803 528429
rect 174803 528377 174815 528429
rect 174815 528377 174845 528429
rect 174869 528377 174879 528429
rect 174879 528377 174925 528429
rect 174629 528375 174685 528377
rect 174709 528375 174765 528377
rect 174789 528375 174845 528377
rect 174869 528375 174925 528377
rect 173969 527885 174025 527887
rect 174049 527885 174105 527887
rect 174129 527885 174185 527887
rect 174209 527885 174265 527887
rect 173969 527833 174015 527885
rect 174015 527833 174025 527885
rect 174049 527833 174079 527885
rect 174079 527833 174091 527885
rect 174091 527833 174105 527885
rect 174129 527833 174143 527885
rect 174143 527833 174155 527885
rect 174155 527833 174185 527885
rect 174209 527833 174219 527885
rect 174219 527833 174265 527885
rect 173969 527831 174025 527833
rect 174049 527831 174105 527833
rect 174129 527831 174185 527833
rect 174209 527831 174265 527833
rect 177787 530061 177843 530063
rect 177867 530061 177923 530063
rect 177947 530061 178003 530063
rect 178027 530061 178083 530063
rect 177787 530009 177833 530061
rect 177833 530009 177843 530061
rect 177867 530009 177897 530061
rect 177897 530009 177909 530061
rect 177909 530009 177923 530061
rect 177947 530009 177961 530061
rect 177961 530009 177973 530061
rect 177973 530009 178003 530061
rect 178027 530009 178037 530061
rect 178037 530009 178083 530061
rect 177787 530007 177843 530009
rect 177867 530007 177923 530009
rect 177947 530007 178003 530009
rect 178027 530007 178083 530009
rect 177787 528973 177843 528975
rect 177867 528973 177923 528975
rect 177947 528973 178003 528975
rect 178027 528973 178083 528975
rect 177787 528921 177833 528973
rect 177833 528921 177843 528973
rect 177867 528921 177897 528973
rect 177897 528921 177909 528973
rect 177909 528921 177923 528973
rect 177947 528921 177961 528973
rect 177961 528921 177973 528973
rect 177973 528921 178003 528973
rect 178027 528921 178037 528973
rect 178037 528921 178083 528973
rect 177787 528919 177843 528921
rect 177867 528919 177923 528921
rect 177947 528919 178003 528921
rect 178027 528919 178083 528921
rect 178447 529517 178503 529519
rect 178527 529517 178583 529519
rect 178607 529517 178663 529519
rect 178687 529517 178743 529519
rect 178447 529465 178493 529517
rect 178493 529465 178503 529517
rect 178527 529465 178557 529517
rect 178557 529465 178569 529517
rect 178569 529465 178583 529517
rect 178607 529465 178621 529517
rect 178621 529465 178633 529517
rect 178633 529465 178663 529517
rect 178687 529465 178697 529517
rect 178697 529465 178743 529517
rect 178447 529463 178503 529465
rect 178527 529463 178583 529465
rect 178607 529463 178663 529465
rect 178687 529463 178743 529465
rect 177787 527885 177843 527887
rect 177867 527885 177923 527887
rect 177947 527885 178003 527887
rect 178027 527885 178083 527887
rect 177787 527833 177833 527885
rect 177833 527833 177843 527885
rect 177867 527833 177897 527885
rect 177897 527833 177909 527885
rect 177909 527833 177923 527885
rect 177947 527833 177961 527885
rect 177961 527833 177973 527885
rect 177973 527833 178003 527885
rect 178027 527833 178037 527885
rect 178037 527833 178083 527885
rect 177787 527831 177843 527833
rect 177867 527831 177923 527833
rect 177947 527831 178003 527833
rect 178027 527831 178083 527833
rect 174629 527341 174685 527343
rect 174709 527341 174765 527343
rect 174789 527341 174845 527343
rect 174869 527341 174925 527343
rect 174629 527289 174675 527341
rect 174675 527289 174685 527341
rect 174709 527289 174739 527341
rect 174739 527289 174751 527341
rect 174751 527289 174765 527341
rect 174789 527289 174803 527341
rect 174803 527289 174815 527341
rect 174815 527289 174845 527341
rect 174869 527289 174879 527341
rect 174879 527289 174925 527341
rect 174629 527287 174685 527289
rect 174709 527287 174765 527289
rect 174789 527287 174845 527289
rect 174869 527287 174925 527289
rect 173969 526797 174025 526799
rect 174049 526797 174105 526799
rect 174129 526797 174185 526799
rect 174209 526797 174265 526799
rect 173969 526745 174015 526797
rect 174015 526745 174025 526797
rect 174049 526745 174079 526797
rect 174079 526745 174091 526797
rect 174091 526745 174105 526797
rect 174129 526745 174143 526797
rect 174143 526745 174155 526797
rect 174155 526745 174185 526797
rect 174209 526745 174219 526797
rect 174219 526745 174265 526797
rect 173969 526743 174025 526745
rect 174049 526743 174105 526745
rect 174129 526743 174185 526745
rect 174209 526743 174265 526745
rect 177787 526797 177843 526799
rect 177867 526797 177923 526799
rect 177947 526797 178003 526799
rect 178027 526797 178083 526799
rect 177787 526745 177833 526797
rect 177833 526745 177843 526797
rect 177867 526745 177897 526797
rect 177897 526745 177909 526797
rect 177909 526745 177923 526797
rect 177947 526745 177961 526797
rect 177961 526745 177973 526797
rect 177973 526745 178003 526797
rect 178027 526745 178037 526797
rect 178037 526745 178083 526797
rect 177787 526743 177843 526745
rect 177867 526743 177923 526745
rect 177947 526743 178003 526745
rect 178027 526743 178083 526745
rect 174629 526253 174685 526255
rect 174709 526253 174765 526255
rect 174789 526253 174845 526255
rect 174869 526253 174925 526255
rect 174629 526201 174675 526253
rect 174675 526201 174685 526253
rect 174709 526201 174739 526253
rect 174739 526201 174751 526253
rect 174751 526201 174765 526253
rect 174789 526201 174803 526253
rect 174803 526201 174815 526253
rect 174815 526201 174845 526253
rect 174869 526201 174879 526253
rect 174879 526201 174925 526253
rect 174629 526199 174685 526201
rect 174709 526199 174765 526201
rect 174789 526199 174845 526201
rect 174869 526199 174925 526201
rect 173969 525709 174025 525711
rect 174049 525709 174105 525711
rect 174129 525709 174185 525711
rect 174209 525709 174265 525711
rect 173969 525657 174015 525709
rect 174015 525657 174025 525709
rect 174049 525657 174079 525709
rect 174079 525657 174091 525709
rect 174091 525657 174105 525709
rect 174129 525657 174143 525709
rect 174143 525657 174155 525709
rect 174155 525657 174185 525709
rect 174209 525657 174219 525709
rect 174219 525657 174265 525709
rect 173969 525655 174025 525657
rect 174049 525655 174105 525657
rect 174129 525655 174185 525657
rect 174209 525655 174265 525657
rect 177787 525709 177843 525711
rect 177867 525709 177923 525711
rect 177947 525709 178003 525711
rect 178027 525709 178083 525711
rect 177787 525657 177833 525709
rect 177833 525657 177843 525709
rect 177867 525657 177897 525709
rect 177897 525657 177909 525709
rect 177909 525657 177923 525709
rect 177947 525657 177961 525709
rect 177961 525657 177973 525709
rect 177973 525657 178003 525709
rect 178027 525657 178037 525709
rect 178037 525657 178083 525709
rect 177787 525655 177843 525657
rect 177867 525655 177923 525657
rect 177947 525655 178003 525657
rect 178027 525655 178083 525657
rect 174629 525165 174685 525167
rect 174709 525165 174765 525167
rect 174789 525165 174845 525167
rect 174869 525165 174925 525167
rect 174629 525113 174675 525165
rect 174675 525113 174685 525165
rect 174709 525113 174739 525165
rect 174739 525113 174751 525165
rect 174751 525113 174765 525165
rect 174789 525113 174803 525165
rect 174803 525113 174815 525165
rect 174815 525113 174845 525165
rect 174869 525113 174879 525165
rect 174879 525113 174925 525165
rect 174629 525111 174685 525113
rect 174709 525111 174765 525113
rect 174789 525111 174845 525113
rect 174869 525111 174925 525113
rect 173969 524621 174025 524623
rect 174049 524621 174105 524623
rect 174129 524621 174185 524623
rect 174209 524621 174265 524623
rect 173969 524569 174015 524621
rect 174015 524569 174025 524621
rect 174049 524569 174079 524621
rect 174079 524569 174091 524621
rect 174091 524569 174105 524621
rect 174129 524569 174143 524621
rect 174143 524569 174155 524621
rect 174155 524569 174185 524621
rect 174209 524569 174219 524621
rect 174219 524569 174265 524621
rect 173969 524567 174025 524569
rect 174049 524567 174105 524569
rect 174129 524567 174185 524569
rect 174209 524567 174265 524569
rect 177787 524621 177843 524623
rect 177867 524621 177923 524623
rect 177947 524621 178003 524623
rect 178027 524621 178083 524623
rect 177787 524569 177833 524621
rect 177833 524569 177843 524621
rect 177867 524569 177897 524621
rect 177897 524569 177909 524621
rect 177909 524569 177923 524621
rect 177947 524569 177961 524621
rect 177961 524569 177973 524621
rect 177973 524569 178003 524621
rect 178027 524569 178037 524621
rect 178037 524569 178083 524621
rect 177787 524567 177843 524569
rect 177867 524567 177923 524569
rect 177947 524567 178003 524569
rect 178027 524567 178083 524569
rect 174629 524077 174685 524079
rect 174709 524077 174765 524079
rect 174789 524077 174845 524079
rect 174869 524077 174925 524079
rect 174629 524025 174675 524077
rect 174675 524025 174685 524077
rect 174709 524025 174739 524077
rect 174739 524025 174751 524077
rect 174751 524025 174765 524077
rect 174789 524025 174803 524077
rect 174803 524025 174815 524077
rect 174815 524025 174845 524077
rect 174869 524025 174879 524077
rect 174879 524025 174925 524077
rect 174629 524023 174685 524025
rect 174709 524023 174765 524025
rect 174789 524023 174845 524025
rect 174869 524023 174925 524025
rect 173969 523533 174025 523535
rect 174049 523533 174105 523535
rect 174129 523533 174185 523535
rect 174209 523533 174265 523535
rect 173969 523481 174015 523533
rect 174015 523481 174025 523533
rect 174049 523481 174079 523533
rect 174079 523481 174091 523533
rect 174091 523481 174105 523533
rect 174129 523481 174143 523533
rect 174143 523481 174155 523533
rect 174155 523481 174185 523533
rect 174209 523481 174219 523533
rect 174219 523481 174265 523533
rect 173969 523479 174025 523481
rect 174049 523479 174105 523481
rect 174129 523479 174185 523481
rect 174209 523479 174265 523481
rect 177787 523533 177843 523535
rect 177867 523533 177923 523535
rect 177947 523533 178003 523535
rect 178027 523533 178083 523535
rect 177787 523481 177833 523533
rect 177833 523481 177843 523533
rect 177867 523481 177897 523533
rect 177897 523481 177909 523533
rect 177909 523481 177923 523533
rect 177947 523481 177961 523533
rect 177961 523481 177973 523533
rect 177973 523481 178003 523533
rect 178027 523481 178037 523533
rect 178037 523481 178083 523533
rect 177787 523479 177843 523481
rect 177867 523479 177923 523481
rect 177947 523479 178003 523481
rect 178027 523479 178083 523481
rect 174629 522989 174685 522991
rect 174709 522989 174765 522991
rect 174789 522989 174845 522991
rect 174869 522989 174925 522991
rect 174629 522937 174675 522989
rect 174675 522937 174685 522989
rect 174709 522937 174739 522989
rect 174739 522937 174751 522989
rect 174751 522937 174765 522989
rect 174789 522937 174803 522989
rect 174803 522937 174815 522989
rect 174815 522937 174845 522989
rect 174869 522937 174879 522989
rect 174879 522937 174925 522989
rect 174629 522935 174685 522937
rect 174709 522935 174765 522937
rect 174789 522935 174845 522937
rect 174869 522935 174925 522937
rect 173969 522445 174025 522447
rect 174049 522445 174105 522447
rect 174129 522445 174185 522447
rect 174209 522445 174265 522447
rect 173969 522393 174015 522445
rect 174015 522393 174025 522445
rect 174049 522393 174079 522445
rect 174079 522393 174091 522445
rect 174091 522393 174105 522445
rect 174129 522393 174143 522445
rect 174143 522393 174155 522445
rect 174155 522393 174185 522445
rect 174209 522393 174219 522445
rect 174219 522393 174265 522445
rect 173969 522391 174025 522393
rect 174049 522391 174105 522393
rect 174129 522391 174185 522393
rect 174209 522391 174265 522393
rect 177787 522445 177843 522447
rect 177867 522445 177923 522447
rect 177947 522445 178003 522447
rect 178027 522445 178083 522447
rect 177787 522393 177833 522445
rect 177833 522393 177843 522445
rect 177867 522393 177897 522445
rect 177897 522393 177909 522445
rect 177909 522393 177923 522445
rect 177947 522393 177961 522445
rect 177961 522393 177973 522445
rect 177973 522393 178003 522445
rect 178027 522393 178037 522445
rect 178037 522393 178083 522445
rect 177787 522391 177843 522393
rect 177867 522391 177923 522393
rect 177947 522391 178003 522393
rect 178027 522391 178083 522393
rect 174629 521901 174685 521903
rect 174709 521901 174765 521903
rect 174789 521901 174845 521903
rect 174869 521901 174925 521903
rect 174629 521849 174675 521901
rect 174675 521849 174685 521901
rect 174709 521849 174739 521901
rect 174739 521849 174751 521901
rect 174751 521849 174765 521901
rect 174789 521849 174803 521901
rect 174803 521849 174815 521901
rect 174815 521849 174845 521901
rect 174869 521849 174879 521901
rect 174879 521849 174925 521901
rect 174629 521847 174685 521849
rect 174709 521847 174765 521849
rect 174789 521847 174845 521849
rect 174869 521847 174925 521849
rect 173969 521357 174025 521359
rect 174049 521357 174105 521359
rect 174129 521357 174185 521359
rect 174209 521357 174265 521359
rect 173969 521305 174015 521357
rect 174015 521305 174025 521357
rect 174049 521305 174079 521357
rect 174079 521305 174091 521357
rect 174091 521305 174105 521357
rect 174129 521305 174143 521357
rect 174143 521305 174155 521357
rect 174155 521305 174185 521357
rect 174209 521305 174219 521357
rect 174219 521305 174265 521357
rect 173969 521303 174025 521305
rect 174049 521303 174105 521305
rect 174129 521303 174185 521305
rect 174209 521303 174265 521305
rect 177787 521357 177843 521359
rect 177867 521357 177923 521359
rect 177947 521357 178003 521359
rect 178027 521357 178083 521359
rect 177787 521305 177833 521357
rect 177833 521305 177843 521357
rect 177867 521305 177897 521357
rect 177897 521305 177909 521357
rect 177909 521305 177923 521357
rect 177947 521305 177961 521357
rect 177961 521305 177973 521357
rect 177973 521305 178003 521357
rect 178027 521305 178037 521357
rect 178037 521305 178083 521357
rect 177787 521303 177843 521305
rect 177867 521303 177923 521305
rect 177947 521303 178003 521305
rect 178027 521303 178083 521305
rect 174629 520813 174685 520815
rect 174709 520813 174765 520815
rect 174789 520813 174845 520815
rect 174869 520813 174925 520815
rect 174629 520761 174675 520813
rect 174675 520761 174685 520813
rect 174709 520761 174739 520813
rect 174739 520761 174751 520813
rect 174751 520761 174765 520813
rect 174789 520761 174803 520813
rect 174803 520761 174815 520813
rect 174815 520761 174845 520813
rect 174869 520761 174879 520813
rect 174879 520761 174925 520813
rect 174629 520759 174685 520761
rect 174709 520759 174765 520761
rect 174789 520759 174845 520761
rect 174869 520759 174925 520761
rect 173969 520269 174025 520271
rect 174049 520269 174105 520271
rect 174129 520269 174185 520271
rect 174209 520269 174265 520271
rect 173969 520217 174015 520269
rect 174015 520217 174025 520269
rect 174049 520217 174079 520269
rect 174079 520217 174091 520269
rect 174091 520217 174105 520269
rect 174129 520217 174143 520269
rect 174143 520217 174155 520269
rect 174155 520217 174185 520269
rect 174209 520217 174219 520269
rect 174219 520217 174265 520269
rect 173969 520215 174025 520217
rect 174049 520215 174105 520217
rect 174129 520215 174185 520217
rect 174209 520215 174265 520217
rect 177787 520269 177843 520271
rect 177867 520269 177923 520271
rect 177947 520269 178003 520271
rect 178027 520269 178083 520271
rect 177787 520217 177833 520269
rect 177833 520217 177843 520269
rect 177867 520217 177897 520269
rect 177897 520217 177909 520269
rect 177909 520217 177923 520269
rect 177947 520217 177961 520269
rect 177961 520217 177973 520269
rect 177973 520217 178003 520269
rect 178027 520217 178037 520269
rect 178037 520217 178083 520269
rect 177787 520215 177843 520217
rect 177867 520215 177923 520217
rect 177947 520215 178003 520217
rect 178027 520215 178083 520217
rect 174629 519725 174685 519727
rect 174709 519725 174765 519727
rect 174789 519725 174845 519727
rect 174869 519725 174925 519727
rect 174629 519673 174675 519725
rect 174675 519673 174685 519725
rect 174709 519673 174739 519725
rect 174739 519673 174751 519725
rect 174751 519673 174765 519725
rect 174789 519673 174803 519725
rect 174803 519673 174815 519725
rect 174815 519673 174845 519725
rect 174869 519673 174879 519725
rect 174879 519673 174925 519725
rect 174629 519671 174685 519673
rect 174709 519671 174765 519673
rect 174789 519671 174845 519673
rect 174869 519671 174925 519673
rect 173969 519181 174025 519183
rect 174049 519181 174105 519183
rect 174129 519181 174185 519183
rect 174209 519181 174265 519183
rect 173969 519129 174015 519181
rect 174015 519129 174025 519181
rect 174049 519129 174079 519181
rect 174079 519129 174091 519181
rect 174091 519129 174105 519181
rect 174129 519129 174143 519181
rect 174143 519129 174155 519181
rect 174155 519129 174185 519181
rect 174209 519129 174219 519181
rect 174219 519129 174265 519181
rect 173969 519127 174025 519129
rect 174049 519127 174105 519129
rect 174129 519127 174185 519129
rect 174209 519127 174265 519129
rect 177787 519181 177843 519183
rect 177867 519181 177923 519183
rect 177947 519181 178003 519183
rect 178027 519181 178083 519183
rect 177787 519129 177833 519181
rect 177833 519129 177843 519181
rect 177867 519129 177897 519181
rect 177897 519129 177909 519181
rect 177909 519129 177923 519181
rect 177947 519129 177961 519181
rect 177961 519129 177973 519181
rect 177973 519129 178003 519181
rect 178027 519129 178037 519181
rect 178037 519129 178083 519181
rect 177787 519127 177843 519129
rect 177867 519127 177923 519129
rect 177947 519127 178003 519129
rect 178027 519127 178083 519129
rect 174629 518637 174685 518639
rect 174709 518637 174765 518639
rect 174789 518637 174845 518639
rect 174869 518637 174925 518639
rect 174629 518585 174675 518637
rect 174675 518585 174685 518637
rect 174709 518585 174739 518637
rect 174739 518585 174751 518637
rect 174751 518585 174765 518637
rect 174789 518585 174803 518637
rect 174803 518585 174815 518637
rect 174815 518585 174845 518637
rect 174869 518585 174879 518637
rect 174879 518585 174925 518637
rect 174629 518583 174685 518585
rect 174709 518583 174765 518585
rect 174789 518583 174845 518585
rect 174869 518583 174925 518585
rect 173969 518093 174025 518095
rect 174049 518093 174105 518095
rect 174129 518093 174185 518095
rect 174209 518093 174265 518095
rect 173969 518041 174015 518093
rect 174015 518041 174025 518093
rect 174049 518041 174079 518093
rect 174079 518041 174091 518093
rect 174091 518041 174105 518093
rect 174129 518041 174143 518093
rect 174143 518041 174155 518093
rect 174155 518041 174185 518093
rect 174209 518041 174219 518093
rect 174219 518041 174265 518093
rect 173969 518039 174025 518041
rect 174049 518039 174105 518041
rect 174129 518039 174185 518041
rect 174209 518039 174265 518041
rect 177787 518093 177843 518095
rect 177867 518093 177923 518095
rect 177947 518093 178003 518095
rect 178027 518093 178083 518095
rect 177787 518041 177833 518093
rect 177833 518041 177843 518093
rect 177867 518041 177897 518093
rect 177897 518041 177909 518093
rect 177909 518041 177923 518093
rect 177947 518041 177961 518093
rect 177961 518041 177973 518093
rect 177973 518041 178003 518093
rect 178027 518041 178037 518093
rect 178037 518041 178083 518093
rect 177787 518039 177843 518041
rect 177867 518039 177923 518041
rect 177947 518039 178003 518041
rect 178027 518039 178083 518041
rect 174629 517549 174685 517551
rect 174709 517549 174765 517551
rect 174789 517549 174845 517551
rect 174869 517549 174925 517551
rect 174629 517497 174675 517549
rect 174675 517497 174685 517549
rect 174709 517497 174739 517549
rect 174739 517497 174751 517549
rect 174751 517497 174765 517549
rect 174789 517497 174803 517549
rect 174803 517497 174815 517549
rect 174815 517497 174845 517549
rect 174869 517497 174879 517549
rect 174879 517497 174925 517549
rect 174629 517495 174685 517497
rect 174709 517495 174765 517497
rect 174789 517495 174845 517497
rect 174869 517495 174925 517497
rect 178447 528429 178503 528431
rect 178527 528429 178583 528431
rect 178607 528429 178663 528431
rect 178687 528429 178743 528431
rect 178447 528377 178493 528429
rect 178493 528377 178503 528429
rect 178527 528377 178557 528429
rect 178557 528377 178569 528429
rect 178569 528377 178583 528429
rect 178607 528377 178621 528429
rect 178621 528377 178633 528429
rect 178633 528377 178663 528429
rect 178687 528377 178697 528429
rect 178697 528377 178743 528429
rect 178447 528375 178503 528377
rect 178527 528375 178583 528377
rect 178607 528375 178663 528377
rect 178687 528375 178743 528377
rect 182265 530605 182321 530607
rect 182345 530605 182401 530607
rect 182425 530605 182481 530607
rect 182505 530605 182561 530607
rect 182265 530553 182311 530605
rect 182311 530553 182321 530605
rect 182345 530553 182375 530605
rect 182375 530553 182387 530605
rect 182387 530553 182401 530605
rect 182425 530553 182439 530605
rect 182439 530553 182451 530605
rect 182451 530553 182481 530605
rect 182505 530553 182515 530605
rect 182515 530553 182561 530605
rect 182265 530551 182321 530553
rect 182345 530551 182401 530553
rect 182425 530551 182481 530553
rect 182505 530551 182561 530553
rect 186083 530605 186139 530607
rect 186163 530605 186219 530607
rect 186243 530605 186299 530607
rect 186323 530605 186379 530607
rect 186083 530553 186129 530605
rect 186129 530553 186139 530605
rect 186163 530553 186193 530605
rect 186193 530553 186205 530605
rect 186205 530553 186219 530605
rect 186243 530553 186257 530605
rect 186257 530553 186269 530605
rect 186269 530553 186299 530605
rect 186323 530553 186333 530605
rect 186333 530553 186379 530605
rect 186083 530551 186139 530553
rect 186163 530551 186219 530553
rect 186243 530551 186299 530553
rect 186323 530551 186379 530553
rect 181605 530061 181661 530063
rect 181685 530061 181741 530063
rect 181765 530061 181821 530063
rect 181845 530061 181901 530063
rect 181605 530009 181651 530061
rect 181651 530009 181661 530061
rect 181685 530009 181715 530061
rect 181715 530009 181727 530061
rect 181727 530009 181741 530061
rect 181765 530009 181779 530061
rect 181779 530009 181791 530061
rect 181791 530009 181821 530061
rect 181845 530009 181855 530061
rect 181855 530009 181901 530061
rect 181605 530007 181661 530009
rect 181685 530007 181741 530009
rect 181765 530007 181821 530009
rect 181845 530007 181901 530009
rect 181605 528973 181661 528975
rect 181685 528973 181741 528975
rect 181765 528973 181821 528975
rect 181845 528973 181901 528975
rect 181605 528921 181651 528973
rect 181651 528921 181661 528973
rect 181685 528921 181715 528973
rect 181715 528921 181727 528973
rect 181727 528921 181741 528973
rect 181765 528921 181779 528973
rect 181779 528921 181791 528973
rect 181791 528921 181821 528973
rect 181845 528921 181855 528973
rect 181855 528921 181901 528973
rect 181605 528919 181661 528921
rect 181685 528919 181741 528921
rect 181765 528919 181821 528921
rect 181845 528919 181901 528921
rect 182265 529517 182321 529519
rect 182345 529517 182401 529519
rect 182425 529517 182481 529519
rect 182505 529517 182561 529519
rect 182265 529465 182311 529517
rect 182311 529465 182321 529517
rect 182345 529465 182375 529517
rect 182375 529465 182387 529517
rect 182387 529465 182401 529517
rect 182425 529465 182439 529517
rect 182439 529465 182451 529517
rect 182451 529465 182481 529517
rect 182505 529465 182515 529517
rect 182515 529465 182561 529517
rect 182265 529463 182321 529465
rect 182345 529463 182401 529465
rect 182425 529463 182481 529465
rect 182505 529463 182561 529465
rect 185423 530061 185479 530063
rect 185503 530061 185559 530063
rect 185583 530061 185639 530063
rect 185663 530061 185719 530063
rect 185423 530009 185469 530061
rect 185469 530009 185479 530061
rect 185503 530009 185533 530061
rect 185533 530009 185545 530061
rect 185545 530009 185559 530061
rect 185583 530009 185597 530061
rect 185597 530009 185609 530061
rect 185609 530009 185639 530061
rect 185663 530009 185673 530061
rect 185673 530009 185719 530061
rect 185423 530007 185479 530009
rect 185503 530007 185559 530009
rect 185583 530007 185639 530009
rect 185663 530007 185719 530009
rect 186083 529517 186139 529519
rect 186163 529517 186219 529519
rect 186243 529517 186299 529519
rect 186323 529517 186379 529519
rect 186083 529465 186129 529517
rect 186129 529465 186139 529517
rect 186163 529465 186193 529517
rect 186193 529465 186205 529517
rect 186205 529465 186219 529517
rect 186243 529465 186257 529517
rect 186257 529465 186269 529517
rect 186269 529465 186299 529517
rect 186323 529465 186333 529517
rect 186333 529465 186379 529517
rect 186083 529463 186139 529465
rect 186163 529463 186219 529465
rect 186243 529463 186299 529465
rect 186323 529463 186379 529465
rect 185423 528973 185479 528975
rect 185503 528973 185559 528975
rect 185583 528973 185639 528975
rect 185663 528973 185719 528975
rect 185423 528921 185469 528973
rect 185469 528921 185479 528973
rect 185503 528921 185533 528973
rect 185533 528921 185545 528973
rect 185545 528921 185559 528973
rect 185583 528921 185597 528973
rect 185597 528921 185609 528973
rect 185609 528921 185639 528973
rect 185663 528921 185673 528973
rect 185673 528921 185719 528973
rect 185423 528919 185479 528921
rect 185503 528919 185559 528921
rect 185583 528919 185639 528921
rect 185663 528919 185719 528921
rect 182265 528429 182321 528431
rect 182345 528429 182401 528431
rect 182425 528429 182481 528431
rect 182505 528429 182561 528431
rect 182265 528377 182311 528429
rect 182311 528377 182321 528429
rect 182345 528377 182375 528429
rect 182375 528377 182387 528429
rect 182387 528377 182401 528429
rect 182425 528377 182439 528429
rect 182439 528377 182451 528429
rect 182451 528377 182481 528429
rect 182505 528377 182515 528429
rect 182515 528377 182561 528429
rect 182265 528375 182321 528377
rect 182345 528375 182401 528377
rect 182425 528375 182481 528377
rect 182505 528375 182561 528377
rect 186083 528429 186139 528431
rect 186163 528429 186219 528431
rect 186243 528429 186299 528431
rect 186323 528429 186379 528431
rect 186083 528377 186129 528429
rect 186129 528377 186139 528429
rect 186163 528377 186193 528429
rect 186193 528377 186205 528429
rect 186205 528377 186219 528429
rect 186243 528377 186257 528429
rect 186257 528377 186269 528429
rect 186269 528377 186299 528429
rect 186323 528377 186333 528429
rect 186333 528377 186379 528429
rect 186083 528375 186139 528377
rect 186163 528375 186219 528377
rect 186243 528375 186299 528377
rect 186323 528375 186379 528377
rect 178447 527341 178503 527343
rect 178527 527341 178583 527343
rect 178607 527341 178663 527343
rect 178687 527341 178743 527343
rect 178447 527289 178493 527341
rect 178493 527289 178503 527341
rect 178527 527289 178557 527341
rect 178557 527289 178569 527341
rect 178569 527289 178583 527341
rect 178607 527289 178621 527341
rect 178621 527289 178633 527341
rect 178633 527289 178663 527341
rect 178687 527289 178697 527341
rect 178697 527289 178743 527341
rect 178447 527287 178503 527289
rect 178527 527287 178583 527289
rect 178607 527287 178663 527289
rect 178687 527287 178743 527289
rect 178447 526253 178503 526255
rect 178527 526253 178583 526255
rect 178607 526253 178663 526255
rect 178687 526253 178743 526255
rect 178447 526201 178493 526253
rect 178493 526201 178503 526253
rect 178527 526201 178557 526253
rect 178557 526201 178569 526253
rect 178569 526201 178583 526253
rect 178607 526201 178621 526253
rect 178621 526201 178633 526253
rect 178633 526201 178663 526253
rect 178687 526201 178697 526253
rect 178697 526201 178743 526253
rect 178447 526199 178503 526201
rect 178527 526199 178583 526201
rect 178607 526199 178663 526201
rect 178687 526199 178743 526201
rect 178447 525165 178503 525167
rect 178527 525165 178583 525167
rect 178607 525165 178663 525167
rect 178687 525165 178743 525167
rect 178447 525113 178493 525165
rect 178493 525113 178503 525165
rect 178527 525113 178557 525165
rect 178557 525113 178569 525165
rect 178569 525113 178583 525165
rect 178607 525113 178621 525165
rect 178621 525113 178633 525165
rect 178633 525113 178663 525165
rect 178687 525113 178697 525165
rect 178697 525113 178743 525165
rect 178447 525111 178503 525113
rect 178527 525111 178583 525113
rect 178607 525111 178663 525113
rect 178687 525111 178743 525113
rect 178447 524077 178503 524079
rect 178527 524077 178583 524079
rect 178607 524077 178663 524079
rect 178687 524077 178743 524079
rect 178447 524025 178493 524077
rect 178493 524025 178503 524077
rect 178527 524025 178557 524077
rect 178557 524025 178569 524077
rect 178569 524025 178583 524077
rect 178607 524025 178621 524077
rect 178621 524025 178633 524077
rect 178633 524025 178663 524077
rect 178687 524025 178697 524077
rect 178697 524025 178743 524077
rect 178447 524023 178503 524025
rect 178527 524023 178583 524025
rect 178607 524023 178663 524025
rect 178687 524023 178743 524025
rect 178447 522989 178503 522991
rect 178527 522989 178583 522991
rect 178607 522989 178663 522991
rect 178687 522989 178743 522991
rect 178447 522937 178493 522989
rect 178493 522937 178503 522989
rect 178527 522937 178557 522989
rect 178557 522937 178569 522989
rect 178569 522937 178583 522989
rect 178607 522937 178621 522989
rect 178621 522937 178633 522989
rect 178633 522937 178663 522989
rect 178687 522937 178697 522989
rect 178697 522937 178743 522989
rect 178447 522935 178503 522937
rect 178527 522935 178583 522937
rect 178607 522935 178663 522937
rect 178687 522935 178743 522937
rect 178447 521901 178503 521903
rect 178527 521901 178583 521903
rect 178607 521901 178663 521903
rect 178687 521901 178743 521903
rect 178447 521849 178493 521901
rect 178493 521849 178503 521901
rect 178527 521849 178557 521901
rect 178557 521849 178569 521901
rect 178569 521849 178583 521901
rect 178607 521849 178621 521901
rect 178621 521849 178633 521901
rect 178633 521849 178663 521901
rect 178687 521849 178697 521901
rect 178697 521849 178743 521901
rect 178447 521847 178503 521849
rect 178527 521847 178583 521849
rect 178607 521847 178663 521849
rect 178687 521847 178743 521849
rect 178447 520813 178503 520815
rect 178527 520813 178583 520815
rect 178607 520813 178663 520815
rect 178687 520813 178743 520815
rect 178447 520761 178493 520813
rect 178493 520761 178503 520813
rect 178527 520761 178557 520813
rect 178557 520761 178569 520813
rect 178569 520761 178583 520813
rect 178607 520761 178621 520813
rect 178621 520761 178633 520813
rect 178633 520761 178663 520813
rect 178687 520761 178697 520813
rect 178697 520761 178743 520813
rect 178447 520759 178503 520761
rect 178527 520759 178583 520761
rect 178607 520759 178663 520761
rect 178687 520759 178743 520761
rect 178447 519725 178503 519727
rect 178527 519725 178583 519727
rect 178607 519725 178663 519727
rect 178687 519725 178743 519727
rect 178447 519673 178493 519725
rect 178493 519673 178503 519725
rect 178527 519673 178557 519725
rect 178557 519673 178569 519725
rect 178569 519673 178583 519725
rect 178607 519673 178621 519725
rect 178621 519673 178633 519725
rect 178633 519673 178663 519725
rect 178687 519673 178697 519725
rect 178697 519673 178743 519725
rect 178447 519671 178503 519673
rect 178527 519671 178583 519673
rect 178607 519671 178663 519673
rect 178687 519671 178743 519673
rect 178447 518637 178503 518639
rect 178527 518637 178583 518639
rect 178607 518637 178663 518639
rect 178687 518637 178743 518639
rect 178447 518585 178493 518637
rect 178493 518585 178503 518637
rect 178527 518585 178557 518637
rect 178557 518585 178569 518637
rect 178569 518585 178583 518637
rect 178607 518585 178621 518637
rect 178621 518585 178633 518637
rect 178633 518585 178663 518637
rect 178687 518585 178697 518637
rect 178697 518585 178743 518637
rect 178447 518583 178503 518585
rect 178527 518583 178583 518585
rect 178607 518583 178663 518585
rect 178687 518583 178743 518585
rect 178447 517549 178503 517551
rect 178527 517549 178583 517551
rect 178607 517549 178663 517551
rect 178687 517549 178743 517551
rect 178447 517497 178493 517549
rect 178493 517497 178503 517549
rect 178527 517497 178557 517549
rect 178557 517497 178569 517549
rect 178569 517497 178583 517549
rect 178607 517497 178621 517549
rect 178621 517497 178633 517549
rect 178633 517497 178663 517549
rect 178687 517497 178697 517549
rect 178697 517497 178743 517549
rect 178447 517495 178503 517497
rect 178527 517495 178583 517497
rect 178607 517495 178663 517497
rect 178687 517495 178743 517497
rect 173969 517005 174025 517007
rect 174049 517005 174105 517007
rect 174129 517005 174185 517007
rect 174209 517005 174265 517007
rect 173969 516953 174015 517005
rect 174015 516953 174025 517005
rect 174049 516953 174079 517005
rect 174079 516953 174091 517005
rect 174091 516953 174105 517005
rect 174129 516953 174143 517005
rect 174143 516953 174155 517005
rect 174155 516953 174185 517005
rect 174209 516953 174219 517005
rect 174219 516953 174265 517005
rect 173969 516951 174025 516953
rect 174049 516951 174105 516953
rect 174129 516951 174185 516953
rect 174209 516951 174265 516953
rect 174629 516461 174685 516463
rect 174709 516461 174765 516463
rect 174789 516461 174845 516463
rect 174869 516461 174925 516463
rect 174629 516409 174675 516461
rect 174675 516409 174685 516461
rect 174709 516409 174739 516461
rect 174739 516409 174751 516461
rect 174751 516409 174765 516461
rect 174789 516409 174803 516461
rect 174803 516409 174815 516461
rect 174815 516409 174845 516461
rect 174869 516409 174879 516461
rect 174879 516409 174925 516461
rect 174629 516407 174685 516409
rect 174709 516407 174765 516409
rect 174789 516407 174845 516409
rect 174869 516407 174925 516409
rect 173969 515917 174025 515919
rect 174049 515917 174105 515919
rect 174129 515917 174185 515919
rect 174209 515917 174265 515919
rect 173969 515865 174015 515917
rect 174015 515865 174025 515917
rect 174049 515865 174079 515917
rect 174079 515865 174091 515917
rect 174091 515865 174105 515917
rect 174129 515865 174143 515917
rect 174143 515865 174155 515917
rect 174155 515865 174185 515917
rect 174209 515865 174219 515917
rect 174219 515865 174265 515917
rect 173969 515863 174025 515865
rect 174049 515863 174105 515865
rect 174129 515863 174185 515865
rect 174209 515863 174265 515865
rect 174629 515373 174685 515375
rect 174709 515373 174765 515375
rect 174789 515373 174845 515375
rect 174869 515373 174925 515375
rect 174629 515321 174675 515373
rect 174675 515321 174685 515373
rect 174709 515321 174739 515373
rect 174739 515321 174751 515373
rect 174751 515321 174765 515373
rect 174789 515321 174803 515373
rect 174803 515321 174815 515373
rect 174815 515321 174845 515373
rect 174869 515321 174879 515373
rect 174879 515321 174925 515373
rect 174629 515319 174685 515321
rect 174709 515319 174765 515321
rect 174789 515319 174845 515321
rect 174869 515319 174925 515321
rect 177787 517005 177843 517007
rect 177867 517005 177923 517007
rect 177947 517005 178003 517007
rect 178027 517005 178083 517007
rect 177787 516953 177833 517005
rect 177833 516953 177843 517005
rect 177867 516953 177897 517005
rect 177897 516953 177909 517005
rect 177909 516953 177923 517005
rect 177947 516953 177961 517005
rect 177961 516953 177973 517005
rect 177973 516953 178003 517005
rect 178027 516953 178037 517005
rect 178037 516953 178083 517005
rect 177787 516951 177843 516953
rect 177867 516951 177923 516953
rect 177947 516951 178003 516953
rect 178027 516951 178083 516953
rect 178447 516461 178503 516463
rect 178527 516461 178583 516463
rect 178607 516461 178663 516463
rect 178687 516461 178743 516463
rect 178447 516409 178493 516461
rect 178493 516409 178503 516461
rect 178527 516409 178557 516461
rect 178557 516409 178569 516461
rect 178569 516409 178583 516461
rect 178607 516409 178621 516461
rect 178621 516409 178633 516461
rect 178633 516409 178663 516461
rect 178687 516409 178697 516461
rect 178697 516409 178743 516461
rect 178447 516407 178503 516409
rect 178527 516407 178583 516409
rect 178607 516407 178663 516409
rect 178687 516407 178743 516409
rect 177787 515917 177843 515919
rect 177867 515917 177923 515919
rect 177947 515917 178003 515919
rect 178027 515917 178083 515919
rect 177787 515865 177833 515917
rect 177833 515865 177843 515917
rect 177867 515865 177897 515917
rect 177897 515865 177909 515917
rect 177909 515865 177923 515917
rect 177947 515865 177961 515917
rect 177961 515865 177973 515917
rect 177973 515865 178003 515917
rect 178027 515865 178037 515917
rect 178037 515865 178083 515917
rect 177787 515863 177843 515865
rect 177867 515863 177923 515865
rect 177947 515863 178003 515865
rect 178027 515863 178083 515865
rect 181605 527885 181661 527887
rect 181685 527885 181741 527887
rect 181765 527885 181821 527887
rect 181845 527885 181901 527887
rect 181605 527833 181651 527885
rect 181651 527833 181661 527885
rect 181685 527833 181715 527885
rect 181715 527833 181727 527885
rect 181727 527833 181741 527885
rect 181765 527833 181779 527885
rect 181779 527833 181791 527885
rect 181791 527833 181821 527885
rect 181845 527833 181855 527885
rect 181855 527833 181901 527885
rect 181605 527831 181661 527833
rect 181685 527831 181741 527833
rect 181765 527831 181821 527833
rect 181845 527831 181901 527833
rect 185423 527885 185479 527887
rect 185503 527885 185559 527887
rect 185583 527885 185639 527887
rect 185663 527885 185719 527887
rect 185423 527833 185469 527885
rect 185469 527833 185479 527885
rect 185503 527833 185533 527885
rect 185533 527833 185545 527885
rect 185545 527833 185559 527885
rect 185583 527833 185597 527885
rect 185597 527833 185609 527885
rect 185609 527833 185639 527885
rect 185663 527833 185673 527885
rect 185673 527833 185719 527885
rect 185423 527831 185479 527833
rect 185503 527831 185559 527833
rect 185583 527831 185639 527833
rect 185663 527831 185719 527833
rect 182265 527341 182321 527343
rect 182345 527341 182401 527343
rect 182425 527341 182481 527343
rect 182505 527341 182561 527343
rect 182265 527289 182311 527341
rect 182311 527289 182321 527341
rect 182345 527289 182375 527341
rect 182375 527289 182387 527341
rect 182387 527289 182401 527341
rect 182425 527289 182439 527341
rect 182439 527289 182451 527341
rect 182451 527289 182481 527341
rect 182505 527289 182515 527341
rect 182515 527289 182561 527341
rect 182265 527287 182321 527289
rect 182345 527287 182401 527289
rect 182425 527287 182481 527289
rect 182505 527287 182561 527289
rect 186083 527341 186139 527343
rect 186163 527341 186219 527343
rect 186243 527341 186299 527343
rect 186323 527341 186379 527343
rect 186083 527289 186129 527341
rect 186129 527289 186139 527341
rect 186163 527289 186193 527341
rect 186193 527289 186205 527341
rect 186205 527289 186219 527341
rect 186243 527289 186257 527341
rect 186257 527289 186269 527341
rect 186269 527289 186299 527341
rect 186323 527289 186333 527341
rect 186333 527289 186379 527341
rect 186083 527287 186139 527289
rect 186163 527287 186219 527289
rect 186243 527287 186299 527289
rect 186323 527287 186379 527289
rect 181605 526797 181661 526799
rect 181685 526797 181741 526799
rect 181765 526797 181821 526799
rect 181845 526797 181901 526799
rect 181605 526745 181651 526797
rect 181651 526745 181661 526797
rect 181685 526745 181715 526797
rect 181715 526745 181727 526797
rect 181727 526745 181741 526797
rect 181765 526745 181779 526797
rect 181779 526745 181791 526797
rect 181791 526745 181821 526797
rect 181845 526745 181855 526797
rect 181855 526745 181901 526797
rect 181605 526743 181661 526745
rect 181685 526743 181741 526745
rect 181765 526743 181821 526745
rect 181845 526743 181901 526745
rect 185423 526797 185479 526799
rect 185503 526797 185559 526799
rect 185583 526797 185639 526799
rect 185663 526797 185719 526799
rect 185423 526745 185469 526797
rect 185469 526745 185479 526797
rect 185503 526745 185533 526797
rect 185533 526745 185545 526797
rect 185545 526745 185559 526797
rect 185583 526745 185597 526797
rect 185597 526745 185609 526797
rect 185609 526745 185639 526797
rect 185663 526745 185673 526797
rect 185673 526745 185719 526797
rect 185423 526743 185479 526745
rect 185503 526743 185559 526745
rect 185583 526743 185639 526745
rect 185663 526743 185719 526745
rect 182265 526253 182321 526255
rect 182345 526253 182401 526255
rect 182425 526253 182481 526255
rect 182505 526253 182561 526255
rect 182265 526201 182311 526253
rect 182311 526201 182321 526253
rect 182345 526201 182375 526253
rect 182375 526201 182387 526253
rect 182387 526201 182401 526253
rect 182425 526201 182439 526253
rect 182439 526201 182451 526253
rect 182451 526201 182481 526253
rect 182505 526201 182515 526253
rect 182515 526201 182561 526253
rect 182265 526199 182321 526201
rect 182345 526199 182401 526201
rect 182425 526199 182481 526201
rect 182505 526199 182561 526201
rect 186083 526253 186139 526255
rect 186163 526253 186219 526255
rect 186243 526253 186299 526255
rect 186323 526253 186379 526255
rect 186083 526201 186129 526253
rect 186129 526201 186139 526253
rect 186163 526201 186193 526253
rect 186193 526201 186205 526253
rect 186205 526201 186219 526253
rect 186243 526201 186257 526253
rect 186257 526201 186269 526253
rect 186269 526201 186299 526253
rect 186323 526201 186333 526253
rect 186333 526201 186379 526253
rect 186083 526199 186139 526201
rect 186163 526199 186219 526201
rect 186243 526199 186299 526201
rect 186323 526199 186379 526201
rect 181605 525709 181661 525711
rect 181685 525709 181741 525711
rect 181765 525709 181821 525711
rect 181845 525709 181901 525711
rect 181605 525657 181651 525709
rect 181651 525657 181661 525709
rect 181685 525657 181715 525709
rect 181715 525657 181727 525709
rect 181727 525657 181741 525709
rect 181765 525657 181779 525709
rect 181779 525657 181791 525709
rect 181791 525657 181821 525709
rect 181845 525657 181855 525709
rect 181855 525657 181901 525709
rect 181605 525655 181661 525657
rect 181685 525655 181741 525657
rect 181765 525655 181821 525657
rect 181845 525655 181901 525657
rect 185423 525709 185479 525711
rect 185503 525709 185559 525711
rect 185583 525709 185639 525711
rect 185663 525709 185719 525711
rect 185423 525657 185469 525709
rect 185469 525657 185479 525709
rect 185503 525657 185533 525709
rect 185533 525657 185545 525709
rect 185545 525657 185559 525709
rect 185583 525657 185597 525709
rect 185597 525657 185609 525709
rect 185609 525657 185639 525709
rect 185663 525657 185673 525709
rect 185673 525657 185719 525709
rect 185423 525655 185479 525657
rect 185503 525655 185559 525657
rect 185583 525655 185639 525657
rect 185663 525655 185719 525657
rect 182265 525165 182321 525167
rect 182345 525165 182401 525167
rect 182425 525165 182481 525167
rect 182505 525165 182561 525167
rect 182265 525113 182311 525165
rect 182311 525113 182321 525165
rect 182345 525113 182375 525165
rect 182375 525113 182387 525165
rect 182387 525113 182401 525165
rect 182425 525113 182439 525165
rect 182439 525113 182451 525165
rect 182451 525113 182481 525165
rect 182505 525113 182515 525165
rect 182515 525113 182561 525165
rect 182265 525111 182321 525113
rect 182345 525111 182401 525113
rect 182425 525111 182481 525113
rect 182505 525111 182561 525113
rect 186083 525165 186139 525167
rect 186163 525165 186219 525167
rect 186243 525165 186299 525167
rect 186323 525165 186379 525167
rect 186083 525113 186129 525165
rect 186129 525113 186139 525165
rect 186163 525113 186193 525165
rect 186193 525113 186205 525165
rect 186205 525113 186219 525165
rect 186243 525113 186257 525165
rect 186257 525113 186269 525165
rect 186269 525113 186299 525165
rect 186323 525113 186333 525165
rect 186333 525113 186379 525165
rect 186083 525111 186139 525113
rect 186163 525111 186219 525113
rect 186243 525111 186299 525113
rect 186323 525111 186379 525113
rect 181605 524621 181661 524623
rect 181685 524621 181741 524623
rect 181765 524621 181821 524623
rect 181845 524621 181901 524623
rect 181605 524569 181651 524621
rect 181651 524569 181661 524621
rect 181685 524569 181715 524621
rect 181715 524569 181727 524621
rect 181727 524569 181741 524621
rect 181765 524569 181779 524621
rect 181779 524569 181791 524621
rect 181791 524569 181821 524621
rect 181845 524569 181855 524621
rect 181855 524569 181901 524621
rect 181605 524567 181661 524569
rect 181685 524567 181741 524569
rect 181765 524567 181821 524569
rect 181845 524567 181901 524569
rect 185423 524621 185479 524623
rect 185503 524621 185559 524623
rect 185583 524621 185639 524623
rect 185663 524621 185719 524623
rect 185423 524569 185469 524621
rect 185469 524569 185479 524621
rect 185503 524569 185533 524621
rect 185533 524569 185545 524621
rect 185545 524569 185559 524621
rect 185583 524569 185597 524621
rect 185597 524569 185609 524621
rect 185609 524569 185639 524621
rect 185663 524569 185673 524621
rect 185673 524569 185719 524621
rect 185423 524567 185479 524569
rect 185503 524567 185559 524569
rect 185583 524567 185639 524569
rect 185663 524567 185719 524569
rect 182265 524077 182321 524079
rect 182345 524077 182401 524079
rect 182425 524077 182481 524079
rect 182505 524077 182561 524079
rect 182265 524025 182311 524077
rect 182311 524025 182321 524077
rect 182345 524025 182375 524077
rect 182375 524025 182387 524077
rect 182387 524025 182401 524077
rect 182425 524025 182439 524077
rect 182439 524025 182451 524077
rect 182451 524025 182481 524077
rect 182505 524025 182515 524077
rect 182515 524025 182561 524077
rect 182265 524023 182321 524025
rect 182345 524023 182401 524025
rect 182425 524023 182481 524025
rect 182505 524023 182561 524025
rect 186083 524077 186139 524079
rect 186163 524077 186219 524079
rect 186243 524077 186299 524079
rect 186323 524077 186379 524079
rect 186083 524025 186129 524077
rect 186129 524025 186139 524077
rect 186163 524025 186193 524077
rect 186193 524025 186205 524077
rect 186205 524025 186219 524077
rect 186243 524025 186257 524077
rect 186257 524025 186269 524077
rect 186269 524025 186299 524077
rect 186323 524025 186333 524077
rect 186333 524025 186379 524077
rect 186083 524023 186139 524025
rect 186163 524023 186219 524025
rect 186243 524023 186299 524025
rect 186323 524023 186379 524025
rect 181605 523533 181661 523535
rect 181685 523533 181741 523535
rect 181765 523533 181821 523535
rect 181845 523533 181901 523535
rect 181605 523481 181651 523533
rect 181651 523481 181661 523533
rect 181685 523481 181715 523533
rect 181715 523481 181727 523533
rect 181727 523481 181741 523533
rect 181765 523481 181779 523533
rect 181779 523481 181791 523533
rect 181791 523481 181821 523533
rect 181845 523481 181855 523533
rect 181855 523481 181901 523533
rect 181605 523479 181661 523481
rect 181685 523479 181741 523481
rect 181765 523479 181821 523481
rect 181845 523479 181901 523481
rect 185423 523533 185479 523535
rect 185503 523533 185559 523535
rect 185583 523533 185639 523535
rect 185663 523533 185719 523535
rect 185423 523481 185469 523533
rect 185469 523481 185479 523533
rect 185503 523481 185533 523533
rect 185533 523481 185545 523533
rect 185545 523481 185559 523533
rect 185583 523481 185597 523533
rect 185597 523481 185609 523533
rect 185609 523481 185639 523533
rect 185663 523481 185673 523533
rect 185673 523481 185719 523533
rect 185423 523479 185479 523481
rect 185503 523479 185559 523481
rect 185583 523479 185639 523481
rect 185663 523479 185719 523481
rect 182265 522989 182321 522991
rect 182345 522989 182401 522991
rect 182425 522989 182481 522991
rect 182505 522989 182561 522991
rect 182265 522937 182311 522989
rect 182311 522937 182321 522989
rect 182345 522937 182375 522989
rect 182375 522937 182387 522989
rect 182387 522937 182401 522989
rect 182425 522937 182439 522989
rect 182439 522937 182451 522989
rect 182451 522937 182481 522989
rect 182505 522937 182515 522989
rect 182515 522937 182561 522989
rect 182265 522935 182321 522937
rect 182345 522935 182401 522937
rect 182425 522935 182481 522937
rect 182505 522935 182561 522937
rect 186083 522989 186139 522991
rect 186163 522989 186219 522991
rect 186243 522989 186299 522991
rect 186323 522989 186379 522991
rect 186083 522937 186129 522989
rect 186129 522937 186139 522989
rect 186163 522937 186193 522989
rect 186193 522937 186205 522989
rect 186205 522937 186219 522989
rect 186243 522937 186257 522989
rect 186257 522937 186269 522989
rect 186269 522937 186299 522989
rect 186323 522937 186333 522989
rect 186333 522937 186379 522989
rect 186083 522935 186139 522937
rect 186163 522935 186219 522937
rect 186243 522935 186299 522937
rect 186323 522935 186379 522937
rect 181605 522445 181661 522447
rect 181685 522445 181741 522447
rect 181765 522445 181821 522447
rect 181845 522445 181901 522447
rect 181605 522393 181651 522445
rect 181651 522393 181661 522445
rect 181685 522393 181715 522445
rect 181715 522393 181727 522445
rect 181727 522393 181741 522445
rect 181765 522393 181779 522445
rect 181779 522393 181791 522445
rect 181791 522393 181821 522445
rect 181845 522393 181855 522445
rect 181855 522393 181901 522445
rect 181605 522391 181661 522393
rect 181685 522391 181741 522393
rect 181765 522391 181821 522393
rect 181845 522391 181901 522393
rect 185423 522445 185479 522447
rect 185503 522445 185559 522447
rect 185583 522445 185639 522447
rect 185663 522445 185719 522447
rect 185423 522393 185469 522445
rect 185469 522393 185479 522445
rect 185503 522393 185533 522445
rect 185533 522393 185545 522445
rect 185545 522393 185559 522445
rect 185583 522393 185597 522445
rect 185597 522393 185609 522445
rect 185609 522393 185639 522445
rect 185663 522393 185673 522445
rect 185673 522393 185719 522445
rect 185423 522391 185479 522393
rect 185503 522391 185559 522393
rect 185583 522391 185639 522393
rect 185663 522391 185719 522393
rect 182265 521901 182321 521903
rect 182345 521901 182401 521903
rect 182425 521901 182481 521903
rect 182505 521901 182561 521903
rect 182265 521849 182311 521901
rect 182311 521849 182321 521901
rect 182345 521849 182375 521901
rect 182375 521849 182387 521901
rect 182387 521849 182401 521901
rect 182425 521849 182439 521901
rect 182439 521849 182451 521901
rect 182451 521849 182481 521901
rect 182505 521849 182515 521901
rect 182515 521849 182561 521901
rect 182265 521847 182321 521849
rect 182345 521847 182401 521849
rect 182425 521847 182481 521849
rect 182505 521847 182561 521849
rect 186083 521901 186139 521903
rect 186163 521901 186219 521903
rect 186243 521901 186299 521903
rect 186323 521901 186379 521903
rect 186083 521849 186129 521901
rect 186129 521849 186139 521901
rect 186163 521849 186193 521901
rect 186193 521849 186205 521901
rect 186205 521849 186219 521901
rect 186243 521849 186257 521901
rect 186257 521849 186269 521901
rect 186269 521849 186299 521901
rect 186323 521849 186333 521901
rect 186333 521849 186379 521901
rect 186083 521847 186139 521849
rect 186163 521847 186219 521849
rect 186243 521847 186299 521849
rect 186323 521847 186379 521849
rect 181605 521357 181661 521359
rect 181685 521357 181741 521359
rect 181765 521357 181821 521359
rect 181845 521357 181901 521359
rect 181605 521305 181651 521357
rect 181651 521305 181661 521357
rect 181685 521305 181715 521357
rect 181715 521305 181727 521357
rect 181727 521305 181741 521357
rect 181765 521305 181779 521357
rect 181779 521305 181791 521357
rect 181791 521305 181821 521357
rect 181845 521305 181855 521357
rect 181855 521305 181901 521357
rect 181605 521303 181661 521305
rect 181685 521303 181741 521305
rect 181765 521303 181821 521305
rect 181845 521303 181901 521305
rect 185423 521357 185479 521359
rect 185503 521357 185559 521359
rect 185583 521357 185639 521359
rect 185663 521357 185719 521359
rect 185423 521305 185469 521357
rect 185469 521305 185479 521357
rect 185503 521305 185533 521357
rect 185533 521305 185545 521357
rect 185545 521305 185559 521357
rect 185583 521305 185597 521357
rect 185597 521305 185609 521357
rect 185609 521305 185639 521357
rect 185663 521305 185673 521357
rect 185673 521305 185719 521357
rect 185423 521303 185479 521305
rect 185503 521303 185559 521305
rect 185583 521303 185639 521305
rect 185663 521303 185719 521305
rect 182265 520813 182321 520815
rect 182345 520813 182401 520815
rect 182425 520813 182481 520815
rect 182505 520813 182561 520815
rect 182265 520761 182311 520813
rect 182311 520761 182321 520813
rect 182345 520761 182375 520813
rect 182375 520761 182387 520813
rect 182387 520761 182401 520813
rect 182425 520761 182439 520813
rect 182439 520761 182451 520813
rect 182451 520761 182481 520813
rect 182505 520761 182515 520813
rect 182515 520761 182561 520813
rect 182265 520759 182321 520761
rect 182345 520759 182401 520761
rect 182425 520759 182481 520761
rect 182505 520759 182561 520761
rect 186083 520813 186139 520815
rect 186163 520813 186219 520815
rect 186243 520813 186299 520815
rect 186323 520813 186379 520815
rect 186083 520761 186129 520813
rect 186129 520761 186139 520813
rect 186163 520761 186193 520813
rect 186193 520761 186205 520813
rect 186205 520761 186219 520813
rect 186243 520761 186257 520813
rect 186257 520761 186269 520813
rect 186269 520761 186299 520813
rect 186323 520761 186333 520813
rect 186333 520761 186379 520813
rect 186083 520759 186139 520761
rect 186163 520759 186219 520761
rect 186243 520759 186299 520761
rect 186323 520759 186379 520761
rect 181605 520269 181661 520271
rect 181685 520269 181741 520271
rect 181765 520269 181821 520271
rect 181845 520269 181901 520271
rect 181605 520217 181651 520269
rect 181651 520217 181661 520269
rect 181685 520217 181715 520269
rect 181715 520217 181727 520269
rect 181727 520217 181741 520269
rect 181765 520217 181779 520269
rect 181779 520217 181791 520269
rect 181791 520217 181821 520269
rect 181845 520217 181855 520269
rect 181855 520217 181901 520269
rect 181605 520215 181661 520217
rect 181685 520215 181741 520217
rect 181765 520215 181821 520217
rect 181845 520215 181901 520217
rect 185423 520269 185479 520271
rect 185503 520269 185559 520271
rect 185583 520269 185639 520271
rect 185663 520269 185719 520271
rect 185423 520217 185469 520269
rect 185469 520217 185479 520269
rect 185503 520217 185533 520269
rect 185533 520217 185545 520269
rect 185545 520217 185559 520269
rect 185583 520217 185597 520269
rect 185597 520217 185609 520269
rect 185609 520217 185639 520269
rect 185663 520217 185673 520269
rect 185673 520217 185719 520269
rect 185423 520215 185479 520217
rect 185503 520215 185559 520217
rect 185583 520215 185639 520217
rect 185663 520215 185719 520217
rect 182265 519725 182321 519727
rect 182345 519725 182401 519727
rect 182425 519725 182481 519727
rect 182505 519725 182561 519727
rect 182265 519673 182311 519725
rect 182311 519673 182321 519725
rect 182345 519673 182375 519725
rect 182375 519673 182387 519725
rect 182387 519673 182401 519725
rect 182425 519673 182439 519725
rect 182439 519673 182451 519725
rect 182451 519673 182481 519725
rect 182505 519673 182515 519725
rect 182515 519673 182561 519725
rect 182265 519671 182321 519673
rect 182345 519671 182401 519673
rect 182425 519671 182481 519673
rect 182505 519671 182561 519673
rect 186083 519725 186139 519727
rect 186163 519725 186219 519727
rect 186243 519725 186299 519727
rect 186323 519725 186379 519727
rect 186083 519673 186129 519725
rect 186129 519673 186139 519725
rect 186163 519673 186193 519725
rect 186193 519673 186205 519725
rect 186205 519673 186219 519725
rect 186243 519673 186257 519725
rect 186257 519673 186269 519725
rect 186269 519673 186299 519725
rect 186323 519673 186333 519725
rect 186333 519673 186379 519725
rect 186083 519671 186139 519673
rect 186163 519671 186219 519673
rect 186243 519671 186299 519673
rect 186323 519671 186379 519673
rect 181605 519181 181661 519183
rect 181685 519181 181741 519183
rect 181765 519181 181821 519183
rect 181845 519181 181901 519183
rect 181605 519129 181651 519181
rect 181651 519129 181661 519181
rect 181685 519129 181715 519181
rect 181715 519129 181727 519181
rect 181727 519129 181741 519181
rect 181765 519129 181779 519181
rect 181779 519129 181791 519181
rect 181791 519129 181821 519181
rect 181845 519129 181855 519181
rect 181855 519129 181901 519181
rect 181605 519127 181661 519129
rect 181685 519127 181741 519129
rect 181765 519127 181821 519129
rect 181845 519127 181901 519129
rect 185423 519181 185479 519183
rect 185503 519181 185559 519183
rect 185583 519181 185639 519183
rect 185663 519181 185719 519183
rect 185423 519129 185469 519181
rect 185469 519129 185479 519181
rect 185503 519129 185533 519181
rect 185533 519129 185545 519181
rect 185545 519129 185559 519181
rect 185583 519129 185597 519181
rect 185597 519129 185609 519181
rect 185609 519129 185639 519181
rect 185663 519129 185673 519181
rect 185673 519129 185719 519181
rect 185423 519127 185479 519129
rect 185503 519127 185559 519129
rect 185583 519127 185639 519129
rect 185663 519127 185719 519129
rect 182265 518637 182321 518639
rect 182345 518637 182401 518639
rect 182425 518637 182481 518639
rect 182505 518637 182561 518639
rect 182265 518585 182311 518637
rect 182311 518585 182321 518637
rect 182345 518585 182375 518637
rect 182375 518585 182387 518637
rect 182387 518585 182401 518637
rect 182425 518585 182439 518637
rect 182439 518585 182451 518637
rect 182451 518585 182481 518637
rect 182505 518585 182515 518637
rect 182515 518585 182561 518637
rect 182265 518583 182321 518585
rect 182345 518583 182401 518585
rect 182425 518583 182481 518585
rect 182505 518583 182561 518585
rect 186083 518637 186139 518639
rect 186163 518637 186219 518639
rect 186243 518637 186299 518639
rect 186323 518637 186379 518639
rect 186083 518585 186129 518637
rect 186129 518585 186139 518637
rect 186163 518585 186193 518637
rect 186193 518585 186205 518637
rect 186205 518585 186219 518637
rect 186243 518585 186257 518637
rect 186257 518585 186269 518637
rect 186269 518585 186299 518637
rect 186323 518585 186333 518637
rect 186333 518585 186379 518637
rect 186083 518583 186139 518585
rect 186163 518583 186219 518585
rect 186243 518583 186299 518585
rect 186323 518583 186379 518585
rect 181605 518093 181661 518095
rect 181685 518093 181741 518095
rect 181765 518093 181821 518095
rect 181845 518093 181901 518095
rect 181605 518041 181651 518093
rect 181651 518041 181661 518093
rect 181685 518041 181715 518093
rect 181715 518041 181727 518093
rect 181727 518041 181741 518093
rect 181765 518041 181779 518093
rect 181779 518041 181791 518093
rect 181791 518041 181821 518093
rect 181845 518041 181855 518093
rect 181855 518041 181901 518093
rect 181605 518039 181661 518041
rect 181685 518039 181741 518041
rect 181765 518039 181821 518041
rect 181845 518039 181901 518041
rect 185423 518093 185479 518095
rect 185503 518093 185559 518095
rect 185583 518093 185639 518095
rect 185663 518093 185719 518095
rect 185423 518041 185469 518093
rect 185469 518041 185479 518093
rect 185503 518041 185533 518093
rect 185533 518041 185545 518093
rect 185545 518041 185559 518093
rect 185583 518041 185597 518093
rect 185597 518041 185609 518093
rect 185609 518041 185639 518093
rect 185663 518041 185673 518093
rect 185673 518041 185719 518093
rect 185423 518039 185479 518041
rect 185503 518039 185559 518041
rect 185583 518039 185639 518041
rect 185663 518039 185719 518041
rect 182265 517549 182321 517551
rect 182345 517549 182401 517551
rect 182425 517549 182481 517551
rect 182505 517549 182561 517551
rect 182265 517497 182311 517549
rect 182311 517497 182321 517549
rect 182345 517497 182375 517549
rect 182375 517497 182387 517549
rect 182387 517497 182401 517549
rect 182425 517497 182439 517549
rect 182439 517497 182451 517549
rect 182451 517497 182481 517549
rect 182505 517497 182515 517549
rect 182515 517497 182561 517549
rect 182265 517495 182321 517497
rect 182345 517495 182401 517497
rect 182425 517495 182481 517497
rect 182505 517495 182561 517497
rect 186083 517549 186139 517551
rect 186163 517549 186219 517551
rect 186243 517549 186299 517551
rect 186323 517549 186379 517551
rect 186083 517497 186129 517549
rect 186129 517497 186139 517549
rect 186163 517497 186193 517549
rect 186193 517497 186205 517549
rect 186205 517497 186219 517549
rect 186243 517497 186257 517549
rect 186257 517497 186269 517549
rect 186269 517497 186299 517549
rect 186323 517497 186333 517549
rect 186333 517497 186379 517549
rect 186083 517495 186139 517497
rect 186163 517495 186219 517497
rect 186243 517495 186299 517497
rect 186323 517495 186379 517497
rect 181605 517005 181661 517007
rect 181685 517005 181741 517007
rect 181765 517005 181821 517007
rect 181845 517005 181901 517007
rect 181605 516953 181651 517005
rect 181651 516953 181661 517005
rect 181685 516953 181715 517005
rect 181715 516953 181727 517005
rect 181727 516953 181741 517005
rect 181765 516953 181779 517005
rect 181779 516953 181791 517005
rect 181791 516953 181821 517005
rect 181845 516953 181855 517005
rect 181855 516953 181901 517005
rect 181605 516951 181661 516953
rect 181685 516951 181741 516953
rect 181765 516951 181821 516953
rect 181845 516951 181901 516953
rect 185423 517005 185479 517007
rect 185503 517005 185559 517007
rect 185583 517005 185639 517007
rect 185663 517005 185719 517007
rect 185423 516953 185469 517005
rect 185469 516953 185479 517005
rect 185503 516953 185533 517005
rect 185533 516953 185545 517005
rect 185545 516953 185559 517005
rect 185583 516953 185597 517005
rect 185597 516953 185609 517005
rect 185609 516953 185639 517005
rect 185663 516953 185673 517005
rect 185673 516953 185719 517005
rect 185423 516951 185479 516953
rect 185503 516951 185559 516953
rect 185583 516951 185639 516953
rect 185663 516951 185719 516953
rect 182265 516461 182321 516463
rect 182345 516461 182401 516463
rect 182425 516461 182481 516463
rect 182505 516461 182561 516463
rect 182265 516409 182311 516461
rect 182311 516409 182321 516461
rect 182345 516409 182375 516461
rect 182375 516409 182387 516461
rect 182387 516409 182401 516461
rect 182425 516409 182439 516461
rect 182439 516409 182451 516461
rect 182451 516409 182481 516461
rect 182505 516409 182515 516461
rect 182515 516409 182561 516461
rect 182265 516407 182321 516409
rect 182345 516407 182401 516409
rect 182425 516407 182481 516409
rect 182505 516407 182561 516409
rect 186083 516461 186139 516463
rect 186163 516461 186219 516463
rect 186243 516461 186299 516463
rect 186323 516461 186379 516463
rect 186083 516409 186129 516461
rect 186129 516409 186139 516461
rect 186163 516409 186193 516461
rect 186193 516409 186205 516461
rect 186205 516409 186219 516461
rect 186243 516409 186257 516461
rect 186257 516409 186269 516461
rect 186269 516409 186299 516461
rect 186323 516409 186333 516461
rect 186333 516409 186379 516461
rect 186083 516407 186139 516409
rect 186163 516407 186219 516409
rect 186243 516407 186299 516409
rect 186323 516407 186379 516409
rect 181605 515917 181661 515919
rect 181685 515917 181741 515919
rect 181765 515917 181821 515919
rect 181845 515917 181901 515919
rect 181605 515865 181651 515917
rect 181651 515865 181661 515917
rect 181685 515865 181715 515917
rect 181715 515865 181727 515917
rect 181727 515865 181741 515917
rect 181765 515865 181779 515917
rect 181779 515865 181791 515917
rect 181791 515865 181821 515917
rect 181845 515865 181855 515917
rect 181855 515865 181901 515917
rect 181605 515863 181661 515865
rect 181685 515863 181741 515865
rect 181765 515863 181821 515865
rect 181845 515863 181901 515865
rect 185423 515917 185479 515919
rect 185503 515917 185559 515919
rect 185583 515917 185639 515919
rect 185663 515917 185719 515919
rect 185423 515865 185469 515917
rect 185469 515865 185479 515917
rect 185503 515865 185533 515917
rect 185533 515865 185545 515917
rect 185545 515865 185559 515917
rect 185583 515865 185597 515917
rect 185597 515865 185609 515917
rect 185609 515865 185639 515917
rect 185663 515865 185673 515917
rect 185673 515865 185719 515917
rect 185423 515863 185479 515865
rect 185503 515863 185559 515865
rect 185583 515863 185639 515865
rect 185663 515863 185719 515865
rect 178447 515373 178503 515375
rect 178527 515373 178583 515375
rect 178607 515373 178663 515375
rect 178687 515373 178743 515375
rect 178447 515321 178493 515373
rect 178493 515321 178503 515373
rect 178527 515321 178557 515373
rect 178557 515321 178569 515373
rect 178569 515321 178583 515373
rect 178607 515321 178621 515373
rect 178621 515321 178633 515373
rect 178633 515321 178663 515373
rect 178687 515321 178697 515373
rect 178697 515321 178743 515373
rect 178447 515319 178503 515321
rect 178527 515319 178583 515321
rect 178607 515319 178663 515321
rect 178687 515319 178743 515321
rect 182265 515373 182321 515375
rect 182345 515373 182401 515375
rect 182425 515373 182481 515375
rect 182505 515373 182561 515375
rect 182265 515321 182311 515373
rect 182311 515321 182321 515373
rect 182345 515321 182375 515373
rect 182375 515321 182387 515373
rect 182387 515321 182401 515373
rect 182425 515321 182439 515373
rect 182439 515321 182451 515373
rect 182451 515321 182481 515373
rect 182505 515321 182515 515373
rect 182515 515321 182561 515373
rect 182265 515319 182321 515321
rect 182345 515319 182401 515321
rect 182425 515319 182481 515321
rect 182505 515319 182561 515321
rect 186083 515373 186139 515375
rect 186163 515373 186219 515375
rect 186243 515373 186299 515375
rect 186323 515373 186379 515375
rect 186083 515321 186129 515373
rect 186129 515321 186139 515373
rect 186163 515321 186193 515373
rect 186193 515321 186205 515373
rect 186205 515321 186219 515373
rect 186243 515321 186257 515373
rect 186257 515321 186269 515373
rect 186269 515321 186299 515373
rect 186323 515321 186333 515373
rect 186333 515321 186379 515373
rect 186083 515319 186139 515321
rect 186163 515319 186219 515321
rect 186243 515319 186299 515321
rect 186323 515319 186379 515321
rect 2000 507000 4000 509000
rect 2000 464000 4000 466000
rect 2000 421000 4000 423000
rect 2000 378000 4000 380000
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 18000 701005 20000 702300
rect 70000 701005 72000 702300
rect 122000 701005 124000 702300
rect 17990 701000 20010 701005
rect 17990 699000 18000 701000
rect 20000 699000 20010 701000
rect 17990 698995 20010 699000
rect 69990 701000 72010 701005
rect 69990 699000 70000 701000
rect 72000 699000 72010 701000
rect 69990 698995 72010 699000
rect 121990 701000 124010 701005
rect 121990 699000 122000 701000
rect 124000 699000 124010 701000
rect 121990 698995 124010 699000
rect -800 684000 1700 685242
rect 2990 684000 5010 684005
rect -800 682000 3000 684000
rect 5000 682000 5010 684000
rect -800 680242 1700 682000
rect 2990 681995 5010 682000
rect 157609 541837 162708 541865
rect 157609 538893 162624 541837
rect 162688 538893 162708 541837
rect 157609 538865 162708 538893
rect 163118 540255 191998 540265
rect 163118 540245 174188 540255
rect 163118 540065 166688 540245
rect 166868 540065 170488 540245
rect 170668 540075 174188 540245
rect 174368 540245 191998 540255
rect 174368 540075 177698 540245
rect 170668 540065 177698 540075
rect 177878 540065 181288 540245
rect 181468 540065 184588 540245
rect 184768 540065 187898 540245
rect 188078 540065 191188 540245
rect 191368 540065 191808 540245
rect 191988 540065 191998 540245
rect 163118 540045 191998 540065
rect 163118 538870 163338 540045
rect 163018 538865 163338 538870
rect 161378 538665 161528 538675
rect 159388 538655 159488 538665
rect 159388 538555 159398 538655
rect 159478 538555 159488 538655
rect 159388 538545 159488 538555
rect 161378 538545 161388 538665
rect 161508 538545 161528 538665
rect 163018 538665 163028 538865
rect 163328 538665 163338 538865
rect 163018 538660 163338 538665
rect 163118 538555 163338 538660
rect 163898 539315 192008 539325
rect 163898 539305 191198 539315
rect 163898 539125 166688 539305
rect 166868 539125 170488 539305
rect 170668 539125 174188 539305
rect 174368 539125 177688 539305
rect 177868 539125 181288 539305
rect 181468 539125 184588 539305
rect 184768 539125 187888 539305
rect 188068 539135 191198 539305
rect 191378 539305 192008 539315
rect 191378 539135 191818 539305
rect 188068 539125 191818 539135
rect 191998 539125 192008 539305
rect 163898 539105 192008 539125
rect 161378 538535 161528 538545
rect 163898 535625 164118 539105
rect 160198 535565 164118 535625
rect 160198 535425 160208 535565
rect 160358 535425 164118 535565
rect 160198 535405 164118 535425
rect 174619 530611 174935 530612
rect 174619 530547 174625 530611
rect 174689 530547 174705 530611
rect 174769 530547 174785 530611
rect 174849 530547 174865 530611
rect 174929 530547 174935 530611
rect 174619 530546 174935 530547
rect 178437 530611 178753 530612
rect 178437 530547 178443 530611
rect 178507 530547 178523 530611
rect 178587 530547 178603 530611
rect 178667 530547 178683 530611
rect 178747 530547 178753 530611
rect 178437 530546 178753 530547
rect 182255 530611 182571 530612
rect 182255 530547 182261 530611
rect 182325 530547 182341 530611
rect 182405 530547 182421 530611
rect 182485 530547 182501 530611
rect 182565 530547 182571 530611
rect 182255 530546 182571 530547
rect 186073 530611 186389 530612
rect 186073 530547 186079 530611
rect 186143 530547 186159 530611
rect 186223 530547 186239 530611
rect 186303 530547 186319 530611
rect 186383 530547 186389 530611
rect 186073 530546 186389 530547
rect 173959 530067 174275 530068
rect 173959 530003 173965 530067
rect 174029 530003 174045 530067
rect 174109 530003 174125 530067
rect 174189 530003 174205 530067
rect 174269 530003 174275 530067
rect 173959 530002 174275 530003
rect 177777 530067 178093 530068
rect 177777 530003 177783 530067
rect 177847 530003 177863 530067
rect 177927 530003 177943 530067
rect 178007 530003 178023 530067
rect 178087 530003 178093 530067
rect 177777 530002 178093 530003
rect 181595 530067 181911 530068
rect 181595 530003 181601 530067
rect 181665 530003 181681 530067
rect 181745 530003 181761 530067
rect 181825 530003 181841 530067
rect 181905 530003 181911 530067
rect 181595 530002 181911 530003
rect 185413 530067 185729 530068
rect 185413 530003 185419 530067
rect 185483 530003 185499 530067
rect 185563 530003 185579 530067
rect 185643 530003 185659 530067
rect 185723 530003 185729 530067
rect 185413 530002 185729 530003
rect 174619 529523 174935 529524
rect 174619 529459 174625 529523
rect 174689 529459 174705 529523
rect 174769 529459 174785 529523
rect 174849 529459 174865 529523
rect 174929 529459 174935 529523
rect 174619 529458 174935 529459
rect 178437 529523 178753 529524
rect 178437 529459 178443 529523
rect 178507 529459 178523 529523
rect 178587 529459 178603 529523
rect 178667 529459 178683 529523
rect 178747 529459 178753 529523
rect 178437 529458 178753 529459
rect 182255 529523 182571 529524
rect 182255 529459 182261 529523
rect 182325 529459 182341 529523
rect 182405 529459 182421 529523
rect 182485 529459 182501 529523
rect 182565 529459 182571 529523
rect 182255 529458 182571 529459
rect 186073 529523 186389 529524
rect 186073 529459 186079 529523
rect 186143 529459 186159 529523
rect 186223 529459 186239 529523
rect 186303 529459 186319 529523
rect 186383 529459 186389 529523
rect 186073 529458 186389 529459
rect 173959 528979 174275 528980
rect 173959 528915 173965 528979
rect 174029 528915 174045 528979
rect 174109 528915 174125 528979
rect 174189 528915 174205 528979
rect 174269 528915 174275 528979
rect 173959 528914 174275 528915
rect 177777 528979 178093 528980
rect 177777 528915 177783 528979
rect 177847 528915 177863 528979
rect 177927 528915 177943 528979
rect 178007 528915 178023 528979
rect 178087 528915 178093 528979
rect 177777 528914 178093 528915
rect 181595 528979 181911 528980
rect 181595 528915 181601 528979
rect 181665 528915 181681 528979
rect 181745 528915 181761 528979
rect 181825 528915 181841 528979
rect 181905 528915 181911 528979
rect 181595 528914 181911 528915
rect 185413 528979 185729 528980
rect 185413 528915 185419 528979
rect 185483 528915 185499 528979
rect 185563 528915 185579 528979
rect 185643 528915 185659 528979
rect 185723 528915 185729 528979
rect 185413 528914 185729 528915
rect 174619 528435 174935 528436
rect 174619 528371 174625 528435
rect 174689 528371 174705 528435
rect 174769 528371 174785 528435
rect 174849 528371 174865 528435
rect 174929 528371 174935 528435
rect 174619 528370 174935 528371
rect 178437 528435 178753 528436
rect 178437 528371 178443 528435
rect 178507 528371 178523 528435
rect 178587 528371 178603 528435
rect 178667 528371 178683 528435
rect 178747 528371 178753 528435
rect 178437 528370 178753 528371
rect 182255 528435 182571 528436
rect 182255 528371 182261 528435
rect 182325 528371 182341 528435
rect 182405 528371 182421 528435
rect 182485 528371 182501 528435
rect 182565 528371 182571 528435
rect 182255 528370 182571 528371
rect 186073 528435 186389 528436
rect 186073 528371 186079 528435
rect 186143 528371 186159 528435
rect 186223 528371 186239 528435
rect 186303 528371 186319 528435
rect 186383 528371 186389 528435
rect 186073 528370 186389 528371
rect 173959 527891 174275 527892
rect 173959 527827 173965 527891
rect 174029 527827 174045 527891
rect 174109 527827 174125 527891
rect 174189 527827 174205 527891
rect 174269 527827 174275 527891
rect 173959 527826 174275 527827
rect 177777 527891 178093 527892
rect 177777 527827 177783 527891
rect 177847 527827 177863 527891
rect 177927 527827 177943 527891
rect 178007 527827 178023 527891
rect 178087 527827 178093 527891
rect 177777 527826 178093 527827
rect 181595 527891 181911 527892
rect 181595 527827 181601 527891
rect 181665 527827 181681 527891
rect 181745 527827 181761 527891
rect 181825 527827 181841 527891
rect 181905 527827 181911 527891
rect 181595 527826 181911 527827
rect 185413 527891 185729 527892
rect 185413 527827 185419 527891
rect 185483 527827 185499 527891
rect 185563 527827 185579 527891
rect 185643 527827 185659 527891
rect 185723 527827 185729 527891
rect 185413 527826 185729 527827
rect 174619 527347 174935 527348
rect 174619 527283 174625 527347
rect 174689 527283 174705 527347
rect 174769 527283 174785 527347
rect 174849 527283 174865 527347
rect 174929 527283 174935 527347
rect 174619 527282 174935 527283
rect 178437 527347 178753 527348
rect 178437 527283 178443 527347
rect 178507 527283 178523 527347
rect 178587 527283 178603 527347
rect 178667 527283 178683 527347
rect 178747 527283 178753 527347
rect 178437 527282 178753 527283
rect 182255 527347 182571 527348
rect 182255 527283 182261 527347
rect 182325 527283 182341 527347
rect 182405 527283 182421 527347
rect 182485 527283 182501 527347
rect 182565 527283 182571 527347
rect 182255 527282 182571 527283
rect 186073 527347 186389 527348
rect 186073 527283 186079 527347
rect 186143 527283 186159 527347
rect 186223 527283 186239 527347
rect 186303 527283 186319 527347
rect 186383 527283 186389 527347
rect 186073 527282 186389 527283
rect 173959 526803 174275 526804
rect 173959 526739 173965 526803
rect 174029 526739 174045 526803
rect 174109 526739 174125 526803
rect 174189 526739 174205 526803
rect 174269 526739 174275 526803
rect 173959 526738 174275 526739
rect 177777 526803 178093 526804
rect 177777 526739 177783 526803
rect 177847 526739 177863 526803
rect 177927 526739 177943 526803
rect 178007 526739 178023 526803
rect 178087 526739 178093 526803
rect 177777 526738 178093 526739
rect 181595 526803 181911 526804
rect 181595 526739 181601 526803
rect 181665 526739 181681 526803
rect 181745 526739 181761 526803
rect 181825 526739 181841 526803
rect 181905 526739 181911 526803
rect 181595 526738 181911 526739
rect 185413 526803 185729 526804
rect 185413 526739 185419 526803
rect 185483 526739 185499 526803
rect 185563 526739 185579 526803
rect 185643 526739 185659 526803
rect 185723 526739 185729 526803
rect 185413 526738 185729 526739
rect 174619 526259 174935 526260
rect 174619 526195 174625 526259
rect 174689 526195 174705 526259
rect 174769 526195 174785 526259
rect 174849 526195 174865 526259
rect 174929 526195 174935 526259
rect 174619 526194 174935 526195
rect 178437 526259 178753 526260
rect 178437 526195 178443 526259
rect 178507 526195 178523 526259
rect 178587 526195 178603 526259
rect 178667 526195 178683 526259
rect 178747 526195 178753 526259
rect 178437 526194 178753 526195
rect 182255 526259 182571 526260
rect 182255 526195 182261 526259
rect 182325 526195 182341 526259
rect 182405 526195 182421 526259
rect 182485 526195 182501 526259
rect 182565 526195 182571 526259
rect 182255 526194 182571 526195
rect 186073 526259 186389 526260
rect 186073 526195 186079 526259
rect 186143 526195 186159 526259
rect 186223 526195 186239 526259
rect 186303 526195 186319 526259
rect 186383 526195 186389 526259
rect 186073 526194 186389 526195
rect 173959 525715 174275 525716
rect 173959 525651 173965 525715
rect 174029 525651 174045 525715
rect 174109 525651 174125 525715
rect 174189 525651 174205 525715
rect 174269 525651 174275 525715
rect 173959 525650 174275 525651
rect 177777 525715 178093 525716
rect 177777 525651 177783 525715
rect 177847 525651 177863 525715
rect 177927 525651 177943 525715
rect 178007 525651 178023 525715
rect 178087 525651 178093 525715
rect 177777 525650 178093 525651
rect 181595 525715 181911 525716
rect 181595 525651 181601 525715
rect 181665 525651 181681 525715
rect 181745 525651 181761 525715
rect 181825 525651 181841 525715
rect 181905 525651 181911 525715
rect 181595 525650 181911 525651
rect 185413 525715 185729 525716
rect 185413 525651 185419 525715
rect 185483 525651 185499 525715
rect 185563 525651 185579 525715
rect 185643 525651 185659 525715
rect 185723 525651 185729 525715
rect 185413 525650 185729 525651
rect 174619 525171 174935 525172
rect 174619 525107 174625 525171
rect 174689 525107 174705 525171
rect 174769 525107 174785 525171
rect 174849 525107 174865 525171
rect 174929 525107 174935 525171
rect 174619 525106 174935 525107
rect 178437 525171 178753 525172
rect 178437 525107 178443 525171
rect 178507 525107 178523 525171
rect 178587 525107 178603 525171
rect 178667 525107 178683 525171
rect 178747 525107 178753 525171
rect 178437 525106 178753 525107
rect 182255 525171 182571 525172
rect 182255 525107 182261 525171
rect 182325 525107 182341 525171
rect 182405 525107 182421 525171
rect 182485 525107 182501 525171
rect 182565 525107 182571 525171
rect 182255 525106 182571 525107
rect 186073 525171 186389 525172
rect 186073 525107 186079 525171
rect 186143 525107 186159 525171
rect 186223 525107 186239 525171
rect 186303 525107 186319 525171
rect 186383 525107 186389 525171
rect 186073 525106 186389 525107
rect 173959 524627 174275 524628
rect 173959 524563 173965 524627
rect 174029 524563 174045 524627
rect 174109 524563 174125 524627
rect 174189 524563 174205 524627
rect 174269 524563 174275 524627
rect 173959 524562 174275 524563
rect 177777 524627 178093 524628
rect 177777 524563 177783 524627
rect 177847 524563 177863 524627
rect 177927 524563 177943 524627
rect 178007 524563 178023 524627
rect 178087 524563 178093 524627
rect 177777 524562 178093 524563
rect 181595 524627 181911 524628
rect 181595 524563 181601 524627
rect 181665 524563 181681 524627
rect 181745 524563 181761 524627
rect 181825 524563 181841 524627
rect 181905 524563 181911 524627
rect 181595 524562 181911 524563
rect 185413 524627 185729 524628
rect 185413 524563 185419 524627
rect 185483 524563 185499 524627
rect 185563 524563 185579 524627
rect 185643 524563 185659 524627
rect 185723 524563 185729 524627
rect 185413 524562 185729 524563
rect 174619 524083 174935 524084
rect 174619 524019 174625 524083
rect 174689 524019 174705 524083
rect 174769 524019 174785 524083
rect 174849 524019 174865 524083
rect 174929 524019 174935 524083
rect 174619 524018 174935 524019
rect 178437 524083 178753 524084
rect 178437 524019 178443 524083
rect 178507 524019 178523 524083
rect 178587 524019 178603 524083
rect 178667 524019 178683 524083
rect 178747 524019 178753 524083
rect 178437 524018 178753 524019
rect 182255 524083 182571 524084
rect 182255 524019 182261 524083
rect 182325 524019 182341 524083
rect 182405 524019 182421 524083
rect 182485 524019 182501 524083
rect 182565 524019 182571 524083
rect 182255 524018 182571 524019
rect 186073 524083 186389 524084
rect 186073 524019 186079 524083
rect 186143 524019 186159 524083
rect 186223 524019 186239 524083
rect 186303 524019 186319 524083
rect 186383 524019 186389 524083
rect 186073 524018 186389 524019
rect 173959 523539 174275 523540
rect 173959 523475 173965 523539
rect 174029 523475 174045 523539
rect 174109 523475 174125 523539
rect 174189 523475 174205 523539
rect 174269 523475 174275 523539
rect 173959 523474 174275 523475
rect 177777 523539 178093 523540
rect 177777 523475 177783 523539
rect 177847 523475 177863 523539
rect 177927 523475 177943 523539
rect 178007 523475 178023 523539
rect 178087 523475 178093 523539
rect 177777 523474 178093 523475
rect 181595 523539 181911 523540
rect 181595 523475 181601 523539
rect 181665 523475 181681 523539
rect 181745 523475 181761 523539
rect 181825 523475 181841 523539
rect 181905 523475 181911 523539
rect 181595 523474 181911 523475
rect 185413 523539 185729 523540
rect 185413 523475 185419 523539
rect 185483 523475 185499 523539
rect 185563 523475 185579 523539
rect 185643 523475 185659 523539
rect 185723 523475 185729 523539
rect 185413 523474 185729 523475
rect 174619 522995 174935 522996
rect 174619 522931 174625 522995
rect 174689 522931 174705 522995
rect 174769 522931 174785 522995
rect 174849 522931 174865 522995
rect 174929 522931 174935 522995
rect 174619 522930 174935 522931
rect 178437 522995 178753 522996
rect 178437 522931 178443 522995
rect 178507 522931 178523 522995
rect 178587 522931 178603 522995
rect 178667 522931 178683 522995
rect 178747 522931 178753 522995
rect 178437 522930 178753 522931
rect 182255 522995 182571 522996
rect 182255 522931 182261 522995
rect 182325 522931 182341 522995
rect 182405 522931 182421 522995
rect 182485 522931 182501 522995
rect 182565 522931 182571 522995
rect 182255 522930 182571 522931
rect 186073 522995 186389 522996
rect 186073 522931 186079 522995
rect 186143 522931 186159 522995
rect 186223 522931 186239 522995
rect 186303 522931 186319 522995
rect 186383 522931 186389 522995
rect 186073 522930 186389 522931
rect 173959 522451 174275 522452
rect 173959 522387 173965 522451
rect 174029 522387 174045 522451
rect 174109 522387 174125 522451
rect 174189 522387 174205 522451
rect 174269 522387 174275 522451
rect 173959 522386 174275 522387
rect 177777 522451 178093 522452
rect 177777 522387 177783 522451
rect 177847 522387 177863 522451
rect 177927 522387 177943 522451
rect 178007 522387 178023 522451
rect 178087 522387 178093 522451
rect 177777 522386 178093 522387
rect 181595 522451 181911 522452
rect 181595 522387 181601 522451
rect 181665 522387 181681 522451
rect 181745 522387 181761 522451
rect 181825 522387 181841 522451
rect 181905 522387 181911 522451
rect 181595 522386 181911 522387
rect 185413 522451 185729 522452
rect 185413 522387 185419 522451
rect 185483 522387 185499 522451
rect 185563 522387 185579 522451
rect 185643 522387 185659 522451
rect 185723 522387 185729 522451
rect 185413 522386 185729 522387
rect 174619 521907 174935 521908
rect 174619 521843 174625 521907
rect 174689 521843 174705 521907
rect 174769 521843 174785 521907
rect 174849 521843 174865 521907
rect 174929 521843 174935 521907
rect 174619 521842 174935 521843
rect 178437 521907 178753 521908
rect 178437 521843 178443 521907
rect 178507 521843 178523 521907
rect 178587 521843 178603 521907
rect 178667 521843 178683 521907
rect 178747 521843 178753 521907
rect 178437 521842 178753 521843
rect 182255 521907 182571 521908
rect 182255 521843 182261 521907
rect 182325 521843 182341 521907
rect 182405 521843 182421 521907
rect 182485 521843 182501 521907
rect 182565 521843 182571 521907
rect 182255 521842 182571 521843
rect 186073 521907 186389 521908
rect 186073 521843 186079 521907
rect 186143 521843 186159 521907
rect 186223 521843 186239 521907
rect 186303 521843 186319 521907
rect 186383 521843 186389 521907
rect 186073 521842 186389 521843
rect 173959 521363 174275 521364
rect 173959 521299 173965 521363
rect 174029 521299 174045 521363
rect 174109 521299 174125 521363
rect 174189 521299 174205 521363
rect 174269 521299 174275 521363
rect 173959 521298 174275 521299
rect 177777 521363 178093 521364
rect 177777 521299 177783 521363
rect 177847 521299 177863 521363
rect 177927 521299 177943 521363
rect 178007 521299 178023 521363
rect 178087 521299 178093 521363
rect 177777 521298 178093 521299
rect 181595 521363 181911 521364
rect 181595 521299 181601 521363
rect 181665 521299 181681 521363
rect 181745 521299 181761 521363
rect 181825 521299 181841 521363
rect 181905 521299 181911 521363
rect 181595 521298 181911 521299
rect 185413 521363 185729 521364
rect 185413 521299 185419 521363
rect 185483 521299 185499 521363
rect 185563 521299 185579 521363
rect 185643 521299 185659 521363
rect 185723 521299 185729 521363
rect 185413 521298 185729 521299
rect 174619 520819 174935 520820
rect 174619 520755 174625 520819
rect 174689 520755 174705 520819
rect 174769 520755 174785 520819
rect 174849 520755 174865 520819
rect 174929 520755 174935 520819
rect 174619 520754 174935 520755
rect 178437 520819 178753 520820
rect 178437 520755 178443 520819
rect 178507 520755 178523 520819
rect 178587 520755 178603 520819
rect 178667 520755 178683 520819
rect 178747 520755 178753 520819
rect 178437 520754 178753 520755
rect 182255 520819 182571 520820
rect 182255 520755 182261 520819
rect 182325 520755 182341 520819
rect 182405 520755 182421 520819
rect 182485 520755 182501 520819
rect 182565 520755 182571 520819
rect 182255 520754 182571 520755
rect 186073 520819 186389 520820
rect 186073 520755 186079 520819
rect 186143 520755 186159 520819
rect 186223 520755 186239 520819
rect 186303 520755 186319 520819
rect 186383 520755 186389 520819
rect 186073 520754 186389 520755
rect 173959 520275 174275 520276
rect 173959 520211 173965 520275
rect 174029 520211 174045 520275
rect 174109 520211 174125 520275
rect 174189 520211 174205 520275
rect 174269 520211 174275 520275
rect 173959 520210 174275 520211
rect 177777 520275 178093 520276
rect 177777 520211 177783 520275
rect 177847 520211 177863 520275
rect 177927 520211 177943 520275
rect 178007 520211 178023 520275
rect 178087 520211 178093 520275
rect 177777 520210 178093 520211
rect 181595 520275 181911 520276
rect 181595 520211 181601 520275
rect 181665 520211 181681 520275
rect 181745 520211 181761 520275
rect 181825 520211 181841 520275
rect 181905 520211 181911 520275
rect 181595 520210 181911 520211
rect 185413 520275 185729 520276
rect 185413 520211 185419 520275
rect 185483 520211 185499 520275
rect 185563 520211 185579 520275
rect 185643 520211 185659 520275
rect 185723 520211 185729 520275
rect 185413 520210 185729 520211
rect 174619 519731 174935 519732
rect 174619 519667 174625 519731
rect 174689 519667 174705 519731
rect 174769 519667 174785 519731
rect 174849 519667 174865 519731
rect 174929 519667 174935 519731
rect 174619 519666 174935 519667
rect 178437 519731 178753 519732
rect 178437 519667 178443 519731
rect 178507 519667 178523 519731
rect 178587 519667 178603 519731
rect 178667 519667 178683 519731
rect 178747 519667 178753 519731
rect 178437 519666 178753 519667
rect 182255 519731 182571 519732
rect 182255 519667 182261 519731
rect 182325 519667 182341 519731
rect 182405 519667 182421 519731
rect 182485 519667 182501 519731
rect 182565 519667 182571 519731
rect 182255 519666 182571 519667
rect 186073 519731 186389 519732
rect 186073 519667 186079 519731
rect 186143 519667 186159 519731
rect 186223 519667 186239 519731
rect 186303 519667 186319 519731
rect 186383 519667 186389 519731
rect 186073 519666 186389 519667
rect 173959 519187 174275 519188
rect 173959 519123 173965 519187
rect 174029 519123 174045 519187
rect 174109 519123 174125 519187
rect 174189 519123 174205 519187
rect 174269 519123 174275 519187
rect 173959 519122 174275 519123
rect 177777 519187 178093 519188
rect 177777 519123 177783 519187
rect 177847 519123 177863 519187
rect 177927 519123 177943 519187
rect 178007 519123 178023 519187
rect 178087 519123 178093 519187
rect 177777 519122 178093 519123
rect 181595 519187 181911 519188
rect 181595 519123 181601 519187
rect 181665 519123 181681 519187
rect 181745 519123 181761 519187
rect 181825 519123 181841 519187
rect 181905 519123 181911 519187
rect 181595 519122 181911 519123
rect 185413 519187 185729 519188
rect 185413 519123 185419 519187
rect 185483 519123 185499 519187
rect 185563 519123 185579 519187
rect 185643 519123 185659 519187
rect 185723 519123 185729 519187
rect 185413 519122 185729 519123
rect 174619 518643 174935 518644
rect 174619 518579 174625 518643
rect 174689 518579 174705 518643
rect 174769 518579 174785 518643
rect 174849 518579 174865 518643
rect 174929 518579 174935 518643
rect 174619 518578 174935 518579
rect 178437 518643 178753 518644
rect 178437 518579 178443 518643
rect 178507 518579 178523 518643
rect 178587 518579 178603 518643
rect 178667 518579 178683 518643
rect 178747 518579 178753 518643
rect 178437 518578 178753 518579
rect 182255 518643 182571 518644
rect 182255 518579 182261 518643
rect 182325 518579 182341 518643
rect 182405 518579 182421 518643
rect 182485 518579 182501 518643
rect 182565 518579 182571 518643
rect 182255 518578 182571 518579
rect 186073 518643 186389 518644
rect 186073 518579 186079 518643
rect 186143 518579 186159 518643
rect 186223 518579 186239 518643
rect 186303 518579 186319 518643
rect 186383 518579 186389 518643
rect 186073 518578 186389 518579
rect 173959 518099 174275 518100
rect 173959 518035 173965 518099
rect 174029 518035 174045 518099
rect 174109 518035 174125 518099
rect 174189 518035 174205 518099
rect 174269 518035 174275 518099
rect 173959 518034 174275 518035
rect 177777 518099 178093 518100
rect 177777 518035 177783 518099
rect 177847 518035 177863 518099
rect 177927 518035 177943 518099
rect 178007 518035 178023 518099
rect 178087 518035 178093 518099
rect 177777 518034 178093 518035
rect 181595 518099 181911 518100
rect 181595 518035 181601 518099
rect 181665 518035 181681 518099
rect 181745 518035 181761 518099
rect 181825 518035 181841 518099
rect 181905 518035 181911 518099
rect 181595 518034 181911 518035
rect 185413 518099 185729 518100
rect 185413 518035 185419 518099
rect 185483 518035 185499 518099
rect 185563 518035 185579 518099
rect 185643 518035 185659 518099
rect 185723 518035 185729 518099
rect 185413 518034 185729 518035
rect 174619 517555 174935 517556
rect 174619 517491 174625 517555
rect 174689 517491 174705 517555
rect 174769 517491 174785 517555
rect 174849 517491 174865 517555
rect 174929 517491 174935 517555
rect 174619 517490 174935 517491
rect 178437 517555 178753 517556
rect 178437 517491 178443 517555
rect 178507 517491 178523 517555
rect 178587 517491 178603 517555
rect 178667 517491 178683 517555
rect 178747 517491 178753 517555
rect 178437 517490 178753 517491
rect 182255 517555 182571 517556
rect 182255 517491 182261 517555
rect 182325 517491 182341 517555
rect 182405 517491 182421 517555
rect 182485 517491 182501 517555
rect 182565 517491 182571 517555
rect 182255 517490 182571 517491
rect 186073 517555 186389 517556
rect 186073 517491 186079 517555
rect 186143 517491 186159 517555
rect 186223 517491 186239 517555
rect 186303 517491 186319 517555
rect 186383 517491 186389 517555
rect 186073 517490 186389 517491
rect 173959 517011 174275 517012
rect 173959 516947 173965 517011
rect 174029 516947 174045 517011
rect 174109 516947 174125 517011
rect 174189 516947 174205 517011
rect 174269 516947 174275 517011
rect 173959 516946 174275 516947
rect 177777 517011 178093 517012
rect 177777 516947 177783 517011
rect 177847 516947 177863 517011
rect 177927 516947 177943 517011
rect 178007 516947 178023 517011
rect 178087 516947 178093 517011
rect 177777 516946 178093 516947
rect 181595 517011 181911 517012
rect 181595 516947 181601 517011
rect 181665 516947 181681 517011
rect 181745 516947 181761 517011
rect 181825 516947 181841 517011
rect 181905 516947 181911 517011
rect 181595 516946 181911 516947
rect 185413 517011 185729 517012
rect 185413 516947 185419 517011
rect 185483 516947 185499 517011
rect 185563 516947 185579 517011
rect 185643 516947 185659 517011
rect 185723 516947 185729 517011
rect 185413 516946 185729 516947
rect 174619 516467 174935 516468
rect 174619 516403 174625 516467
rect 174689 516403 174705 516467
rect 174769 516403 174785 516467
rect 174849 516403 174865 516467
rect 174929 516403 174935 516467
rect 174619 516402 174935 516403
rect 178437 516467 178753 516468
rect 178437 516403 178443 516467
rect 178507 516403 178523 516467
rect 178587 516403 178603 516467
rect 178667 516403 178683 516467
rect 178747 516403 178753 516467
rect 178437 516402 178753 516403
rect 182255 516467 182571 516468
rect 182255 516403 182261 516467
rect 182325 516403 182341 516467
rect 182405 516403 182421 516467
rect 182485 516403 182501 516467
rect 182565 516403 182571 516467
rect 182255 516402 182571 516403
rect 186073 516467 186389 516468
rect 186073 516403 186079 516467
rect 186143 516403 186159 516467
rect 186223 516403 186239 516467
rect 186303 516403 186319 516467
rect 186383 516403 186389 516467
rect 186073 516402 186389 516403
rect 173959 515923 174275 515924
rect 173959 515859 173965 515923
rect 174029 515859 174045 515923
rect 174109 515859 174125 515923
rect 174189 515859 174205 515923
rect 174269 515859 174275 515923
rect 173959 515858 174275 515859
rect 177777 515923 178093 515924
rect 177777 515859 177783 515923
rect 177847 515859 177863 515923
rect 177927 515859 177943 515923
rect 178007 515859 178023 515923
rect 178087 515859 178093 515923
rect 177777 515858 178093 515859
rect 181595 515923 181911 515924
rect 181595 515859 181601 515923
rect 181665 515859 181681 515923
rect 181745 515859 181761 515923
rect 181825 515859 181841 515923
rect 181905 515859 181911 515923
rect 181595 515858 181911 515859
rect 185413 515923 185729 515924
rect 185413 515859 185419 515923
rect 185483 515859 185499 515923
rect 185563 515859 185579 515923
rect 185643 515859 185659 515923
rect 185723 515859 185729 515923
rect 185413 515858 185729 515859
rect 174619 515379 174935 515380
rect 174619 515315 174625 515379
rect 174689 515315 174705 515379
rect 174769 515315 174785 515379
rect 174849 515315 174865 515379
rect 174929 515315 174935 515379
rect 174619 515314 174935 515315
rect 178437 515379 178753 515380
rect 178437 515315 178443 515379
rect 178507 515315 178523 515379
rect 178587 515315 178603 515379
rect 178667 515315 178683 515379
rect 178747 515315 178753 515379
rect 178437 515314 178753 515315
rect 182255 515379 182571 515380
rect 182255 515315 182261 515379
rect 182325 515315 182341 515379
rect 182405 515315 182421 515379
rect 182485 515315 182501 515379
rect 182565 515315 182571 515379
rect 182255 515314 182571 515315
rect 186073 515379 186389 515380
rect 186073 515315 186079 515379
rect 186143 515315 186159 515379
rect 186223 515315 186239 515379
rect 186303 515315 186319 515379
rect 186383 515315 186389 515379
rect 186073 515314 186389 515315
rect 1990 509000 4010 509005
rect 1000 508200 2000 509000
rect 400 508096 2000 508200
rect -800 507984 2000 508096
rect 400 507800 2000 507984
rect 1000 507000 2000 507800
rect 4000 507000 4010 509000
rect 1990 506995 4010 507000
rect 1990 466000 4010 466005
rect 1000 465000 2000 466000
rect 400 464874 2000 465000
rect -800 464762 2000 464874
rect 400 464600 2000 464762
rect 1000 464000 2000 464600
rect 4000 464000 4010 466000
rect 1990 463995 4010 464000
rect 1990 423000 4010 423005
rect 1000 421700 2000 423000
rect 400 421652 2000 421700
rect -800 421540 2000 421652
rect 400 421000 2000 421540
rect 4000 421000 4010 423000
rect 1990 420995 4010 421000
rect 1990 380000 4010 380005
rect 1000 378700 2000 380000
rect 400 378430 2000 378700
rect -800 378318 2000 378430
rect 400 378000 2000 378318
rect 4000 378000 4010 380000
rect 1990 377995 4010 378000
<< via3 >>
rect 162624 538893 162688 541837
rect 159398 538555 159478 538655
rect 161388 538545 161508 538665
rect 174625 530607 174689 530611
rect 174625 530551 174629 530607
rect 174629 530551 174685 530607
rect 174685 530551 174689 530607
rect 174625 530547 174689 530551
rect 174705 530607 174769 530611
rect 174705 530551 174709 530607
rect 174709 530551 174765 530607
rect 174765 530551 174769 530607
rect 174705 530547 174769 530551
rect 174785 530607 174849 530611
rect 174785 530551 174789 530607
rect 174789 530551 174845 530607
rect 174845 530551 174849 530607
rect 174785 530547 174849 530551
rect 174865 530607 174929 530611
rect 174865 530551 174869 530607
rect 174869 530551 174925 530607
rect 174925 530551 174929 530607
rect 174865 530547 174929 530551
rect 178443 530607 178507 530611
rect 178443 530551 178447 530607
rect 178447 530551 178503 530607
rect 178503 530551 178507 530607
rect 178443 530547 178507 530551
rect 178523 530607 178587 530611
rect 178523 530551 178527 530607
rect 178527 530551 178583 530607
rect 178583 530551 178587 530607
rect 178523 530547 178587 530551
rect 178603 530607 178667 530611
rect 178603 530551 178607 530607
rect 178607 530551 178663 530607
rect 178663 530551 178667 530607
rect 178603 530547 178667 530551
rect 178683 530607 178747 530611
rect 178683 530551 178687 530607
rect 178687 530551 178743 530607
rect 178743 530551 178747 530607
rect 178683 530547 178747 530551
rect 182261 530607 182325 530611
rect 182261 530551 182265 530607
rect 182265 530551 182321 530607
rect 182321 530551 182325 530607
rect 182261 530547 182325 530551
rect 182341 530607 182405 530611
rect 182341 530551 182345 530607
rect 182345 530551 182401 530607
rect 182401 530551 182405 530607
rect 182341 530547 182405 530551
rect 182421 530607 182485 530611
rect 182421 530551 182425 530607
rect 182425 530551 182481 530607
rect 182481 530551 182485 530607
rect 182421 530547 182485 530551
rect 182501 530607 182565 530611
rect 182501 530551 182505 530607
rect 182505 530551 182561 530607
rect 182561 530551 182565 530607
rect 182501 530547 182565 530551
rect 186079 530607 186143 530611
rect 186079 530551 186083 530607
rect 186083 530551 186139 530607
rect 186139 530551 186143 530607
rect 186079 530547 186143 530551
rect 186159 530607 186223 530611
rect 186159 530551 186163 530607
rect 186163 530551 186219 530607
rect 186219 530551 186223 530607
rect 186159 530547 186223 530551
rect 186239 530607 186303 530611
rect 186239 530551 186243 530607
rect 186243 530551 186299 530607
rect 186299 530551 186303 530607
rect 186239 530547 186303 530551
rect 186319 530607 186383 530611
rect 186319 530551 186323 530607
rect 186323 530551 186379 530607
rect 186379 530551 186383 530607
rect 186319 530547 186383 530551
rect 173965 530063 174029 530067
rect 173965 530007 173969 530063
rect 173969 530007 174025 530063
rect 174025 530007 174029 530063
rect 173965 530003 174029 530007
rect 174045 530063 174109 530067
rect 174045 530007 174049 530063
rect 174049 530007 174105 530063
rect 174105 530007 174109 530063
rect 174045 530003 174109 530007
rect 174125 530063 174189 530067
rect 174125 530007 174129 530063
rect 174129 530007 174185 530063
rect 174185 530007 174189 530063
rect 174125 530003 174189 530007
rect 174205 530063 174269 530067
rect 174205 530007 174209 530063
rect 174209 530007 174265 530063
rect 174265 530007 174269 530063
rect 174205 530003 174269 530007
rect 177783 530063 177847 530067
rect 177783 530007 177787 530063
rect 177787 530007 177843 530063
rect 177843 530007 177847 530063
rect 177783 530003 177847 530007
rect 177863 530063 177927 530067
rect 177863 530007 177867 530063
rect 177867 530007 177923 530063
rect 177923 530007 177927 530063
rect 177863 530003 177927 530007
rect 177943 530063 178007 530067
rect 177943 530007 177947 530063
rect 177947 530007 178003 530063
rect 178003 530007 178007 530063
rect 177943 530003 178007 530007
rect 178023 530063 178087 530067
rect 178023 530007 178027 530063
rect 178027 530007 178083 530063
rect 178083 530007 178087 530063
rect 178023 530003 178087 530007
rect 181601 530063 181665 530067
rect 181601 530007 181605 530063
rect 181605 530007 181661 530063
rect 181661 530007 181665 530063
rect 181601 530003 181665 530007
rect 181681 530063 181745 530067
rect 181681 530007 181685 530063
rect 181685 530007 181741 530063
rect 181741 530007 181745 530063
rect 181681 530003 181745 530007
rect 181761 530063 181825 530067
rect 181761 530007 181765 530063
rect 181765 530007 181821 530063
rect 181821 530007 181825 530063
rect 181761 530003 181825 530007
rect 181841 530063 181905 530067
rect 181841 530007 181845 530063
rect 181845 530007 181901 530063
rect 181901 530007 181905 530063
rect 181841 530003 181905 530007
rect 185419 530063 185483 530067
rect 185419 530007 185423 530063
rect 185423 530007 185479 530063
rect 185479 530007 185483 530063
rect 185419 530003 185483 530007
rect 185499 530063 185563 530067
rect 185499 530007 185503 530063
rect 185503 530007 185559 530063
rect 185559 530007 185563 530063
rect 185499 530003 185563 530007
rect 185579 530063 185643 530067
rect 185579 530007 185583 530063
rect 185583 530007 185639 530063
rect 185639 530007 185643 530063
rect 185579 530003 185643 530007
rect 185659 530063 185723 530067
rect 185659 530007 185663 530063
rect 185663 530007 185719 530063
rect 185719 530007 185723 530063
rect 185659 530003 185723 530007
rect 174625 529519 174689 529523
rect 174625 529463 174629 529519
rect 174629 529463 174685 529519
rect 174685 529463 174689 529519
rect 174625 529459 174689 529463
rect 174705 529519 174769 529523
rect 174705 529463 174709 529519
rect 174709 529463 174765 529519
rect 174765 529463 174769 529519
rect 174705 529459 174769 529463
rect 174785 529519 174849 529523
rect 174785 529463 174789 529519
rect 174789 529463 174845 529519
rect 174845 529463 174849 529519
rect 174785 529459 174849 529463
rect 174865 529519 174929 529523
rect 174865 529463 174869 529519
rect 174869 529463 174925 529519
rect 174925 529463 174929 529519
rect 174865 529459 174929 529463
rect 178443 529519 178507 529523
rect 178443 529463 178447 529519
rect 178447 529463 178503 529519
rect 178503 529463 178507 529519
rect 178443 529459 178507 529463
rect 178523 529519 178587 529523
rect 178523 529463 178527 529519
rect 178527 529463 178583 529519
rect 178583 529463 178587 529519
rect 178523 529459 178587 529463
rect 178603 529519 178667 529523
rect 178603 529463 178607 529519
rect 178607 529463 178663 529519
rect 178663 529463 178667 529519
rect 178603 529459 178667 529463
rect 178683 529519 178747 529523
rect 178683 529463 178687 529519
rect 178687 529463 178743 529519
rect 178743 529463 178747 529519
rect 178683 529459 178747 529463
rect 182261 529519 182325 529523
rect 182261 529463 182265 529519
rect 182265 529463 182321 529519
rect 182321 529463 182325 529519
rect 182261 529459 182325 529463
rect 182341 529519 182405 529523
rect 182341 529463 182345 529519
rect 182345 529463 182401 529519
rect 182401 529463 182405 529519
rect 182341 529459 182405 529463
rect 182421 529519 182485 529523
rect 182421 529463 182425 529519
rect 182425 529463 182481 529519
rect 182481 529463 182485 529519
rect 182421 529459 182485 529463
rect 182501 529519 182565 529523
rect 182501 529463 182505 529519
rect 182505 529463 182561 529519
rect 182561 529463 182565 529519
rect 182501 529459 182565 529463
rect 186079 529519 186143 529523
rect 186079 529463 186083 529519
rect 186083 529463 186139 529519
rect 186139 529463 186143 529519
rect 186079 529459 186143 529463
rect 186159 529519 186223 529523
rect 186159 529463 186163 529519
rect 186163 529463 186219 529519
rect 186219 529463 186223 529519
rect 186159 529459 186223 529463
rect 186239 529519 186303 529523
rect 186239 529463 186243 529519
rect 186243 529463 186299 529519
rect 186299 529463 186303 529519
rect 186239 529459 186303 529463
rect 186319 529519 186383 529523
rect 186319 529463 186323 529519
rect 186323 529463 186379 529519
rect 186379 529463 186383 529519
rect 186319 529459 186383 529463
rect 173965 528975 174029 528979
rect 173965 528919 173969 528975
rect 173969 528919 174025 528975
rect 174025 528919 174029 528975
rect 173965 528915 174029 528919
rect 174045 528975 174109 528979
rect 174045 528919 174049 528975
rect 174049 528919 174105 528975
rect 174105 528919 174109 528975
rect 174045 528915 174109 528919
rect 174125 528975 174189 528979
rect 174125 528919 174129 528975
rect 174129 528919 174185 528975
rect 174185 528919 174189 528975
rect 174125 528915 174189 528919
rect 174205 528975 174269 528979
rect 174205 528919 174209 528975
rect 174209 528919 174265 528975
rect 174265 528919 174269 528975
rect 174205 528915 174269 528919
rect 177783 528975 177847 528979
rect 177783 528919 177787 528975
rect 177787 528919 177843 528975
rect 177843 528919 177847 528975
rect 177783 528915 177847 528919
rect 177863 528975 177927 528979
rect 177863 528919 177867 528975
rect 177867 528919 177923 528975
rect 177923 528919 177927 528975
rect 177863 528915 177927 528919
rect 177943 528975 178007 528979
rect 177943 528919 177947 528975
rect 177947 528919 178003 528975
rect 178003 528919 178007 528975
rect 177943 528915 178007 528919
rect 178023 528975 178087 528979
rect 178023 528919 178027 528975
rect 178027 528919 178083 528975
rect 178083 528919 178087 528975
rect 178023 528915 178087 528919
rect 181601 528975 181665 528979
rect 181601 528919 181605 528975
rect 181605 528919 181661 528975
rect 181661 528919 181665 528975
rect 181601 528915 181665 528919
rect 181681 528975 181745 528979
rect 181681 528919 181685 528975
rect 181685 528919 181741 528975
rect 181741 528919 181745 528975
rect 181681 528915 181745 528919
rect 181761 528975 181825 528979
rect 181761 528919 181765 528975
rect 181765 528919 181821 528975
rect 181821 528919 181825 528975
rect 181761 528915 181825 528919
rect 181841 528975 181905 528979
rect 181841 528919 181845 528975
rect 181845 528919 181901 528975
rect 181901 528919 181905 528975
rect 181841 528915 181905 528919
rect 185419 528975 185483 528979
rect 185419 528919 185423 528975
rect 185423 528919 185479 528975
rect 185479 528919 185483 528975
rect 185419 528915 185483 528919
rect 185499 528975 185563 528979
rect 185499 528919 185503 528975
rect 185503 528919 185559 528975
rect 185559 528919 185563 528975
rect 185499 528915 185563 528919
rect 185579 528975 185643 528979
rect 185579 528919 185583 528975
rect 185583 528919 185639 528975
rect 185639 528919 185643 528975
rect 185579 528915 185643 528919
rect 185659 528975 185723 528979
rect 185659 528919 185663 528975
rect 185663 528919 185719 528975
rect 185719 528919 185723 528975
rect 185659 528915 185723 528919
rect 174625 528431 174689 528435
rect 174625 528375 174629 528431
rect 174629 528375 174685 528431
rect 174685 528375 174689 528431
rect 174625 528371 174689 528375
rect 174705 528431 174769 528435
rect 174705 528375 174709 528431
rect 174709 528375 174765 528431
rect 174765 528375 174769 528431
rect 174705 528371 174769 528375
rect 174785 528431 174849 528435
rect 174785 528375 174789 528431
rect 174789 528375 174845 528431
rect 174845 528375 174849 528431
rect 174785 528371 174849 528375
rect 174865 528431 174929 528435
rect 174865 528375 174869 528431
rect 174869 528375 174925 528431
rect 174925 528375 174929 528431
rect 174865 528371 174929 528375
rect 178443 528431 178507 528435
rect 178443 528375 178447 528431
rect 178447 528375 178503 528431
rect 178503 528375 178507 528431
rect 178443 528371 178507 528375
rect 178523 528431 178587 528435
rect 178523 528375 178527 528431
rect 178527 528375 178583 528431
rect 178583 528375 178587 528431
rect 178523 528371 178587 528375
rect 178603 528431 178667 528435
rect 178603 528375 178607 528431
rect 178607 528375 178663 528431
rect 178663 528375 178667 528431
rect 178603 528371 178667 528375
rect 178683 528431 178747 528435
rect 178683 528375 178687 528431
rect 178687 528375 178743 528431
rect 178743 528375 178747 528431
rect 178683 528371 178747 528375
rect 182261 528431 182325 528435
rect 182261 528375 182265 528431
rect 182265 528375 182321 528431
rect 182321 528375 182325 528431
rect 182261 528371 182325 528375
rect 182341 528431 182405 528435
rect 182341 528375 182345 528431
rect 182345 528375 182401 528431
rect 182401 528375 182405 528431
rect 182341 528371 182405 528375
rect 182421 528431 182485 528435
rect 182421 528375 182425 528431
rect 182425 528375 182481 528431
rect 182481 528375 182485 528431
rect 182421 528371 182485 528375
rect 182501 528431 182565 528435
rect 182501 528375 182505 528431
rect 182505 528375 182561 528431
rect 182561 528375 182565 528431
rect 182501 528371 182565 528375
rect 186079 528431 186143 528435
rect 186079 528375 186083 528431
rect 186083 528375 186139 528431
rect 186139 528375 186143 528431
rect 186079 528371 186143 528375
rect 186159 528431 186223 528435
rect 186159 528375 186163 528431
rect 186163 528375 186219 528431
rect 186219 528375 186223 528431
rect 186159 528371 186223 528375
rect 186239 528431 186303 528435
rect 186239 528375 186243 528431
rect 186243 528375 186299 528431
rect 186299 528375 186303 528431
rect 186239 528371 186303 528375
rect 186319 528431 186383 528435
rect 186319 528375 186323 528431
rect 186323 528375 186379 528431
rect 186379 528375 186383 528431
rect 186319 528371 186383 528375
rect 173965 527887 174029 527891
rect 173965 527831 173969 527887
rect 173969 527831 174025 527887
rect 174025 527831 174029 527887
rect 173965 527827 174029 527831
rect 174045 527887 174109 527891
rect 174045 527831 174049 527887
rect 174049 527831 174105 527887
rect 174105 527831 174109 527887
rect 174045 527827 174109 527831
rect 174125 527887 174189 527891
rect 174125 527831 174129 527887
rect 174129 527831 174185 527887
rect 174185 527831 174189 527887
rect 174125 527827 174189 527831
rect 174205 527887 174269 527891
rect 174205 527831 174209 527887
rect 174209 527831 174265 527887
rect 174265 527831 174269 527887
rect 174205 527827 174269 527831
rect 177783 527887 177847 527891
rect 177783 527831 177787 527887
rect 177787 527831 177843 527887
rect 177843 527831 177847 527887
rect 177783 527827 177847 527831
rect 177863 527887 177927 527891
rect 177863 527831 177867 527887
rect 177867 527831 177923 527887
rect 177923 527831 177927 527887
rect 177863 527827 177927 527831
rect 177943 527887 178007 527891
rect 177943 527831 177947 527887
rect 177947 527831 178003 527887
rect 178003 527831 178007 527887
rect 177943 527827 178007 527831
rect 178023 527887 178087 527891
rect 178023 527831 178027 527887
rect 178027 527831 178083 527887
rect 178083 527831 178087 527887
rect 178023 527827 178087 527831
rect 181601 527887 181665 527891
rect 181601 527831 181605 527887
rect 181605 527831 181661 527887
rect 181661 527831 181665 527887
rect 181601 527827 181665 527831
rect 181681 527887 181745 527891
rect 181681 527831 181685 527887
rect 181685 527831 181741 527887
rect 181741 527831 181745 527887
rect 181681 527827 181745 527831
rect 181761 527887 181825 527891
rect 181761 527831 181765 527887
rect 181765 527831 181821 527887
rect 181821 527831 181825 527887
rect 181761 527827 181825 527831
rect 181841 527887 181905 527891
rect 181841 527831 181845 527887
rect 181845 527831 181901 527887
rect 181901 527831 181905 527887
rect 181841 527827 181905 527831
rect 185419 527887 185483 527891
rect 185419 527831 185423 527887
rect 185423 527831 185479 527887
rect 185479 527831 185483 527887
rect 185419 527827 185483 527831
rect 185499 527887 185563 527891
rect 185499 527831 185503 527887
rect 185503 527831 185559 527887
rect 185559 527831 185563 527887
rect 185499 527827 185563 527831
rect 185579 527887 185643 527891
rect 185579 527831 185583 527887
rect 185583 527831 185639 527887
rect 185639 527831 185643 527887
rect 185579 527827 185643 527831
rect 185659 527887 185723 527891
rect 185659 527831 185663 527887
rect 185663 527831 185719 527887
rect 185719 527831 185723 527887
rect 185659 527827 185723 527831
rect 174625 527343 174689 527347
rect 174625 527287 174629 527343
rect 174629 527287 174685 527343
rect 174685 527287 174689 527343
rect 174625 527283 174689 527287
rect 174705 527343 174769 527347
rect 174705 527287 174709 527343
rect 174709 527287 174765 527343
rect 174765 527287 174769 527343
rect 174705 527283 174769 527287
rect 174785 527343 174849 527347
rect 174785 527287 174789 527343
rect 174789 527287 174845 527343
rect 174845 527287 174849 527343
rect 174785 527283 174849 527287
rect 174865 527343 174929 527347
rect 174865 527287 174869 527343
rect 174869 527287 174925 527343
rect 174925 527287 174929 527343
rect 174865 527283 174929 527287
rect 178443 527343 178507 527347
rect 178443 527287 178447 527343
rect 178447 527287 178503 527343
rect 178503 527287 178507 527343
rect 178443 527283 178507 527287
rect 178523 527343 178587 527347
rect 178523 527287 178527 527343
rect 178527 527287 178583 527343
rect 178583 527287 178587 527343
rect 178523 527283 178587 527287
rect 178603 527343 178667 527347
rect 178603 527287 178607 527343
rect 178607 527287 178663 527343
rect 178663 527287 178667 527343
rect 178603 527283 178667 527287
rect 178683 527343 178747 527347
rect 178683 527287 178687 527343
rect 178687 527287 178743 527343
rect 178743 527287 178747 527343
rect 178683 527283 178747 527287
rect 182261 527343 182325 527347
rect 182261 527287 182265 527343
rect 182265 527287 182321 527343
rect 182321 527287 182325 527343
rect 182261 527283 182325 527287
rect 182341 527343 182405 527347
rect 182341 527287 182345 527343
rect 182345 527287 182401 527343
rect 182401 527287 182405 527343
rect 182341 527283 182405 527287
rect 182421 527343 182485 527347
rect 182421 527287 182425 527343
rect 182425 527287 182481 527343
rect 182481 527287 182485 527343
rect 182421 527283 182485 527287
rect 182501 527343 182565 527347
rect 182501 527287 182505 527343
rect 182505 527287 182561 527343
rect 182561 527287 182565 527343
rect 182501 527283 182565 527287
rect 186079 527343 186143 527347
rect 186079 527287 186083 527343
rect 186083 527287 186139 527343
rect 186139 527287 186143 527343
rect 186079 527283 186143 527287
rect 186159 527343 186223 527347
rect 186159 527287 186163 527343
rect 186163 527287 186219 527343
rect 186219 527287 186223 527343
rect 186159 527283 186223 527287
rect 186239 527343 186303 527347
rect 186239 527287 186243 527343
rect 186243 527287 186299 527343
rect 186299 527287 186303 527343
rect 186239 527283 186303 527287
rect 186319 527343 186383 527347
rect 186319 527287 186323 527343
rect 186323 527287 186379 527343
rect 186379 527287 186383 527343
rect 186319 527283 186383 527287
rect 173965 526799 174029 526803
rect 173965 526743 173969 526799
rect 173969 526743 174025 526799
rect 174025 526743 174029 526799
rect 173965 526739 174029 526743
rect 174045 526799 174109 526803
rect 174045 526743 174049 526799
rect 174049 526743 174105 526799
rect 174105 526743 174109 526799
rect 174045 526739 174109 526743
rect 174125 526799 174189 526803
rect 174125 526743 174129 526799
rect 174129 526743 174185 526799
rect 174185 526743 174189 526799
rect 174125 526739 174189 526743
rect 174205 526799 174269 526803
rect 174205 526743 174209 526799
rect 174209 526743 174265 526799
rect 174265 526743 174269 526799
rect 174205 526739 174269 526743
rect 177783 526799 177847 526803
rect 177783 526743 177787 526799
rect 177787 526743 177843 526799
rect 177843 526743 177847 526799
rect 177783 526739 177847 526743
rect 177863 526799 177927 526803
rect 177863 526743 177867 526799
rect 177867 526743 177923 526799
rect 177923 526743 177927 526799
rect 177863 526739 177927 526743
rect 177943 526799 178007 526803
rect 177943 526743 177947 526799
rect 177947 526743 178003 526799
rect 178003 526743 178007 526799
rect 177943 526739 178007 526743
rect 178023 526799 178087 526803
rect 178023 526743 178027 526799
rect 178027 526743 178083 526799
rect 178083 526743 178087 526799
rect 178023 526739 178087 526743
rect 181601 526799 181665 526803
rect 181601 526743 181605 526799
rect 181605 526743 181661 526799
rect 181661 526743 181665 526799
rect 181601 526739 181665 526743
rect 181681 526799 181745 526803
rect 181681 526743 181685 526799
rect 181685 526743 181741 526799
rect 181741 526743 181745 526799
rect 181681 526739 181745 526743
rect 181761 526799 181825 526803
rect 181761 526743 181765 526799
rect 181765 526743 181821 526799
rect 181821 526743 181825 526799
rect 181761 526739 181825 526743
rect 181841 526799 181905 526803
rect 181841 526743 181845 526799
rect 181845 526743 181901 526799
rect 181901 526743 181905 526799
rect 181841 526739 181905 526743
rect 185419 526799 185483 526803
rect 185419 526743 185423 526799
rect 185423 526743 185479 526799
rect 185479 526743 185483 526799
rect 185419 526739 185483 526743
rect 185499 526799 185563 526803
rect 185499 526743 185503 526799
rect 185503 526743 185559 526799
rect 185559 526743 185563 526799
rect 185499 526739 185563 526743
rect 185579 526799 185643 526803
rect 185579 526743 185583 526799
rect 185583 526743 185639 526799
rect 185639 526743 185643 526799
rect 185579 526739 185643 526743
rect 185659 526799 185723 526803
rect 185659 526743 185663 526799
rect 185663 526743 185719 526799
rect 185719 526743 185723 526799
rect 185659 526739 185723 526743
rect 174625 526255 174689 526259
rect 174625 526199 174629 526255
rect 174629 526199 174685 526255
rect 174685 526199 174689 526255
rect 174625 526195 174689 526199
rect 174705 526255 174769 526259
rect 174705 526199 174709 526255
rect 174709 526199 174765 526255
rect 174765 526199 174769 526255
rect 174705 526195 174769 526199
rect 174785 526255 174849 526259
rect 174785 526199 174789 526255
rect 174789 526199 174845 526255
rect 174845 526199 174849 526255
rect 174785 526195 174849 526199
rect 174865 526255 174929 526259
rect 174865 526199 174869 526255
rect 174869 526199 174925 526255
rect 174925 526199 174929 526255
rect 174865 526195 174929 526199
rect 178443 526255 178507 526259
rect 178443 526199 178447 526255
rect 178447 526199 178503 526255
rect 178503 526199 178507 526255
rect 178443 526195 178507 526199
rect 178523 526255 178587 526259
rect 178523 526199 178527 526255
rect 178527 526199 178583 526255
rect 178583 526199 178587 526255
rect 178523 526195 178587 526199
rect 178603 526255 178667 526259
rect 178603 526199 178607 526255
rect 178607 526199 178663 526255
rect 178663 526199 178667 526255
rect 178603 526195 178667 526199
rect 178683 526255 178747 526259
rect 178683 526199 178687 526255
rect 178687 526199 178743 526255
rect 178743 526199 178747 526255
rect 178683 526195 178747 526199
rect 182261 526255 182325 526259
rect 182261 526199 182265 526255
rect 182265 526199 182321 526255
rect 182321 526199 182325 526255
rect 182261 526195 182325 526199
rect 182341 526255 182405 526259
rect 182341 526199 182345 526255
rect 182345 526199 182401 526255
rect 182401 526199 182405 526255
rect 182341 526195 182405 526199
rect 182421 526255 182485 526259
rect 182421 526199 182425 526255
rect 182425 526199 182481 526255
rect 182481 526199 182485 526255
rect 182421 526195 182485 526199
rect 182501 526255 182565 526259
rect 182501 526199 182505 526255
rect 182505 526199 182561 526255
rect 182561 526199 182565 526255
rect 182501 526195 182565 526199
rect 186079 526255 186143 526259
rect 186079 526199 186083 526255
rect 186083 526199 186139 526255
rect 186139 526199 186143 526255
rect 186079 526195 186143 526199
rect 186159 526255 186223 526259
rect 186159 526199 186163 526255
rect 186163 526199 186219 526255
rect 186219 526199 186223 526255
rect 186159 526195 186223 526199
rect 186239 526255 186303 526259
rect 186239 526199 186243 526255
rect 186243 526199 186299 526255
rect 186299 526199 186303 526255
rect 186239 526195 186303 526199
rect 186319 526255 186383 526259
rect 186319 526199 186323 526255
rect 186323 526199 186379 526255
rect 186379 526199 186383 526255
rect 186319 526195 186383 526199
rect 173965 525711 174029 525715
rect 173965 525655 173969 525711
rect 173969 525655 174025 525711
rect 174025 525655 174029 525711
rect 173965 525651 174029 525655
rect 174045 525711 174109 525715
rect 174045 525655 174049 525711
rect 174049 525655 174105 525711
rect 174105 525655 174109 525711
rect 174045 525651 174109 525655
rect 174125 525711 174189 525715
rect 174125 525655 174129 525711
rect 174129 525655 174185 525711
rect 174185 525655 174189 525711
rect 174125 525651 174189 525655
rect 174205 525711 174269 525715
rect 174205 525655 174209 525711
rect 174209 525655 174265 525711
rect 174265 525655 174269 525711
rect 174205 525651 174269 525655
rect 177783 525711 177847 525715
rect 177783 525655 177787 525711
rect 177787 525655 177843 525711
rect 177843 525655 177847 525711
rect 177783 525651 177847 525655
rect 177863 525711 177927 525715
rect 177863 525655 177867 525711
rect 177867 525655 177923 525711
rect 177923 525655 177927 525711
rect 177863 525651 177927 525655
rect 177943 525711 178007 525715
rect 177943 525655 177947 525711
rect 177947 525655 178003 525711
rect 178003 525655 178007 525711
rect 177943 525651 178007 525655
rect 178023 525711 178087 525715
rect 178023 525655 178027 525711
rect 178027 525655 178083 525711
rect 178083 525655 178087 525711
rect 178023 525651 178087 525655
rect 181601 525711 181665 525715
rect 181601 525655 181605 525711
rect 181605 525655 181661 525711
rect 181661 525655 181665 525711
rect 181601 525651 181665 525655
rect 181681 525711 181745 525715
rect 181681 525655 181685 525711
rect 181685 525655 181741 525711
rect 181741 525655 181745 525711
rect 181681 525651 181745 525655
rect 181761 525711 181825 525715
rect 181761 525655 181765 525711
rect 181765 525655 181821 525711
rect 181821 525655 181825 525711
rect 181761 525651 181825 525655
rect 181841 525711 181905 525715
rect 181841 525655 181845 525711
rect 181845 525655 181901 525711
rect 181901 525655 181905 525711
rect 181841 525651 181905 525655
rect 185419 525711 185483 525715
rect 185419 525655 185423 525711
rect 185423 525655 185479 525711
rect 185479 525655 185483 525711
rect 185419 525651 185483 525655
rect 185499 525711 185563 525715
rect 185499 525655 185503 525711
rect 185503 525655 185559 525711
rect 185559 525655 185563 525711
rect 185499 525651 185563 525655
rect 185579 525711 185643 525715
rect 185579 525655 185583 525711
rect 185583 525655 185639 525711
rect 185639 525655 185643 525711
rect 185579 525651 185643 525655
rect 185659 525711 185723 525715
rect 185659 525655 185663 525711
rect 185663 525655 185719 525711
rect 185719 525655 185723 525711
rect 185659 525651 185723 525655
rect 174625 525167 174689 525171
rect 174625 525111 174629 525167
rect 174629 525111 174685 525167
rect 174685 525111 174689 525167
rect 174625 525107 174689 525111
rect 174705 525167 174769 525171
rect 174705 525111 174709 525167
rect 174709 525111 174765 525167
rect 174765 525111 174769 525167
rect 174705 525107 174769 525111
rect 174785 525167 174849 525171
rect 174785 525111 174789 525167
rect 174789 525111 174845 525167
rect 174845 525111 174849 525167
rect 174785 525107 174849 525111
rect 174865 525167 174929 525171
rect 174865 525111 174869 525167
rect 174869 525111 174925 525167
rect 174925 525111 174929 525167
rect 174865 525107 174929 525111
rect 178443 525167 178507 525171
rect 178443 525111 178447 525167
rect 178447 525111 178503 525167
rect 178503 525111 178507 525167
rect 178443 525107 178507 525111
rect 178523 525167 178587 525171
rect 178523 525111 178527 525167
rect 178527 525111 178583 525167
rect 178583 525111 178587 525167
rect 178523 525107 178587 525111
rect 178603 525167 178667 525171
rect 178603 525111 178607 525167
rect 178607 525111 178663 525167
rect 178663 525111 178667 525167
rect 178603 525107 178667 525111
rect 178683 525167 178747 525171
rect 178683 525111 178687 525167
rect 178687 525111 178743 525167
rect 178743 525111 178747 525167
rect 178683 525107 178747 525111
rect 182261 525167 182325 525171
rect 182261 525111 182265 525167
rect 182265 525111 182321 525167
rect 182321 525111 182325 525167
rect 182261 525107 182325 525111
rect 182341 525167 182405 525171
rect 182341 525111 182345 525167
rect 182345 525111 182401 525167
rect 182401 525111 182405 525167
rect 182341 525107 182405 525111
rect 182421 525167 182485 525171
rect 182421 525111 182425 525167
rect 182425 525111 182481 525167
rect 182481 525111 182485 525167
rect 182421 525107 182485 525111
rect 182501 525167 182565 525171
rect 182501 525111 182505 525167
rect 182505 525111 182561 525167
rect 182561 525111 182565 525167
rect 182501 525107 182565 525111
rect 186079 525167 186143 525171
rect 186079 525111 186083 525167
rect 186083 525111 186139 525167
rect 186139 525111 186143 525167
rect 186079 525107 186143 525111
rect 186159 525167 186223 525171
rect 186159 525111 186163 525167
rect 186163 525111 186219 525167
rect 186219 525111 186223 525167
rect 186159 525107 186223 525111
rect 186239 525167 186303 525171
rect 186239 525111 186243 525167
rect 186243 525111 186299 525167
rect 186299 525111 186303 525167
rect 186239 525107 186303 525111
rect 186319 525167 186383 525171
rect 186319 525111 186323 525167
rect 186323 525111 186379 525167
rect 186379 525111 186383 525167
rect 186319 525107 186383 525111
rect 173965 524623 174029 524627
rect 173965 524567 173969 524623
rect 173969 524567 174025 524623
rect 174025 524567 174029 524623
rect 173965 524563 174029 524567
rect 174045 524623 174109 524627
rect 174045 524567 174049 524623
rect 174049 524567 174105 524623
rect 174105 524567 174109 524623
rect 174045 524563 174109 524567
rect 174125 524623 174189 524627
rect 174125 524567 174129 524623
rect 174129 524567 174185 524623
rect 174185 524567 174189 524623
rect 174125 524563 174189 524567
rect 174205 524623 174269 524627
rect 174205 524567 174209 524623
rect 174209 524567 174265 524623
rect 174265 524567 174269 524623
rect 174205 524563 174269 524567
rect 177783 524623 177847 524627
rect 177783 524567 177787 524623
rect 177787 524567 177843 524623
rect 177843 524567 177847 524623
rect 177783 524563 177847 524567
rect 177863 524623 177927 524627
rect 177863 524567 177867 524623
rect 177867 524567 177923 524623
rect 177923 524567 177927 524623
rect 177863 524563 177927 524567
rect 177943 524623 178007 524627
rect 177943 524567 177947 524623
rect 177947 524567 178003 524623
rect 178003 524567 178007 524623
rect 177943 524563 178007 524567
rect 178023 524623 178087 524627
rect 178023 524567 178027 524623
rect 178027 524567 178083 524623
rect 178083 524567 178087 524623
rect 178023 524563 178087 524567
rect 181601 524623 181665 524627
rect 181601 524567 181605 524623
rect 181605 524567 181661 524623
rect 181661 524567 181665 524623
rect 181601 524563 181665 524567
rect 181681 524623 181745 524627
rect 181681 524567 181685 524623
rect 181685 524567 181741 524623
rect 181741 524567 181745 524623
rect 181681 524563 181745 524567
rect 181761 524623 181825 524627
rect 181761 524567 181765 524623
rect 181765 524567 181821 524623
rect 181821 524567 181825 524623
rect 181761 524563 181825 524567
rect 181841 524623 181905 524627
rect 181841 524567 181845 524623
rect 181845 524567 181901 524623
rect 181901 524567 181905 524623
rect 181841 524563 181905 524567
rect 185419 524623 185483 524627
rect 185419 524567 185423 524623
rect 185423 524567 185479 524623
rect 185479 524567 185483 524623
rect 185419 524563 185483 524567
rect 185499 524623 185563 524627
rect 185499 524567 185503 524623
rect 185503 524567 185559 524623
rect 185559 524567 185563 524623
rect 185499 524563 185563 524567
rect 185579 524623 185643 524627
rect 185579 524567 185583 524623
rect 185583 524567 185639 524623
rect 185639 524567 185643 524623
rect 185579 524563 185643 524567
rect 185659 524623 185723 524627
rect 185659 524567 185663 524623
rect 185663 524567 185719 524623
rect 185719 524567 185723 524623
rect 185659 524563 185723 524567
rect 174625 524079 174689 524083
rect 174625 524023 174629 524079
rect 174629 524023 174685 524079
rect 174685 524023 174689 524079
rect 174625 524019 174689 524023
rect 174705 524079 174769 524083
rect 174705 524023 174709 524079
rect 174709 524023 174765 524079
rect 174765 524023 174769 524079
rect 174705 524019 174769 524023
rect 174785 524079 174849 524083
rect 174785 524023 174789 524079
rect 174789 524023 174845 524079
rect 174845 524023 174849 524079
rect 174785 524019 174849 524023
rect 174865 524079 174929 524083
rect 174865 524023 174869 524079
rect 174869 524023 174925 524079
rect 174925 524023 174929 524079
rect 174865 524019 174929 524023
rect 178443 524079 178507 524083
rect 178443 524023 178447 524079
rect 178447 524023 178503 524079
rect 178503 524023 178507 524079
rect 178443 524019 178507 524023
rect 178523 524079 178587 524083
rect 178523 524023 178527 524079
rect 178527 524023 178583 524079
rect 178583 524023 178587 524079
rect 178523 524019 178587 524023
rect 178603 524079 178667 524083
rect 178603 524023 178607 524079
rect 178607 524023 178663 524079
rect 178663 524023 178667 524079
rect 178603 524019 178667 524023
rect 178683 524079 178747 524083
rect 178683 524023 178687 524079
rect 178687 524023 178743 524079
rect 178743 524023 178747 524079
rect 178683 524019 178747 524023
rect 182261 524079 182325 524083
rect 182261 524023 182265 524079
rect 182265 524023 182321 524079
rect 182321 524023 182325 524079
rect 182261 524019 182325 524023
rect 182341 524079 182405 524083
rect 182341 524023 182345 524079
rect 182345 524023 182401 524079
rect 182401 524023 182405 524079
rect 182341 524019 182405 524023
rect 182421 524079 182485 524083
rect 182421 524023 182425 524079
rect 182425 524023 182481 524079
rect 182481 524023 182485 524079
rect 182421 524019 182485 524023
rect 182501 524079 182565 524083
rect 182501 524023 182505 524079
rect 182505 524023 182561 524079
rect 182561 524023 182565 524079
rect 182501 524019 182565 524023
rect 186079 524079 186143 524083
rect 186079 524023 186083 524079
rect 186083 524023 186139 524079
rect 186139 524023 186143 524079
rect 186079 524019 186143 524023
rect 186159 524079 186223 524083
rect 186159 524023 186163 524079
rect 186163 524023 186219 524079
rect 186219 524023 186223 524079
rect 186159 524019 186223 524023
rect 186239 524079 186303 524083
rect 186239 524023 186243 524079
rect 186243 524023 186299 524079
rect 186299 524023 186303 524079
rect 186239 524019 186303 524023
rect 186319 524079 186383 524083
rect 186319 524023 186323 524079
rect 186323 524023 186379 524079
rect 186379 524023 186383 524079
rect 186319 524019 186383 524023
rect 173965 523535 174029 523539
rect 173965 523479 173969 523535
rect 173969 523479 174025 523535
rect 174025 523479 174029 523535
rect 173965 523475 174029 523479
rect 174045 523535 174109 523539
rect 174045 523479 174049 523535
rect 174049 523479 174105 523535
rect 174105 523479 174109 523535
rect 174045 523475 174109 523479
rect 174125 523535 174189 523539
rect 174125 523479 174129 523535
rect 174129 523479 174185 523535
rect 174185 523479 174189 523535
rect 174125 523475 174189 523479
rect 174205 523535 174269 523539
rect 174205 523479 174209 523535
rect 174209 523479 174265 523535
rect 174265 523479 174269 523535
rect 174205 523475 174269 523479
rect 177783 523535 177847 523539
rect 177783 523479 177787 523535
rect 177787 523479 177843 523535
rect 177843 523479 177847 523535
rect 177783 523475 177847 523479
rect 177863 523535 177927 523539
rect 177863 523479 177867 523535
rect 177867 523479 177923 523535
rect 177923 523479 177927 523535
rect 177863 523475 177927 523479
rect 177943 523535 178007 523539
rect 177943 523479 177947 523535
rect 177947 523479 178003 523535
rect 178003 523479 178007 523535
rect 177943 523475 178007 523479
rect 178023 523535 178087 523539
rect 178023 523479 178027 523535
rect 178027 523479 178083 523535
rect 178083 523479 178087 523535
rect 178023 523475 178087 523479
rect 181601 523535 181665 523539
rect 181601 523479 181605 523535
rect 181605 523479 181661 523535
rect 181661 523479 181665 523535
rect 181601 523475 181665 523479
rect 181681 523535 181745 523539
rect 181681 523479 181685 523535
rect 181685 523479 181741 523535
rect 181741 523479 181745 523535
rect 181681 523475 181745 523479
rect 181761 523535 181825 523539
rect 181761 523479 181765 523535
rect 181765 523479 181821 523535
rect 181821 523479 181825 523535
rect 181761 523475 181825 523479
rect 181841 523535 181905 523539
rect 181841 523479 181845 523535
rect 181845 523479 181901 523535
rect 181901 523479 181905 523535
rect 181841 523475 181905 523479
rect 185419 523535 185483 523539
rect 185419 523479 185423 523535
rect 185423 523479 185479 523535
rect 185479 523479 185483 523535
rect 185419 523475 185483 523479
rect 185499 523535 185563 523539
rect 185499 523479 185503 523535
rect 185503 523479 185559 523535
rect 185559 523479 185563 523535
rect 185499 523475 185563 523479
rect 185579 523535 185643 523539
rect 185579 523479 185583 523535
rect 185583 523479 185639 523535
rect 185639 523479 185643 523535
rect 185579 523475 185643 523479
rect 185659 523535 185723 523539
rect 185659 523479 185663 523535
rect 185663 523479 185719 523535
rect 185719 523479 185723 523535
rect 185659 523475 185723 523479
rect 174625 522991 174689 522995
rect 174625 522935 174629 522991
rect 174629 522935 174685 522991
rect 174685 522935 174689 522991
rect 174625 522931 174689 522935
rect 174705 522991 174769 522995
rect 174705 522935 174709 522991
rect 174709 522935 174765 522991
rect 174765 522935 174769 522991
rect 174705 522931 174769 522935
rect 174785 522991 174849 522995
rect 174785 522935 174789 522991
rect 174789 522935 174845 522991
rect 174845 522935 174849 522991
rect 174785 522931 174849 522935
rect 174865 522991 174929 522995
rect 174865 522935 174869 522991
rect 174869 522935 174925 522991
rect 174925 522935 174929 522991
rect 174865 522931 174929 522935
rect 178443 522991 178507 522995
rect 178443 522935 178447 522991
rect 178447 522935 178503 522991
rect 178503 522935 178507 522991
rect 178443 522931 178507 522935
rect 178523 522991 178587 522995
rect 178523 522935 178527 522991
rect 178527 522935 178583 522991
rect 178583 522935 178587 522991
rect 178523 522931 178587 522935
rect 178603 522991 178667 522995
rect 178603 522935 178607 522991
rect 178607 522935 178663 522991
rect 178663 522935 178667 522991
rect 178603 522931 178667 522935
rect 178683 522991 178747 522995
rect 178683 522935 178687 522991
rect 178687 522935 178743 522991
rect 178743 522935 178747 522991
rect 178683 522931 178747 522935
rect 182261 522991 182325 522995
rect 182261 522935 182265 522991
rect 182265 522935 182321 522991
rect 182321 522935 182325 522991
rect 182261 522931 182325 522935
rect 182341 522991 182405 522995
rect 182341 522935 182345 522991
rect 182345 522935 182401 522991
rect 182401 522935 182405 522991
rect 182341 522931 182405 522935
rect 182421 522991 182485 522995
rect 182421 522935 182425 522991
rect 182425 522935 182481 522991
rect 182481 522935 182485 522991
rect 182421 522931 182485 522935
rect 182501 522991 182565 522995
rect 182501 522935 182505 522991
rect 182505 522935 182561 522991
rect 182561 522935 182565 522991
rect 182501 522931 182565 522935
rect 186079 522991 186143 522995
rect 186079 522935 186083 522991
rect 186083 522935 186139 522991
rect 186139 522935 186143 522991
rect 186079 522931 186143 522935
rect 186159 522991 186223 522995
rect 186159 522935 186163 522991
rect 186163 522935 186219 522991
rect 186219 522935 186223 522991
rect 186159 522931 186223 522935
rect 186239 522991 186303 522995
rect 186239 522935 186243 522991
rect 186243 522935 186299 522991
rect 186299 522935 186303 522991
rect 186239 522931 186303 522935
rect 186319 522991 186383 522995
rect 186319 522935 186323 522991
rect 186323 522935 186379 522991
rect 186379 522935 186383 522991
rect 186319 522931 186383 522935
rect 173965 522447 174029 522451
rect 173965 522391 173969 522447
rect 173969 522391 174025 522447
rect 174025 522391 174029 522447
rect 173965 522387 174029 522391
rect 174045 522447 174109 522451
rect 174045 522391 174049 522447
rect 174049 522391 174105 522447
rect 174105 522391 174109 522447
rect 174045 522387 174109 522391
rect 174125 522447 174189 522451
rect 174125 522391 174129 522447
rect 174129 522391 174185 522447
rect 174185 522391 174189 522447
rect 174125 522387 174189 522391
rect 174205 522447 174269 522451
rect 174205 522391 174209 522447
rect 174209 522391 174265 522447
rect 174265 522391 174269 522447
rect 174205 522387 174269 522391
rect 177783 522447 177847 522451
rect 177783 522391 177787 522447
rect 177787 522391 177843 522447
rect 177843 522391 177847 522447
rect 177783 522387 177847 522391
rect 177863 522447 177927 522451
rect 177863 522391 177867 522447
rect 177867 522391 177923 522447
rect 177923 522391 177927 522447
rect 177863 522387 177927 522391
rect 177943 522447 178007 522451
rect 177943 522391 177947 522447
rect 177947 522391 178003 522447
rect 178003 522391 178007 522447
rect 177943 522387 178007 522391
rect 178023 522447 178087 522451
rect 178023 522391 178027 522447
rect 178027 522391 178083 522447
rect 178083 522391 178087 522447
rect 178023 522387 178087 522391
rect 181601 522447 181665 522451
rect 181601 522391 181605 522447
rect 181605 522391 181661 522447
rect 181661 522391 181665 522447
rect 181601 522387 181665 522391
rect 181681 522447 181745 522451
rect 181681 522391 181685 522447
rect 181685 522391 181741 522447
rect 181741 522391 181745 522447
rect 181681 522387 181745 522391
rect 181761 522447 181825 522451
rect 181761 522391 181765 522447
rect 181765 522391 181821 522447
rect 181821 522391 181825 522447
rect 181761 522387 181825 522391
rect 181841 522447 181905 522451
rect 181841 522391 181845 522447
rect 181845 522391 181901 522447
rect 181901 522391 181905 522447
rect 181841 522387 181905 522391
rect 185419 522447 185483 522451
rect 185419 522391 185423 522447
rect 185423 522391 185479 522447
rect 185479 522391 185483 522447
rect 185419 522387 185483 522391
rect 185499 522447 185563 522451
rect 185499 522391 185503 522447
rect 185503 522391 185559 522447
rect 185559 522391 185563 522447
rect 185499 522387 185563 522391
rect 185579 522447 185643 522451
rect 185579 522391 185583 522447
rect 185583 522391 185639 522447
rect 185639 522391 185643 522447
rect 185579 522387 185643 522391
rect 185659 522447 185723 522451
rect 185659 522391 185663 522447
rect 185663 522391 185719 522447
rect 185719 522391 185723 522447
rect 185659 522387 185723 522391
rect 174625 521903 174689 521907
rect 174625 521847 174629 521903
rect 174629 521847 174685 521903
rect 174685 521847 174689 521903
rect 174625 521843 174689 521847
rect 174705 521903 174769 521907
rect 174705 521847 174709 521903
rect 174709 521847 174765 521903
rect 174765 521847 174769 521903
rect 174705 521843 174769 521847
rect 174785 521903 174849 521907
rect 174785 521847 174789 521903
rect 174789 521847 174845 521903
rect 174845 521847 174849 521903
rect 174785 521843 174849 521847
rect 174865 521903 174929 521907
rect 174865 521847 174869 521903
rect 174869 521847 174925 521903
rect 174925 521847 174929 521903
rect 174865 521843 174929 521847
rect 178443 521903 178507 521907
rect 178443 521847 178447 521903
rect 178447 521847 178503 521903
rect 178503 521847 178507 521903
rect 178443 521843 178507 521847
rect 178523 521903 178587 521907
rect 178523 521847 178527 521903
rect 178527 521847 178583 521903
rect 178583 521847 178587 521903
rect 178523 521843 178587 521847
rect 178603 521903 178667 521907
rect 178603 521847 178607 521903
rect 178607 521847 178663 521903
rect 178663 521847 178667 521903
rect 178603 521843 178667 521847
rect 178683 521903 178747 521907
rect 178683 521847 178687 521903
rect 178687 521847 178743 521903
rect 178743 521847 178747 521903
rect 178683 521843 178747 521847
rect 182261 521903 182325 521907
rect 182261 521847 182265 521903
rect 182265 521847 182321 521903
rect 182321 521847 182325 521903
rect 182261 521843 182325 521847
rect 182341 521903 182405 521907
rect 182341 521847 182345 521903
rect 182345 521847 182401 521903
rect 182401 521847 182405 521903
rect 182341 521843 182405 521847
rect 182421 521903 182485 521907
rect 182421 521847 182425 521903
rect 182425 521847 182481 521903
rect 182481 521847 182485 521903
rect 182421 521843 182485 521847
rect 182501 521903 182565 521907
rect 182501 521847 182505 521903
rect 182505 521847 182561 521903
rect 182561 521847 182565 521903
rect 182501 521843 182565 521847
rect 186079 521903 186143 521907
rect 186079 521847 186083 521903
rect 186083 521847 186139 521903
rect 186139 521847 186143 521903
rect 186079 521843 186143 521847
rect 186159 521903 186223 521907
rect 186159 521847 186163 521903
rect 186163 521847 186219 521903
rect 186219 521847 186223 521903
rect 186159 521843 186223 521847
rect 186239 521903 186303 521907
rect 186239 521847 186243 521903
rect 186243 521847 186299 521903
rect 186299 521847 186303 521903
rect 186239 521843 186303 521847
rect 186319 521903 186383 521907
rect 186319 521847 186323 521903
rect 186323 521847 186379 521903
rect 186379 521847 186383 521903
rect 186319 521843 186383 521847
rect 173965 521359 174029 521363
rect 173965 521303 173969 521359
rect 173969 521303 174025 521359
rect 174025 521303 174029 521359
rect 173965 521299 174029 521303
rect 174045 521359 174109 521363
rect 174045 521303 174049 521359
rect 174049 521303 174105 521359
rect 174105 521303 174109 521359
rect 174045 521299 174109 521303
rect 174125 521359 174189 521363
rect 174125 521303 174129 521359
rect 174129 521303 174185 521359
rect 174185 521303 174189 521359
rect 174125 521299 174189 521303
rect 174205 521359 174269 521363
rect 174205 521303 174209 521359
rect 174209 521303 174265 521359
rect 174265 521303 174269 521359
rect 174205 521299 174269 521303
rect 177783 521359 177847 521363
rect 177783 521303 177787 521359
rect 177787 521303 177843 521359
rect 177843 521303 177847 521359
rect 177783 521299 177847 521303
rect 177863 521359 177927 521363
rect 177863 521303 177867 521359
rect 177867 521303 177923 521359
rect 177923 521303 177927 521359
rect 177863 521299 177927 521303
rect 177943 521359 178007 521363
rect 177943 521303 177947 521359
rect 177947 521303 178003 521359
rect 178003 521303 178007 521359
rect 177943 521299 178007 521303
rect 178023 521359 178087 521363
rect 178023 521303 178027 521359
rect 178027 521303 178083 521359
rect 178083 521303 178087 521359
rect 178023 521299 178087 521303
rect 181601 521359 181665 521363
rect 181601 521303 181605 521359
rect 181605 521303 181661 521359
rect 181661 521303 181665 521359
rect 181601 521299 181665 521303
rect 181681 521359 181745 521363
rect 181681 521303 181685 521359
rect 181685 521303 181741 521359
rect 181741 521303 181745 521359
rect 181681 521299 181745 521303
rect 181761 521359 181825 521363
rect 181761 521303 181765 521359
rect 181765 521303 181821 521359
rect 181821 521303 181825 521359
rect 181761 521299 181825 521303
rect 181841 521359 181905 521363
rect 181841 521303 181845 521359
rect 181845 521303 181901 521359
rect 181901 521303 181905 521359
rect 181841 521299 181905 521303
rect 185419 521359 185483 521363
rect 185419 521303 185423 521359
rect 185423 521303 185479 521359
rect 185479 521303 185483 521359
rect 185419 521299 185483 521303
rect 185499 521359 185563 521363
rect 185499 521303 185503 521359
rect 185503 521303 185559 521359
rect 185559 521303 185563 521359
rect 185499 521299 185563 521303
rect 185579 521359 185643 521363
rect 185579 521303 185583 521359
rect 185583 521303 185639 521359
rect 185639 521303 185643 521359
rect 185579 521299 185643 521303
rect 185659 521359 185723 521363
rect 185659 521303 185663 521359
rect 185663 521303 185719 521359
rect 185719 521303 185723 521359
rect 185659 521299 185723 521303
rect 174625 520815 174689 520819
rect 174625 520759 174629 520815
rect 174629 520759 174685 520815
rect 174685 520759 174689 520815
rect 174625 520755 174689 520759
rect 174705 520815 174769 520819
rect 174705 520759 174709 520815
rect 174709 520759 174765 520815
rect 174765 520759 174769 520815
rect 174705 520755 174769 520759
rect 174785 520815 174849 520819
rect 174785 520759 174789 520815
rect 174789 520759 174845 520815
rect 174845 520759 174849 520815
rect 174785 520755 174849 520759
rect 174865 520815 174929 520819
rect 174865 520759 174869 520815
rect 174869 520759 174925 520815
rect 174925 520759 174929 520815
rect 174865 520755 174929 520759
rect 178443 520815 178507 520819
rect 178443 520759 178447 520815
rect 178447 520759 178503 520815
rect 178503 520759 178507 520815
rect 178443 520755 178507 520759
rect 178523 520815 178587 520819
rect 178523 520759 178527 520815
rect 178527 520759 178583 520815
rect 178583 520759 178587 520815
rect 178523 520755 178587 520759
rect 178603 520815 178667 520819
rect 178603 520759 178607 520815
rect 178607 520759 178663 520815
rect 178663 520759 178667 520815
rect 178603 520755 178667 520759
rect 178683 520815 178747 520819
rect 178683 520759 178687 520815
rect 178687 520759 178743 520815
rect 178743 520759 178747 520815
rect 178683 520755 178747 520759
rect 182261 520815 182325 520819
rect 182261 520759 182265 520815
rect 182265 520759 182321 520815
rect 182321 520759 182325 520815
rect 182261 520755 182325 520759
rect 182341 520815 182405 520819
rect 182341 520759 182345 520815
rect 182345 520759 182401 520815
rect 182401 520759 182405 520815
rect 182341 520755 182405 520759
rect 182421 520815 182485 520819
rect 182421 520759 182425 520815
rect 182425 520759 182481 520815
rect 182481 520759 182485 520815
rect 182421 520755 182485 520759
rect 182501 520815 182565 520819
rect 182501 520759 182505 520815
rect 182505 520759 182561 520815
rect 182561 520759 182565 520815
rect 182501 520755 182565 520759
rect 186079 520815 186143 520819
rect 186079 520759 186083 520815
rect 186083 520759 186139 520815
rect 186139 520759 186143 520815
rect 186079 520755 186143 520759
rect 186159 520815 186223 520819
rect 186159 520759 186163 520815
rect 186163 520759 186219 520815
rect 186219 520759 186223 520815
rect 186159 520755 186223 520759
rect 186239 520815 186303 520819
rect 186239 520759 186243 520815
rect 186243 520759 186299 520815
rect 186299 520759 186303 520815
rect 186239 520755 186303 520759
rect 186319 520815 186383 520819
rect 186319 520759 186323 520815
rect 186323 520759 186379 520815
rect 186379 520759 186383 520815
rect 186319 520755 186383 520759
rect 173965 520271 174029 520275
rect 173965 520215 173969 520271
rect 173969 520215 174025 520271
rect 174025 520215 174029 520271
rect 173965 520211 174029 520215
rect 174045 520271 174109 520275
rect 174045 520215 174049 520271
rect 174049 520215 174105 520271
rect 174105 520215 174109 520271
rect 174045 520211 174109 520215
rect 174125 520271 174189 520275
rect 174125 520215 174129 520271
rect 174129 520215 174185 520271
rect 174185 520215 174189 520271
rect 174125 520211 174189 520215
rect 174205 520271 174269 520275
rect 174205 520215 174209 520271
rect 174209 520215 174265 520271
rect 174265 520215 174269 520271
rect 174205 520211 174269 520215
rect 177783 520271 177847 520275
rect 177783 520215 177787 520271
rect 177787 520215 177843 520271
rect 177843 520215 177847 520271
rect 177783 520211 177847 520215
rect 177863 520271 177927 520275
rect 177863 520215 177867 520271
rect 177867 520215 177923 520271
rect 177923 520215 177927 520271
rect 177863 520211 177927 520215
rect 177943 520271 178007 520275
rect 177943 520215 177947 520271
rect 177947 520215 178003 520271
rect 178003 520215 178007 520271
rect 177943 520211 178007 520215
rect 178023 520271 178087 520275
rect 178023 520215 178027 520271
rect 178027 520215 178083 520271
rect 178083 520215 178087 520271
rect 178023 520211 178087 520215
rect 181601 520271 181665 520275
rect 181601 520215 181605 520271
rect 181605 520215 181661 520271
rect 181661 520215 181665 520271
rect 181601 520211 181665 520215
rect 181681 520271 181745 520275
rect 181681 520215 181685 520271
rect 181685 520215 181741 520271
rect 181741 520215 181745 520271
rect 181681 520211 181745 520215
rect 181761 520271 181825 520275
rect 181761 520215 181765 520271
rect 181765 520215 181821 520271
rect 181821 520215 181825 520271
rect 181761 520211 181825 520215
rect 181841 520271 181905 520275
rect 181841 520215 181845 520271
rect 181845 520215 181901 520271
rect 181901 520215 181905 520271
rect 181841 520211 181905 520215
rect 185419 520271 185483 520275
rect 185419 520215 185423 520271
rect 185423 520215 185479 520271
rect 185479 520215 185483 520271
rect 185419 520211 185483 520215
rect 185499 520271 185563 520275
rect 185499 520215 185503 520271
rect 185503 520215 185559 520271
rect 185559 520215 185563 520271
rect 185499 520211 185563 520215
rect 185579 520271 185643 520275
rect 185579 520215 185583 520271
rect 185583 520215 185639 520271
rect 185639 520215 185643 520271
rect 185579 520211 185643 520215
rect 185659 520271 185723 520275
rect 185659 520215 185663 520271
rect 185663 520215 185719 520271
rect 185719 520215 185723 520271
rect 185659 520211 185723 520215
rect 174625 519727 174689 519731
rect 174625 519671 174629 519727
rect 174629 519671 174685 519727
rect 174685 519671 174689 519727
rect 174625 519667 174689 519671
rect 174705 519727 174769 519731
rect 174705 519671 174709 519727
rect 174709 519671 174765 519727
rect 174765 519671 174769 519727
rect 174705 519667 174769 519671
rect 174785 519727 174849 519731
rect 174785 519671 174789 519727
rect 174789 519671 174845 519727
rect 174845 519671 174849 519727
rect 174785 519667 174849 519671
rect 174865 519727 174929 519731
rect 174865 519671 174869 519727
rect 174869 519671 174925 519727
rect 174925 519671 174929 519727
rect 174865 519667 174929 519671
rect 178443 519727 178507 519731
rect 178443 519671 178447 519727
rect 178447 519671 178503 519727
rect 178503 519671 178507 519727
rect 178443 519667 178507 519671
rect 178523 519727 178587 519731
rect 178523 519671 178527 519727
rect 178527 519671 178583 519727
rect 178583 519671 178587 519727
rect 178523 519667 178587 519671
rect 178603 519727 178667 519731
rect 178603 519671 178607 519727
rect 178607 519671 178663 519727
rect 178663 519671 178667 519727
rect 178603 519667 178667 519671
rect 178683 519727 178747 519731
rect 178683 519671 178687 519727
rect 178687 519671 178743 519727
rect 178743 519671 178747 519727
rect 178683 519667 178747 519671
rect 182261 519727 182325 519731
rect 182261 519671 182265 519727
rect 182265 519671 182321 519727
rect 182321 519671 182325 519727
rect 182261 519667 182325 519671
rect 182341 519727 182405 519731
rect 182341 519671 182345 519727
rect 182345 519671 182401 519727
rect 182401 519671 182405 519727
rect 182341 519667 182405 519671
rect 182421 519727 182485 519731
rect 182421 519671 182425 519727
rect 182425 519671 182481 519727
rect 182481 519671 182485 519727
rect 182421 519667 182485 519671
rect 182501 519727 182565 519731
rect 182501 519671 182505 519727
rect 182505 519671 182561 519727
rect 182561 519671 182565 519727
rect 182501 519667 182565 519671
rect 186079 519727 186143 519731
rect 186079 519671 186083 519727
rect 186083 519671 186139 519727
rect 186139 519671 186143 519727
rect 186079 519667 186143 519671
rect 186159 519727 186223 519731
rect 186159 519671 186163 519727
rect 186163 519671 186219 519727
rect 186219 519671 186223 519727
rect 186159 519667 186223 519671
rect 186239 519727 186303 519731
rect 186239 519671 186243 519727
rect 186243 519671 186299 519727
rect 186299 519671 186303 519727
rect 186239 519667 186303 519671
rect 186319 519727 186383 519731
rect 186319 519671 186323 519727
rect 186323 519671 186379 519727
rect 186379 519671 186383 519727
rect 186319 519667 186383 519671
rect 173965 519183 174029 519187
rect 173965 519127 173969 519183
rect 173969 519127 174025 519183
rect 174025 519127 174029 519183
rect 173965 519123 174029 519127
rect 174045 519183 174109 519187
rect 174045 519127 174049 519183
rect 174049 519127 174105 519183
rect 174105 519127 174109 519183
rect 174045 519123 174109 519127
rect 174125 519183 174189 519187
rect 174125 519127 174129 519183
rect 174129 519127 174185 519183
rect 174185 519127 174189 519183
rect 174125 519123 174189 519127
rect 174205 519183 174269 519187
rect 174205 519127 174209 519183
rect 174209 519127 174265 519183
rect 174265 519127 174269 519183
rect 174205 519123 174269 519127
rect 177783 519183 177847 519187
rect 177783 519127 177787 519183
rect 177787 519127 177843 519183
rect 177843 519127 177847 519183
rect 177783 519123 177847 519127
rect 177863 519183 177927 519187
rect 177863 519127 177867 519183
rect 177867 519127 177923 519183
rect 177923 519127 177927 519183
rect 177863 519123 177927 519127
rect 177943 519183 178007 519187
rect 177943 519127 177947 519183
rect 177947 519127 178003 519183
rect 178003 519127 178007 519183
rect 177943 519123 178007 519127
rect 178023 519183 178087 519187
rect 178023 519127 178027 519183
rect 178027 519127 178083 519183
rect 178083 519127 178087 519183
rect 178023 519123 178087 519127
rect 181601 519183 181665 519187
rect 181601 519127 181605 519183
rect 181605 519127 181661 519183
rect 181661 519127 181665 519183
rect 181601 519123 181665 519127
rect 181681 519183 181745 519187
rect 181681 519127 181685 519183
rect 181685 519127 181741 519183
rect 181741 519127 181745 519183
rect 181681 519123 181745 519127
rect 181761 519183 181825 519187
rect 181761 519127 181765 519183
rect 181765 519127 181821 519183
rect 181821 519127 181825 519183
rect 181761 519123 181825 519127
rect 181841 519183 181905 519187
rect 181841 519127 181845 519183
rect 181845 519127 181901 519183
rect 181901 519127 181905 519183
rect 181841 519123 181905 519127
rect 185419 519183 185483 519187
rect 185419 519127 185423 519183
rect 185423 519127 185479 519183
rect 185479 519127 185483 519183
rect 185419 519123 185483 519127
rect 185499 519183 185563 519187
rect 185499 519127 185503 519183
rect 185503 519127 185559 519183
rect 185559 519127 185563 519183
rect 185499 519123 185563 519127
rect 185579 519183 185643 519187
rect 185579 519127 185583 519183
rect 185583 519127 185639 519183
rect 185639 519127 185643 519183
rect 185579 519123 185643 519127
rect 185659 519183 185723 519187
rect 185659 519127 185663 519183
rect 185663 519127 185719 519183
rect 185719 519127 185723 519183
rect 185659 519123 185723 519127
rect 174625 518639 174689 518643
rect 174625 518583 174629 518639
rect 174629 518583 174685 518639
rect 174685 518583 174689 518639
rect 174625 518579 174689 518583
rect 174705 518639 174769 518643
rect 174705 518583 174709 518639
rect 174709 518583 174765 518639
rect 174765 518583 174769 518639
rect 174705 518579 174769 518583
rect 174785 518639 174849 518643
rect 174785 518583 174789 518639
rect 174789 518583 174845 518639
rect 174845 518583 174849 518639
rect 174785 518579 174849 518583
rect 174865 518639 174929 518643
rect 174865 518583 174869 518639
rect 174869 518583 174925 518639
rect 174925 518583 174929 518639
rect 174865 518579 174929 518583
rect 178443 518639 178507 518643
rect 178443 518583 178447 518639
rect 178447 518583 178503 518639
rect 178503 518583 178507 518639
rect 178443 518579 178507 518583
rect 178523 518639 178587 518643
rect 178523 518583 178527 518639
rect 178527 518583 178583 518639
rect 178583 518583 178587 518639
rect 178523 518579 178587 518583
rect 178603 518639 178667 518643
rect 178603 518583 178607 518639
rect 178607 518583 178663 518639
rect 178663 518583 178667 518639
rect 178603 518579 178667 518583
rect 178683 518639 178747 518643
rect 178683 518583 178687 518639
rect 178687 518583 178743 518639
rect 178743 518583 178747 518639
rect 178683 518579 178747 518583
rect 182261 518639 182325 518643
rect 182261 518583 182265 518639
rect 182265 518583 182321 518639
rect 182321 518583 182325 518639
rect 182261 518579 182325 518583
rect 182341 518639 182405 518643
rect 182341 518583 182345 518639
rect 182345 518583 182401 518639
rect 182401 518583 182405 518639
rect 182341 518579 182405 518583
rect 182421 518639 182485 518643
rect 182421 518583 182425 518639
rect 182425 518583 182481 518639
rect 182481 518583 182485 518639
rect 182421 518579 182485 518583
rect 182501 518639 182565 518643
rect 182501 518583 182505 518639
rect 182505 518583 182561 518639
rect 182561 518583 182565 518639
rect 182501 518579 182565 518583
rect 186079 518639 186143 518643
rect 186079 518583 186083 518639
rect 186083 518583 186139 518639
rect 186139 518583 186143 518639
rect 186079 518579 186143 518583
rect 186159 518639 186223 518643
rect 186159 518583 186163 518639
rect 186163 518583 186219 518639
rect 186219 518583 186223 518639
rect 186159 518579 186223 518583
rect 186239 518639 186303 518643
rect 186239 518583 186243 518639
rect 186243 518583 186299 518639
rect 186299 518583 186303 518639
rect 186239 518579 186303 518583
rect 186319 518639 186383 518643
rect 186319 518583 186323 518639
rect 186323 518583 186379 518639
rect 186379 518583 186383 518639
rect 186319 518579 186383 518583
rect 173965 518095 174029 518099
rect 173965 518039 173969 518095
rect 173969 518039 174025 518095
rect 174025 518039 174029 518095
rect 173965 518035 174029 518039
rect 174045 518095 174109 518099
rect 174045 518039 174049 518095
rect 174049 518039 174105 518095
rect 174105 518039 174109 518095
rect 174045 518035 174109 518039
rect 174125 518095 174189 518099
rect 174125 518039 174129 518095
rect 174129 518039 174185 518095
rect 174185 518039 174189 518095
rect 174125 518035 174189 518039
rect 174205 518095 174269 518099
rect 174205 518039 174209 518095
rect 174209 518039 174265 518095
rect 174265 518039 174269 518095
rect 174205 518035 174269 518039
rect 177783 518095 177847 518099
rect 177783 518039 177787 518095
rect 177787 518039 177843 518095
rect 177843 518039 177847 518095
rect 177783 518035 177847 518039
rect 177863 518095 177927 518099
rect 177863 518039 177867 518095
rect 177867 518039 177923 518095
rect 177923 518039 177927 518095
rect 177863 518035 177927 518039
rect 177943 518095 178007 518099
rect 177943 518039 177947 518095
rect 177947 518039 178003 518095
rect 178003 518039 178007 518095
rect 177943 518035 178007 518039
rect 178023 518095 178087 518099
rect 178023 518039 178027 518095
rect 178027 518039 178083 518095
rect 178083 518039 178087 518095
rect 178023 518035 178087 518039
rect 181601 518095 181665 518099
rect 181601 518039 181605 518095
rect 181605 518039 181661 518095
rect 181661 518039 181665 518095
rect 181601 518035 181665 518039
rect 181681 518095 181745 518099
rect 181681 518039 181685 518095
rect 181685 518039 181741 518095
rect 181741 518039 181745 518095
rect 181681 518035 181745 518039
rect 181761 518095 181825 518099
rect 181761 518039 181765 518095
rect 181765 518039 181821 518095
rect 181821 518039 181825 518095
rect 181761 518035 181825 518039
rect 181841 518095 181905 518099
rect 181841 518039 181845 518095
rect 181845 518039 181901 518095
rect 181901 518039 181905 518095
rect 181841 518035 181905 518039
rect 185419 518095 185483 518099
rect 185419 518039 185423 518095
rect 185423 518039 185479 518095
rect 185479 518039 185483 518095
rect 185419 518035 185483 518039
rect 185499 518095 185563 518099
rect 185499 518039 185503 518095
rect 185503 518039 185559 518095
rect 185559 518039 185563 518095
rect 185499 518035 185563 518039
rect 185579 518095 185643 518099
rect 185579 518039 185583 518095
rect 185583 518039 185639 518095
rect 185639 518039 185643 518095
rect 185579 518035 185643 518039
rect 185659 518095 185723 518099
rect 185659 518039 185663 518095
rect 185663 518039 185719 518095
rect 185719 518039 185723 518095
rect 185659 518035 185723 518039
rect 174625 517551 174689 517555
rect 174625 517495 174629 517551
rect 174629 517495 174685 517551
rect 174685 517495 174689 517551
rect 174625 517491 174689 517495
rect 174705 517551 174769 517555
rect 174705 517495 174709 517551
rect 174709 517495 174765 517551
rect 174765 517495 174769 517551
rect 174705 517491 174769 517495
rect 174785 517551 174849 517555
rect 174785 517495 174789 517551
rect 174789 517495 174845 517551
rect 174845 517495 174849 517551
rect 174785 517491 174849 517495
rect 174865 517551 174929 517555
rect 174865 517495 174869 517551
rect 174869 517495 174925 517551
rect 174925 517495 174929 517551
rect 174865 517491 174929 517495
rect 178443 517551 178507 517555
rect 178443 517495 178447 517551
rect 178447 517495 178503 517551
rect 178503 517495 178507 517551
rect 178443 517491 178507 517495
rect 178523 517551 178587 517555
rect 178523 517495 178527 517551
rect 178527 517495 178583 517551
rect 178583 517495 178587 517551
rect 178523 517491 178587 517495
rect 178603 517551 178667 517555
rect 178603 517495 178607 517551
rect 178607 517495 178663 517551
rect 178663 517495 178667 517551
rect 178603 517491 178667 517495
rect 178683 517551 178747 517555
rect 178683 517495 178687 517551
rect 178687 517495 178743 517551
rect 178743 517495 178747 517551
rect 178683 517491 178747 517495
rect 182261 517551 182325 517555
rect 182261 517495 182265 517551
rect 182265 517495 182321 517551
rect 182321 517495 182325 517551
rect 182261 517491 182325 517495
rect 182341 517551 182405 517555
rect 182341 517495 182345 517551
rect 182345 517495 182401 517551
rect 182401 517495 182405 517551
rect 182341 517491 182405 517495
rect 182421 517551 182485 517555
rect 182421 517495 182425 517551
rect 182425 517495 182481 517551
rect 182481 517495 182485 517551
rect 182421 517491 182485 517495
rect 182501 517551 182565 517555
rect 182501 517495 182505 517551
rect 182505 517495 182561 517551
rect 182561 517495 182565 517551
rect 182501 517491 182565 517495
rect 186079 517551 186143 517555
rect 186079 517495 186083 517551
rect 186083 517495 186139 517551
rect 186139 517495 186143 517551
rect 186079 517491 186143 517495
rect 186159 517551 186223 517555
rect 186159 517495 186163 517551
rect 186163 517495 186219 517551
rect 186219 517495 186223 517551
rect 186159 517491 186223 517495
rect 186239 517551 186303 517555
rect 186239 517495 186243 517551
rect 186243 517495 186299 517551
rect 186299 517495 186303 517551
rect 186239 517491 186303 517495
rect 186319 517551 186383 517555
rect 186319 517495 186323 517551
rect 186323 517495 186379 517551
rect 186379 517495 186383 517551
rect 186319 517491 186383 517495
rect 173965 517007 174029 517011
rect 173965 516951 173969 517007
rect 173969 516951 174025 517007
rect 174025 516951 174029 517007
rect 173965 516947 174029 516951
rect 174045 517007 174109 517011
rect 174045 516951 174049 517007
rect 174049 516951 174105 517007
rect 174105 516951 174109 517007
rect 174045 516947 174109 516951
rect 174125 517007 174189 517011
rect 174125 516951 174129 517007
rect 174129 516951 174185 517007
rect 174185 516951 174189 517007
rect 174125 516947 174189 516951
rect 174205 517007 174269 517011
rect 174205 516951 174209 517007
rect 174209 516951 174265 517007
rect 174265 516951 174269 517007
rect 174205 516947 174269 516951
rect 177783 517007 177847 517011
rect 177783 516951 177787 517007
rect 177787 516951 177843 517007
rect 177843 516951 177847 517007
rect 177783 516947 177847 516951
rect 177863 517007 177927 517011
rect 177863 516951 177867 517007
rect 177867 516951 177923 517007
rect 177923 516951 177927 517007
rect 177863 516947 177927 516951
rect 177943 517007 178007 517011
rect 177943 516951 177947 517007
rect 177947 516951 178003 517007
rect 178003 516951 178007 517007
rect 177943 516947 178007 516951
rect 178023 517007 178087 517011
rect 178023 516951 178027 517007
rect 178027 516951 178083 517007
rect 178083 516951 178087 517007
rect 178023 516947 178087 516951
rect 181601 517007 181665 517011
rect 181601 516951 181605 517007
rect 181605 516951 181661 517007
rect 181661 516951 181665 517007
rect 181601 516947 181665 516951
rect 181681 517007 181745 517011
rect 181681 516951 181685 517007
rect 181685 516951 181741 517007
rect 181741 516951 181745 517007
rect 181681 516947 181745 516951
rect 181761 517007 181825 517011
rect 181761 516951 181765 517007
rect 181765 516951 181821 517007
rect 181821 516951 181825 517007
rect 181761 516947 181825 516951
rect 181841 517007 181905 517011
rect 181841 516951 181845 517007
rect 181845 516951 181901 517007
rect 181901 516951 181905 517007
rect 181841 516947 181905 516951
rect 185419 517007 185483 517011
rect 185419 516951 185423 517007
rect 185423 516951 185479 517007
rect 185479 516951 185483 517007
rect 185419 516947 185483 516951
rect 185499 517007 185563 517011
rect 185499 516951 185503 517007
rect 185503 516951 185559 517007
rect 185559 516951 185563 517007
rect 185499 516947 185563 516951
rect 185579 517007 185643 517011
rect 185579 516951 185583 517007
rect 185583 516951 185639 517007
rect 185639 516951 185643 517007
rect 185579 516947 185643 516951
rect 185659 517007 185723 517011
rect 185659 516951 185663 517007
rect 185663 516951 185719 517007
rect 185719 516951 185723 517007
rect 185659 516947 185723 516951
rect 174625 516463 174689 516467
rect 174625 516407 174629 516463
rect 174629 516407 174685 516463
rect 174685 516407 174689 516463
rect 174625 516403 174689 516407
rect 174705 516463 174769 516467
rect 174705 516407 174709 516463
rect 174709 516407 174765 516463
rect 174765 516407 174769 516463
rect 174705 516403 174769 516407
rect 174785 516463 174849 516467
rect 174785 516407 174789 516463
rect 174789 516407 174845 516463
rect 174845 516407 174849 516463
rect 174785 516403 174849 516407
rect 174865 516463 174929 516467
rect 174865 516407 174869 516463
rect 174869 516407 174925 516463
rect 174925 516407 174929 516463
rect 174865 516403 174929 516407
rect 178443 516463 178507 516467
rect 178443 516407 178447 516463
rect 178447 516407 178503 516463
rect 178503 516407 178507 516463
rect 178443 516403 178507 516407
rect 178523 516463 178587 516467
rect 178523 516407 178527 516463
rect 178527 516407 178583 516463
rect 178583 516407 178587 516463
rect 178523 516403 178587 516407
rect 178603 516463 178667 516467
rect 178603 516407 178607 516463
rect 178607 516407 178663 516463
rect 178663 516407 178667 516463
rect 178603 516403 178667 516407
rect 178683 516463 178747 516467
rect 178683 516407 178687 516463
rect 178687 516407 178743 516463
rect 178743 516407 178747 516463
rect 178683 516403 178747 516407
rect 182261 516463 182325 516467
rect 182261 516407 182265 516463
rect 182265 516407 182321 516463
rect 182321 516407 182325 516463
rect 182261 516403 182325 516407
rect 182341 516463 182405 516467
rect 182341 516407 182345 516463
rect 182345 516407 182401 516463
rect 182401 516407 182405 516463
rect 182341 516403 182405 516407
rect 182421 516463 182485 516467
rect 182421 516407 182425 516463
rect 182425 516407 182481 516463
rect 182481 516407 182485 516463
rect 182421 516403 182485 516407
rect 182501 516463 182565 516467
rect 182501 516407 182505 516463
rect 182505 516407 182561 516463
rect 182561 516407 182565 516463
rect 182501 516403 182565 516407
rect 186079 516463 186143 516467
rect 186079 516407 186083 516463
rect 186083 516407 186139 516463
rect 186139 516407 186143 516463
rect 186079 516403 186143 516407
rect 186159 516463 186223 516467
rect 186159 516407 186163 516463
rect 186163 516407 186219 516463
rect 186219 516407 186223 516463
rect 186159 516403 186223 516407
rect 186239 516463 186303 516467
rect 186239 516407 186243 516463
rect 186243 516407 186299 516463
rect 186299 516407 186303 516463
rect 186239 516403 186303 516407
rect 186319 516463 186383 516467
rect 186319 516407 186323 516463
rect 186323 516407 186379 516463
rect 186379 516407 186383 516463
rect 186319 516403 186383 516407
rect 173965 515919 174029 515923
rect 173965 515863 173969 515919
rect 173969 515863 174025 515919
rect 174025 515863 174029 515919
rect 173965 515859 174029 515863
rect 174045 515919 174109 515923
rect 174045 515863 174049 515919
rect 174049 515863 174105 515919
rect 174105 515863 174109 515919
rect 174045 515859 174109 515863
rect 174125 515919 174189 515923
rect 174125 515863 174129 515919
rect 174129 515863 174185 515919
rect 174185 515863 174189 515919
rect 174125 515859 174189 515863
rect 174205 515919 174269 515923
rect 174205 515863 174209 515919
rect 174209 515863 174265 515919
rect 174265 515863 174269 515919
rect 174205 515859 174269 515863
rect 177783 515919 177847 515923
rect 177783 515863 177787 515919
rect 177787 515863 177843 515919
rect 177843 515863 177847 515919
rect 177783 515859 177847 515863
rect 177863 515919 177927 515923
rect 177863 515863 177867 515919
rect 177867 515863 177923 515919
rect 177923 515863 177927 515919
rect 177863 515859 177927 515863
rect 177943 515919 178007 515923
rect 177943 515863 177947 515919
rect 177947 515863 178003 515919
rect 178003 515863 178007 515919
rect 177943 515859 178007 515863
rect 178023 515919 178087 515923
rect 178023 515863 178027 515919
rect 178027 515863 178083 515919
rect 178083 515863 178087 515919
rect 178023 515859 178087 515863
rect 181601 515919 181665 515923
rect 181601 515863 181605 515919
rect 181605 515863 181661 515919
rect 181661 515863 181665 515919
rect 181601 515859 181665 515863
rect 181681 515919 181745 515923
rect 181681 515863 181685 515919
rect 181685 515863 181741 515919
rect 181741 515863 181745 515919
rect 181681 515859 181745 515863
rect 181761 515919 181825 515923
rect 181761 515863 181765 515919
rect 181765 515863 181821 515919
rect 181821 515863 181825 515919
rect 181761 515859 181825 515863
rect 181841 515919 181905 515923
rect 181841 515863 181845 515919
rect 181845 515863 181901 515919
rect 181901 515863 181905 515919
rect 181841 515859 181905 515863
rect 185419 515919 185483 515923
rect 185419 515863 185423 515919
rect 185423 515863 185479 515919
rect 185479 515863 185483 515919
rect 185419 515859 185483 515863
rect 185499 515919 185563 515923
rect 185499 515863 185503 515919
rect 185503 515863 185559 515919
rect 185559 515863 185563 515919
rect 185499 515859 185563 515863
rect 185579 515919 185643 515923
rect 185579 515863 185583 515919
rect 185583 515863 185639 515919
rect 185639 515863 185643 515919
rect 185579 515859 185643 515863
rect 185659 515919 185723 515923
rect 185659 515863 185663 515919
rect 185663 515863 185719 515919
rect 185719 515863 185723 515919
rect 185659 515859 185723 515863
rect 174625 515375 174689 515379
rect 174625 515319 174629 515375
rect 174629 515319 174685 515375
rect 174685 515319 174689 515375
rect 174625 515315 174689 515319
rect 174705 515375 174769 515379
rect 174705 515319 174709 515375
rect 174709 515319 174765 515375
rect 174765 515319 174769 515375
rect 174705 515315 174769 515319
rect 174785 515375 174849 515379
rect 174785 515319 174789 515375
rect 174789 515319 174845 515375
rect 174845 515319 174849 515375
rect 174785 515315 174849 515319
rect 174865 515375 174929 515379
rect 174865 515319 174869 515375
rect 174869 515319 174925 515375
rect 174925 515319 174929 515375
rect 174865 515315 174929 515319
rect 178443 515375 178507 515379
rect 178443 515319 178447 515375
rect 178447 515319 178503 515375
rect 178503 515319 178507 515375
rect 178443 515315 178507 515319
rect 178523 515375 178587 515379
rect 178523 515319 178527 515375
rect 178527 515319 178583 515375
rect 178583 515319 178587 515375
rect 178523 515315 178587 515319
rect 178603 515375 178667 515379
rect 178603 515319 178607 515375
rect 178607 515319 178663 515375
rect 178663 515319 178667 515375
rect 178603 515315 178667 515319
rect 178683 515375 178747 515379
rect 178683 515319 178687 515375
rect 178687 515319 178743 515375
rect 178743 515319 178747 515375
rect 178683 515315 178747 515319
rect 182261 515375 182325 515379
rect 182261 515319 182265 515375
rect 182265 515319 182321 515375
rect 182321 515319 182325 515375
rect 182261 515315 182325 515319
rect 182341 515375 182405 515379
rect 182341 515319 182345 515375
rect 182345 515319 182401 515375
rect 182401 515319 182405 515375
rect 182341 515315 182405 515319
rect 182421 515375 182485 515379
rect 182421 515319 182425 515375
rect 182425 515319 182481 515375
rect 182481 515319 182485 515375
rect 182421 515315 182485 515319
rect 182501 515375 182565 515379
rect 182501 515319 182505 515375
rect 182505 515319 182561 515375
rect 182561 515319 182565 515375
rect 182501 515315 182565 515319
rect 186079 515375 186143 515379
rect 186079 515319 186083 515375
rect 186083 515319 186139 515375
rect 186139 515319 186143 515375
rect 186079 515315 186143 515319
rect 186159 515375 186223 515379
rect 186159 515319 186163 515375
rect 186163 515319 186219 515375
rect 186219 515319 186223 515375
rect 186159 515315 186223 515319
rect 186239 515375 186303 515379
rect 186239 515319 186243 515375
rect 186243 515319 186299 515375
rect 186299 515319 186303 515375
rect 186239 515315 186303 515319
rect 186319 515375 186383 515379
rect 186319 515319 186323 515375
rect 186323 515319 186379 515375
rect 186379 515319 186383 515375
rect 186319 515315 186383 515319
<< mimcap >>
rect 157709 541725 162509 541765
rect 157709 539005 157749 541725
rect 162469 539005 162509 541725
rect 157709 538965 162509 539005
<< mimcapcontact >>
rect 157749 539005 162469 541725
<< metal4 >>
rect 162608 541837 162704 541853
rect 157748 541725 162470 541726
rect 157748 539005 157749 541725
rect 162469 539005 162470 541725
rect 157748 539004 162470 539005
rect 159388 538655 159488 539004
rect 162608 538893 162624 541837
rect 162688 539080 162704 541837
rect 162688 538893 162763 539080
rect 162608 538877 162763 538893
rect 162628 538805 162763 538877
rect 159388 538555 159398 538655
rect 159478 538555 159488 538655
rect 159388 538545 159488 538555
rect 161378 538715 162763 538805
rect 161378 538665 161528 538715
rect 161378 538545 161388 538665
rect 161508 538545 161528 538665
rect 161378 538535 161528 538545
rect 173957 530067 174277 530627
rect 173957 530003 173965 530067
rect 174029 530003 174045 530067
rect 174109 530003 174125 530067
rect 174189 530003 174205 530067
rect 174269 530003 174277 530067
rect 173957 528979 174277 530003
rect 173957 528915 173965 528979
rect 174029 528915 174045 528979
rect 174109 528915 174125 528979
rect 174189 528915 174205 528979
rect 174269 528915 174277 528979
rect 173957 528793 174277 528915
rect 173957 528557 173999 528793
rect 174235 528557 174277 528793
rect 173957 527891 174277 528557
rect 173957 527827 173965 527891
rect 174029 527827 174045 527891
rect 174109 527827 174125 527891
rect 174189 527827 174205 527891
rect 174269 527827 174277 527891
rect 173957 526803 174277 527827
rect 173957 526739 173965 526803
rect 174029 526739 174045 526803
rect 174109 526739 174125 526803
rect 174189 526739 174205 526803
rect 174269 526739 174277 526803
rect 173957 525715 174277 526739
rect 173957 525651 173965 525715
rect 174029 525651 174045 525715
rect 174109 525651 174125 525715
rect 174189 525651 174205 525715
rect 174269 525651 174277 525715
rect 173957 524985 174277 525651
rect 173957 524749 173999 524985
rect 174235 524749 174277 524985
rect 173957 524627 174277 524749
rect 173957 524563 173965 524627
rect 174029 524563 174045 524627
rect 174109 524563 174125 524627
rect 174189 524563 174205 524627
rect 174269 524563 174277 524627
rect 173957 523539 174277 524563
rect 173957 523475 173965 523539
rect 174029 523475 174045 523539
rect 174109 523475 174125 523539
rect 174189 523475 174205 523539
rect 174269 523475 174277 523539
rect 173957 522451 174277 523475
rect 173957 522387 173965 522451
rect 174029 522387 174045 522451
rect 174109 522387 174125 522451
rect 174189 522387 174205 522451
rect 174269 522387 174277 522451
rect 173957 521363 174277 522387
rect 173957 521299 173965 521363
rect 174029 521299 174045 521363
rect 174109 521299 174125 521363
rect 174189 521299 174205 521363
rect 174269 521299 174277 521363
rect 173957 521177 174277 521299
rect 173957 520941 173999 521177
rect 174235 520941 174277 521177
rect 173957 520275 174277 520941
rect 173957 520211 173965 520275
rect 174029 520211 174045 520275
rect 174109 520211 174125 520275
rect 174189 520211 174205 520275
rect 174269 520211 174277 520275
rect 173957 519187 174277 520211
rect 173957 519123 173965 519187
rect 174029 519123 174045 519187
rect 174109 519123 174125 519187
rect 174189 519123 174205 519187
rect 174269 519123 174277 519187
rect 173957 518099 174277 519123
rect 173957 518035 173965 518099
rect 174029 518035 174045 518099
rect 174109 518035 174125 518099
rect 174189 518035 174205 518099
rect 174269 518035 174277 518099
rect 173957 517369 174277 518035
rect 173957 517133 173999 517369
rect 174235 517133 174277 517369
rect 173957 517011 174277 517133
rect 173957 516947 173965 517011
rect 174029 516947 174045 517011
rect 174109 516947 174125 517011
rect 174189 516947 174205 517011
rect 174269 516947 174277 517011
rect 173957 515923 174277 516947
rect 173957 515859 173965 515923
rect 174029 515859 174045 515923
rect 174109 515859 174125 515923
rect 174189 515859 174205 515923
rect 174269 515859 174277 515923
rect 173957 515299 174277 515859
rect 174617 530611 174937 530627
rect 174617 530547 174625 530611
rect 174689 530547 174705 530611
rect 174769 530547 174785 530611
rect 174849 530547 174865 530611
rect 174929 530547 174937 530611
rect 174617 529523 174937 530547
rect 174617 529459 174625 529523
rect 174689 529459 174705 529523
rect 174769 529459 174785 529523
rect 174849 529459 174865 529523
rect 174929 529459 174937 529523
rect 174617 528435 174937 529459
rect 174617 528371 174625 528435
rect 174689 528371 174705 528435
rect 174769 528371 174785 528435
rect 174849 528371 174865 528435
rect 174929 528371 174937 528435
rect 174617 528133 174937 528371
rect 174617 527897 174659 528133
rect 174895 527897 174937 528133
rect 174617 527347 174937 527897
rect 174617 527283 174625 527347
rect 174689 527283 174705 527347
rect 174769 527283 174785 527347
rect 174849 527283 174865 527347
rect 174929 527283 174937 527347
rect 174617 526259 174937 527283
rect 174617 526195 174625 526259
rect 174689 526195 174705 526259
rect 174769 526195 174785 526259
rect 174849 526195 174865 526259
rect 174929 526195 174937 526259
rect 174617 525171 174937 526195
rect 174617 525107 174625 525171
rect 174689 525107 174705 525171
rect 174769 525107 174785 525171
rect 174849 525107 174865 525171
rect 174929 525107 174937 525171
rect 174617 524325 174937 525107
rect 174617 524089 174659 524325
rect 174895 524089 174937 524325
rect 174617 524083 174937 524089
rect 174617 524019 174625 524083
rect 174689 524019 174705 524083
rect 174769 524019 174785 524083
rect 174849 524019 174865 524083
rect 174929 524019 174937 524083
rect 174617 522995 174937 524019
rect 174617 522931 174625 522995
rect 174689 522931 174705 522995
rect 174769 522931 174785 522995
rect 174849 522931 174865 522995
rect 174929 522931 174937 522995
rect 174617 521907 174937 522931
rect 174617 521843 174625 521907
rect 174689 521843 174705 521907
rect 174769 521843 174785 521907
rect 174849 521843 174865 521907
rect 174929 521843 174937 521907
rect 174617 520819 174937 521843
rect 174617 520755 174625 520819
rect 174689 520755 174705 520819
rect 174769 520755 174785 520819
rect 174849 520755 174865 520819
rect 174929 520755 174937 520819
rect 174617 520517 174937 520755
rect 174617 520281 174659 520517
rect 174895 520281 174937 520517
rect 174617 519731 174937 520281
rect 174617 519667 174625 519731
rect 174689 519667 174705 519731
rect 174769 519667 174785 519731
rect 174849 519667 174865 519731
rect 174929 519667 174937 519731
rect 174617 518643 174937 519667
rect 174617 518579 174625 518643
rect 174689 518579 174705 518643
rect 174769 518579 174785 518643
rect 174849 518579 174865 518643
rect 174929 518579 174937 518643
rect 174617 517555 174937 518579
rect 174617 517491 174625 517555
rect 174689 517491 174705 517555
rect 174769 517491 174785 517555
rect 174849 517491 174865 517555
rect 174929 517491 174937 517555
rect 174617 516709 174937 517491
rect 174617 516473 174659 516709
rect 174895 516473 174937 516709
rect 174617 516467 174937 516473
rect 174617 516403 174625 516467
rect 174689 516403 174705 516467
rect 174769 516403 174785 516467
rect 174849 516403 174865 516467
rect 174929 516403 174937 516467
rect 174617 515379 174937 516403
rect 174617 515315 174625 515379
rect 174689 515315 174705 515379
rect 174769 515315 174785 515379
rect 174849 515315 174865 515379
rect 174929 515315 174937 515379
rect 174617 515299 174937 515315
rect 177775 530067 178095 530627
rect 177775 530003 177783 530067
rect 177847 530003 177863 530067
rect 177927 530003 177943 530067
rect 178007 530003 178023 530067
rect 178087 530003 178095 530067
rect 177775 528979 178095 530003
rect 177775 528915 177783 528979
rect 177847 528915 177863 528979
rect 177927 528915 177943 528979
rect 178007 528915 178023 528979
rect 178087 528915 178095 528979
rect 177775 528793 178095 528915
rect 177775 528557 177817 528793
rect 178053 528557 178095 528793
rect 177775 527891 178095 528557
rect 177775 527827 177783 527891
rect 177847 527827 177863 527891
rect 177927 527827 177943 527891
rect 178007 527827 178023 527891
rect 178087 527827 178095 527891
rect 177775 526803 178095 527827
rect 177775 526739 177783 526803
rect 177847 526739 177863 526803
rect 177927 526739 177943 526803
rect 178007 526739 178023 526803
rect 178087 526739 178095 526803
rect 177775 525715 178095 526739
rect 177775 525651 177783 525715
rect 177847 525651 177863 525715
rect 177927 525651 177943 525715
rect 178007 525651 178023 525715
rect 178087 525651 178095 525715
rect 177775 524985 178095 525651
rect 177775 524749 177817 524985
rect 178053 524749 178095 524985
rect 177775 524627 178095 524749
rect 177775 524563 177783 524627
rect 177847 524563 177863 524627
rect 177927 524563 177943 524627
rect 178007 524563 178023 524627
rect 178087 524563 178095 524627
rect 177775 523539 178095 524563
rect 177775 523475 177783 523539
rect 177847 523475 177863 523539
rect 177927 523475 177943 523539
rect 178007 523475 178023 523539
rect 178087 523475 178095 523539
rect 177775 522451 178095 523475
rect 177775 522387 177783 522451
rect 177847 522387 177863 522451
rect 177927 522387 177943 522451
rect 178007 522387 178023 522451
rect 178087 522387 178095 522451
rect 177775 521363 178095 522387
rect 177775 521299 177783 521363
rect 177847 521299 177863 521363
rect 177927 521299 177943 521363
rect 178007 521299 178023 521363
rect 178087 521299 178095 521363
rect 177775 521177 178095 521299
rect 177775 520941 177817 521177
rect 178053 520941 178095 521177
rect 177775 520275 178095 520941
rect 177775 520211 177783 520275
rect 177847 520211 177863 520275
rect 177927 520211 177943 520275
rect 178007 520211 178023 520275
rect 178087 520211 178095 520275
rect 177775 519187 178095 520211
rect 177775 519123 177783 519187
rect 177847 519123 177863 519187
rect 177927 519123 177943 519187
rect 178007 519123 178023 519187
rect 178087 519123 178095 519187
rect 177775 518099 178095 519123
rect 177775 518035 177783 518099
rect 177847 518035 177863 518099
rect 177927 518035 177943 518099
rect 178007 518035 178023 518099
rect 178087 518035 178095 518099
rect 177775 517369 178095 518035
rect 177775 517133 177817 517369
rect 178053 517133 178095 517369
rect 177775 517011 178095 517133
rect 177775 516947 177783 517011
rect 177847 516947 177863 517011
rect 177927 516947 177943 517011
rect 178007 516947 178023 517011
rect 178087 516947 178095 517011
rect 177775 515923 178095 516947
rect 177775 515859 177783 515923
rect 177847 515859 177863 515923
rect 177927 515859 177943 515923
rect 178007 515859 178023 515923
rect 178087 515859 178095 515923
rect 177775 515299 178095 515859
rect 178435 530611 178755 530627
rect 178435 530547 178443 530611
rect 178507 530547 178523 530611
rect 178587 530547 178603 530611
rect 178667 530547 178683 530611
rect 178747 530547 178755 530611
rect 178435 529523 178755 530547
rect 178435 529459 178443 529523
rect 178507 529459 178523 529523
rect 178587 529459 178603 529523
rect 178667 529459 178683 529523
rect 178747 529459 178755 529523
rect 178435 528435 178755 529459
rect 178435 528371 178443 528435
rect 178507 528371 178523 528435
rect 178587 528371 178603 528435
rect 178667 528371 178683 528435
rect 178747 528371 178755 528435
rect 178435 528133 178755 528371
rect 178435 527897 178477 528133
rect 178713 527897 178755 528133
rect 178435 527347 178755 527897
rect 178435 527283 178443 527347
rect 178507 527283 178523 527347
rect 178587 527283 178603 527347
rect 178667 527283 178683 527347
rect 178747 527283 178755 527347
rect 178435 526259 178755 527283
rect 178435 526195 178443 526259
rect 178507 526195 178523 526259
rect 178587 526195 178603 526259
rect 178667 526195 178683 526259
rect 178747 526195 178755 526259
rect 178435 525171 178755 526195
rect 178435 525107 178443 525171
rect 178507 525107 178523 525171
rect 178587 525107 178603 525171
rect 178667 525107 178683 525171
rect 178747 525107 178755 525171
rect 178435 524325 178755 525107
rect 178435 524089 178477 524325
rect 178713 524089 178755 524325
rect 178435 524083 178755 524089
rect 178435 524019 178443 524083
rect 178507 524019 178523 524083
rect 178587 524019 178603 524083
rect 178667 524019 178683 524083
rect 178747 524019 178755 524083
rect 178435 522995 178755 524019
rect 178435 522931 178443 522995
rect 178507 522931 178523 522995
rect 178587 522931 178603 522995
rect 178667 522931 178683 522995
rect 178747 522931 178755 522995
rect 178435 521907 178755 522931
rect 178435 521843 178443 521907
rect 178507 521843 178523 521907
rect 178587 521843 178603 521907
rect 178667 521843 178683 521907
rect 178747 521843 178755 521907
rect 178435 520819 178755 521843
rect 178435 520755 178443 520819
rect 178507 520755 178523 520819
rect 178587 520755 178603 520819
rect 178667 520755 178683 520819
rect 178747 520755 178755 520819
rect 178435 520517 178755 520755
rect 178435 520281 178477 520517
rect 178713 520281 178755 520517
rect 178435 519731 178755 520281
rect 178435 519667 178443 519731
rect 178507 519667 178523 519731
rect 178587 519667 178603 519731
rect 178667 519667 178683 519731
rect 178747 519667 178755 519731
rect 178435 518643 178755 519667
rect 178435 518579 178443 518643
rect 178507 518579 178523 518643
rect 178587 518579 178603 518643
rect 178667 518579 178683 518643
rect 178747 518579 178755 518643
rect 178435 517555 178755 518579
rect 178435 517491 178443 517555
rect 178507 517491 178523 517555
rect 178587 517491 178603 517555
rect 178667 517491 178683 517555
rect 178747 517491 178755 517555
rect 178435 516709 178755 517491
rect 178435 516473 178477 516709
rect 178713 516473 178755 516709
rect 178435 516467 178755 516473
rect 178435 516403 178443 516467
rect 178507 516403 178523 516467
rect 178587 516403 178603 516467
rect 178667 516403 178683 516467
rect 178747 516403 178755 516467
rect 178435 515379 178755 516403
rect 178435 515315 178443 515379
rect 178507 515315 178523 515379
rect 178587 515315 178603 515379
rect 178667 515315 178683 515379
rect 178747 515315 178755 515379
rect 178435 515299 178755 515315
rect 181593 530067 181913 530627
rect 181593 530003 181601 530067
rect 181665 530003 181681 530067
rect 181745 530003 181761 530067
rect 181825 530003 181841 530067
rect 181905 530003 181913 530067
rect 181593 528979 181913 530003
rect 181593 528915 181601 528979
rect 181665 528915 181681 528979
rect 181745 528915 181761 528979
rect 181825 528915 181841 528979
rect 181905 528915 181913 528979
rect 181593 528793 181913 528915
rect 181593 528557 181635 528793
rect 181871 528557 181913 528793
rect 181593 527891 181913 528557
rect 181593 527827 181601 527891
rect 181665 527827 181681 527891
rect 181745 527827 181761 527891
rect 181825 527827 181841 527891
rect 181905 527827 181913 527891
rect 181593 526803 181913 527827
rect 181593 526739 181601 526803
rect 181665 526739 181681 526803
rect 181745 526739 181761 526803
rect 181825 526739 181841 526803
rect 181905 526739 181913 526803
rect 181593 525715 181913 526739
rect 181593 525651 181601 525715
rect 181665 525651 181681 525715
rect 181745 525651 181761 525715
rect 181825 525651 181841 525715
rect 181905 525651 181913 525715
rect 181593 524985 181913 525651
rect 181593 524749 181635 524985
rect 181871 524749 181913 524985
rect 181593 524627 181913 524749
rect 181593 524563 181601 524627
rect 181665 524563 181681 524627
rect 181745 524563 181761 524627
rect 181825 524563 181841 524627
rect 181905 524563 181913 524627
rect 181593 523539 181913 524563
rect 181593 523475 181601 523539
rect 181665 523475 181681 523539
rect 181745 523475 181761 523539
rect 181825 523475 181841 523539
rect 181905 523475 181913 523539
rect 181593 522451 181913 523475
rect 181593 522387 181601 522451
rect 181665 522387 181681 522451
rect 181745 522387 181761 522451
rect 181825 522387 181841 522451
rect 181905 522387 181913 522451
rect 181593 521363 181913 522387
rect 181593 521299 181601 521363
rect 181665 521299 181681 521363
rect 181745 521299 181761 521363
rect 181825 521299 181841 521363
rect 181905 521299 181913 521363
rect 181593 521177 181913 521299
rect 181593 520941 181635 521177
rect 181871 520941 181913 521177
rect 181593 520275 181913 520941
rect 181593 520211 181601 520275
rect 181665 520211 181681 520275
rect 181745 520211 181761 520275
rect 181825 520211 181841 520275
rect 181905 520211 181913 520275
rect 181593 519187 181913 520211
rect 181593 519123 181601 519187
rect 181665 519123 181681 519187
rect 181745 519123 181761 519187
rect 181825 519123 181841 519187
rect 181905 519123 181913 519187
rect 181593 518099 181913 519123
rect 181593 518035 181601 518099
rect 181665 518035 181681 518099
rect 181745 518035 181761 518099
rect 181825 518035 181841 518099
rect 181905 518035 181913 518099
rect 181593 517369 181913 518035
rect 181593 517133 181635 517369
rect 181871 517133 181913 517369
rect 181593 517011 181913 517133
rect 181593 516947 181601 517011
rect 181665 516947 181681 517011
rect 181745 516947 181761 517011
rect 181825 516947 181841 517011
rect 181905 516947 181913 517011
rect 181593 515923 181913 516947
rect 181593 515859 181601 515923
rect 181665 515859 181681 515923
rect 181745 515859 181761 515923
rect 181825 515859 181841 515923
rect 181905 515859 181913 515923
rect 181593 515299 181913 515859
rect 182253 530611 182573 530627
rect 182253 530547 182261 530611
rect 182325 530547 182341 530611
rect 182405 530547 182421 530611
rect 182485 530547 182501 530611
rect 182565 530547 182573 530611
rect 182253 529523 182573 530547
rect 182253 529459 182261 529523
rect 182325 529459 182341 529523
rect 182405 529459 182421 529523
rect 182485 529459 182501 529523
rect 182565 529459 182573 529523
rect 182253 528435 182573 529459
rect 182253 528371 182261 528435
rect 182325 528371 182341 528435
rect 182405 528371 182421 528435
rect 182485 528371 182501 528435
rect 182565 528371 182573 528435
rect 182253 528133 182573 528371
rect 182253 527897 182295 528133
rect 182531 527897 182573 528133
rect 182253 527347 182573 527897
rect 182253 527283 182261 527347
rect 182325 527283 182341 527347
rect 182405 527283 182421 527347
rect 182485 527283 182501 527347
rect 182565 527283 182573 527347
rect 182253 526259 182573 527283
rect 182253 526195 182261 526259
rect 182325 526195 182341 526259
rect 182405 526195 182421 526259
rect 182485 526195 182501 526259
rect 182565 526195 182573 526259
rect 182253 525171 182573 526195
rect 182253 525107 182261 525171
rect 182325 525107 182341 525171
rect 182405 525107 182421 525171
rect 182485 525107 182501 525171
rect 182565 525107 182573 525171
rect 182253 524325 182573 525107
rect 182253 524089 182295 524325
rect 182531 524089 182573 524325
rect 182253 524083 182573 524089
rect 182253 524019 182261 524083
rect 182325 524019 182341 524083
rect 182405 524019 182421 524083
rect 182485 524019 182501 524083
rect 182565 524019 182573 524083
rect 182253 522995 182573 524019
rect 182253 522931 182261 522995
rect 182325 522931 182341 522995
rect 182405 522931 182421 522995
rect 182485 522931 182501 522995
rect 182565 522931 182573 522995
rect 182253 521907 182573 522931
rect 182253 521843 182261 521907
rect 182325 521843 182341 521907
rect 182405 521843 182421 521907
rect 182485 521843 182501 521907
rect 182565 521843 182573 521907
rect 182253 520819 182573 521843
rect 182253 520755 182261 520819
rect 182325 520755 182341 520819
rect 182405 520755 182421 520819
rect 182485 520755 182501 520819
rect 182565 520755 182573 520819
rect 182253 520517 182573 520755
rect 182253 520281 182295 520517
rect 182531 520281 182573 520517
rect 182253 519731 182573 520281
rect 182253 519667 182261 519731
rect 182325 519667 182341 519731
rect 182405 519667 182421 519731
rect 182485 519667 182501 519731
rect 182565 519667 182573 519731
rect 182253 518643 182573 519667
rect 182253 518579 182261 518643
rect 182325 518579 182341 518643
rect 182405 518579 182421 518643
rect 182485 518579 182501 518643
rect 182565 518579 182573 518643
rect 182253 517555 182573 518579
rect 182253 517491 182261 517555
rect 182325 517491 182341 517555
rect 182405 517491 182421 517555
rect 182485 517491 182501 517555
rect 182565 517491 182573 517555
rect 182253 516709 182573 517491
rect 182253 516473 182295 516709
rect 182531 516473 182573 516709
rect 182253 516467 182573 516473
rect 182253 516403 182261 516467
rect 182325 516403 182341 516467
rect 182405 516403 182421 516467
rect 182485 516403 182501 516467
rect 182565 516403 182573 516467
rect 182253 515379 182573 516403
rect 182253 515315 182261 515379
rect 182325 515315 182341 515379
rect 182405 515315 182421 515379
rect 182485 515315 182501 515379
rect 182565 515315 182573 515379
rect 182253 515299 182573 515315
rect 185411 530067 185731 530627
rect 185411 530003 185419 530067
rect 185483 530003 185499 530067
rect 185563 530003 185579 530067
rect 185643 530003 185659 530067
rect 185723 530003 185731 530067
rect 185411 528979 185731 530003
rect 185411 528915 185419 528979
rect 185483 528915 185499 528979
rect 185563 528915 185579 528979
rect 185643 528915 185659 528979
rect 185723 528915 185731 528979
rect 185411 528793 185731 528915
rect 185411 528557 185453 528793
rect 185689 528557 185731 528793
rect 185411 527891 185731 528557
rect 185411 527827 185419 527891
rect 185483 527827 185499 527891
rect 185563 527827 185579 527891
rect 185643 527827 185659 527891
rect 185723 527827 185731 527891
rect 185411 526803 185731 527827
rect 185411 526739 185419 526803
rect 185483 526739 185499 526803
rect 185563 526739 185579 526803
rect 185643 526739 185659 526803
rect 185723 526739 185731 526803
rect 185411 525715 185731 526739
rect 185411 525651 185419 525715
rect 185483 525651 185499 525715
rect 185563 525651 185579 525715
rect 185643 525651 185659 525715
rect 185723 525651 185731 525715
rect 185411 524985 185731 525651
rect 185411 524749 185453 524985
rect 185689 524749 185731 524985
rect 185411 524627 185731 524749
rect 185411 524563 185419 524627
rect 185483 524563 185499 524627
rect 185563 524563 185579 524627
rect 185643 524563 185659 524627
rect 185723 524563 185731 524627
rect 185411 523539 185731 524563
rect 185411 523475 185419 523539
rect 185483 523475 185499 523539
rect 185563 523475 185579 523539
rect 185643 523475 185659 523539
rect 185723 523475 185731 523539
rect 185411 522451 185731 523475
rect 185411 522387 185419 522451
rect 185483 522387 185499 522451
rect 185563 522387 185579 522451
rect 185643 522387 185659 522451
rect 185723 522387 185731 522451
rect 185411 521363 185731 522387
rect 185411 521299 185419 521363
rect 185483 521299 185499 521363
rect 185563 521299 185579 521363
rect 185643 521299 185659 521363
rect 185723 521299 185731 521363
rect 185411 521177 185731 521299
rect 185411 520941 185453 521177
rect 185689 520941 185731 521177
rect 185411 520275 185731 520941
rect 185411 520211 185419 520275
rect 185483 520211 185499 520275
rect 185563 520211 185579 520275
rect 185643 520211 185659 520275
rect 185723 520211 185731 520275
rect 185411 519187 185731 520211
rect 185411 519123 185419 519187
rect 185483 519123 185499 519187
rect 185563 519123 185579 519187
rect 185643 519123 185659 519187
rect 185723 519123 185731 519187
rect 185411 518099 185731 519123
rect 185411 518035 185419 518099
rect 185483 518035 185499 518099
rect 185563 518035 185579 518099
rect 185643 518035 185659 518099
rect 185723 518035 185731 518099
rect 185411 517369 185731 518035
rect 185411 517133 185453 517369
rect 185689 517133 185731 517369
rect 185411 517011 185731 517133
rect 185411 516947 185419 517011
rect 185483 516947 185499 517011
rect 185563 516947 185579 517011
rect 185643 516947 185659 517011
rect 185723 516947 185731 517011
rect 185411 515923 185731 516947
rect 185411 515859 185419 515923
rect 185483 515859 185499 515923
rect 185563 515859 185579 515923
rect 185643 515859 185659 515923
rect 185723 515859 185731 515923
rect 185411 515299 185731 515859
rect 186071 530611 186391 530627
rect 186071 530547 186079 530611
rect 186143 530547 186159 530611
rect 186223 530547 186239 530611
rect 186303 530547 186319 530611
rect 186383 530547 186391 530611
rect 186071 529523 186391 530547
rect 186071 529459 186079 529523
rect 186143 529459 186159 529523
rect 186223 529459 186239 529523
rect 186303 529459 186319 529523
rect 186383 529459 186391 529523
rect 186071 528435 186391 529459
rect 186071 528371 186079 528435
rect 186143 528371 186159 528435
rect 186223 528371 186239 528435
rect 186303 528371 186319 528435
rect 186383 528371 186391 528435
rect 186071 528133 186391 528371
rect 186071 527897 186113 528133
rect 186349 527897 186391 528133
rect 186071 527347 186391 527897
rect 186071 527283 186079 527347
rect 186143 527283 186159 527347
rect 186223 527283 186239 527347
rect 186303 527283 186319 527347
rect 186383 527283 186391 527347
rect 186071 526259 186391 527283
rect 186071 526195 186079 526259
rect 186143 526195 186159 526259
rect 186223 526195 186239 526259
rect 186303 526195 186319 526259
rect 186383 526195 186391 526259
rect 186071 525171 186391 526195
rect 186071 525107 186079 525171
rect 186143 525107 186159 525171
rect 186223 525107 186239 525171
rect 186303 525107 186319 525171
rect 186383 525107 186391 525171
rect 186071 524325 186391 525107
rect 186071 524089 186113 524325
rect 186349 524089 186391 524325
rect 186071 524083 186391 524089
rect 186071 524019 186079 524083
rect 186143 524019 186159 524083
rect 186223 524019 186239 524083
rect 186303 524019 186319 524083
rect 186383 524019 186391 524083
rect 186071 522995 186391 524019
rect 186071 522931 186079 522995
rect 186143 522931 186159 522995
rect 186223 522931 186239 522995
rect 186303 522931 186319 522995
rect 186383 522931 186391 522995
rect 186071 521907 186391 522931
rect 186071 521843 186079 521907
rect 186143 521843 186159 521907
rect 186223 521843 186239 521907
rect 186303 521843 186319 521907
rect 186383 521843 186391 521907
rect 186071 520819 186391 521843
rect 186071 520755 186079 520819
rect 186143 520755 186159 520819
rect 186223 520755 186239 520819
rect 186303 520755 186319 520819
rect 186383 520755 186391 520819
rect 186071 520517 186391 520755
rect 186071 520281 186113 520517
rect 186349 520281 186391 520517
rect 186071 519731 186391 520281
rect 186071 519667 186079 519731
rect 186143 519667 186159 519731
rect 186223 519667 186239 519731
rect 186303 519667 186319 519731
rect 186383 519667 186391 519731
rect 186071 518643 186391 519667
rect 186071 518579 186079 518643
rect 186143 518579 186159 518643
rect 186223 518579 186239 518643
rect 186303 518579 186319 518643
rect 186383 518579 186391 518643
rect 186071 517555 186391 518579
rect 186071 517491 186079 517555
rect 186143 517491 186159 517555
rect 186223 517491 186239 517555
rect 186303 517491 186319 517555
rect 186383 517491 186391 517555
rect 186071 516709 186391 517491
rect 186071 516473 186113 516709
rect 186349 516473 186391 516709
rect 186071 516467 186391 516473
rect 186071 516403 186079 516467
rect 186143 516403 186159 516467
rect 186223 516403 186239 516467
rect 186303 516403 186319 516467
rect 186383 516403 186391 516467
rect 186071 515379 186391 516403
rect 186071 515315 186079 515379
rect 186143 515315 186159 515379
rect 186223 515315 186239 515379
rect 186303 515315 186319 515379
rect 186383 515315 186391 515379
rect 186071 515299 186391 515315
<< via4 >>
rect 173999 528557 174235 528793
rect 173999 524749 174235 524985
rect 173999 520941 174235 521177
rect 173999 517133 174235 517369
rect 174659 527897 174895 528133
rect 174659 524089 174895 524325
rect 174659 520281 174895 520517
rect 174659 516473 174895 516709
rect 177817 528557 178053 528793
rect 177817 524749 178053 524985
rect 177817 520941 178053 521177
rect 177817 517133 178053 517369
rect 178477 527897 178713 528133
rect 178477 524089 178713 524325
rect 178477 520281 178713 520517
rect 178477 516473 178713 516709
rect 181635 528557 181871 528793
rect 181635 524749 181871 524985
rect 181635 520941 181871 521177
rect 181635 517133 181871 517369
rect 182295 527897 182531 528133
rect 182295 524089 182531 524325
rect 182295 520281 182531 520517
rect 182295 516473 182531 516709
rect 185453 528557 185689 528793
rect 185453 524749 185689 524985
rect 185453 520941 185689 521177
rect 185453 517133 185689 517369
rect 186113 527897 186349 528133
rect 186113 524089 186349 524325
rect 186113 520281 186349 520517
rect 186113 516473 186349 516709
<< metal5 >>
rect 172160 528793 187528 528835
rect 172160 528557 173999 528793
rect 174235 528557 177817 528793
rect 178053 528557 181635 528793
rect 181871 528557 185453 528793
rect 185689 528557 187528 528793
rect 172160 528515 187528 528557
rect 172160 528133 187528 528175
rect 172160 527897 174659 528133
rect 174895 527897 178477 528133
rect 178713 527897 182295 528133
rect 182531 527897 186113 528133
rect 186349 527897 187528 528133
rect 172160 527855 187528 527897
rect 172160 524985 187528 525027
rect 172160 524749 173999 524985
rect 174235 524749 177817 524985
rect 178053 524749 181635 524985
rect 181871 524749 185453 524985
rect 185689 524749 187528 524985
rect 172160 524707 187528 524749
rect 172160 524325 187528 524367
rect 172160 524089 174659 524325
rect 174895 524089 178477 524325
rect 178713 524089 182295 524325
rect 182531 524089 186113 524325
rect 186349 524089 187528 524325
rect 172160 524047 187528 524089
rect 172160 521177 187528 521219
rect 172160 520941 173999 521177
rect 174235 520941 177817 521177
rect 178053 520941 181635 521177
rect 181871 520941 185453 521177
rect 185689 520941 187528 521177
rect 172160 520899 187528 520941
rect 172160 520517 187528 520559
rect 172160 520281 174659 520517
rect 174895 520281 178477 520517
rect 178713 520281 182295 520517
rect 182531 520281 186113 520517
rect 186349 520281 187528 520517
rect 172160 520239 187528 520281
rect 172160 517369 187528 517411
rect 172160 517133 173999 517369
rect 174235 517133 177817 517369
rect 178053 517133 181635 517369
rect 181871 517133 185453 517369
rect 185689 517133 187528 517369
rect 172160 517091 187528 517133
rect 172160 516709 187528 516751
rect 172160 516473 174659 516709
rect 174895 516473 178477 516709
rect 178713 516473 182295 516709
rect 182531 516473 186113 516709
rect 186349 516473 187528 516709
rect 172160 516431 187528 516473
<< res0p35 >>
rect 164314 536431 164388 537519
rect 164632 536431 164706 537519
rect 164950 536431 165024 537519
rect 165268 536431 165342 537519
rect 165586 536431 165660 537519
rect 165904 536431 165978 537519
rect 166222 536431 166296 537519
rect 166540 536431 166614 537519
rect 168086 536431 168160 537519
rect 168404 536431 168478 537519
rect 168722 536431 168796 537519
rect 169040 536431 169114 537519
rect 171822 536431 171896 537519
rect 172140 536431 172214 537519
rect 175340 536431 175414 537519
rect 178940 536991 179014 537519
rect 182240 537271 182314 537519
rect 185540 537411 185614 537519
rect 188840 537315 188914 537519
rect 164284 534091 164358 535179
rect 164602 534091 164676 535179
rect 164920 534091 164994 535179
rect 165238 534091 165312 535179
rect 165556 534091 165630 535179
rect 165874 534091 165948 535179
rect 166192 534091 166266 535179
rect 166510 534091 166584 535179
<< labels >>
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 reset
port 64 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 sdi
port 63 nsew signal input
flabel metal3 s -800 464762 480 464874 0 FreeSans 1120 0 0 0 sclk
port 62 nsew signal input
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 ss
port 61 nsew signal input
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 ib
port 37 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 inp
port 46 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 inn
port 45 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 out
port 44 nsew signal bidirectional
flabel metal1 193000 521000 195000 523000 0 FreeSans 1600 0 0 0 gnd_spi
port 71 nsew
flabel metal1 193000 524000 195000 526000 0 FreeSans 1600 0 0 0 vd_spi
port 73 nsew
flabel space 163528 542565 163728 542755 0 FreeSans 1600 0 0 0 dpga_flat_0.inp
flabel metal2 186228 513055 186428 513245 0 FreeSans 1600 0 0 0 dpga_flat_0.reset
flabel metal2 181908 513095 182108 513285 0 FreeSans 1600 0 0 0 dpga_flat_0.sdi
flabel metal1 192428 539115 192628 539315 0 FreeSans 1600 0 0 0 dpga_flat_0.vd
flabel metal1 192428 540055 192628 540255 0 FreeSans 1600 0 0 0 dpga_flat_0.gnd
flabel metal1 178178 542715 178378 542915 0 FreeSans 1600 0 0 0 dpga_flat_0.inn
flabel metal1 163528 542755 163728 542955 0 FreeSans 1600 0 0 0 dpga_flat_0.inp
flabel metal1 156798 536765 156998 536965 0 FreeSans 1600 0 0 0 dpga_flat_0.out
flabel metal1 163028 533115 163228 533315 0 FreeSans 1600 0 0 0 dpga_flat_0.ib
flabel metal1 192428 522875 192628 523065 0 FreeSans 1600 0 0 0 dpga_flat_0.gndd
flabel metal2 177578 513095 177778 513285 0 FreeSans 1600 0 0 0 dpga_flat_0.sclk
flabel metal2 173248 513095 173448 513285 0 FreeSans 1600 0 0 0 dpga_flat_0.ss
flabel metal1 192428 523395 192628 523585 0 FreeSans 1600 0 0 0 dpga_flat_0.vpwr
flabel metal1 190920 522967 191010 522985 0 FreeSans 1600 0 0 0 dpga_flat_0.vgnd
flabel metal4 174617 515299 174937 530627 0 FreeSans 1920 90 0 0 dpga_flat_0.sr_0.VGND
flabel metal4 178435 515299 178755 530627 0 FreeSans 1920 90 0 0 dpga_flat_0.sr_0.VGND
flabel metal4 182253 515299 182573 530627 0 FreeSans 1920 90 0 0 dpga_flat_0.sr_0.VGND
flabel metal4 186071 515299 186391 530627 0 FreeSans 1920 90 0 0 dpga_flat_0.sr_0.VGND
flabel metal5 172160 527855 187528 528175 0 FreeSans 2560 0 0 0 dpga_flat_0.sr_0.VGND
flabel metal5 172160 524047 187528 524367 0 FreeSans 2560 0 0 0 dpga_flat_0.sr_0.VGND
flabel metal5 172160 520239 187528 520559 0 FreeSans 2560 0 0 0 dpga_flat_0.sr_0.VGND
flabel metal5 172160 516431 187528 516751 0 FreeSans 2560 0 0 0 dpga_flat_0.sr_0.VGND
flabel metal4 173957 515299 174277 530627 0 FreeSans 1920 90 0 0 dpga_flat_0.sr_0.VPWR
flabel metal4 177775 515299 178095 530627 0 FreeSans 1920 90 0 0 dpga_flat_0.sr_0.VPWR
flabel metal4 181593 515299 181913 530627 0 FreeSans 1920 90 0 0 dpga_flat_0.sr_0.VPWR
flabel metal4 185411 515299 185731 530627 0 FreeSans 1920 90 0 0 dpga_flat_0.sr_0.VPWR
flabel metal5 172160 528515 187528 528835 0 FreeSans 2560 0 0 0 dpga_flat_0.sr_0.VPWR
flabel metal5 172160 524707 187528 525027 0 FreeSans 2560 0 0 0 dpga_flat_0.sr_0.VPWR
flabel metal5 172160 520899 187528 521219 0 FreeSans 2560 0 0 0 dpga_flat_0.sr_0.VPWR
flabel metal5 172160 517091 187528 517411 0 FreeSans 2560 0 0 0 dpga_flat_0.sr_0.VPWR
flabel metal2 172410 531955 172466 532755 0 FreeSans 224 90 0 0 dpga_flat_0.sr_0.data[0]
flabel metal2 174526 531955 174582 532755 0 FreeSans 224 90 0 0 dpga_flat_0.sr_0.data[1]
flabel metal2 176642 531955 176698 532755 0 FreeSans 224 90 0 0 dpga_flat_0.sr_0.data[2]
flabel metal2 178758 531955 178814 532755 0 FreeSans 224 90 0 0 dpga_flat_0.sr_0.data[3]
flabel metal2 180874 531955 180930 532755 0 FreeSans 224 90 0 0 dpga_flat_0.sr_0.data[4]
flabel metal2 182990 531955 183046 532755 0 FreeSans 224 90 0 0 dpga_flat_0.sr_0.data[5]
flabel metal2 185106 531955 185162 532755 0 FreeSans 224 90 0 0 dpga_flat_0.sr_0.data[6]
flabel metal2 187222 531955 187278 532755 0 FreeSans 224 90 0 0 dpga_flat_0.sr_0.data[7]
flabel metal2 186302 513099 186358 513899 0 FreeSans 224 90 0 0 dpga_flat_0.sr_0.reset
flabel metal2 177654 513099 177710 513899 0 FreeSans 224 90 0 0 dpga_flat_0.sr_0.sclk
flabel metal2 181978 513099 182034 513899 0 FreeSans 224 90 0 0 dpga_flat_0.sr_0.sdi
flabel metal2 173330 513099 173386 513899 0 FreeSans 224 90 0 0 dpga_flat_0.sr_0.ss
rlabel metal1 179844 515347 179844 515347 0 dpga_flat_0.sr_0.VGND
rlabel metal1 179844 515891 179844 515891 0 dpga_flat_0.sr_0.VPWR
rlabel metal1 176624 529797 176624 529797 0 dpga_flat_0.sr_0._00_
rlabel metal1 178372 530137 178372 530137 0 dpga_flat_0.sr_0._01_
rlabel metal2 179890 529593 179890 529593 0 dpga_flat_0.sr_0._02_
rlabel metal1 181178 529797 181178 529797 0 dpga_flat_0.sr_0._03_
rlabel metal1 180718 528709 180718 528709 0 dpga_flat_0.sr_0._04_
rlabel metal1 176854 530273 176854 530273 0 dpga_flat_0.sr_0._05_
rlabel metal2 176394 528369 176394 528369 0 dpga_flat_0.sr_0._06_
rlabel metal1 175888 529049 175888 529049 0 dpga_flat_0.sr_0._07_
rlabel metal1 177130 528505 177130 528505 0 dpga_flat_0.sr_0._08_
rlabel metal1 178234 529865 178234 529865 0 dpga_flat_0.sr_0._09_
rlabel metal1 178786 530341 178786 530341 0 dpga_flat_0.sr_0._10_
rlabel metal1 179982 530137 179982 530137 0 dpga_flat_0.sr_0._11_
rlabel metal1 182328 530205 182328 530205 0 dpga_flat_0.sr_0._12_
rlabel metal1 180396 528641 180396 528641 0 dpga_flat_0.sr_0._13_
rlabel metal2 177682 529049 177682 529049 0 dpga_flat_0.sr_0.clknet_0_sclk
rlabel metal1 176164 529049 176164 529049 0 dpga_flat_0.sr_0.clknet_1_0__leaf_sclk
rlabel metal2 180534 528879 180534 528879 0 dpga_flat_0.sr_0.clknet_1_1__leaf_sclk
rlabel metal2 172438 531201 172438 531201 0 dpga_flat_0.sr_0.data[0]
rlabel metal2 174554 531201 174554 531201 0 dpga_flat_0.sr_0.data[1]
rlabel metal2 176670 531796 176670 531796 0 dpga_flat_0.sr_0.data[2]
rlabel metal2 178786 531796 178786 531796 0 dpga_flat_0.sr_0.data[3]
rlabel metal2 180902 530963 180902 530963 0 dpga_flat_0.sr_0.data[4]
rlabel metal2 183018 531235 183018 531235 0 dpga_flat_0.sr_0.data[5]
rlabel metal2 185134 531235 185134 531235 0 dpga_flat_0.sr_0.data[6]
rlabel metal1 176893 529729 176893 529729 0 dpga_flat_0.sr_0.net1
rlabel metal1 182098 530341 182098 530341 0 dpga_flat_0.sr_0.net10
rlabel metal2 187250 531728 187250 531728 0 dpga_flat_0.sr_0.net11
rlabel metal1 175428 529593 175428 529593 0 dpga_flat_0.sr_0.net12
rlabel metal1 177176 528641 177176 528641 0 dpga_flat_0.sr_0.net13
rlabel metal1 176256 528641 176256 528641 0 dpga_flat_0.sr_0.net14
rlabel metal1 179338 528063 179338 528063 0 dpga_flat_0.sr_0.net15
rlabel metal1 182052 530273 182052 530273 0 dpga_flat_0.sr_0.net16
rlabel metal2 177682 529899 177682 529899 0 dpga_flat_0.sr_0.net17
rlabel metal1 181730 515789 181730 515789 0 dpga_flat_0.sr_0.net2
rlabel metal1 174462 529185 174462 529185 0 dpga_flat_0.sr_0.net3
rlabel metal2 174830 530069 174830 530069 0 dpga_flat_0.sr_0.net4
rlabel metal2 176762 528403 176762 528403 0 dpga_flat_0.sr_0.net5
rlabel metal2 178234 529321 178234 529321 0 dpga_flat_0.sr_0.net6
rlabel metal1 177958 529763 177958 529763 0 dpga_flat_0.sr_0.net7
rlabel metal1 178970 529933 178970 529933 0 dpga_flat_0.sr_0.net8
rlabel metal1 182604 529797 182604 529797 0 dpga_flat_0.sr_0.net9
rlabel metal2 186514 514650 186514 514650 0 dpga_flat_0.sr_0.reset
rlabel metal2 177682 515609 177682 515609 0 dpga_flat_0.sr_0.sclk
rlabel metal1 182236 515585 182236 515585 0 dpga_flat_0.sr_0.sdi
rlabel metal1 173450 515517 173450 515517 0 dpga_flat_0.sr_0.ss
flabel metal1 173065 530562 173099 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_9.VGND
flabel metal1 173065 530018 173099 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_9.VPWR
flabel nwell 173065 530018 173099 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_9.VPB
flabel pwell 173065 530562 173099 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_9.VNB
rlabel comment 173036 530579 173036 530579 2 dpga_flat_0.sr_0.FILLER_0_0_9.decap_12
flabel metal1 172513 529474 172547 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_3.VGND
flabel metal1 172513 530018 172547 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_3.VPWR
flabel nwell 172513 530018 172547 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_3.VPB
flabel pwell 172513 529474 172547 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_3.VNB
rlabel comment 172484 529491 172484 529491 4 dpga_flat_0.sr_0.FILLER_0_1_3.decap_12
flabel metal1 173617 529474 173651 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_15.VGND
flabel metal1 173617 530018 173651 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_15.VPWR
flabel nwell 173617 530018 173651 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_15.VPB
flabel pwell 173617 529474 173651 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_15.VNB
rlabel comment 173588 529491 173588 529491 4 dpga_flat_0.sr_0.FILLER_0_1_15.decap_12
flabel metal1 172237 530018 172271 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_0_Left_28.VPWR
flabel metal1 172237 530562 172271 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_0_Left_28.VGND
flabel nwell 172237 530018 172271 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_0_Left_28.VPB
flabel pwell 172237 530562 172271 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_0_Left_28.VNB
rlabel comment 172208 530579 172208 530579 2 dpga_flat_0.sr_0.PHY_EDGE_ROW_0_Left_28.decap_3
rlabel metal1 172208 530531 172484 530627 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_0_Left_28.VGND
rlabel metal1 172208 529987 172484 530083 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_0_Left_28.VPWR
flabel metal1 172237 530018 172271 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_1_Left_29.VPWR
flabel metal1 172237 529474 172271 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_1_Left_29.VGND
flabel nwell 172237 530018 172271 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_1_Left_29.VPB
flabel pwell 172237 529474 172271 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_1_Left_29.VNB
rlabel comment 172208 529491 172208 529491 4 dpga_flat_0.sr_0.PHY_EDGE_ROW_1_Left_29.decap_3
rlabel metal1 172208 529443 172484 529539 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_1_Left_29.VGND
rlabel metal1 172208 529987 172484 530083 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_1_Left_29.VPWR
flabel locali 172605 530256 172639 530290 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output4.X
flabel locali 172881 530392 172915 530426 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output4.A
flabel locali 172513 530392 172547 530426 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output4.X
flabel locali 172881 530324 172915 530358 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output4.A
flabel locali 172513 530324 172547 530358 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output4.X
flabel metal1 172973 530562 173007 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output4.VGND
flabel metal1 172973 530018 173007 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output4.VPWR
flabel nwell 172973 530018 173007 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output4.VPB
flabel pwell 172973 530562 173007 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output4.VNB
rlabel comment 173036 530579 173036 530579 8 dpga_flat_0.sr_0.output4.clkbuf_4
rlabel metal1 172484 530531 173036 530627 5 dpga_flat_0.sr_0.output4.VGND
rlabel metal1 172484 529987 173036 530083 5 dpga_flat_0.sr_0.output4.VPWR
flabel metal1 174169 530018 174203 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_21.VPWR
flabel metal1 174169 530562 174203 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_21.VGND
flabel nwell 174169 530018 174203 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_21.VPB
flabel pwell 174169 530562 174203 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_21.VNB
rlabel comment 174140 530579 174140 530579 2 dpga_flat_0.sr_0.FILLER_0_0_21.decap_6
rlabel metal1 174140 530531 174692 530627 5 dpga_flat_0.sr_0.FILLER_0_0_21.VGND
rlabel metal1 174140 529987 174692 530083 5 dpga_flat_0.sr_0.FILLER_0_0_21.VPWR
flabel metal1 174714 530022 174750 530052 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_27.VPWR
flabel metal1 174714 530563 174750 530592 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_27.VGND
flabel nwell 174723 530028 174743 530045 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_27.VPB
flabel pwell 174720 530568 174744 530590 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_27.VNB
rlabel comment 174692 530579 174692 530579 2 dpga_flat_0.sr_0.FILLER_0_0_27.fill_1
rlabel metal1 174692 530531 174784 530627 5 dpga_flat_0.sr_0.FILLER_0_0_27.VGND
rlabel metal1 174692 529987 174784 530083 5 dpga_flat_0.sr_0.FILLER_0_0_27.VPWR
flabel metal1 175450 530022 175486 530052 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_35.VPWR
flabel metal1 175450 530563 175486 530592 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_35.VGND
flabel nwell 175459 530028 175479 530045 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_35.VPB
flabel pwell 175456 530568 175480 530590 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_35.VNB
rlabel comment 175428 530579 175428 530579 2 dpga_flat_0.sr_0.FILLER_0_0_35.fill_1
rlabel metal1 175428 530531 175520 530627 5 dpga_flat_0.sr_0.FILLER_0_0_35.VGND
rlabel metal1 175428 529987 175520 530083 5 dpga_flat_0.sr_0.FILLER_0_0_35.VPWR
flabel metal1 174714 530018 174750 530048 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_27.VPWR
flabel metal1 174714 529478 174750 529507 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_27.VGND
flabel nwell 174723 530025 174743 530042 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_27.VPB
flabel pwell 174720 529480 174744 529502 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_27.VNB
rlabel comment 174692 529491 174692 529491 4 dpga_flat_0.sr_0.FILLER_0_1_27.fill_1
rlabel metal1 174692 529443 174784 529539 1 dpga_flat_0.sr_0.FILLER_0_1_27.VGND
rlabel metal1 174692 529987 174784 530083 1 dpga_flat_0.sr_0.FILLER_0_1_27.VPWR
flabel metal1 174806 530026 174859 530055 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_56.VPWR
flabel metal1 174805 530559 174856 530597 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_56.VGND
rlabel comment 174784 530579 174784 530579 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_56.tapvpwrvgnd_1
rlabel metal1 174784 530531 174876 530627 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_56.VGND
rlabel metal1 174784 529987 174876 530083 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_56.VPWR
flabel locali 175550 530120 175584 530154 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._28_.Q
flabel locali 175550 530188 175584 530222 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._28_.Q
flabel locali 175550 530256 175584 530290 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._28_.Q
flabel locali 175550 530460 175584 530494 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._28_.Q
flabel locali 175845 530392 175879 530426 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._28_.RESET_B
flabel locali 177021 530256 177055 530290 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._28_.D
flabel locali 177296 530256 177330 530290 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._28_.CLK
flabel locali 177296 530324 177330 530358 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._28_.CLK
flabel locali 175845 530324 175879 530358 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._28_.RESET_B
flabel metal1 177297 530562 177331 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._28_.VGND
flabel metal1 177297 530018 177331 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._28_.VPWR
flabel nwell 177297 530018 177331 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._28_.VPB
flabel pwell 177297 530562 177331 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._28_.VNB
rlabel comment 177360 530579 177360 530579 8 dpga_flat_0.sr_0._28_.dfrtp_1
rlabel locali 175831 530372 175879 530452 5 dpga_flat_0.sr_0._28_.RESET_B
rlabel locali 175831 530298 175939 530372 5 dpga_flat_0.sr_0._28_.RESET_B
rlabel metal1 175833 530423 175891 530432 5 dpga_flat_0.sr_0._28_.RESET_B
rlabel metal1 175893 530323 175951 530386 5 dpga_flat_0.sr_0._28_.RESET_B
rlabel metal1 175833 530386 175951 530395 5 dpga_flat_0.sr_0._28_.RESET_B
rlabel metal1 176481 530386 176611 530395 5 dpga_flat_0.sr_0._28_.RESET_B
rlabel metal1 175833 530395 176611 530423 5 dpga_flat_0.sr_0._28_.RESET_B
rlabel metal1 176481 530423 176611 530432 5 dpga_flat_0.sr_0._28_.RESET_B
rlabel metal1 175520 530531 177360 530627 5 dpga_flat_0.sr_0._28_.VGND
rlabel metal1 175520 529987 177360 530083 5 dpga_flat_0.sr_0._28_.VPWR
flabel locali 177296 529916 177330 529950 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._30_.Q
flabel locali 177296 529848 177330 529882 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._30_.Q
flabel locali 177296 529780 177330 529814 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._30_.Q
flabel locali 177296 529576 177330 529610 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._30_.Q
flabel locali 177001 529644 177035 529678 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._30_.RESET_B
flabel locali 175825 529780 175859 529814 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._30_.D
flabel locali 175550 529780 175584 529814 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._30_.CLK
flabel locali 175550 529712 175584 529746 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._30_.CLK
flabel locali 177001 529712 177035 529746 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._30_.RESET_B
flabel metal1 175549 529474 175583 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._30_.VGND
flabel metal1 175549 530018 175583 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._30_.VPWR
flabel nwell 175549 530018 175583 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._30_.VPB
flabel pwell 175549 529474 175583 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._30_.VNB
rlabel comment 175520 529491 175520 529491 4 dpga_flat_0.sr_0._30_.dfrtp_1
rlabel locali 177001 529618 177049 529698 1 dpga_flat_0.sr_0._30_.RESET_B
rlabel locali 176941 529698 177049 529772 1 dpga_flat_0.sr_0._30_.RESET_B
rlabel metal1 176989 529638 177047 529647 1 dpga_flat_0.sr_0._30_.RESET_B
rlabel metal1 176929 529684 176987 529747 1 dpga_flat_0.sr_0._30_.RESET_B
rlabel metal1 176929 529675 177047 529684 1 dpga_flat_0.sr_0._30_.RESET_B
rlabel metal1 176269 529675 176399 529684 1 dpga_flat_0.sr_0._30_.RESET_B
rlabel metal1 176269 529647 177047 529675 1 dpga_flat_0.sr_0._30_.RESET_B
rlabel metal1 176269 529638 176399 529647 1 dpga_flat_0.sr_0._30_.RESET_B
rlabel metal1 175520 529443 177360 529539 1 dpga_flat_0.sr_0._30_.VGND
rlabel metal1 175520 529987 177360 530083 1 dpga_flat_0.sr_0._30_.VPWR
flabel locali 174813 529712 174847 529746 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold1.A
flabel locali 175461 529644 175495 529678 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold1.X
flabel locali 174813 529780 174847 529814 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold1.A
flabel locali 175461 529576 175495 529610 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold1.X
flabel locali 174905 529712 174939 529746 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold1.A
flabel locali 174905 529780 174939 529814 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold1.A
flabel locali 175461 529916 175495 529950 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold1.X
flabel locali 175461 529780 175495 529814 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold1.X
flabel locali 175461 529848 175495 529882 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold1.X
flabel locali 175461 529712 175495 529746 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold1.X
flabel nwell 174813 530018 174847 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold1.VPB
flabel pwell 174813 529474 174847 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold1.VNB
flabel metal1 174813 529474 174847 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold1.VGND
flabel metal1 174813 530018 174847 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold1.VPWR
rlabel comment 174784 529491 174784 529491 4 dpga_flat_0.sr_0.hold1.dlygate4sd3_1
rlabel metal1 174784 529443 175520 529539 1 dpga_flat_0.sr_0.hold1.VGND
rlabel metal1 174784 529987 175520 530083 1 dpga_flat_0.sr_0.hold1.VPWR
flabel locali 174997 530256 175031 530290 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output5.X
flabel locali 175273 530392 175307 530426 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output5.A
flabel locali 174905 530392 174939 530426 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output5.X
flabel locali 175273 530324 175307 530358 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output5.A
flabel locali 174905 530324 174939 530358 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output5.X
flabel metal1 175365 530562 175399 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output5.VGND
flabel metal1 175365 530018 175399 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output5.VPWR
flabel nwell 175365 530018 175399 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output5.VPB
flabel pwell 175365 530562 175399 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output5.VNB
rlabel comment 175428 530579 175428 530579 8 dpga_flat_0.sr_0.output5.clkbuf_4
rlabel metal1 174876 530531 175428 530627 5 dpga_flat_0.sr_0.output5.VGND
rlabel metal1 174876 529987 175428 530083 5 dpga_flat_0.sr_0.output5.VPWR
flabel metal1 177472 530561 177525 530593 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_57.VGND
flabel metal1 177473 530018 177525 530049 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_57.VPWR
flabel nwell 177480 530026 177514 530044 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_57.VPB
flabel pwell 177483 530567 177515 530589 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_57.VNB
rlabel comment 177452 530579 177452 530579 2 dpga_flat_0.sr_0.FILLER_0_0_57.fill_2
rlabel metal1 177452 530531 177636 530627 5 dpga_flat_0.sr_0.FILLER_0_0_57.VGND
rlabel metal1 177452 529987 177636 530083 5 dpga_flat_0.sr_0.FILLER_0_0_57.VPWR
flabel metal1 177474 530018 177510 530048 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_57.VPWR
flabel metal1 177474 529478 177510 529507 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_57.VGND
flabel nwell 177483 530025 177503 530042 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_57.VPB
flabel pwell 177480 529480 177504 529502 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_57.VNB
rlabel comment 177452 529491 177452 529491 4 dpga_flat_0.sr_0.FILLER_0_1_57.fill_1
rlabel metal1 177452 529443 177544 529539 1 dpga_flat_0.sr_0.FILLER_0_1_57.VGND
rlabel metal1 177452 529987 177544 530083 1 dpga_flat_0.sr_0.FILLER_0_1_57.VPWR
flabel metal1 177382 530026 177435 530055 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_57.VPWR
flabel metal1 177381 530559 177432 530597 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_57.VGND
rlabel comment 177360 530579 177360 530579 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_57.tapvpwrvgnd_1
rlabel metal1 177360 530531 177452 530627 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_57.VGND
rlabel metal1 177360 529987 177452 530083 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_57.VPWR
flabel metal1 177382 530015 177435 530044 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_1_61.VPWR
flabel metal1 177381 529473 177432 529511 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_1_61.VGND
rlabel comment 177360 529491 177360 529491 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_1_61.tapvpwrvgnd_1
rlabel metal1 177360 529443 177452 529539 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_1_61.VGND
rlabel metal1 177360 529987 177452 530083 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_1_61.VPWR
flabel metal1 178308 529474 178342 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._18_.VGND
flabel metal1 178308 530018 178342 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._18_.VPWR
flabel locali 177664 529780 177698 529814 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._18_.S
flabel locali 177756 529780 177790 529814 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._18_.S
flabel locali 177848 529644 177882 529678 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._18_.A1
flabel locali 177848 529712 177882 529746 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._18_.A1
flabel locali 177940 529712 177974 529746 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._18_.A0
flabel locali 178308 529576 178342 529610 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._18_.X
flabel locali 178308 529848 178342 529882 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._18_.X
flabel locali 178308 529916 178342 529950 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._18_.X
flabel nwell 178264 530018 178298 530052 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._18_.VPB
flabel pwell 178254 529474 178288 529508 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._18_.VNB
rlabel comment 178372 529491 178372 529491 6 dpga_flat_0.sr_0._18_.mux2_1
rlabel metal1 177544 529443 178372 529539 1 dpga_flat_0.sr_0._18_.VGND
rlabel metal1 177544 529987 178372 530083 1 dpga_flat_0.sr_0._18_.VPWR
flabel locali 178309 530324 178343 530358 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold6.A
flabel locali 177661 530392 177695 530426 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold6.X
flabel locali 178309 530256 178343 530290 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold6.A
flabel locali 177661 530460 177695 530494 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold6.X
flabel locali 178217 530324 178251 530358 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold6.A
flabel locali 178217 530256 178251 530290 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold6.A
flabel locali 177661 530120 177695 530154 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold6.X
flabel locali 177661 530256 177695 530290 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold6.X
flabel locali 177661 530188 177695 530222 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold6.X
flabel locali 177661 530324 177695 530358 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold6.X
flabel nwell 178309 530018 178343 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold6.VPB
flabel pwell 178309 530562 178343 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold6.VNB
flabel metal1 178309 530562 178343 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold6.VGND
flabel metal1 178309 530018 178343 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold6.VPWR
rlabel comment 178372 530579 178372 530579 8 dpga_flat_0.sr_0.hold6.dlygate4sd3_1
rlabel metal1 177636 530531 178372 530627 5 dpga_flat_0.sr_0.hold6.VGND
rlabel metal1 177636 529987 178372 530083 5 dpga_flat_0.sr_0.hold6.VPWR
flabel metal1 179772 530561 179825 530593 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_82.VGND
flabel metal1 179773 530018 179825 530049 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_82.VPWR
flabel nwell 179780 530026 179814 530044 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_82.VPB
flabel pwell 179783 530567 179815 530589 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_82.VNB
rlabel comment 179752 530579 179752 530579 2 dpga_flat_0.sr_0.FILLER_0_0_82.fill_2
rlabel metal1 179752 530531 179936 530627 5 dpga_flat_0.sr_0.FILLER_0_0_82.VGND
rlabel metal1 179752 529987 179936 530083 5 dpga_flat_0.sr_0.FILLER_0_0_82.VPWR
flabel metal1 178585 530562 178619 530596 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._21_.VGND
flabel metal1 178585 530018 178619 530052 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._21_.VPWR
flabel locali 178401 530460 178435 530494 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._21_.X
flabel locali 178401 530188 178435 530222 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._21_.X
flabel locali 178401 530120 178435 530154 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._21_.X
flabel locali 178585 530324 178619 530358 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._21_.A
flabel nwell 178585 530018 178619 530052 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._21_.VPB
flabel pwell 178585 530562 178619 530596 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._21_.VNB
rlabel comment 178372 530579 178372 530579 2 dpga_flat_0.sr_0._21_.clkbuf_1
rlabel metal1 178372 530531 178648 530627 5 dpga_flat_0.sr_0._21_.VGND
rlabel metal1 178372 529987 178648 530083 5 dpga_flat_0.sr_0._21_.VPWR
flabel locali 178402 529916 178436 529950 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._32_.Q
flabel locali 178402 529848 178436 529882 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._32_.Q
flabel locali 178402 529780 178436 529814 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._32_.Q
flabel locali 178402 529576 178436 529610 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._32_.Q
flabel locali 178697 529644 178731 529678 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._32_.RESET_B
flabel locali 179873 529780 179907 529814 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._32_.D
flabel locali 180148 529780 180182 529814 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._32_.CLK
flabel locali 180148 529712 180182 529746 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._32_.CLK
flabel locali 178697 529712 178731 529746 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._32_.RESET_B
flabel metal1 180149 529474 180183 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._32_.VGND
flabel metal1 180149 530018 180183 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._32_.VPWR
flabel nwell 180149 530018 180183 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._32_.VPB
flabel pwell 180149 529474 180183 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._32_.VNB
rlabel comment 180212 529491 180212 529491 6 dpga_flat_0.sr_0._32_.dfrtp_1
rlabel locali 178683 529618 178731 529698 1 dpga_flat_0.sr_0._32_.RESET_B
rlabel locali 178683 529698 178791 529772 1 dpga_flat_0.sr_0._32_.RESET_B
rlabel metal1 178685 529638 178743 529647 1 dpga_flat_0.sr_0._32_.RESET_B
rlabel metal1 178745 529684 178803 529747 1 dpga_flat_0.sr_0._32_.RESET_B
rlabel metal1 178685 529675 178803 529684 1 dpga_flat_0.sr_0._32_.RESET_B
rlabel metal1 179333 529675 179463 529684 1 dpga_flat_0.sr_0._32_.RESET_B
rlabel metal1 178685 529647 179463 529675 1 dpga_flat_0.sr_0._32_.RESET_B
rlabel metal1 179333 529638 179463 529647 1 dpga_flat_0.sr_0._32_.RESET_B
rlabel metal1 178372 529443 180212 529539 1 dpga_flat_0.sr_0._32_.VGND
rlabel metal1 178372 529987 180212 530083 1 dpga_flat_0.sr_0._32_.VPWR
flabel locali 179597 530256 179631 530290 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output6.X
flabel locali 179321 530392 179355 530426 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output6.A
flabel locali 179689 530392 179723 530426 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output6.X
flabel locali 179321 530324 179355 530358 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output6.A
flabel locali 179689 530324 179723 530358 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output6.X
flabel metal1 179229 530562 179263 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output6.VGND
flabel metal1 179229 530018 179263 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output6.VPWR
flabel nwell 179229 530018 179263 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output6.VPB
flabel pwell 179229 530562 179263 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output6.VNB
rlabel comment 179200 530579 179200 530579 2 dpga_flat_0.sr_0.output6.clkbuf_4
rlabel metal1 179200 530531 179752 530627 5 dpga_flat_0.sr_0.output6.VGND
rlabel metal1 179200 529987 179752 530083 5 dpga_flat_0.sr_0.output6.VPWR
flabel locali 178769 530256 178803 530290 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output7.X
flabel locali 179045 530392 179079 530426 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output7.A
flabel locali 178677 530392 178711 530426 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output7.X
flabel locali 179045 530324 179079 530358 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output7.A
flabel locali 178677 530324 178711 530358 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output7.X
flabel metal1 179137 530562 179171 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output7.VGND
flabel metal1 179137 530018 179171 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output7.VPWR
flabel nwell 179137 530018 179171 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output7.VPB
flabel pwell 179137 530562 179171 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output7.VNB
rlabel comment 179200 530579 179200 530579 8 dpga_flat_0.sr_0.output7.clkbuf_4
rlabel metal1 178648 530531 179200 530627 5 dpga_flat_0.sr_0.output7.VGND
rlabel metal1 178648 529987 179200 530083 5 dpga_flat_0.sr_0.output7.VPWR
flabel metal1 180048 530561 180101 530593 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_85.VGND
flabel metal1 180049 530018 180101 530049 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_85.VPWR
flabel nwell 180056 530026 180090 530044 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_85.VPB
flabel pwell 180059 530567 180091 530589 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_85.VNB
rlabel comment 180028 530579 180028 530579 2 dpga_flat_0.sr_0.FILLER_0_0_85.fill_2
rlabel metal1 180028 530531 180212 530627 5 dpga_flat_0.sr_0.FILLER_0_0_85.VGND
rlabel metal1 180028 529987 180212 530083 5 dpga_flat_0.sr_0.FILLER_0_0_85.VPWR
flabel metal1 181062 530022 181098 530052 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_96.VPWR
flabel metal1 181062 530563 181098 530592 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_96.VGND
flabel nwell 181071 530028 181091 530045 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_96.VPB
flabel pwell 181068 530568 181092 530590 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_96.VNB
rlabel comment 181040 530579 181040 530579 2 dpga_flat_0.sr_0.FILLER_0_0_96.fill_1
rlabel metal1 181040 530531 181132 530627 5 dpga_flat_0.sr_0.FILLER_0_0_96.VGND
rlabel metal1 181040 529987 181132 530083 5 dpga_flat_0.sr_0.FILLER_0_0_96.VPWR
flabel metal1 179958 530026 180011 530055 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_58.VPWR
flabel metal1 179957 530559 180008 530597 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_58.VGND
rlabel comment 179936 530579 179936 530579 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_58.tapvpwrvgnd_1
rlabel metal1 179936 530531 180028 530627 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_58.VGND
rlabel metal1 179936 529987 180028 530083 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_58.VPWR
flabel metal1 180242 530562 180276 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._22_.VGND
flabel metal1 180242 530018 180276 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._22_.VPWR
flabel locali 180886 530256 180920 530290 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._22_.S
flabel locali 180794 530256 180828 530290 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._22_.S
flabel locali 180702 530392 180736 530426 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._22_.A1
flabel locali 180702 530324 180736 530358 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._22_.A1
flabel locali 180610 530324 180644 530358 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._22_.A0
flabel locali 180242 530460 180276 530494 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._22_.X
flabel locali 180242 530188 180276 530222 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._22_.X
flabel locali 180242 530120 180276 530154 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._22_.X
flabel nwell 180286 530018 180320 530052 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._22_.VPB
flabel pwell 180296 530562 180330 530596 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._22_.VNB
rlabel comment 180212 530579 180212 530579 2 dpga_flat_0.sr_0._22_.mux2_1
rlabel metal1 180212 530531 181040 530627 5 dpga_flat_0.sr_0._22_.VGND
rlabel metal1 180212 529987 181040 530083 5 dpga_flat_0.sr_0._22_.VPWR
flabel metal1 181896 530562 181930 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._24_.VGND
flabel metal1 181896 530018 181930 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._24_.VPWR
flabel locali 181252 530256 181286 530290 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._24_.S
flabel locali 181344 530256 181378 530290 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._24_.S
flabel locali 181436 530392 181470 530426 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._24_.A1
flabel locali 181436 530324 181470 530358 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._24_.A1
flabel locali 181528 530324 181562 530358 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._24_.A0
flabel locali 181896 530460 181930 530494 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._24_.X
flabel locali 181896 530188 181930 530222 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._24_.X
flabel locali 181896 530120 181930 530154 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._24_.X
flabel nwell 181852 530018 181886 530052 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._24_.VPB
flabel pwell 181842 530562 181876 530596 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._24_.VNB
rlabel comment 181960 530579 181960 530579 8 dpga_flat_0.sr_0._24_.mux2_1
rlabel metal1 181132 530531 181960 530627 5 dpga_flat_0.sr_0._24_.VGND
rlabel metal1 181132 529987 181960 530083 5 dpga_flat_0.sr_0._24_.VPWR
flabel locali 181988 529916 182022 529950 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._33_.Q
flabel locali 181988 529848 182022 529882 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._33_.Q
flabel locali 181988 529780 182022 529814 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._33_.Q
flabel locali 181988 529576 182022 529610 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._33_.Q
flabel locali 181693 529644 181727 529678 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._33_.RESET_B
flabel locali 180517 529780 180551 529814 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._33_.D
flabel locali 180242 529780 180276 529814 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._33_.CLK
flabel locali 180242 529712 180276 529746 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._33_.CLK
flabel locali 181693 529712 181727 529746 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._33_.RESET_B
flabel metal1 180241 529474 180275 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._33_.VGND
flabel metal1 180241 530018 180275 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._33_.VPWR
flabel nwell 180241 530018 180275 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._33_.VPB
flabel pwell 180241 529474 180275 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._33_.VNB
rlabel comment 180212 529491 180212 529491 4 dpga_flat_0.sr_0._33_.dfrtp_1
rlabel locali 181693 529618 181741 529698 1 dpga_flat_0.sr_0._33_.RESET_B
rlabel locali 181633 529698 181741 529772 1 dpga_flat_0.sr_0._33_.RESET_B
rlabel metal1 181681 529638 181739 529647 1 dpga_flat_0.sr_0._33_.RESET_B
rlabel metal1 181621 529684 181679 529747 1 dpga_flat_0.sr_0._33_.RESET_B
rlabel metal1 181621 529675 181739 529684 1 dpga_flat_0.sr_0._33_.RESET_B
rlabel metal1 180961 529675 181091 529684 1 dpga_flat_0.sr_0._33_.RESET_B
rlabel metal1 180961 529647 181739 529675 1 dpga_flat_0.sr_0._33_.RESET_B
rlabel metal1 180961 529638 181091 529647 1 dpga_flat_0.sr_0._33_.RESET_B
rlabel metal1 180212 529443 182052 529539 1 dpga_flat_0.sr_0._33_.VGND
rlabel metal1 180212 529987 182052 530083 1 dpga_flat_0.sr_0._33_.VPWR
flabel locali 182357 530256 182391 530290 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output8.X
flabel locali 182081 530392 182115 530426 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output8.A
flabel locali 182449 530392 182483 530426 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output8.X
flabel locali 182081 530324 182115 530358 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output8.A
flabel locali 182449 530324 182483 530358 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output8.X
flabel metal1 181989 530562 182023 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output8.VGND
flabel metal1 181989 530018 182023 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output8.VPWR
flabel nwell 181989 530018 182023 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output8.VPB
flabel pwell 181989 530562 182023 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output8.VNB
rlabel comment 181960 530579 181960 530579 2 dpga_flat_0.sr_0.output8.clkbuf_4
rlabel metal1 181960 530531 182512 530627 5 dpga_flat_0.sr_0.output8.VGND
rlabel metal1 181960 529987 182512 530083 5 dpga_flat_0.sr_0.output8.VPWR
flabel locali 183277 529712 183311 529746 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold5.A
flabel locali 182629 529644 182663 529678 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold5.X
flabel locali 183277 529780 183311 529814 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold5.A
flabel locali 182629 529576 182663 529610 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold5.X
flabel locali 183185 529712 183219 529746 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold5.A
flabel locali 183185 529780 183219 529814 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold5.A
flabel locali 182629 529916 182663 529950 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold5.X
flabel locali 182629 529780 182663 529814 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold5.X
flabel locali 182629 529848 182663 529882 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold5.X
flabel locali 182629 529712 182663 529746 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold5.X
flabel nwell 183277 530018 183311 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold5.VPB
flabel pwell 183277 529474 183311 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold5.VNB
flabel metal1 183277 529474 183311 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold5.VGND
flabel metal1 183277 530018 183311 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold5.VPWR
rlabel comment 183340 529491 183340 529491 6 dpga_flat_0.sr_0.hold5.dlygate4sd3_1
rlabel metal1 182604 529443 183340 529539 1 dpga_flat_0.sr_0.hold5.VGND
rlabel metal1 182604 529987 183340 530083 1 dpga_flat_0.sr_0.hold5.VPWR
flabel metal1 182534 530015 182587 530044 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_1_62.VPWR
flabel metal1 182533 529473 182584 529511 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_1_62.VGND
rlabel comment 182512 529491 182512 529491 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_1_62.tapvpwrvgnd_1
rlabel metal1 182512 529443 182604 529539 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_1_62.VGND
rlabel metal1 182512 529987 182604 530083 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_1_62.VPWR
flabel metal1 182534 530026 182587 530055 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_59.VPWR
flabel metal1 182533 530559 182584 530597 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_59.VGND
rlabel comment 182512 530579 182512 530579 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_59.tapvpwrvgnd_1
rlabel metal1 182512 530531 182604 530627 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_59.VGND
rlabel metal1 182512 529987 182604 530083 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_59.VPWR
flabel metal1 182442 530018 182478 530048 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_111.VPWR
flabel metal1 182442 529478 182478 529507 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_111.VGND
flabel nwell 182451 530025 182471 530042 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_111.VPB
flabel pwell 182448 529480 182472 529502 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_111.VNB
rlabel comment 182420 529491 182420 529491 4 dpga_flat_0.sr_0.FILLER_0_1_111.fill_1
rlabel metal1 182420 529443 182512 529539 1 dpga_flat_0.sr_0.FILLER_0_1_111.VGND
rlabel metal1 182420 529987 182512 530083 1 dpga_flat_0.sr_0.FILLER_0_1_111.VPWR
flabel metal1 182081 529474 182115 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_107.VGND
flabel metal1 182081 530018 182115 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_107.VPWR
flabel nwell 182081 530018 182115 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_107.VPB
flabel pwell 182081 529474 182115 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_107.VNB
rlabel comment 182052 529491 182052 529491 4 dpga_flat_0.sr_0.FILLER_0_1_107.decap_4
rlabel metal1 182052 529443 182420 529539 1 dpga_flat_0.sr_0.FILLER_0_1_107.VGND
rlabel metal1 182052 529987 182420 530083 1 dpga_flat_0.sr_0.FILLER_0_1_107.VPWR
flabel metal1 182633 530562 182667 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_113.VGND
flabel metal1 182633 530018 182667 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_113.VPWR
flabel nwell 182633 530018 182667 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_113.VPB
flabel pwell 182633 530562 182667 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_113.VNB
rlabel comment 182604 530579 182604 530579 2 dpga_flat_0.sr_0.FILLER_0_0_113.decap_4
rlabel metal1 182604 530531 182972 530627 5 dpga_flat_0.sr_0.FILLER_0_0_113.VGND
rlabel metal1 182604 529987 182972 530083 5 dpga_flat_0.sr_0.FILLER_0_0_113.VPWR
flabel locali 183461 530256 183495 530290 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output9.X
flabel locali 183185 530392 183219 530426 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output9.A
flabel locali 183553 530392 183587 530426 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output9.X
flabel locali 183185 530324 183219 530358 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output9.A
flabel locali 183553 530324 183587 530358 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output9.X
flabel metal1 183093 530562 183127 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output9.VGND
flabel metal1 183093 530018 183127 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output9.VPWR
flabel nwell 183093 530018 183127 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output9.VPB
flabel pwell 183093 530562 183127 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output9.VNB
rlabel comment 183064 530579 183064 530579 2 dpga_flat_0.sr_0.output9.clkbuf_4
rlabel metal1 183064 530531 183616 530627 5 dpga_flat_0.sr_0.output9.VGND
rlabel metal1 183064 529987 183616 530083 5 dpga_flat_0.sr_0.output9.VPWR
flabel metal1 182994 530022 183030 530052 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_117.VPWR
flabel metal1 182994 530563 183030 530592 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_117.VGND
flabel nwell 183003 530028 183023 530045 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_117.VPB
flabel pwell 183000 530568 183024 530590 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_117.VNB
rlabel comment 182972 530579 182972 530579 2 dpga_flat_0.sr_0.FILLER_0_0_117.fill_1
rlabel metal1 182972 530531 183064 530627 5 dpga_flat_0.sr_0.FILLER_0_0_117.VGND
rlabel metal1 182972 529987 183064 530083 5 dpga_flat_0.sr_0.FILLER_0_0_117.VPWR
flabel metal1 183369 529474 183403 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_121.VGND
flabel metal1 183369 530018 183403 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_121.VPWR
flabel nwell 183369 530018 183403 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_121.VPB
flabel pwell 183369 529474 183403 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_121.VNB
rlabel comment 183340 529491 183340 529491 4 dpga_flat_0.sr_0.FILLER_0_1_121.decap_12
flabel metal1 183645 530562 183679 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_124.VGND
flabel metal1 183645 530018 183679 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_124.VPWR
flabel nwell 183645 530018 183679 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_124.VPB
flabel pwell 183645 530562 183679 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_124.VNB
rlabel comment 183616 530579 183616 530579 2 dpga_flat_0.sr_0.FILLER_0_0_124.decap_12
flabel metal1 184749 530562 184783 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_136.VGND
flabel metal1 184749 530018 184783 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_136.VPWR
flabel nwell 184749 530018 184783 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_136.VPB
flabel pwell 184749 530562 184783 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_136.VNB
rlabel comment 184720 530579 184720 530579 2 dpga_flat_0.sr_0.FILLER_0_0_136.decap_4
rlabel metal1 184720 530531 185088 530627 5 dpga_flat_0.sr_0.FILLER_0_0_136.VGND
rlabel metal1 184720 529987 185088 530083 5 dpga_flat_0.sr_0.FILLER_0_0_136.VPWR
flabel metal1 184473 529474 184507 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_133.VGND
flabel metal1 184473 530018 184507 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_133.VPWR
flabel nwell 184473 530018 184507 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_133.VPB
flabel pwell 184473 529474 184507 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_133.VNB
rlabel comment 184444 529491 184444 529491 4 dpga_flat_0.sr_0.FILLER_0_1_133.decap_12
flabel metal1 185577 529474 185611 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_145.VGND
flabel metal1 185577 530018 185611 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_145.VPWR
flabel nwell 185577 530018 185611 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_145.VPB
flabel pwell 185577 529474 185611 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_145.VNB
rlabel comment 185548 529491 185548 529491 4 dpga_flat_0.sr_0.FILLER_0_1_145.decap_12
flabel metal1 185110 530026 185163 530055 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_60.VPWR
flabel metal1 185109 530559 185160 530597 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_60.VGND
rlabel comment 185088 530579 185088 530579 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_60.tapvpwrvgnd_1
rlabel metal1 185088 530531 185180 530627 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_60.VGND
rlabel metal1 185088 529987 185180 530083 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_60.VPWR
flabel locali 185577 530256 185611 530290 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output10.X
flabel locali 185301 530392 185335 530426 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output10.A
flabel locali 185669 530392 185703 530426 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output10.X
flabel locali 185301 530324 185335 530358 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output10.A
flabel locali 185669 530324 185703 530358 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output10.X
flabel metal1 185209 530562 185243 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output10.VGND
flabel metal1 185209 530018 185243 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output10.VPWR
flabel nwell 185209 530018 185243 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output10.VPB
flabel pwell 185209 530562 185243 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output10.VNB
rlabel comment 185180 530579 185180 530579 2 dpga_flat_0.sr_0.output10.clkbuf_4
rlabel metal1 185180 530531 185732 530627 5 dpga_flat_0.sr_0.output10.VGND
rlabel metal1 185180 529987 185732 530083 5 dpga_flat_0.sr_0.output10.VPWR
flabel metal1 185761 530562 185795 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_147.VGND
flabel metal1 185761 530018 185795 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_147.VPWR
flabel nwell 185761 530018 185795 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_147.VPB
flabel pwell 185761 530562 185795 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_147.VNB
rlabel comment 185732 530579 185732 530579 2 dpga_flat_0.sr_0.FILLER_0_0_147.decap_12
flabel metal1 186858 530022 186894 530052 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_159.VPWR
flabel metal1 186858 530563 186894 530592 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_159.VGND
flabel nwell 186867 530028 186887 530045 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_159.VPB
flabel pwell 186864 530568 186888 530590 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_159.VNB
rlabel comment 186836 530579 186836 530579 2 dpga_flat_0.sr_0.FILLER_0_0_159.fill_1
rlabel metal1 186836 530531 186928 530627 5 dpga_flat_0.sr_0.FILLER_0_0_159.VGND
rlabel metal1 186836 529987 186928 530083 5 dpga_flat_0.sr_0.FILLER_0_0_159.VPWR
flabel metal1 186681 530018 186715 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_157.VPWR
flabel metal1 186681 529474 186715 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_157.VGND
flabel nwell 186681 530018 186715 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_157.VPB
flabel pwell 186681 529474 186715 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_157.VNB
rlabel comment 186652 529491 186652 529491 4 dpga_flat_0.sr_0.FILLER_0_1_157.decap_6
rlabel metal1 186652 529443 187204 529539 1 dpga_flat_0.sr_0.FILLER_0_1_157.VGND
rlabel metal1 186652 529987 187204 530083 1 dpga_flat_0.sr_0.FILLER_0_1_157.VPWR
flabel metal1 187417 530018 187451 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_0_Right_0.VPWR
flabel metal1 187417 530562 187451 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_0_Right_0.VGND
flabel nwell 187417 530018 187451 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_0_Right_0.VPB
flabel pwell 187417 530562 187451 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_0_Right_0.VNB
rlabel comment 187480 530579 187480 530579 8 dpga_flat_0.sr_0.PHY_EDGE_ROW_0_Right_0.decap_3
rlabel metal1 187204 530531 187480 530627 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_0_Right_0.VGND
rlabel metal1 187204 529987 187480 530083 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_0_Right_0.VPWR
flabel metal1 187417 530018 187451 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_1_Right_1.VPWR
flabel metal1 187417 529474 187451 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_1_Right_1.VGND
flabel nwell 187417 530018 187451 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_1_Right_1.VPB
flabel pwell 187417 529474 187451 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_1_Right_1.VNB
rlabel comment 187480 529491 187480 529491 6 dpga_flat_0.sr_0.PHY_EDGE_ROW_1_Right_1.decap_3
rlabel metal1 187204 529443 187480 529539 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_1_Right_1.VGND
rlabel metal1 187204 529987 187480 530083 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_1_Right_1.VPWR
flabel locali 187122 530256 187156 530290 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.sr_11.LO
flabel locali 186995 530320 187029 530354 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.sr_11.HI
flabel nwell 186957 530018 186991 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.sr_11.VPB
flabel pwell 186957 530562 186991 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.sr_11.VNB
flabel metal1 186957 530562 186991 530596 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.sr_11.VGND
flabel metal1 186957 530018 186991 530052 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.sr_11.VPWR
rlabel comment 186928 530579 186928 530579 2 dpga_flat_0.sr_0.sr_11.conb_1
flabel comment 186973 530306 186973 530306 0 FreeSans 200 90 0 0 dpga_flat_0.sr_0.sr_11.resistive_li1_ok
flabel comment 187161 530306 187161 530306 0 FreeSans 200 90 0 0 dpga_flat_0.sr_0.sr_11.resistive_li1_ok
flabel comment 187114 530321 187114 530321 0 FreeSans 200 90 0 0 dpga_flat_0.sr_0.sr_11.no_jumper_check
flabel comment 187011 530321 187011 530321 0 FreeSans 200 90 0 0 dpga_flat_0.sr_0.sr_11.no_jumper_check
rlabel metal1 186928 530531 187204 530627 5 dpga_flat_0.sr_0.sr_11.VGND
rlabel metal1 186928 529987 187204 530083 5 dpga_flat_0.sr_0.sr_11.VPWR
flabel metal1 172513 529474 172547 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_3.VGND
flabel metal1 172513 528930 172547 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_3.VPWR
flabel nwell 172513 528930 172547 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_3.VPB
flabel pwell 172513 529474 172547 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_3.VNB
rlabel comment 172484 529491 172484 529491 2 dpga_flat_0.sr_0.FILLER_0_2_3.decap_12
flabel metal1 173617 529474 173651 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_15.VGND
flabel metal1 173617 528930 173651 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_15.VPWR
flabel nwell 173617 528930 173651 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_15.VPB
flabel pwell 173617 529474 173651 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_15.VNB
rlabel comment 173588 529491 173588 529491 2 dpga_flat_0.sr_0.FILLER_0_2_15.decap_12
flabel metal1 172237 528930 172271 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_2_Left_30.VPWR
flabel metal1 172237 529474 172271 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_2_Left_30.VGND
flabel nwell 172237 528930 172271 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_2_Left_30.VPB
flabel pwell 172237 529474 172271 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_2_Left_30.VNB
rlabel comment 172208 529491 172208 529491 2 dpga_flat_0.sr_0.PHY_EDGE_ROW_2_Left_30.decap_3
rlabel metal1 172208 529443 172484 529539 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_2_Left_30.VGND
rlabel metal1 172208 528899 172484 528995 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_2_Left_30.VPWR
flabel metal1 174714 528934 174750 528964 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_27.VPWR
flabel metal1 174714 529475 174750 529504 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_27.VGND
flabel nwell 174723 528940 174743 528957 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_27.VPB
flabel pwell 174720 529480 174744 529502 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_27.VNB
rlabel comment 174692 529491 174692 529491 2 dpga_flat_0.sr_0.FILLER_0_2_27.fill_1
rlabel metal1 174692 529443 174784 529539 5 dpga_flat_0.sr_0.FILLER_0_2_27.VGND
rlabel metal1 174692 528899 174784 528995 5 dpga_flat_0.sr_0.FILLER_0_2_27.VPWR
flabel metal1 174896 529473 174949 529505 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_29.VGND
flabel metal1 174897 528930 174949 528961 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_29.VPWR
flabel nwell 174904 528938 174938 528956 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_29.VPB
flabel pwell 174907 529479 174939 529501 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_29.VNB
rlabel comment 174876 529491 174876 529491 2 dpga_flat_0.sr_0.FILLER_0_2_29.fill_2
rlabel metal1 174876 529443 175060 529539 5 dpga_flat_0.sr_0.FILLER_0_2_29.VGND
rlabel metal1 174876 528899 175060 528995 5 dpga_flat_0.sr_0.FILLER_0_2_29.VPWR
flabel metal1 174806 528938 174859 528967 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_2_63.VPWR
flabel metal1 174805 529471 174856 529509 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_2_63.VGND
rlabel comment 174784 529491 174784 529491 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_2_63.tapvpwrvgnd_1
rlabel metal1 174784 529443 174876 529539 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_2_63.VGND
rlabel metal1 174784 528899 174876 528995 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_2_63.VPWR
flabel metal1 175824 529474 175858 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._14_.VGND
flabel metal1 175824 528930 175858 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._14_.VPWR
flabel locali 175180 529168 175214 529202 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._14_.S
flabel locali 175272 529168 175306 529202 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._14_.S
flabel locali 175364 529304 175398 529338 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._14_.A1
flabel locali 175364 529236 175398 529270 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._14_.A1
flabel locali 175456 529236 175490 529270 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._14_.A0
flabel locali 175824 529372 175858 529406 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._14_.X
flabel locali 175824 529100 175858 529134 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._14_.X
flabel locali 175824 529032 175858 529066 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._14_.X
flabel nwell 175780 528930 175814 528964 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._14_.VPB
flabel pwell 175770 529474 175804 529508 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._14_.VNB
rlabel comment 175888 529491 175888 529491 8 dpga_flat_0.sr_0._14_.mux2_1
rlabel metal1 175060 529443 175888 529539 5 dpga_flat_0.sr_0._14_.VGND
rlabel metal1 175060 528899 175888 528995 5 dpga_flat_0.sr_0._14_.VPWR
flabel locali 176101 529168 176135 529202 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_0__f_sclk.X
flabel locali 176009 529168 176043 529202 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_0__f_sclk.X
flabel locali 176009 529236 176043 529270 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_0__f_sclk.X
flabel locali 176101 529236 176135 529270 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_0__f_sclk.X
flabel locali 176101 529304 176135 529338 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_0__f_sclk.X
flabel locali 176009 529304 176043 529338 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_0__f_sclk.X
flabel locali 177665 529304 177699 529338 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_0__f_sclk.A
flabel locali 177665 529236 177699 529270 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_0__f_sclk.A
flabel pwell 177665 529474 177699 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_0__f_sclk.VNB
flabel pwell 177682 529491 177682 529491 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_0__f_sclk.VNB
flabel nwell 177665 528930 177699 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_0__f_sclk.VPB
flabel nwell 177682 528947 177682 528947 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_0__f_sclk.VPB
flabel metal1 177665 529474 177699 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_0__f_sclk.VGND
flabel metal1 177665 528930 177699 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_0__f_sclk.VPWR
rlabel comment 177728 529491 177728 529491 8 dpga_flat_0.sr_0.clkbuf_1_0__f_sclk.clkbuf_16
rlabel metal1 175888 529443 177728 529539 5 dpga_flat_0.sr_0.clkbuf_1_0__f_sclk.VGND
rlabel metal1 175888 528899 177728 528995 5 dpga_flat_0.sr_0.clkbuf_1_0__f_sclk.VPWR
flabel locali 179504 529032 179538 529066 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._31_.Q
flabel locali 179504 529100 179538 529134 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._31_.Q
flabel locali 179504 529168 179538 529202 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._31_.Q
flabel locali 179504 529372 179538 529406 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._31_.Q
flabel locali 179209 529304 179243 529338 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._31_.RESET_B
flabel locali 178033 529168 178067 529202 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._31_.D
flabel locali 177758 529168 177792 529202 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._31_.CLK
flabel locali 177758 529236 177792 529270 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._31_.CLK
flabel locali 179209 529236 179243 529270 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._31_.RESET_B
flabel metal1 177757 529474 177791 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._31_.VGND
flabel metal1 177757 528930 177791 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._31_.VPWR
flabel nwell 177757 528930 177791 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._31_.VPB
flabel pwell 177757 529474 177791 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._31_.VNB
rlabel comment 177728 529491 177728 529491 2 dpga_flat_0.sr_0._31_.dfrtp_1
rlabel locali 179209 529284 179257 529364 5 dpga_flat_0.sr_0._31_.RESET_B
rlabel locali 179149 529210 179257 529284 5 dpga_flat_0.sr_0._31_.RESET_B
rlabel metal1 179197 529335 179255 529344 5 dpga_flat_0.sr_0._31_.RESET_B
rlabel metal1 179137 529235 179195 529298 5 dpga_flat_0.sr_0._31_.RESET_B
rlabel metal1 179137 529298 179255 529307 5 dpga_flat_0.sr_0._31_.RESET_B
rlabel metal1 178477 529298 178607 529307 5 dpga_flat_0.sr_0._31_.RESET_B
rlabel metal1 178477 529307 179255 529335 5 dpga_flat_0.sr_0._31_.RESET_B
rlabel metal1 178477 529335 178607 529344 5 dpga_flat_0.sr_0._31_.RESET_B
rlabel metal1 177728 529443 179568 529539 5 dpga_flat_0.sr_0._31_.VGND
rlabel metal1 177728 528899 179568 528995 5 dpga_flat_0.sr_0._31_.VPWR
flabel metal1 179590 528934 179626 528964 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_80.VPWR
flabel metal1 179590 529475 179626 529504 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_80.VGND
flabel nwell 179599 528940 179619 528957 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_80.VPB
flabel pwell 179596 529480 179620 529502 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_80.VNB
rlabel comment 179568 529491 179568 529491 2 dpga_flat_0.sr_0.FILLER_0_2_80.fill_1
rlabel metal1 179568 529443 179660 529539 5 dpga_flat_0.sr_0.FILLER_0_2_80.VGND
rlabel metal1 179568 528899 179660 528995 5 dpga_flat_0.sr_0.FILLER_0_2_80.VPWR
flabel metal1 179689 529474 179723 529508 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._23_.VGND
flabel metal1 179689 528930 179723 528964 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._23_.VPWR
flabel locali 179873 529372 179907 529406 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._23_.X
flabel locali 179873 529100 179907 529134 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._23_.X
flabel locali 179873 529032 179907 529066 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._23_.X
flabel locali 179689 529236 179723 529270 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._23_.A
flabel nwell 179689 528930 179723 528964 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._23_.VPB
flabel pwell 179689 529474 179723 529508 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._23_.VNB
rlabel comment 179936 529491 179936 529491 8 dpga_flat_0.sr_0._23_.clkbuf_1
rlabel metal1 179660 529443 179936 529539 5 dpga_flat_0.sr_0._23_.VGND
rlabel metal1 179660 528899 179936 528995 5 dpga_flat_0.sr_0._23_.VPWR
flabel metal1 180057 528930 180091 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_85.VPWR
flabel metal1 180057 529474 180091 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_85.VGND
flabel nwell 180057 528930 180091 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_85.VPB
flabel pwell 180057 529474 180091 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_85.VNB
rlabel comment 180028 529491 180028 529491 2 dpga_flat_0.sr_0.FILLER_0_2_85.decap_6
rlabel metal1 180028 529443 180580 529539 5 dpga_flat_0.sr_0.FILLER_0_2_85.VGND
rlabel metal1 180028 528899 180580 528995 5 dpga_flat_0.sr_0.FILLER_0_2_85.VPWR
flabel metal1 180602 528934 180638 528964 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_91.VPWR
flabel metal1 180602 529475 180638 529504 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_91.VGND
flabel nwell 180611 528940 180631 528957 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_91.VPB
flabel pwell 180608 529480 180632 529502 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_91.VNB
rlabel comment 180580 529491 180580 529491 2 dpga_flat_0.sr_0.FILLER_0_2_91.fill_1
rlabel metal1 180580 529443 180672 529539 5 dpga_flat_0.sr_0.FILLER_0_2_91.VGND
rlabel metal1 180580 528899 180672 528995 5 dpga_flat_0.sr_0.FILLER_0_2_91.VPWR
flabel metal1 179958 528938 180011 528967 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_2_64.VPWR
flabel metal1 179957 529471 180008 529509 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_2_64.VGND
rlabel comment 179936 529491 179936 529491 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_2_64.tapvpwrvgnd_1
rlabel metal1 179936 529443 180028 529539 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_2_64.VGND
rlabel metal1 179936 528899 180028 528995 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_2_64.VPWR
flabel locali 182265 529168 182299 529202 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_1__f_sclk.X
flabel locali 182357 529168 182391 529202 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_1__f_sclk.X
flabel locali 182357 529236 182391 529270 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_1__f_sclk.X
flabel locali 182265 529236 182299 529270 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_1__f_sclk.X
flabel locali 182265 529304 182299 529338 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_1__f_sclk.X
flabel locali 182357 529304 182391 529338 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_1__f_sclk.X
flabel locali 180701 529304 180735 529338 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_1__f_sclk.A
flabel locali 180701 529236 180735 529270 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_1__f_sclk.A
flabel pwell 180701 529474 180735 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_1__f_sclk.VNB
flabel pwell 180718 529491 180718 529491 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_1__f_sclk.VNB
flabel nwell 180701 528930 180735 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_1__f_sclk.VPB
flabel nwell 180718 528947 180718 528947 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_1__f_sclk.VPB
flabel metal1 180701 529474 180735 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_1__f_sclk.VGND
flabel metal1 180701 528930 180735 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_1__f_sclk.VPWR
rlabel comment 180672 529491 180672 529491 2 dpga_flat_0.sr_0.clkbuf_1_1__f_sclk.clkbuf_16
rlabel metal1 180672 529443 182512 529539 5 dpga_flat_0.sr_0.clkbuf_1_1__f_sclk.VGND
rlabel metal1 180672 528899 182512 528995 5 dpga_flat_0.sr_0.clkbuf_1_1__f_sclk.VPWR
flabel metal1 182817 529474 182851 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_115.VGND
flabel metal1 182817 528930 182851 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_115.VPWR
flabel nwell 182817 528930 182851 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_115.VPB
flabel pwell 182817 529474 182851 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_115.VNB
rlabel comment 182788 529491 182788 529491 2 dpga_flat_0.sr_0.FILLER_0_2_115.decap_12
flabel metal1 182725 529474 182759 529508 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._25_.VGND
flabel metal1 182725 528930 182759 528964 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._25_.VPWR
flabel locali 182541 529372 182575 529406 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._25_.X
flabel locali 182541 529100 182575 529134 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._25_.X
flabel locali 182541 529032 182575 529066 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._25_.X
flabel locali 182725 529236 182759 529270 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._25_.A
flabel nwell 182725 528930 182759 528964 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._25_.VPB
flabel pwell 182725 529474 182759 529508 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._25_.VNB
rlabel comment 182512 529491 182512 529491 2 dpga_flat_0.sr_0._25_.clkbuf_1
rlabel metal1 182512 529443 182788 529539 5 dpga_flat_0.sr_0._25_.VGND
rlabel metal1 182512 528899 182788 528995 5 dpga_flat_0.sr_0._25_.VPWR
flabel metal1 183921 529474 183955 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_127.VGND
flabel metal1 183921 528930 183955 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_127.VPWR
flabel nwell 183921 528930 183955 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_127.VPB
flabel pwell 183921 529474 183955 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_127.VNB
rlabel comment 183892 529491 183892 529491 2 dpga_flat_0.sr_0.FILLER_0_2_127.decap_12
flabel metal1 185018 528934 185054 528964 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_139.VPWR
flabel metal1 185018 529475 185054 529504 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_139.VGND
flabel nwell 185027 528940 185047 528957 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_139.VPB
flabel pwell 185024 529480 185048 529502 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_139.VNB
rlabel comment 184996 529491 184996 529491 2 dpga_flat_0.sr_0.FILLER_0_2_139.fill_1
rlabel metal1 184996 529443 185088 529539 5 dpga_flat_0.sr_0.FILLER_0_2_139.VGND
rlabel metal1 184996 528899 185088 528995 5 dpga_flat_0.sr_0.FILLER_0_2_139.VPWR
flabel metal1 185209 529474 185243 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_141.VGND
flabel metal1 185209 528930 185243 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_141.VPWR
flabel nwell 185209 528930 185243 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_141.VPB
flabel pwell 185209 529474 185243 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_141.VNB
rlabel comment 185180 529491 185180 529491 2 dpga_flat_0.sr_0.FILLER_0_2_141.decap_12
flabel metal1 185110 528938 185163 528967 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_2_65.VPWR
flabel metal1 185109 529471 185160 529509 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_2_65.VGND
rlabel comment 185088 529491 185088 529491 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_2_65.tapvpwrvgnd_1
rlabel metal1 185088 529443 185180 529539 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_2_65.VGND
rlabel metal1 185088 528899 185180 528995 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_2_65.VPWR
flabel metal1 186313 528930 186347 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_153.VPWR
flabel metal1 186313 529474 186347 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_153.VGND
flabel nwell 186313 528930 186347 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_153.VPB
flabel pwell 186313 529474 186347 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_153.VNB
rlabel comment 186284 529491 186284 529491 2 dpga_flat_0.sr_0.FILLER_0_2_153.decap_8
rlabel metal1 186284 529443 187020 529539 5 dpga_flat_0.sr_0.FILLER_0_2_153.VGND
rlabel metal1 186284 528899 187020 528995 5 dpga_flat_0.sr_0.FILLER_0_2_153.VPWR
flabel metal1 187040 529473 187093 529505 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_161.VGND
flabel metal1 187041 528930 187093 528961 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_161.VPWR
flabel nwell 187048 528938 187082 528956 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_161.VPB
flabel pwell 187051 529479 187083 529501 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_161.VNB
rlabel comment 187020 529491 187020 529491 2 dpga_flat_0.sr_0.FILLER_0_2_161.fill_2
rlabel metal1 187020 529443 187204 529539 5 dpga_flat_0.sr_0.FILLER_0_2_161.VGND
rlabel metal1 187020 528899 187204 528995 5 dpga_flat_0.sr_0.FILLER_0_2_161.VPWR
flabel metal1 187417 528930 187451 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_2_Right_2.VPWR
flabel metal1 187417 529474 187451 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_2_Right_2.VGND
flabel nwell 187417 528930 187451 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_2_Right_2.VPB
flabel pwell 187417 529474 187451 529508 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_2_Right_2.VNB
rlabel comment 187480 529491 187480 529491 8 dpga_flat_0.sr_0.PHY_EDGE_ROW_2_Right_2.decap_3
rlabel metal1 187204 529443 187480 529539 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_2_Right_2.VGND
rlabel metal1 187204 528899 187480 528995 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_2_Right_2.VPWR
flabel metal1 172513 528386 172547 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_3.VGND
flabel metal1 172513 528930 172547 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_3.VPWR
flabel nwell 172513 528930 172547 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_3.VPB
flabel pwell 172513 528386 172547 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_3.VNB
rlabel comment 172484 528403 172484 528403 4 dpga_flat_0.sr_0.FILLER_0_3_3.decap_12
flabel metal1 173617 528386 173651 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_15.VGND
flabel metal1 173617 528930 173651 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_15.VPWR
flabel nwell 173617 528930 173651 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_15.VPB
flabel pwell 173617 528386 173651 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_15.VNB
rlabel comment 173588 528403 173588 528403 4 dpga_flat_0.sr_0.FILLER_0_3_15.decap_12
flabel metal1 172237 528930 172271 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_3_Left_31.VPWR
flabel metal1 172237 528386 172271 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_3_Left_31.VGND
flabel nwell 172237 528930 172271 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_3_Left_31.VPB
flabel pwell 172237 528386 172271 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_3_Left_31.VNB
rlabel comment 172208 528403 172208 528403 4 dpga_flat_0.sr_0.PHY_EDGE_ROW_3_Left_31.decap_3
rlabel metal1 172208 528355 172484 528451 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_3_Left_31.VGND
rlabel metal1 172208 528899 172484 528995 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_3_Left_31.VPWR
flabel metal1 174721 528386 174755 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_27.VGND
flabel metal1 174721 528930 174755 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_27.VPWR
flabel nwell 174721 528930 174755 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_27.VPB
flabel pwell 174721 528386 174755 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_27.VNB
rlabel comment 174692 528403 174692 528403 4 dpga_flat_0.sr_0.FILLER_0_3_27.decap_12
flabel metal1 175818 528930 175854 528960 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_39.VPWR
flabel metal1 175818 528390 175854 528419 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_39.VGND
flabel nwell 175827 528937 175847 528954 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_39.VPB
flabel pwell 175824 528392 175848 528414 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_39.VNB
rlabel comment 175796 528403 175796 528403 4 dpga_flat_0.sr_0.FILLER_0_3_39.fill_1
rlabel metal1 175796 528355 175888 528451 1 dpga_flat_0.sr_0.FILLER_0_3_39.VGND
rlabel metal1 175796 528899 175888 528995 1 dpga_flat_0.sr_0.FILLER_0_3_39.VPWR
flabel metal1 175917 528386 175951 528420 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._15_.VGND
flabel metal1 175917 528930 175951 528964 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._15_.VPWR
flabel locali 176101 528488 176135 528522 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._15_.X
flabel locali 176101 528760 176135 528794 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._15_.X
flabel locali 176101 528828 176135 528862 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._15_.X
flabel locali 175917 528624 175951 528658 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._15_.A
flabel nwell 175917 528930 175951 528964 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._15_.VPB
flabel pwell 175917 528386 175951 528420 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._15_.VNB
rlabel comment 176164 528403 176164 528403 6 dpga_flat_0.sr_0._15_.clkbuf_1
rlabel metal1 175888 528355 176164 528451 1 dpga_flat_0.sr_0._15_.VGND
rlabel metal1 175888 528899 176164 528995 1 dpga_flat_0.sr_0._15_.VPWR
flabel metal1 177290 528930 177326 528960 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_55.VPWR
flabel metal1 177290 528390 177326 528419 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_55.VGND
flabel nwell 177299 528937 177319 528954 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_55.VPB
flabel pwell 177296 528392 177320 528414 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_55.VNB
rlabel comment 177268 528403 177268 528403 4 dpga_flat_0.sr_0.FILLER_0_3_55.fill_1
rlabel metal1 177268 528355 177360 528451 1 dpga_flat_0.sr_0.FILLER_0_3_55.VGND
rlabel metal1 177268 528899 177360 528995 1 dpga_flat_0.sr_0.FILLER_0_3_55.VPWR
flabel metal1 177382 528927 177435 528956 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_3_66.VPWR
flabel metal1 177381 528385 177432 528423 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_3_66.VGND
rlabel comment 177360 528403 177360 528403 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_3_66.tapvpwrvgnd_1
rlabel metal1 177360 528355 177452 528451 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_3_66.VGND
rlabel metal1 177360 528899 177452 528995 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_3_66.VPWR
flabel metal1 177204 528386 177238 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._16_.VGND
flabel metal1 177204 528930 177238 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._16_.VPWR
flabel locali 176560 528692 176594 528726 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._16_.S
flabel locali 176652 528692 176686 528726 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._16_.S
flabel locali 176744 528556 176778 528590 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._16_.A1
flabel locali 176744 528624 176778 528658 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._16_.A1
flabel locali 176836 528624 176870 528658 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._16_.A0
flabel locali 177204 528488 177238 528522 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._16_.X
flabel locali 177204 528760 177238 528794 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._16_.X
flabel locali 177204 528828 177238 528862 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._16_.X
flabel nwell 177160 528930 177194 528964 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._16_.VPB
flabel pwell 177150 528386 177184 528420 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._16_.VNB
rlabel comment 177268 528403 177268 528403 6 dpga_flat_0.sr_0._16_.mux2_1
rlabel metal1 176440 528355 177268 528451 1 dpga_flat_0.sr_0._16_.VGND
rlabel metal1 176440 528899 177268 528995 1 dpga_flat_0.sr_0._16_.VPWR
flabel metal1 176193 528386 176227 528420 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._17_.VGND
flabel metal1 176193 528930 176227 528964 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._17_.VPWR
flabel locali 176377 528488 176411 528522 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._17_.X
flabel locali 176377 528760 176411 528794 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._17_.X
flabel locali 176377 528828 176411 528862 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._17_.X
flabel locali 176193 528624 176227 528658 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._17_.A
flabel nwell 176193 528930 176227 528964 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._17_.VPB
flabel pwell 176193 528386 176227 528420 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._17_.VNB
rlabel comment 176440 528403 176440 528403 6 dpga_flat_0.sr_0._17_.clkbuf_1
rlabel metal1 176164 528355 176440 528451 1 dpga_flat_0.sr_0._17_.VGND
rlabel metal1 176164 528899 176440 528995 1 dpga_flat_0.sr_0._17_.VPWR
flabel locali 178125 528624 178159 528658 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold2.A
flabel locali 177477 528556 177511 528590 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold2.X
flabel locali 178125 528692 178159 528726 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold2.A
flabel locali 177477 528488 177511 528522 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold2.X
flabel locali 178033 528624 178067 528658 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold2.A
flabel locali 178033 528692 178067 528726 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold2.A
flabel locali 177477 528828 177511 528862 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold2.X
flabel locali 177477 528692 177511 528726 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold2.X
flabel locali 177477 528760 177511 528794 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold2.X
flabel locali 177477 528624 177511 528658 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold2.X
flabel nwell 178125 528930 178159 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold2.VPB
flabel pwell 178125 528386 178159 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold2.VNB
flabel metal1 178125 528386 178159 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold2.VGND
flabel metal1 178125 528930 178159 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold2.VPWR
rlabel comment 178188 528403 178188 528403 6 dpga_flat_0.sr_0.hold2.dlygate4sd3_1
rlabel metal1 177452 528355 178188 528451 1 dpga_flat_0.sr_0.hold2.VGND
rlabel metal1 177452 528899 178188 528995 1 dpga_flat_0.sr_0.hold2.VPWR
flabel metal1 178208 528389 178261 528421 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_65.VGND
flabel metal1 178209 528933 178261 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_65.VPWR
flabel nwell 178216 528938 178250 528956 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_65.VPB
flabel pwell 178219 528393 178251 528415 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_65.VNB
rlabel comment 178188 528403 178188 528403 4 dpga_flat_0.sr_0.FILLER_0_3_65.fill_2
rlabel metal1 178188 528355 178372 528451 1 dpga_flat_0.sr_0.FILLER_0_3_65.VGND
rlabel metal1 178188 528899 178372 528995 1 dpga_flat_0.sr_0.FILLER_0_3_65.VPWR
flabel locali 179965 528692 179999 528726 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_0_sclk.X
flabel locali 180057 528692 180091 528726 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_0_sclk.X
flabel locali 180057 528624 180091 528658 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_0_sclk.X
flabel locali 179965 528624 179999 528658 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_0_sclk.X
flabel locali 179965 528556 179999 528590 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_0_sclk.X
flabel locali 180057 528556 180091 528590 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_0_sclk.X
flabel locali 178401 528556 178435 528590 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_0_sclk.A
flabel locali 178401 528624 178435 528658 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_0_sclk.A
flabel pwell 178401 528386 178435 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_0_sclk.VNB
flabel pwell 178418 528403 178418 528403 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_0_sclk.VNB
flabel nwell 178401 528930 178435 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_0_sclk.VPB
flabel nwell 178418 528947 178418 528947 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_0_sclk.VPB
flabel metal1 178401 528386 178435 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_0_sclk.VGND
flabel metal1 178401 528930 178435 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_0_sclk.VPWR
rlabel comment 178372 528403 178372 528403 4 dpga_flat_0.sr_0.clkbuf_0_sclk.clkbuf_16
rlabel metal1 178372 528355 180212 528451 1 dpga_flat_0.sr_0.clkbuf_0_sclk.VGND
rlabel metal1 178372 528899 180212 528995 1 dpga_flat_0.sr_0.clkbuf_0_sclk.VPWR
flabel metal1 180241 528386 180275 528420 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._27_.VGND
flabel metal1 180241 528930 180275 528964 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._27_.VPWR
flabel locali 180425 528488 180459 528522 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._27_.X
flabel locali 180425 528760 180459 528794 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._27_.X
flabel locali 180425 528828 180459 528862 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._27_.X
flabel locali 180241 528624 180275 528658 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._27_.A
flabel nwell 180241 528930 180275 528964 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._27_.VPB
flabel pwell 180241 528386 180275 528420 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._27_.VNB
rlabel comment 180488 528403 180488 528403 6 dpga_flat_0.sr_0._27_.clkbuf_1
rlabel metal1 180212 528355 180488 528451 1 dpga_flat_0.sr_0._27_.VGND
rlabel metal1 180212 528899 180488 528995 1 dpga_flat_0.sr_0._27_.VPWR
flabel locali 182264 528828 182298 528862 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._34_.Q
flabel locali 182264 528760 182298 528794 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._34_.Q
flabel locali 182264 528692 182298 528726 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._34_.Q
flabel locali 182264 528488 182298 528522 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._34_.Q
flabel locali 181969 528556 182003 528590 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._34_.RESET_B
flabel locali 180793 528692 180827 528726 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._34_.D
flabel locali 180518 528692 180552 528726 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._34_.CLK
flabel locali 180518 528624 180552 528658 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._34_.CLK
flabel locali 181969 528624 182003 528658 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._34_.RESET_B
flabel metal1 180517 528386 180551 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._34_.VGND
flabel metal1 180517 528930 180551 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._34_.VPWR
flabel nwell 180517 528930 180551 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._34_.VPB
flabel pwell 180517 528386 180551 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._34_.VNB
rlabel comment 180488 528403 180488 528403 4 dpga_flat_0.sr_0._34_.dfrtp_1
rlabel locali 181969 528530 182017 528610 1 dpga_flat_0.sr_0._34_.RESET_B
rlabel locali 181909 528610 182017 528684 1 dpga_flat_0.sr_0._34_.RESET_B
rlabel metal1 181957 528550 182015 528559 1 dpga_flat_0.sr_0._34_.RESET_B
rlabel metal1 181897 528596 181955 528659 1 dpga_flat_0.sr_0._34_.RESET_B
rlabel metal1 181897 528587 182015 528596 1 dpga_flat_0.sr_0._34_.RESET_B
rlabel metal1 181237 528587 181367 528596 1 dpga_flat_0.sr_0._34_.RESET_B
rlabel metal1 181237 528559 182015 528587 1 dpga_flat_0.sr_0._34_.RESET_B
rlabel metal1 181237 528550 181367 528559 1 dpga_flat_0.sr_0._34_.RESET_B
rlabel metal1 180488 528355 182328 528451 1 dpga_flat_0.sr_0._34_.VGND
rlabel metal1 180488 528899 182328 528995 1 dpga_flat_0.sr_0._34_.VPWR
flabel metal1 182348 528389 182401 528421 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_110.VGND
flabel metal1 182349 528933 182401 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_110.VPWR
flabel nwell 182356 528938 182390 528956 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_110.VPB
flabel pwell 182359 528393 182391 528415 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_110.VNB
rlabel comment 182328 528403 182328 528403 4 dpga_flat_0.sr_0.FILLER_0_3_110.fill_2
rlabel metal1 182328 528355 182512 528451 1 dpga_flat_0.sr_0.FILLER_0_3_110.VGND
rlabel metal1 182328 528899 182512 528995 1 dpga_flat_0.sr_0.FILLER_0_3_110.VPWR
flabel metal1 182633 528386 182667 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_113.VGND
flabel metal1 182633 528930 182667 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_113.VPWR
flabel nwell 182633 528930 182667 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_113.VPB
flabel pwell 182633 528386 182667 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_113.VNB
rlabel comment 182604 528403 182604 528403 4 dpga_flat_0.sr_0.FILLER_0_3_113.decap_12
flabel metal1 183737 528386 183771 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_125.VGND
flabel metal1 183737 528930 183771 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_125.VPWR
flabel nwell 183737 528930 183771 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_125.VPB
flabel pwell 183737 528386 183771 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_125.VNB
rlabel comment 183708 528403 183708 528403 4 dpga_flat_0.sr_0.FILLER_0_3_125.decap_12
flabel metal1 182534 528927 182587 528956 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_3_67.VPWR
flabel metal1 182533 528385 182584 528423 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_3_67.VGND
rlabel comment 182512 528403 182512 528403 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_3_67.tapvpwrvgnd_1
rlabel metal1 182512 528355 182604 528451 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_3_67.VGND
rlabel metal1 182512 528899 182604 528995 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_3_67.VPWR
flabel metal1 184841 528386 184875 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_137.VGND
flabel metal1 184841 528930 184875 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_137.VPWR
flabel nwell 184841 528930 184875 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_137.VPB
flabel pwell 184841 528386 184875 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_137.VNB
rlabel comment 184812 528403 184812 528403 4 dpga_flat_0.sr_0.FILLER_0_3_137.decap_12
flabel metal1 185945 528386 185979 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_149.VGND
flabel metal1 185945 528930 185979 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_149.VPWR
flabel nwell 185945 528930 185979 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_149.VPB
flabel pwell 185945 528386 185979 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_149.VNB
rlabel comment 185916 528403 185916 528403 4 dpga_flat_0.sr_0.FILLER_0_3_149.decap_12
flabel metal1 187040 528389 187093 528421 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_161.VGND
flabel metal1 187041 528933 187093 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_161.VPWR
flabel nwell 187048 528938 187082 528956 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_161.VPB
flabel pwell 187051 528393 187083 528415 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_161.VNB
rlabel comment 187020 528403 187020 528403 4 dpga_flat_0.sr_0.FILLER_0_3_161.fill_2
rlabel metal1 187020 528355 187204 528451 1 dpga_flat_0.sr_0.FILLER_0_3_161.VGND
rlabel metal1 187020 528899 187204 528995 1 dpga_flat_0.sr_0.FILLER_0_3_161.VPWR
flabel metal1 187417 528930 187451 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_3_Right_3.VPWR
flabel metal1 187417 528386 187451 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_3_Right_3.VGND
flabel nwell 187417 528930 187451 528964 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_3_Right_3.VPB
flabel pwell 187417 528386 187451 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_3_Right_3.VNB
rlabel comment 187480 528403 187480 528403 6 dpga_flat_0.sr_0.PHY_EDGE_ROW_3_Right_3.decap_3
rlabel metal1 187204 528355 187480 528451 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_3_Right_3.VGND
rlabel metal1 187204 528899 187480 528995 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_3_Right_3.VPWR
flabel metal1 172513 528386 172547 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_3.VGND
flabel metal1 172513 527842 172547 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_3.VPWR
flabel nwell 172513 527842 172547 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_3.VPB
flabel pwell 172513 528386 172547 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_3.VNB
rlabel comment 172484 528403 172484 528403 2 dpga_flat_0.sr_0.FILLER_0_4_3.decap_12
flabel metal1 173617 528386 173651 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_15.VGND
flabel metal1 173617 527842 173651 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_15.VPWR
flabel nwell 173617 527842 173651 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_15.VPB
flabel pwell 173617 528386 173651 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_15.VNB
rlabel comment 173588 528403 173588 528403 2 dpga_flat_0.sr_0.FILLER_0_4_15.decap_12
flabel metal1 172237 527842 172271 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_4_Left_32.VPWR
flabel metal1 172237 528386 172271 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_4_Left_32.VGND
flabel nwell 172237 527842 172271 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_4_Left_32.VPB
flabel pwell 172237 528386 172271 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_4_Left_32.VNB
rlabel comment 172208 528403 172208 528403 2 dpga_flat_0.sr_0.PHY_EDGE_ROW_4_Left_32.decap_3
rlabel metal1 172208 528355 172484 528451 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_4_Left_32.VGND
rlabel metal1 172208 527811 172484 527907 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_4_Left_32.VPWR
flabel metal1 174714 527846 174750 527876 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_27.VPWR
flabel metal1 174714 528387 174750 528416 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_27.VGND
flabel nwell 174723 527852 174743 527869 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_27.VPB
flabel pwell 174720 528392 174744 528414 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_27.VNB
rlabel comment 174692 528403 174692 528403 2 dpga_flat_0.sr_0.FILLER_0_4_27.fill_1
rlabel metal1 174692 528355 174784 528451 5 dpga_flat_0.sr_0.FILLER_0_4_27.VGND
rlabel metal1 174692 527811 174784 527907 5 dpga_flat_0.sr_0.FILLER_0_4_27.VPWR
flabel metal1 174905 528386 174939 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_29.VGND
flabel metal1 174905 527842 174939 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_29.VPWR
flabel nwell 174905 527842 174939 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_29.VPB
flabel pwell 174905 528386 174939 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_29.VNB
rlabel comment 174876 528403 174876 528403 2 dpga_flat_0.sr_0.FILLER_0_4_29.decap_12
flabel metal1 176002 527846 176038 527876 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_41.VPWR
flabel metal1 176002 528387 176038 528416 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_41.VGND
flabel nwell 176011 527852 176031 527869 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_41.VPB
flabel pwell 176008 528392 176032 528414 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_41.VNB
rlabel comment 175980 528403 175980 528403 2 dpga_flat_0.sr_0.FILLER_0_4_41.fill_1
rlabel metal1 175980 528355 176072 528451 5 dpga_flat_0.sr_0.FILLER_0_4_41.VGND
rlabel metal1 175980 527811 176072 527907 5 dpga_flat_0.sr_0.FILLER_0_4_41.VPWR
flabel metal1 174806 527850 174859 527879 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_4_68.VPWR
flabel metal1 174805 528383 174856 528421 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_4_68.VGND
rlabel comment 174784 528403 174784 528403 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_4_68.tapvpwrvgnd_1
rlabel metal1 174784 528355 174876 528451 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_4_68.VGND
rlabel metal1 174784 527811 174876 527907 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_4_68.VPWR
flabel metal1 178125 528386 178159 528420 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._19_.VGND
flabel metal1 178125 527842 178159 527876 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._19_.VPWR
flabel locali 177941 528284 177975 528318 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._19_.X
flabel locali 177941 528012 177975 528046 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._19_.X
flabel locali 177941 527944 177975 527978 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._19_.X
flabel locali 178125 528148 178159 528182 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._19_.A
flabel nwell 178125 527842 178159 527876 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._19_.VPB
flabel pwell 178125 528386 178159 528420 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._19_.VNB
rlabel comment 177912 528403 177912 528403 2 dpga_flat_0.sr_0._19_.clkbuf_1
rlabel metal1 177912 528355 178188 528451 5 dpga_flat_0.sr_0._19_.VGND
rlabel metal1 177912 527811 178188 527907 5 dpga_flat_0.sr_0._19_.VPWR
flabel locali 177848 527944 177882 527978 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._29_.Q
flabel locali 177848 528012 177882 528046 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._29_.Q
flabel locali 177848 528080 177882 528114 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._29_.Q
flabel locali 177848 528284 177882 528318 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._29_.Q
flabel locali 177553 528216 177587 528250 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._29_.RESET_B
flabel locali 176377 528080 176411 528114 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._29_.D
flabel locali 176102 528080 176136 528114 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._29_.CLK
flabel locali 176102 528148 176136 528182 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._29_.CLK
flabel locali 177553 528148 177587 528182 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._29_.RESET_B
flabel metal1 176101 528386 176135 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._29_.VGND
flabel metal1 176101 527842 176135 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._29_.VPWR
flabel nwell 176101 527842 176135 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._29_.VPB
flabel pwell 176101 528386 176135 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._29_.VNB
rlabel comment 176072 528403 176072 528403 2 dpga_flat_0.sr_0._29_.dfrtp_1
rlabel locali 177553 528196 177601 528276 5 dpga_flat_0.sr_0._29_.RESET_B
rlabel locali 177493 528122 177601 528196 5 dpga_flat_0.sr_0._29_.RESET_B
rlabel metal1 177541 528247 177599 528256 5 dpga_flat_0.sr_0._29_.RESET_B
rlabel metal1 177481 528147 177539 528210 5 dpga_flat_0.sr_0._29_.RESET_B
rlabel metal1 177481 528210 177599 528219 5 dpga_flat_0.sr_0._29_.RESET_B
rlabel metal1 176821 528210 176951 528219 5 dpga_flat_0.sr_0._29_.RESET_B
rlabel metal1 176821 528219 177599 528247 5 dpga_flat_0.sr_0._29_.RESET_B
rlabel metal1 176821 528247 176951 528256 5 dpga_flat_0.sr_0._29_.RESET_B
rlabel metal1 176072 528355 177912 528451 5 dpga_flat_0.sr_0._29_.VGND
rlabel metal1 176072 527811 177912 527907 5 dpga_flat_0.sr_0._29_.VPWR
flabel metal1 178217 527842 178251 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_65.VPWR
flabel metal1 178217 528386 178251 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_65.VGND
flabel nwell 178217 527842 178251 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_65.VPB
flabel pwell 178217 528386 178251 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_65.VNB
rlabel comment 178188 528403 178188 528403 2 dpga_flat_0.sr_0.FILLER_0_4_65.decap_8
rlabel metal1 178188 528355 178924 528451 5 dpga_flat_0.sr_0.FILLER_0_4_65.VGND
rlabel metal1 178188 527811 178924 527907 5 dpga_flat_0.sr_0.FILLER_0_4_65.VPWR
flabel metal1 179772 528385 179825 528417 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_82.VGND
flabel metal1 179773 527842 179825 527873 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_82.VPWR
flabel nwell 179780 527850 179814 527868 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_82.VPB
flabel pwell 179783 528391 179815 528413 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_82.VNB
rlabel comment 179752 528403 179752 528403 2 dpga_flat_0.sr_0.FILLER_0_4_82.fill_2
rlabel metal1 179752 528355 179936 528451 5 dpga_flat_0.sr_0.FILLER_0_4_82.VGND
rlabel metal1 179752 527811 179936 527907 5 dpga_flat_0.sr_0.FILLER_0_4_82.VPWR
flabel metal1 178954 528386 178988 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._20_.VGND
flabel metal1 178954 527842 178988 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._20_.VPWR
flabel locali 179598 528080 179632 528114 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._20_.S
flabel locali 179506 528080 179540 528114 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._20_.S
flabel locali 179414 528216 179448 528250 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._20_.A1
flabel locali 179414 528148 179448 528182 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._20_.A1
flabel locali 179322 528148 179356 528182 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._20_.A0
flabel locali 178954 528284 178988 528318 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._20_.X
flabel locali 178954 528012 178988 528046 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._20_.X
flabel locali 178954 527944 178988 527978 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._20_.X
flabel nwell 178998 527842 179032 527876 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._20_.VPB
flabel pwell 179008 528386 179042 528420 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._20_.VNB
rlabel comment 178924 528403 178924 528403 2 dpga_flat_0.sr_0._20_.mux2_1
rlabel metal1 178924 528355 179752 528451 5 dpga_flat_0.sr_0._20_.VGND
rlabel metal1 178924 527811 179752 527907 5 dpga_flat_0.sr_0._20_.VPWR
flabel metal1 180057 527842 180091 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_85.VPWR
flabel metal1 180057 528386 180091 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_85.VGND
flabel nwell 180057 527842 180091 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_85.VPB
flabel pwell 180057 528386 180091 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_85.VNB
rlabel comment 180028 528403 180028 528403 2 dpga_flat_0.sr_0.FILLER_0_4_85.decap_8
rlabel metal1 180028 528355 180764 528451 5 dpga_flat_0.sr_0.FILLER_0_4_85.VGND
rlabel metal1 180028 527811 180764 527907 5 dpga_flat_0.sr_0.FILLER_0_4_85.VPWR
flabel metal1 180784 528385 180837 528417 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_93.VGND
flabel metal1 180785 527842 180837 527873 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_93.VPWR
flabel nwell 180792 527850 180826 527868 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_93.VPB
flabel pwell 180795 528391 180827 528413 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_93.VNB
rlabel comment 180764 528403 180764 528403 2 dpga_flat_0.sr_0.FILLER_0_4_93.fill_2
rlabel metal1 180764 528355 180948 528451 5 dpga_flat_0.sr_0.FILLER_0_4_93.VGND
rlabel metal1 180764 527811 180948 527907 5 dpga_flat_0.sr_0.FILLER_0_4_93.VPWR
flabel metal1 181805 528386 181839 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_104.VGND
flabel metal1 181805 527842 181839 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_104.VPWR
flabel nwell 181805 527842 181839 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_104.VPB
flabel pwell 181805 528386 181839 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_104.VNB
rlabel comment 181776 528403 181776 528403 2 dpga_flat_0.sr_0.FILLER_0_4_104.decap_12
flabel metal1 179958 527850 180011 527879 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_4_69.VPWR
flabel metal1 179957 528383 180008 528421 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_4_69.VGND
rlabel comment 179936 528403 179936 528403 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_4_69.tapvpwrvgnd_1
rlabel metal1 179936 528355 180028 528451 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_4_69.VGND
rlabel metal1 179936 527811 180028 527907 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_4_69.VPWR
flabel metal1 180978 528386 181012 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._26_.VGND
flabel metal1 180978 527842 181012 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._26_.VPWR
flabel locali 181622 528080 181656 528114 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._26_.S
flabel locali 181530 528080 181564 528114 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._26_.S
flabel locali 181438 528216 181472 528250 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._26_.A1
flabel locali 181438 528148 181472 528182 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._26_.A1
flabel locali 181346 528148 181380 528182 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._26_.A0
flabel locali 180978 528284 181012 528318 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._26_.X
flabel locali 180978 528012 181012 528046 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._26_.X
flabel locali 180978 527944 181012 527978 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._26_.X
flabel nwell 181022 527842 181056 527876 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._26_.VPB
flabel pwell 181032 528386 181066 528420 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._26_.VNB
rlabel comment 180948 528403 180948 528403 2 dpga_flat_0.sr_0._26_.mux2_1
rlabel metal1 180948 528355 181776 528451 5 dpga_flat_0.sr_0._26_.VGND
rlabel metal1 180948 527811 181776 527907 5 dpga_flat_0.sr_0._26_.VPWR
flabel metal1 182909 528386 182943 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_116.VGND
flabel metal1 182909 527842 182943 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_116.VPWR
flabel nwell 182909 527842 182943 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_116.VPB
flabel pwell 182909 528386 182943 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_116.VNB
rlabel comment 182880 528403 182880 528403 2 dpga_flat_0.sr_0.FILLER_0_4_116.decap_12
flabel metal1 184013 528386 184047 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_128.VGND
flabel metal1 184013 527842 184047 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_128.VPWR
flabel nwell 184013 527842 184047 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_128.VPB
flabel pwell 184013 528386 184047 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_128.VNB
rlabel comment 183984 528403 183984 528403 2 dpga_flat_0.sr_0.FILLER_0_4_128.decap_12
flabel metal1 185209 528386 185243 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_141.VGND
flabel metal1 185209 527842 185243 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_141.VPWR
flabel nwell 185209 527842 185243 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_141.VPB
flabel pwell 185209 528386 185243 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_141.VNB
rlabel comment 185180 528403 185180 528403 2 dpga_flat_0.sr_0.FILLER_0_4_141.decap_12
flabel metal1 185110 527850 185163 527879 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_4_70.VPWR
flabel metal1 185109 528383 185160 528421 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_4_70.VGND
rlabel comment 185088 528403 185088 528403 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_4_70.tapvpwrvgnd_1
rlabel metal1 185088 528355 185180 528451 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_4_70.VGND
rlabel metal1 185088 527811 185180 527907 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_4_70.VPWR
flabel metal1 186313 527842 186347 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_153.VPWR
flabel metal1 186313 528386 186347 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_153.VGND
flabel nwell 186313 527842 186347 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_153.VPB
flabel pwell 186313 528386 186347 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_153.VNB
rlabel comment 186284 528403 186284 528403 2 dpga_flat_0.sr_0.FILLER_0_4_153.decap_8
rlabel metal1 186284 528355 187020 528451 5 dpga_flat_0.sr_0.FILLER_0_4_153.VGND
rlabel metal1 186284 527811 187020 527907 5 dpga_flat_0.sr_0.FILLER_0_4_153.VPWR
flabel metal1 187040 528385 187093 528417 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_161.VGND
flabel metal1 187041 527842 187093 527873 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_161.VPWR
flabel nwell 187048 527850 187082 527868 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_161.VPB
flabel pwell 187051 528391 187083 528413 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_161.VNB
rlabel comment 187020 528403 187020 528403 2 dpga_flat_0.sr_0.FILLER_0_4_161.fill_2
rlabel metal1 187020 528355 187204 528451 5 dpga_flat_0.sr_0.FILLER_0_4_161.VGND
rlabel metal1 187020 527811 187204 527907 5 dpga_flat_0.sr_0.FILLER_0_4_161.VPWR
flabel metal1 187417 527842 187451 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_4_Right_4.VPWR
flabel metal1 187417 528386 187451 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_4_Right_4.VGND
flabel nwell 187417 527842 187451 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_4_Right_4.VPB
flabel pwell 187417 528386 187451 528420 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_4_Right_4.VNB
rlabel comment 187480 528403 187480 528403 8 dpga_flat_0.sr_0.PHY_EDGE_ROW_4_Right_4.decap_3
rlabel metal1 187204 528355 187480 528451 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_4_Right_4.VGND
rlabel metal1 187204 527811 187480 527907 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_4_Right_4.VPWR
flabel metal1 172513 527298 172547 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_3.VGND
flabel metal1 172513 527842 172547 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_3.VPWR
flabel nwell 172513 527842 172547 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_3.VPB
flabel pwell 172513 527298 172547 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_3.VNB
rlabel comment 172484 527315 172484 527315 4 dpga_flat_0.sr_0.FILLER_0_5_3.decap_12
flabel metal1 173617 527298 173651 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_15.VGND
flabel metal1 173617 527842 173651 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_15.VPWR
flabel nwell 173617 527842 173651 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_15.VPB
flabel pwell 173617 527298 173651 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_15.VNB
rlabel comment 173588 527315 173588 527315 4 dpga_flat_0.sr_0.FILLER_0_5_15.decap_12
flabel metal1 172237 527842 172271 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_5_Left_33.VPWR
flabel metal1 172237 527298 172271 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_5_Left_33.VGND
flabel nwell 172237 527842 172271 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_5_Left_33.VPB
flabel pwell 172237 527298 172271 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_5_Left_33.VNB
rlabel comment 172208 527315 172208 527315 4 dpga_flat_0.sr_0.PHY_EDGE_ROW_5_Left_33.decap_3
rlabel metal1 172208 527267 172484 527363 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_5_Left_33.VGND
rlabel metal1 172208 527811 172484 527907 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_5_Left_33.VPWR
flabel metal1 174721 527298 174755 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_27.VGND
flabel metal1 174721 527842 174755 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_27.VPWR
flabel nwell 174721 527842 174755 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_27.VPB
flabel pwell 174721 527298 174755 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_27.VNB
rlabel comment 174692 527315 174692 527315 4 dpga_flat_0.sr_0.FILLER_0_5_27.decap_12
flabel metal1 175825 527842 175859 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_39.VPWR
flabel metal1 175825 527298 175859 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_39.VGND
flabel nwell 175825 527842 175859 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_39.VPB
flabel pwell 175825 527298 175859 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_39.VNB
rlabel comment 175796 527315 175796 527315 4 dpga_flat_0.sr_0.FILLER_0_5_39.decap_6
rlabel metal1 175796 527267 176348 527363 1 dpga_flat_0.sr_0.FILLER_0_5_39.VGND
rlabel metal1 175796 527811 176348 527907 1 dpga_flat_0.sr_0.FILLER_0_5_39.VPWR
flabel metal1 177113 527842 177147 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_53.VPWR
flabel metal1 177113 527298 177147 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_53.VGND
flabel nwell 177113 527842 177147 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_53.VPB
flabel pwell 177113 527298 177147 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_53.VNB
rlabel comment 177084 527315 177084 527315 4 dpga_flat_0.sr_0.FILLER_0_5_53.decap_3
rlabel metal1 177084 527267 177360 527363 1 dpga_flat_0.sr_0.FILLER_0_5_53.VGND
rlabel metal1 177084 527811 177360 527907 1 dpga_flat_0.sr_0.FILLER_0_5_53.VPWR
flabel metal1 177481 527298 177515 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_57.VGND
flabel metal1 177481 527842 177515 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_57.VPWR
flabel nwell 177481 527842 177515 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_57.VPB
flabel pwell 177481 527298 177515 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_57.VNB
rlabel comment 177452 527315 177452 527315 4 dpga_flat_0.sr_0.FILLER_0_5_57.decap_12
flabel metal1 177382 527839 177435 527868 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_5_71.VPWR
flabel metal1 177381 527297 177432 527335 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_5_71.VGND
rlabel comment 177360 527315 177360 527315 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_5_71.tapvpwrvgnd_1
rlabel metal1 177360 527267 177452 527363 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_5_71.VGND
rlabel metal1 177360 527811 177452 527907 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_5_71.VPWR
flabel locali 177021 527536 177055 527570 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold3.A
flabel locali 176373 527468 176407 527502 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold3.X
flabel locali 177021 527604 177055 527638 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold3.A
flabel locali 176373 527400 176407 527434 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold3.X
flabel locali 176929 527536 176963 527570 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold3.A
flabel locali 176929 527604 176963 527638 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold3.A
flabel locali 176373 527740 176407 527774 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold3.X
flabel locali 176373 527604 176407 527638 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold3.X
flabel locali 176373 527672 176407 527706 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold3.X
flabel locali 176373 527536 176407 527570 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold3.X
flabel nwell 177021 527842 177055 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold3.VPB
flabel pwell 177021 527298 177055 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold3.VNB
flabel metal1 177021 527298 177055 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold3.VGND
flabel metal1 177021 527842 177055 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold3.VPWR
rlabel comment 177084 527315 177084 527315 6 dpga_flat_0.sr_0.hold3.dlygate4sd3_1
rlabel metal1 176348 527267 177084 527363 1 dpga_flat_0.sr_0.hold3.VGND
rlabel metal1 176348 527811 177084 527907 1 dpga_flat_0.sr_0.hold3.VPWR
flabel metal1 178585 527298 178619 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_69.VGND
flabel metal1 178585 527842 178619 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_69.VPWR
flabel nwell 178585 527842 178619 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_69.VPB
flabel pwell 178585 527298 178619 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_69.VNB
rlabel comment 178556 527315 178556 527315 4 dpga_flat_0.sr_0.FILLER_0_5_69.decap_4
rlabel metal1 178556 527267 178924 527363 1 dpga_flat_0.sr_0.FILLER_0_5_69.VGND
rlabel metal1 178556 527811 178924 527907 1 dpga_flat_0.sr_0.FILLER_0_5_69.VPWR
flabel metal1 179689 527298 179723 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_81.VGND
flabel metal1 179689 527842 179723 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_81.VPWR
flabel nwell 179689 527842 179723 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_81.VPB
flabel pwell 179689 527298 179723 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_81.VNB
rlabel comment 179660 527315 179660 527315 4 dpga_flat_0.sr_0.FILLER_0_5_81.decap_12
flabel locali 179597 527536 179631 527570 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold4.A
flabel locali 178949 527468 178983 527502 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold4.X
flabel locali 179597 527604 179631 527638 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold4.A
flabel locali 178949 527400 178983 527434 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold4.X
flabel locali 179505 527536 179539 527570 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold4.A
flabel locali 179505 527604 179539 527638 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold4.A
flabel locali 178949 527740 178983 527774 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold4.X
flabel locali 178949 527604 178983 527638 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold4.X
flabel locali 178949 527672 178983 527706 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold4.X
flabel locali 178949 527536 178983 527570 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold4.X
flabel nwell 179597 527842 179631 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold4.VPB
flabel pwell 179597 527298 179631 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold4.VNB
flabel metal1 179597 527298 179631 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold4.VGND
flabel metal1 179597 527842 179631 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold4.VPWR
rlabel comment 179660 527315 179660 527315 6 dpga_flat_0.sr_0.hold4.dlygate4sd3_1
rlabel metal1 178924 527267 179660 527363 1 dpga_flat_0.sr_0.hold4.VGND
rlabel metal1 178924 527811 179660 527907 1 dpga_flat_0.sr_0.hold4.VPWR
flabel metal1 180793 527298 180827 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_93.VGND
flabel metal1 180793 527842 180827 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_93.VPWR
flabel nwell 180793 527842 180827 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_93.VPB
flabel pwell 180793 527298 180827 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_93.VNB
rlabel comment 180764 527315 180764 527315 4 dpga_flat_0.sr_0.FILLER_0_5_93.decap_12
flabel metal1 181897 527842 181931 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_105.VPWR
flabel metal1 181897 527298 181931 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_105.VGND
flabel nwell 181897 527842 181931 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_105.VPB
flabel pwell 181897 527298 181931 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_105.VNB
rlabel comment 181868 527315 181868 527315 4 dpga_flat_0.sr_0.FILLER_0_5_105.decap_6
rlabel metal1 181868 527267 182420 527363 1 dpga_flat_0.sr_0.FILLER_0_5_105.VGND
rlabel metal1 181868 527811 182420 527907 1 dpga_flat_0.sr_0.FILLER_0_5_105.VPWR
flabel metal1 182442 527842 182478 527872 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_111.VPWR
flabel metal1 182442 527302 182478 527331 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_111.VGND
flabel nwell 182451 527849 182471 527866 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_111.VPB
flabel pwell 182448 527304 182472 527326 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_111.VNB
rlabel comment 182420 527315 182420 527315 4 dpga_flat_0.sr_0.FILLER_0_5_111.fill_1
rlabel metal1 182420 527267 182512 527363 1 dpga_flat_0.sr_0.FILLER_0_5_111.VGND
rlabel metal1 182420 527811 182512 527907 1 dpga_flat_0.sr_0.FILLER_0_5_111.VPWR
flabel metal1 182633 527298 182667 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_113.VGND
flabel metal1 182633 527842 182667 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_113.VPWR
flabel nwell 182633 527842 182667 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_113.VPB
flabel pwell 182633 527298 182667 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_113.VNB
rlabel comment 182604 527315 182604 527315 4 dpga_flat_0.sr_0.FILLER_0_5_113.decap_12
flabel metal1 183737 527298 183771 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_125.VGND
flabel metal1 183737 527842 183771 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_125.VPWR
flabel nwell 183737 527842 183771 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_125.VPB
flabel pwell 183737 527298 183771 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_125.VNB
rlabel comment 183708 527315 183708 527315 4 dpga_flat_0.sr_0.FILLER_0_5_125.decap_12
flabel metal1 182534 527839 182587 527868 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_5_72.VPWR
flabel metal1 182533 527297 182584 527335 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_5_72.VGND
rlabel comment 182512 527315 182512 527315 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_5_72.tapvpwrvgnd_1
rlabel metal1 182512 527267 182604 527363 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_5_72.VGND
rlabel metal1 182512 527811 182604 527907 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_5_72.VPWR
flabel metal1 184841 527298 184875 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_137.VGND
flabel metal1 184841 527842 184875 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_137.VPWR
flabel nwell 184841 527842 184875 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_137.VPB
flabel pwell 184841 527298 184875 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_137.VNB
rlabel comment 184812 527315 184812 527315 4 dpga_flat_0.sr_0.FILLER_0_5_137.decap_12
flabel metal1 185945 527298 185979 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_149.VGND
flabel metal1 185945 527842 185979 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_149.VPWR
flabel nwell 185945 527842 185979 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_149.VPB
flabel pwell 185945 527298 185979 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_149.VNB
rlabel comment 185916 527315 185916 527315 4 dpga_flat_0.sr_0.FILLER_0_5_149.decap_12
flabel metal1 187040 527301 187093 527333 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_161.VGND
flabel metal1 187041 527845 187093 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_161.VPWR
flabel nwell 187048 527850 187082 527868 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_161.VPB
flabel pwell 187051 527305 187083 527327 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_161.VNB
rlabel comment 187020 527315 187020 527315 4 dpga_flat_0.sr_0.FILLER_0_5_161.fill_2
rlabel metal1 187020 527267 187204 527363 1 dpga_flat_0.sr_0.FILLER_0_5_161.VGND
rlabel metal1 187020 527811 187204 527907 1 dpga_flat_0.sr_0.FILLER_0_5_161.VPWR
flabel metal1 187417 527842 187451 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_5_Right_5.VPWR
flabel metal1 187417 527298 187451 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_5_Right_5.VGND
flabel nwell 187417 527842 187451 527876 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_5_Right_5.VPB
flabel pwell 187417 527298 187451 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_5_Right_5.VNB
rlabel comment 187480 527315 187480 527315 6 dpga_flat_0.sr_0.PHY_EDGE_ROW_5_Right_5.decap_3
rlabel metal1 187204 527267 187480 527363 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_5_Right_5.VGND
rlabel metal1 187204 527811 187480 527907 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_5_Right_5.VPWR
flabel metal1 172513 527298 172547 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_3.VGND
flabel metal1 172513 526754 172547 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_3.VPWR
flabel nwell 172513 526754 172547 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_3.VPB
flabel pwell 172513 527298 172547 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_3.VNB
rlabel comment 172484 527315 172484 527315 2 dpga_flat_0.sr_0.FILLER_0_6_3.decap_12
flabel metal1 173617 527298 173651 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_15.VGND
flabel metal1 173617 526754 173651 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_15.VPWR
flabel nwell 173617 526754 173651 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_15.VPB
flabel pwell 173617 527298 173651 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_15.VNB
rlabel comment 173588 527315 173588 527315 2 dpga_flat_0.sr_0.FILLER_0_6_15.decap_12
flabel metal1 172513 526210 172547 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_3.VGND
flabel metal1 172513 526754 172547 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_3.VPWR
flabel nwell 172513 526754 172547 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_3.VPB
flabel pwell 172513 526210 172547 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_3.VNB
rlabel comment 172484 526227 172484 526227 4 dpga_flat_0.sr_0.FILLER_0_7_3.decap_12
flabel metal1 173617 526210 173651 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_15.VGND
flabel metal1 173617 526754 173651 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_15.VPWR
flabel nwell 173617 526754 173651 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_15.VPB
flabel pwell 173617 526210 173651 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_15.VNB
rlabel comment 173588 526227 173588 526227 4 dpga_flat_0.sr_0.FILLER_0_7_15.decap_12
flabel metal1 172237 526754 172271 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_6_Left_34.VPWR
flabel metal1 172237 527298 172271 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_6_Left_34.VGND
flabel nwell 172237 526754 172271 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_6_Left_34.VPB
flabel pwell 172237 527298 172271 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_6_Left_34.VNB
rlabel comment 172208 527315 172208 527315 2 dpga_flat_0.sr_0.PHY_EDGE_ROW_6_Left_34.decap_3
rlabel metal1 172208 527267 172484 527363 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_6_Left_34.VGND
rlabel metal1 172208 526723 172484 526819 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_6_Left_34.VPWR
flabel metal1 172237 526754 172271 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_7_Left_35.VPWR
flabel metal1 172237 526210 172271 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_7_Left_35.VGND
flabel nwell 172237 526754 172271 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_7_Left_35.VPB
flabel pwell 172237 526210 172271 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_7_Left_35.VNB
rlabel comment 172208 526227 172208 526227 4 dpga_flat_0.sr_0.PHY_EDGE_ROW_7_Left_35.decap_3
rlabel metal1 172208 526179 172484 526275 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_7_Left_35.VGND
rlabel metal1 172208 526723 172484 526819 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_7_Left_35.VPWR
flabel metal1 174714 526758 174750 526788 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_27.VPWR
flabel metal1 174714 527299 174750 527328 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_27.VGND
flabel nwell 174723 526764 174743 526781 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_27.VPB
flabel pwell 174720 527304 174744 527326 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_27.VNB
rlabel comment 174692 527315 174692 527315 2 dpga_flat_0.sr_0.FILLER_0_6_27.fill_1
rlabel metal1 174692 527267 174784 527363 5 dpga_flat_0.sr_0.FILLER_0_6_27.VGND
rlabel metal1 174692 526723 174784 526819 5 dpga_flat_0.sr_0.FILLER_0_6_27.VPWR
flabel metal1 174905 527298 174939 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_29.VGND
flabel metal1 174905 526754 174939 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_29.VPWR
flabel nwell 174905 526754 174939 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_29.VPB
flabel pwell 174905 527298 174939 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_29.VNB
rlabel comment 174876 527315 174876 527315 2 dpga_flat_0.sr_0.FILLER_0_6_29.decap_12
flabel metal1 176009 527298 176043 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_41.VGND
flabel metal1 176009 526754 176043 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_41.VPWR
flabel nwell 176009 526754 176043 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_41.VPB
flabel pwell 176009 527298 176043 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_41.VNB
rlabel comment 175980 527315 175980 527315 2 dpga_flat_0.sr_0.FILLER_0_6_41.decap_12
flabel metal1 174721 526210 174755 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_27.VGND
flabel metal1 174721 526754 174755 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_27.VPWR
flabel nwell 174721 526754 174755 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_27.VPB
flabel pwell 174721 526210 174755 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_27.VNB
rlabel comment 174692 526227 174692 526227 4 dpga_flat_0.sr_0.FILLER_0_7_27.decap_12
flabel metal1 175825 526210 175859 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_39.VGND
flabel metal1 175825 526754 175859 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_39.VPWR
flabel nwell 175825 526754 175859 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_39.VPB
flabel pwell 175825 526210 175859 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_39.VNB
rlabel comment 175796 526227 175796 526227 4 dpga_flat_0.sr_0.FILLER_0_7_39.decap_12
flabel metal1 174806 526762 174859 526791 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_6_73.VPWR
flabel metal1 174805 527295 174856 527333 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_6_73.VGND
rlabel comment 174784 527315 174784 527315 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_6_73.tapvpwrvgnd_1
rlabel metal1 174784 527267 174876 527363 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_6_73.VGND
rlabel metal1 174784 526723 174876 526819 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_6_73.VPWR
flabel metal1 177113 527298 177147 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_53.VGND
flabel metal1 177113 526754 177147 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_53.VPWR
flabel nwell 177113 526754 177147 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_53.VPB
flabel pwell 177113 527298 177147 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_53.VNB
rlabel comment 177084 527315 177084 527315 2 dpga_flat_0.sr_0.FILLER_0_6_53.decap_12
flabel metal1 176929 526210 176963 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_51.VGND
flabel metal1 176929 526754 176963 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_51.VPWR
flabel nwell 176929 526754 176963 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_51.VPB
flabel pwell 176929 526210 176963 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_51.VNB
rlabel comment 176900 526227 176900 526227 4 dpga_flat_0.sr_0.FILLER_0_7_51.decap_4
rlabel metal1 176900 526179 177268 526275 1 dpga_flat_0.sr_0.FILLER_0_7_51.VGND
rlabel metal1 176900 526723 177268 526819 1 dpga_flat_0.sr_0.FILLER_0_7_51.VPWR
flabel metal1 177290 526754 177326 526784 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_55.VPWR
flabel metal1 177290 526214 177326 526243 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_55.VGND
flabel nwell 177299 526761 177319 526778 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_55.VPB
flabel pwell 177296 526216 177320 526238 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_55.VNB
rlabel comment 177268 526227 177268 526227 4 dpga_flat_0.sr_0.FILLER_0_7_55.fill_1
rlabel metal1 177268 526179 177360 526275 1 dpga_flat_0.sr_0.FILLER_0_7_55.VGND
rlabel metal1 177268 526723 177360 526819 1 dpga_flat_0.sr_0.FILLER_0_7_55.VPWR
flabel metal1 177481 526210 177515 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_57.VGND
flabel metal1 177481 526754 177515 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_57.VPWR
flabel nwell 177481 526754 177515 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_57.VPB
flabel pwell 177481 526210 177515 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_57.VNB
rlabel comment 177452 526227 177452 526227 4 dpga_flat_0.sr_0.FILLER_0_7_57.decap_12
flabel metal1 177382 526751 177435 526780 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_7_76.VPWR
flabel metal1 177381 526209 177432 526247 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_7_76.VGND
rlabel comment 177360 526227 177360 526227 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_7_76.tapvpwrvgnd_1
rlabel metal1 177360 526179 177452 526275 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_7_76.VGND
rlabel metal1 177360 526723 177452 526819 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_7_76.VPWR
flabel metal1 178217 527298 178251 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_65.VGND
flabel metal1 178217 526754 178251 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_65.VPWR
flabel nwell 178217 526754 178251 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_65.VPB
flabel pwell 178217 527298 178251 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_65.VNB
rlabel comment 178188 527315 178188 527315 2 dpga_flat_0.sr_0.FILLER_0_6_65.decap_12
flabel metal1 179321 526754 179355 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_77.VPWR
flabel metal1 179321 527298 179355 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_77.VGND
flabel nwell 179321 526754 179355 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_77.VPB
flabel pwell 179321 527298 179355 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_77.VNB
rlabel comment 179292 527315 179292 527315 2 dpga_flat_0.sr_0.FILLER_0_6_77.decap_6
rlabel metal1 179292 527267 179844 527363 5 dpga_flat_0.sr_0.FILLER_0_6_77.VGND
rlabel metal1 179292 526723 179844 526819 5 dpga_flat_0.sr_0.FILLER_0_6_77.VPWR
flabel metal1 179866 526758 179902 526788 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_83.VPWR
flabel metal1 179866 527299 179902 527328 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_83.VGND
flabel nwell 179875 526764 179895 526781 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_83.VPB
flabel pwell 179872 527304 179896 527326 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_83.VNB
rlabel comment 179844 527315 179844 527315 2 dpga_flat_0.sr_0.FILLER_0_6_83.fill_1
rlabel metal1 179844 527267 179936 527363 5 dpga_flat_0.sr_0.FILLER_0_6_83.VGND
rlabel metal1 179844 526723 179936 526819 5 dpga_flat_0.sr_0.FILLER_0_6_83.VPWR
flabel metal1 178585 526210 178619 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_69.VGND
flabel metal1 178585 526754 178619 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_69.VPWR
flabel nwell 178585 526754 178619 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_69.VPB
flabel pwell 178585 526210 178619 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_69.VNB
rlabel comment 178556 526227 178556 526227 4 dpga_flat_0.sr_0.FILLER_0_7_69.decap_12
flabel metal1 179689 526210 179723 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_81.VGND
flabel metal1 179689 526754 179723 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_81.VPWR
flabel nwell 179689 526754 179723 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_81.VPB
flabel pwell 179689 526210 179723 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_81.VNB
rlabel comment 179660 526227 179660 526227 4 dpga_flat_0.sr_0.FILLER_0_7_81.decap_12
flabel metal1 180057 527298 180091 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_85.VGND
flabel metal1 180057 526754 180091 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_85.VPWR
flabel nwell 180057 526754 180091 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_85.VPB
flabel pwell 180057 527298 180091 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_85.VNB
rlabel comment 180028 527315 180028 527315 2 dpga_flat_0.sr_0.FILLER_0_6_85.decap_12
flabel metal1 181161 527298 181195 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_97.VGND
flabel metal1 181161 526754 181195 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_97.VPWR
flabel nwell 181161 526754 181195 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_97.VPB
flabel pwell 181161 527298 181195 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_97.VNB
rlabel comment 181132 527315 181132 527315 2 dpga_flat_0.sr_0.FILLER_0_6_97.decap_12
flabel metal1 180793 526210 180827 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_93.VGND
flabel metal1 180793 526754 180827 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_93.VPWR
flabel nwell 180793 526754 180827 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_93.VPB
flabel pwell 180793 526210 180827 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_93.VNB
rlabel comment 180764 526227 180764 526227 4 dpga_flat_0.sr_0.FILLER_0_7_93.decap_12
flabel metal1 179958 526762 180011 526791 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_6_74.VPWR
flabel metal1 179957 527295 180008 527333 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_6_74.VGND
rlabel comment 179936 527315 179936 527315 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_6_74.tapvpwrvgnd_1
rlabel metal1 179936 527267 180028 527363 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_6_74.VGND
rlabel metal1 179936 526723 180028 526819 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_6_74.VPWR
flabel metal1 182265 527298 182299 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_109.VGND
flabel metal1 182265 526754 182299 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_109.VPWR
flabel nwell 182265 526754 182299 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_109.VPB
flabel pwell 182265 527298 182299 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_109.VNB
rlabel comment 182236 527315 182236 527315 2 dpga_flat_0.sr_0.FILLER_0_6_109.decap_12
flabel metal1 183369 527298 183403 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_121.VGND
flabel metal1 183369 526754 183403 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_121.VPWR
flabel nwell 183369 526754 183403 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_121.VPB
flabel pwell 183369 527298 183403 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_121.VNB
rlabel comment 183340 527315 183340 527315 2 dpga_flat_0.sr_0.FILLER_0_6_121.decap_12
flabel metal1 181897 526754 181931 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_105.VPWR
flabel metal1 181897 526210 181931 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_105.VGND
flabel nwell 181897 526754 181931 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_105.VPB
flabel pwell 181897 526210 181931 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_105.VNB
rlabel comment 181868 526227 181868 526227 4 dpga_flat_0.sr_0.FILLER_0_7_105.decap_6
rlabel metal1 181868 526179 182420 526275 1 dpga_flat_0.sr_0.FILLER_0_7_105.VGND
rlabel metal1 181868 526723 182420 526819 1 dpga_flat_0.sr_0.FILLER_0_7_105.VPWR
flabel metal1 182442 526754 182478 526784 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_111.VPWR
flabel metal1 182442 526214 182478 526243 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_111.VGND
flabel nwell 182451 526761 182471 526778 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_111.VPB
flabel pwell 182448 526216 182472 526238 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_111.VNB
rlabel comment 182420 526227 182420 526227 4 dpga_flat_0.sr_0.FILLER_0_7_111.fill_1
rlabel metal1 182420 526179 182512 526275 1 dpga_flat_0.sr_0.FILLER_0_7_111.VGND
rlabel metal1 182420 526723 182512 526819 1 dpga_flat_0.sr_0.FILLER_0_7_111.VPWR
flabel metal1 182633 526210 182667 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_113.VGND
flabel metal1 182633 526754 182667 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_113.VPWR
flabel nwell 182633 526754 182667 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_113.VPB
flabel pwell 182633 526210 182667 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_113.VNB
rlabel comment 182604 526227 182604 526227 4 dpga_flat_0.sr_0.FILLER_0_7_113.decap_12
flabel metal1 183737 526210 183771 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_125.VGND
flabel metal1 183737 526754 183771 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_125.VPWR
flabel nwell 183737 526754 183771 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_125.VPB
flabel pwell 183737 526210 183771 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_125.VNB
rlabel comment 183708 526227 183708 526227 4 dpga_flat_0.sr_0.FILLER_0_7_125.decap_12
flabel metal1 182534 526751 182587 526780 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_7_77.VPWR
flabel metal1 182533 526209 182584 526247 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_7_77.VGND
rlabel comment 182512 526227 182512 526227 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_7_77.tapvpwrvgnd_1
rlabel metal1 182512 526179 182604 526275 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_7_77.VGND
rlabel metal1 182512 526723 182604 526819 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_7_77.VPWR
flabel metal1 184473 526754 184507 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_133.VPWR
flabel metal1 184473 527298 184507 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_133.VGND
flabel nwell 184473 526754 184507 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_133.VPB
flabel pwell 184473 527298 184507 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_133.VNB
rlabel comment 184444 527315 184444 527315 2 dpga_flat_0.sr_0.FILLER_0_6_133.decap_6
rlabel metal1 184444 527267 184996 527363 5 dpga_flat_0.sr_0.FILLER_0_6_133.VGND
rlabel metal1 184444 526723 184996 526819 5 dpga_flat_0.sr_0.FILLER_0_6_133.VPWR
flabel metal1 185018 526758 185054 526788 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_139.VPWR
flabel metal1 185018 527299 185054 527328 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_139.VGND
flabel nwell 185027 526764 185047 526781 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_139.VPB
flabel pwell 185024 527304 185048 527326 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_139.VNB
rlabel comment 184996 527315 184996 527315 2 dpga_flat_0.sr_0.FILLER_0_6_139.fill_1
rlabel metal1 184996 527267 185088 527363 5 dpga_flat_0.sr_0.FILLER_0_6_139.VGND
rlabel metal1 184996 526723 185088 526819 5 dpga_flat_0.sr_0.FILLER_0_6_139.VPWR
flabel metal1 185209 527298 185243 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_141.VGND
flabel metal1 185209 526754 185243 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_141.VPWR
flabel nwell 185209 526754 185243 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_141.VPB
flabel pwell 185209 527298 185243 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_141.VNB
rlabel comment 185180 527315 185180 527315 2 dpga_flat_0.sr_0.FILLER_0_6_141.decap_12
flabel metal1 184841 526210 184875 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_137.VGND
flabel metal1 184841 526754 184875 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_137.VPWR
flabel nwell 184841 526754 184875 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_137.VPB
flabel pwell 184841 526210 184875 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_137.VNB
rlabel comment 184812 526227 184812 526227 4 dpga_flat_0.sr_0.FILLER_0_7_137.decap_12
flabel metal1 185110 526762 185163 526791 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_6_75.VPWR
flabel metal1 185109 527295 185160 527333 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_6_75.VGND
rlabel comment 185088 527315 185088 527315 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_6_75.tapvpwrvgnd_1
rlabel metal1 185088 527267 185180 527363 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_6_75.VGND
rlabel metal1 185088 526723 185180 526819 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_6_75.VPWR
flabel metal1 186313 526754 186347 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_153.VPWR
flabel metal1 186313 527298 186347 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_153.VGND
flabel nwell 186313 526754 186347 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_153.VPB
flabel pwell 186313 527298 186347 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_153.VNB
rlabel comment 186284 527315 186284 527315 2 dpga_flat_0.sr_0.FILLER_0_6_153.decap_8
rlabel metal1 186284 527267 187020 527363 5 dpga_flat_0.sr_0.FILLER_0_6_153.VGND
rlabel metal1 186284 526723 187020 526819 5 dpga_flat_0.sr_0.FILLER_0_6_153.VPWR
flabel metal1 187040 527297 187093 527329 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_161.VGND
flabel metal1 187041 526754 187093 526785 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_161.VPWR
flabel nwell 187048 526762 187082 526780 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_161.VPB
flabel pwell 187051 527303 187083 527325 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_161.VNB
rlabel comment 187020 527315 187020 527315 2 dpga_flat_0.sr_0.FILLER_0_6_161.fill_2
rlabel metal1 187020 527267 187204 527363 5 dpga_flat_0.sr_0.FILLER_0_6_161.VGND
rlabel metal1 187020 526723 187204 526819 5 dpga_flat_0.sr_0.FILLER_0_6_161.VPWR
flabel metal1 185945 526210 185979 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_149.VGND
flabel metal1 185945 526754 185979 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_149.VPWR
flabel nwell 185945 526754 185979 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_149.VPB
flabel pwell 185945 526210 185979 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_149.VNB
rlabel comment 185916 526227 185916 526227 4 dpga_flat_0.sr_0.FILLER_0_7_149.decap_12
flabel metal1 187040 526213 187093 526245 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_161.VGND
flabel metal1 187041 526757 187093 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_161.VPWR
flabel nwell 187048 526762 187082 526780 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_161.VPB
flabel pwell 187051 526217 187083 526239 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_161.VNB
rlabel comment 187020 526227 187020 526227 4 dpga_flat_0.sr_0.FILLER_0_7_161.fill_2
rlabel metal1 187020 526179 187204 526275 1 dpga_flat_0.sr_0.FILLER_0_7_161.VGND
rlabel metal1 187020 526723 187204 526819 1 dpga_flat_0.sr_0.FILLER_0_7_161.VPWR
flabel metal1 187417 526754 187451 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_6_Right_6.VPWR
flabel metal1 187417 527298 187451 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_6_Right_6.VGND
flabel nwell 187417 526754 187451 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_6_Right_6.VPB
flabel pwell 187417 527298 187451 527332 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_6_Right_6.VNB
rlabel comment 187480 527315 187480 527315 8 dpga_flat_0.sr_0.PHY_EDGE_ROW_6_Right_6.decap_3
rlabel metal1 187204 527267 187480 527363 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_6_Right_6.VGND
rlabel metal1 187204 526723 187480 526819 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_6_Right_6.VPWR
flabel metal1 187417 526754 187451 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_7_Right_7.VPWR
flabel metal1 187417 526210 187451 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_7_Right_7.VGND
flabel nwell 187417 526754 187451 526788 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_7_Right_7.VPB
flabel pwell 187417 526210 187451 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_7_Right_7.VNB
rlabel comment 187480 526227 187480 526227 6 dpga_flat_0.sr_0.PHY_EDGE_ROW_7_Right_7.decap_3
rlabel metal1 187204 526179 187480 526275 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_7_Right_7.VGND
rlabel metal1 187204 526723 187480 526819 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_7_Right_7.VPWR
flabel metal1 172513 526210 172547 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_3.VGND
flabel metal1 172513 525666 172547 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_3.VPWR
flabel nwell 172513 525666 172547 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_3.VPB
flabel pwell 172513 526210 172547 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_3.VNB
rlabel comment 172484 526227 172484 526227 2 dpga_flat_0.sr_0.FILLER_0_8_3.decap_12
flabel metal1 173617 526210 173651 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_15.VGND
flabel metal1 173617 525666 173651 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_15.VPWR
flabel nwell 173617 525666 173651 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_15.VPB
flabel pwell 173617 526210 173651 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_15.VNB
rlabel comment 173588 526227 173588 526227 2 dpga_flat_0.sr_0.FILLER_0_8_15.decap_12
flabel metal1 172237 525666 172271 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_8_Left_36.VPWR
flabel metal1 172237 526210 172271 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_8_Left_36.VGND
flabel nwell 172237 525666 172271 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_8_Left_36.VPB
flabel pwell 172237 526210 172271 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_8_Left_36.VNB
rlabel comment 172208 526227 172208 526227 2 dpga_flat_0.sr_0.PHY_EDGE_ROW_8_Left_36.decap_3
rlabel metal1 172208 526179 172484 526275 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_8_Left_36.VGND
rlabel metal1 172208 525635 172484 525731 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_8_Left_36.VPWR
flabel metal1 174714 525670 174750 525700 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_27.VPWR
flabel metal1 174714 526211 174750 526240 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_27.VGND
flabel nwell 174723 525676 174743 525693 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_27.VPB
flabel pwell 174720 526216 174744 526238 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_27.VNB
rlabel comment 174692 526227 174692 526227 2 dpga_flat_0.sr_0.FILLER_0_8_27.fill_1
rlabel metal1 174692 526179 174784 526275 5 dpga_flat_0.sr_0.FILLER_0_8_27.VGND
rlabel metal1 174692 525635 174784 525731 5 dpga_flat_0.sr_0.FILLER_0_8_27.VPWR
flabel metal1 174905 526210 174939 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_29.VGND
flabel metal1 174905 525666 174939 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_29.VPWR
flabel nwell 174905 525666 174939 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_29.VPB
flabel pwell 174905 526210 174939 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_29.VNB
rlabel comment 174876 526227 174876 526227 2 dpga_flat_0.sr_0.FILLER_0_8_29.decap_12
flabel metal1 176009 526210 176043 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_41.VGND
flabel metal1 176009 525666 176043 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_41.VPWR
flabel nwell 176009 525666 176043 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_41.VPB
flabel pwell 176009 526210 176043 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_41.VNB
rlabel comment 175980 526227 175980 526227 2 dpga_flat_0.sr_0.FILLER_0_8_41.decap_12
flabel metal1 174806 525674 174859 525703 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_8_78.VPWR
flabel metal1 174805 526207 174856 526245 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_8_78.VGND
rlabel comment 174784 526227 174784 526227 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_8_78.tapvpwrvgnd_1
rlabel metal1 174784 526179 174876 526275 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_8_78.VGND
rlabel metal1 174784 525635 174876 525731 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_8_78.VPWR
flabel metal1 177113 526210 177147 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_53.VGND
flabel metal1 177113 525666 177147 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_53.VPWR
flabel nwell 177113 525666 177147 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_53.VPB
flabel pwell 177113 526210 177147 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_53.VNB
rlabel comment 177084 526227 177084 526227 2 dpga_flat_0.sr_0.FILLER_0_8_53.decap_12
flabel metal1 178217 526210 178251 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_65.VGND
flabel metal1 178217 525666 178251 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_65.VPWR
flabel nwell 178217 525666 178251 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_65.VPB
flabel pwell 178217 526210 178251 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_65.VNB
rlabel comment 178188 526227 178188 526227 2 dpga_flat_0.sr_0.FILLER_0_8_65.decap_12
flabel metal1 179321 525666 179355 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_77.VPWR
flabel metal1 179321 526210 179355 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_77.VGND
flabel nwell 179321 525666 179355 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_77.VPB
flabel pwell 179321 526210 179355 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_77.VNB
rlabel comment 179292 526227 179292 526227 2 dpga_flat_0.sr_0.FILLER_0_8_77.decap_6
rlabel metal1 179292 526179 179844 526275 5 dpga_flat_0.sr_0.FILLER_0_8_77.VGND
rlabel metal1 179292 525635 179844 525731 5 dpga_flat_0.sr_0.FILLER_0_8_77.VPWR
flabel metal1 179866 525670 179902 525700 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_83.VPWR
flabel metal1 179866 526211 179902 526240 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_83.VGND
flabel nwell 179875 525676 179895 525693 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_83.VPB
flabel pwell 179872 526216 179896 526238 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_83.VNB
rlabel comment 179844 526227 179844 526227 2 dpga_flat_0.sr_0.FILLER_0_8_83.fill_1
rlabel metal1 179844 526179 179936 526275 5 dpga_flat_0.sr_0.FILLER_0_8_83.VGND
rlabel metal1 179844 525635 179936 525731 5 dpga_flat_0.sr_0.FILLER_0_8_83.VPWR
flabel metal1 180057 526210 180091 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_85.VGND
flabel metal1 180057 525666 180091 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_85.VPWR
flabel nwell 180057 525666 180091 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_85.VPB
flabel pwell 180057 526210 180091 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_85.VNB
rlabel comment 180028 526227 180028 526227 2 dpga_flat_0.sr_0.FILLER_0_8_85.decap_12
flabel metal1 181161 526210 181195 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_97.VGND
flabel metal1 181161 525666 181195 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_97.VPWR
flabel nwell 181161 525666 181195 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_97.VPB
flabel pwell 181161 526210 181195 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_97.VNB
rlabel comment 181132 526227 181132 526227 2 dpga_flat_0.sr_0.FILLER_0_8_97.decap_12
flabel metal1 179958 525674 180011 525703 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_8_79.VPWR
flabel metal1 179957 526207 180008 526245 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_8_79.VGND
rlabel comment 179936 526227 179936 526227 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_8_79.tapvpwrvgnd_1
rlabel metal1 179936 526179 180028 526275 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_8_79.VGND
rlabel metal1 179936 525635 180028 525731 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_8_79.VPWR
flabel metal1 182265 526210 182299 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_109.VGND
flabel metal1 182265 525666 182299 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_109.VPWR
flabel nwell 182265 525666 182299 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_109.VPB
flabel pwell 182265 526210 182299 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_109.VNB
rlabel comment 182236 526227 182236 526227 2 dpga_flat_0.sr_0.FILLER_0_8_109.decap_12
flabel metal1 183369 526210 183403 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_121.VGND
flabel metal1 183369 525666 183403 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_121.VPWR
flabel nwell 183369 525666 183403 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_121.VPB
flabel pwell 183369 526210 183403 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_121.VNB
rlabel comment 183340 526227 183340 526227 2 dpga_flat_0.sr_0.FILLER_0_8_121.decap_12
flabel metal1 184473 525666 184507 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_133.VPWR
flabel metal1 184473 526210 184507 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_133.VGND
flabel nwell 184473 525666 184507 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_133.VPB
flabel pwell 184473 526210 184507 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_133.VNB
rlabel comment 184444 526227 184444 526227 2 dpga_flat_0.sr_0.FILLER_0_8_133.decap_6
rlabel metal1 184444 526179 184996 526275 5 dpga_flat_0.sr_0.FILLER_0_8_133.VGND
rlabel metal1 184444 525635 184996 525731 5 dpga_flat_0.sr_0.FILLER_0_8_133.VPWR
flabel metal1 185018 525670 185054 525700 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_139.VPWR
flabel metal1 185018 526211 185054 526240 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_139.VGND
flabel nwell 185027 525676 185047 525693 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_139.VPB
flabel pwell 185024 526216 185048 526238 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_139.VNB
rlabel comment 184996 526227 184996 526227 2 dpga_flat_0.sr_0.FILLER_0_8_139.fill_1
rlabel metal1 184996 526179 185088 526275 5 dpga_flat_0.sr_0.FILLER_0_8_139.VGND
rlabel metal1 184996 525635 185088 525731 5 dpga_flat_0.sr_0.FILLER_0_8_139.VPWR
flabel metal1 185209 526210 185243 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_141.VGND
flabel metal1 185209 525666 185243 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_141.VPWR
flabel nwell 185209 525666 185243 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_141.VPB
flabel pwell 185209 526210 185243 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_141.VNB
rlabel comment 185180 526227 185180 526227 2 dpga_flat_0.sr_0.FILLER_0_8_141.decap_12
flabel metal1 185110 525674 185163 525703 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_8_80.VPWR
flabel metal1 185109 526207 185160 526245 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_8_80.VGND
rlabel comment 185088 526227 185088 526227 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_8_80.tapvpwrvgnd_1
rlabel metal1 185088 526179 185180 526275 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_8_80.VGND
rlabel metal1 185088 525635 185180 525731 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_8_80.VPWR
flabel metal1 186313 525666 186347 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_153.VPWR
flabel metal1 186313 526210 186347 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_153.VGND
flabel nwell 186313 525666 186347 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_153.VPB
flabel pwell 186313 526210 186347 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_153.VNB
rlabel comment 186284 526227 186284 526227 2 dpga_flat_0.sr_0.FILLER_0_8_153.decap_8
rlabel metal1 186284 526179 187020 526275 5 dpga_flat_0.sr_0.FILLER_0_8_153.VGND
rlabel metal1 186284 525635 187020 525731 5 dpga_flat_0.sr_0.FILLER_0_8_153.VPWR
flabel metal1 187040 526209 187093 526241 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_161.VGND
flabel metal1 187041 525666 187093 525697 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_161.VPWR
flabel nwell 187048 525674 187082 525692 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_161.VPB
flabel pwell 187051 526215 187083 526237 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_161.VNB
rlabel comment 187020 526227 187020 526227 2 dpga_flat_0.sr_0.FILLER_0_8_161.fill_2
rlabel metal1 187020 526179 187204 526275 5 dpga_flat_0.sr_0.FILLER_0_8_161.VGND
rlabel metal1 187020 525635 187204 525731 5 dpga_flat_0.sr_0.FILLER_0_8_161.VPWR
flabel metal1 187417 525666 187451 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_8_Right_8.VPWR
flabel metal1 187417 526210 187451 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_8_Right_8.VGND
flabel nwell 187417 525666 187451 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_8_Right_8.VPB
flabel pwell 187417 526210 187451 526244 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_8_Right_8.VNB
rlabel comment 187480 526227 187480 526227 8 dpga_flat_0.sr_0.PHY_EDGE_ROW_8_Right_8.decap_3
rlabel metal1 187204 526179 187480 526275 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_8_Right_8.VGND
rlabel metal1 187204 525635 187480 525731 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_8_Right_8.VPWR
flabel metal1 172513 525122 172547 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_3.VGND
flabel metal1 172513 525666 172547 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_3.VPWR
flabel nwell 172513 525666 172547 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_3.VPB
flabel pwell 172513 525122 172547 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_3.VNB
rlabel comment 172484 525139 172484 525139 4 dpga_flat_0.sr_0.FILLER_0_9_3.decap_12
flabel metal1 173617 525122 173651 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_15.VGND
flabel metal1 173617 525666 173651 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_15.VPWR
flabel nwell 173617 525666 173651 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_15.VPB
flabel pwell 173617 525122 173651 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_15.VNB
rlabel comment 173588 525139 173588 525139 4 dpga_flat_0.sr_0.FILLER_0_9_15.decap_12
flabel metal1 172237 525666 172271 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_9_Left_37.VPWR
flabel metal1 172237 525122 172271 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_9_Left_37.VGND
flabel nwell 172237 525666 172271 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_9_Left_37.VPB
flabel pwell 172237 525122 172271 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_9_Left_37.VNB
rlabel comment 172208 525139 172208 525139 4 dpga_flat_0.sr_0.PHY_EDGE_ROW_9_Left_37.decap_3
rlabel metal1 172208 525091 172484 525187 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_9_Left_37.VGND
rlabel metal1 172208 525635 172484 525731 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_9_Left_37.VPWR
flabel metal1 174721 525122 174755 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_27.VGND
flabel metal1 174721 525666 174755 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_27.VPWR
flabel nwell 174721 525666 174755 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_27.VPB
flabel pwell 174721 525122 174755 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_27.VNB
rlabel comment 174692 525139 174692 525139 4 dpga_flat_0.sr_0.FILLER_0_9_27.decap_12
flabel metal1 175825 525122 175859 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_39.VGND
flabel metal1 175825 525666 175859 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_39.VPWR
flabel nwell 175825 525666 175859 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_39.VPB
flabel pwell 175825 525122 175859 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_39.VNB
rlabel comment 175796 525139 175796 525139 4 dpga_flat_0.sr_0.FILLER_0_9_39.decap_12
flabel metal1 176929 525122 176963 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_51.VGND
flabel metal1 176929 525666 176963 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_51.VPWR
flabel nwell 176929 525666 176963 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_51.VPB
flabel pwell 176929 525122 176963 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_51.VNB
rlabel comment 176900 525139 176900 525139 4 dpga_flat_0.sr_0.FILLER_0_9_51.decap_4
rlabel metal1 176900 525091 177268 525187 1 dpga_flat_0.sr_0.FILLER_0_9_51.VGND
rlabel metal1 176900 525635 177268 525731 1 dpga_flat_0.sr_0.FILLER_0_9_51.VPWR
flabel metal1 177290 525666 177326 525696 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_55.VPWR
flabel metal1 177290 525126 177326 525155 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_55.VGND
flabel nwell 177299 525673 177319 525690 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_55.VPB
flabel pwell 177296 525128 177320 525150 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_55.VNB
rlabel comment 177268 525139 177268 525139 4 dpga_flat_0.sr_0.FILLER_0_9_55.fill_1
rlabel metal1 177268 525091 177360 525187 1 dpga_flat_0.sr_0.FILLER_0_9_55.VGND
rlabel metal1 177268 525635 177360 525731 1 dpga_flat_0.sr_0.FILLER_0_9_55.VPWR
flabel metal1 177481 525122 177515 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_57.VGND
flabel metal1 177481 525666 177515 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_57.VPWR
flabel nwell 177481 525666 177515 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_57.VPB
flabel pwell 177481 525122 177515 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_57.VNB
rlabel comment 177452 525139 177452 525139 4 dpga_flat_0.sr_0.FILLER_0_9_57.decap_12
flabel metal1 177382 525663 177435 525692 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_9_81.VPWR
flabel metal1 177381 525121 177432 525159 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_9_81.VGND
rlabel comment 177360 525139 177360 525139 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_9_81.tapvpwrvgnd_1
rlabel metal1 177360 525091 177452 525187 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_9_81.VGND
rlabel metal1 177360 525635 177452 525731 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_9_81.VPWR
flabel metal1 178585 525122 178619 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_69.VGND
flabel metal1 178585 525666 178619 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_69.VPWR
flabel nwell 178585 525666 178619 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_69.VPB
flabel pwell 178585 525122 178619 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_69.VNB
rlabel comment 178556 525139 178556 525139 4 dpga_flat_0.sr_0.FILLER_0_9_69.decap_12
flabel metal1 179689 525122 179723 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_81.VGND
flabel metal1 179689 525666 179723 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_81.VPWR
flabel nwell 179689 525666 179723 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_81.VPB
flabel pwell 179689 525122 179723 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_81.VNB
rlabel comment 179660 525139 179660 525139 4 dpga_flat_0.sr_0.FILLER_0_9_81.decap_12
flabel metal1 180793 525122 180827 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_93.VGND
flabel metal1 180793 525666 180827 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_93.VPWR
flabel nwell 180793 525666 180827 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_93.VPB
flabel pwell 180793 525122 180827 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_93.VNB
rlabel comment 180764 525139 180764 525139 4 dpga_flat_0.sr_0.FILLER_0_9_93.decap_12
flabel metal1 181897 525666 181931 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_105.VPWR
flabel metal1 181897 525122 181931 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_105.VGND
flabel nwell 181897 525666 181931 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_105.VPB
flabel pwell 181897 525122 181931 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_105.VNB
rlabel comment 181868 525139 181868 525139 4 dpga_flat_0.sr_0.FILLER_0_9_105.decap_6
rlabel metal1 181868 525091 182420 525187 1 dpga_flat_0.sr_0.FILLER_0_9_105.VGND
rlabel metal1 181868 525635 182420 525731 1 dpga_flat_0.sr_0.FILLER_0_9_105.VPWR
flabel metal1 182442 525666 182478 525696 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_111.VPWR
flabel metal1 182442 525126 182478 525155 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_111.VGND
flabel nwell 182451 525673 182471 525690 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_111.VPB
flabel pwell 182448 525128 182472 525150 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_111.VNB
rlabel comment 182420 525139 182420 525139 4 dpga_flat_0.sr_0.FILLER_0_9_111.fill_1
rlabel metal1 182420 525091 182512 525187 1 dpga_flat_0.sr_0.FILLER_0_9_111.VGND
rlabel metal1 182420 525635 182512 525731 1 dpga_flat_0.sr_0.FILLER_0_9_111.VPWR
flabel metal1 182633 525122 182667 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_113.VGND
flabel metal1 182633 525666 182667 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_113.VPWR
flabel nwell 182633 525666 182667 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_113.VPB
flabel pwell 182633 525122 182667 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_113.VNB
rlabel comment 182604 525139 182604 525139 4 dpga_flat_0.sr_0.FILLER_0_9_113.decap_12
flabel metal1 183737 525122 183771 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_125.VGND
flabel metal1 183737 525666 183771 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_125.VPWR
flabel nwell 183737 525666 183771 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_125.VPB
flabel pwell 183737 525122 183771 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_125.VNB
rlabel comment 183708 525139 183708 525139 4 dpga_flat_0.sr_0.FILLER_0_9_125.decap_12
flabel metal1 182534 525663 182587 525692 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_9_82.VPWR
flabel metal1 182533 525121 182584 525159 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_9_82.VGND
rlabel comment 182512 525139 182512 525139 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_9_82.tapvpwrvgnd_1
rlabel metal1 182512 525091 182604 525187 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_9_82.VGND
rlabel metal1 182512 525635 182604 525731 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_9_82.VPWR
flabel metal1 184841 525122 184875 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_137.VGND
flabel metal1 184841 525666 184875 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_137.VPWR
flabel nwell 184841 525666 184875 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_137.VPB
flabel pwell 184841 525122 184875 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_137.VNB
rlabel comment 184812 525139 184812 525139 4 dpga_flat_0.sr_0.FILLER_0_9_137.decap_12
flabel metal1 185945 525122 185979 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_149.VGND
flabel metal1 185945 525666 185979 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_149.VPWR
flabel nwell 185945 525666 185979 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_149.VPB
flabel pwell 185945 525122 185979 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_149.VNB
rlabel comment 185916 525139 185916 525139 4 dpga_flat_0.sr_0.FILLER_0_9_149.decap_12
flabel metal1 187040 525125 187093 525157 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_161.VGND
flabel metal1 187041 525669 187093 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_161.VPWR
flabel nwell 187048 525674 187082 525692 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_161.VPB
flabel pwell 187051 525129 187083 525151 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_161.VNB
rlabel comment 187020 525139 187020 525139 4 dpga_flat_0.sr_0.FILLER_0_9_161.fill_2
rlabel metal1 187020 525091 187204 525187 1 dpga_flat_0.sr_0.FILLER_0_9_161.VGND
rlabel metal1 187020 525635 187204 525731 1 dpga_flat_0.sr_0.FILLER_0_9_161.VPWR
flabel metal1 187417 525666 187451 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_9_Right_9.VPWR
flabel metal1 187417 525122 187451 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_9_Right_9.VGND
flabel nwell 187417 525666 187451 525700 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_9_Right_9.VPB
flabel pwell 187417 525122 187451 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_9_Right_9.VNB
rlabel comment 187480 525139 187480 525139 6 dpga_flat_0.sr_0.PHY_EDGE_ROW_9_Right_9.decap_3
rlabel metal1 187204 525091 187480 525187 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_9_Right_9.VGND
rlabel metal1 187204 525635 187480 525731 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_9_Right_9.VPWR
flabel metal1 172513 525122 172547 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_3.VGND
flabel metal1 172513 524578 172547 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_3.VPWR
flabel nwell 172513 524578 172547 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_3.VPB
flabel pwell 172513 525122 172547 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_3.VNB
rlabel comment 172484 525139 172484 525139 2 dpga_flat_0.sr_0.FILLER_0_10_3.decap_12
flabel metal1 173617 525122 173651 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_15.VGND
flabel metal1 173617 524578 173651 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_15.VPWR
flabel nwell 173617 524578 173651 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_15.VPB
flabel pwell 173617 525122 173651 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_15.VNB
rlabel comment 173588 525139 173588 525139 2 dpga_flat_0.sr_0.FILLER_0_10_15.decap_12
flabel metal1 172237 524578 172271 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_10_Left_38.VPWR
flabel metal1 172237 525122 172271 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_10_Left_38.VGND
flabel nwell 172237 524578 172271 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_10_Left_38.VPB
flabel pwell 172237 525122 172271 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_10_Left_38.VNB
rlabel comment 172208 525139 172208 525139 2 dpga_flat_0.sr_0.PHY_EDGE_ROW_10_Left_38.decap_3
rlabel metal1 172208 525091 172484 525187 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_10_Left_38.VGND
rlabel metal1 172208 524547 172484 524643 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_10_Left_38.VPWR
flabel metal1 174714 524582 174750 524612 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_27.VPWR
flabel metal1 174714 525123 174750 525152 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_27.VGND
flabel nwell 174723 524588 174743 524605 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_27.VPB
flabel pwell 174720 525128 174744 525150 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_27.VNB
rlabel comment 174692 525139 174692 525139 2 dpga_flat_0.sr_0.FILLER_0_10_27.fill_1
rlabel metal1 174692 525091 174784 525187 5 dpga_flat_0.sr_0.FILLER_0_10_27.VGND
rlabel metal1 174692 524547 174784 524643 5 dpga_flat_0.sr_0.FILLER_0_10_27.VPWR
flabel metal1 174905 525122 174939 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_29.VGND
flabel metal1 174905 524578 174939 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_29.VPWR
flabel nwell 174905 524578 174939 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_29.VPB
flabel pwell 174905 525122 174939 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_29.VNB
rlabel comment 174876 525139 174876 525139 2 dpga_flat_0.sr_0.FILLER_0_10_29.decap_12
flabel metal1 176009 525122 176043 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_41.VGND
flabel metal1 176009 524578 176043 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_41.VPWR
flabel nwell 176009 524578 176043 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_41.VPB
flabel pwell 176009 525122 176043 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_41.VNB
rlabel comment 175980 525139 175980 525139 2 dpga_flat_0.sr_0.FILLER_0_10_41.decap_12
flabel metal1 174806 524586 174859 524615 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_10_83.VPWR
flabel metal1 174805 525119 174856 525157 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_10_83.VGND
rlabel comment 174784 525139 174784 525139 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_10_83.tapvpwrvgnd_1
rlabel metal1 174784 525091 174876 525187 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_10_83.VGND
rlabel metal1 174784 524547 174876 524643 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_10_83.VPWR
flabel metal1 177113 525122 177147 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_53.VGND
flabel metal1 177113 524578 177147 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_53.VPWR
flabel nwell 177113 524578 177147 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_53.VPB
flabel pwell 177113 525122 177147 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_53.VNB
rlabel comment 177084 525139 177084 525139 2 dpga_flat_0.sr_0.FILLER_0_10_53.decap_12
flabel metal1 178217 525122 178251 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_65.VGND
flabel metal1 178217 524578 178251 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_65.VPWR
flabel nwell 178217 524578 178251 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_65.VPB
flabel pwell 178217 525122 178251 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_65.VNB
rlabel comment 178188 525139 178188 525139 2 dpga_flat_0.sr_0.FILLER_0_10_65.decap_12
flabel metal1 179321 524578 179355 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_77.VPWR
flabel metal1 179321 525122 179355 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_77.VGND
flabel nwell 179321 524578 179355 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_77.VPB
flabel pwell 179321 525122 179355 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_77.VNB
rlabel comment 179292 525139 179292 525139 2 dpga_flat_0.sr_0.FILLER_0_10_77.decap_6
rlabel metal1 179292 525091 179844 525187 5 dpga_flat_0.sr_0.FILLER_0_10_77.VGND
rlabel metal1 179292 524547 179844 524643 5 dpga_flat_0.sr_0.FILLER_0_10_77.VPWR
flabel metal1 179866 524582 179902 524612 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_83.VPWR
flabel metal1 179866 525123 179902 525152 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_83.VGND
flabel nwell 179875 524588 179895 524605 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_83.VPB
flabel pwell 179872 525128 179896 525150 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_83.VNB
rlabel comment 179844 525139 179844 525139 2 dpga_flat_0.sr_0.FILLER_0_10_83.fill_1
rlabel metal1 179844 525091 179936 525187 5 dpga_flat_0.sr_0.FILLER_0_10_83.VGND
rlabel metal1 179844 524547 179936 524643 5 dpga_flat_0.sr_0.FILLER_0_10_83.VPWR
flabel metal1 180057 525122 180091 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_85.VGND
flabel metal1 180057 524578 180091 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_85.VPWR
flabel nwell 180057 524578 180091 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_85.VPB
flabel pwell 180057 525122 180091 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_85.VNB
rlabel comment 180028 525139 180028 525139 2 dpga_flat_0.sr_0.FILLER_0_10_85.decap_12
flabel metal1 181161 525122 181195 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_97.VGND
flabel metal1 181161 524578 181195 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_97.VPWR
flabel nwell 181161 524578 181195 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_97.VPB
flabel pwell 181161 525122 181195 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_97.VNB
rlabel comment 181132 525139 181132 525139 2 dpga_flat_0.sr_0.FILLER_0_10_97.decap_12
flabel metal1 179958 524586 180011 524615 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_10_84.VPWR
flabel metal1 179957 525119 180008 525157 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_10_84.VGND
rlabel comment 179936 525139 179936 525139 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_10_84.tapvpwrvgnd_1
rlabel metal1 179936 525091 180028 525187 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_10_84.VGND
rlabel metal1 179936 524547 180028 524643 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_10_84.VPWR
flabel metal1 182265 525122 182299 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_109.VGND
flabel metal1 182265 524578 182299 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_109.VPWR
flabel nwell 182265 524578 182299 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_109.VPB
flabel pwell 182265 525122 182299 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_109.VNB
rlabel comment 182236 525139 182236 525139 2 dpga_flat_0.sr_0.FILLER_0_10_109.decap_12
flabel metal1 183369 525122 183403 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_121.VGND
flabel metal1 183369 524578 183403 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_121.VPWR
flabel nwell 183369 524578 183403 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_121.VPB
flabel pwell 183369 525122 183403 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_121.VNB
rlabel comment 183340 525139 183340 525139 2 dpga_flat_0.sr_0.FILLER_0_10_121.decap_12
flabel metal1 184473 524578 184507 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_133.VPWR
flabel metal1 184473 525122 184507 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_133.VGND
flabel nwell 184473 524578 184507 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_133.VPB
flabel pwell 184473 525122 184507 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_133.VNB
rlabel comment 184444 525139 184444 525139 2 dpga_flat_0.sr_0.FILLER_0_10_133.decap_6
rlabel metal1 184444 525091 184996 525187 5 dpga_flat_0.sr_0.FILLER_0_10_133.VGND
rlabel metal1 184444 524547 184996 524643 5 dpga_flat_0.sr_0.FILLER_0_10_133.VPWR
flabel metal1 185018 524582 185054 524612 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_139.VPWR
flabel metal1 185018 525123 185054 525152 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_139.VGND
flabel nwell 185027 524588 185047 524605 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_139.VPB
flabel pwell 185024 525128 185048 525150 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_139.VNB
rlabel comment 184996 525139 184996 525139 2 dpga_flat_0.sr_0.FILLER_0_10_139.fill_1
rlabel metal1 184996 525091 185088 525187 5 dpga_flat_0.sr_0.FILLER_0_10_139.VGND
rlabel metal1 184996 524547 185088 524643 5 dpga_flat_0.sr_0.FILLER_0_10_139.VPWR
flabel metal1 185209 525122 185243 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_141.VGND
flabel metal1 185209 524578 185243 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_141.VPWR
flabel nwell 185209 524578 185243 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_141.VPB
flabel pwell 185209 525122 185243 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_141.VNB
rlabel comment 185180 525139 185180 525139 2 dpga_flat_0.sr_0.FILLER_0_10_141.decap_12
flabel metal1 185110 524586 185163 524615 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_10_85.VPWR
flabel metal1 185109 525119 185160 525157 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_10_85.VGND
rlabel comment 185088 525139 185088 525139 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_10_85.tapvpwrvgnd_1
rlabel metal1 185088 525091 185180 525187 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_10_85.VGND
rlabel metal1 185088 524547 185180 524643 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_10_85.VPWR
flabel metal1 186313 524578 186347 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_153.VPWR
flabel metal1 186313 525122 186347 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_153.VGND
flabel nwell 186313 524578 186347 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_153.VPB
flabel pwell 186313 525122 186347 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_153.VNB
rlabel comment 186284 525139 186284 525139 2 dpga_flat_0.sr_0.FILLER_0_10_153.decap_8
rlabel metal1 186284 525091 187020 525187 5 dpga_flat_0.sr_0.FILLER_0_10_153.VGND
rlabel metal1 186284 524547 187020 524643 5 dpga_flat_0.sr_0.FILLER_0_10_153.VPWR
flabel metal1 187040 525121 187093 525153 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_161.VGND
flabel metal1 187041 524578 187093 524609 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_161.VPWR
flabel nwell 187048 524586 187082 524604 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_161.VPB
flabel pwell 187051 525127 187083 525149 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_161.VNB
rlabel comment 187020 525139 187020 525139 2 dpga_flat_0.sr_0.FILLER_0_10_161.fill_2
rlabel metal1 187020 525091 187204 525187 5 dpga_flat_0.sr_0.FILLER_0_10_161.VGND
rlabel metal1 187020 524547 187204 524643 5 dpga_flat_0.sr_0.FILLER_0_10_161.VPWR
flabel metal1 187417 524578 187451 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_10_Right_10.VPWR
flabel metal1 187417 525122 187451 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_10_Right_10.VGND
flabel nwell 187417 524578 187451 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_10_Right_10.VPB
flabel pwell 187417 525122 187451 525156 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_10_Right_10.VNB
rlabel comment 187480 525139 187480 525139 8 dpga_flat_0.sr_0.PHY_EDGE_ROW_10_Right_10.decap_3
rlabel metal1 187204 525091 187480 525187 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_10_Right_10.VGND
rlabel metal1 187204 524547 187480 524643 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_10_Right_10.VPWR
flabel metal1 172513 524034 172547 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_3.VGND
flabel metal1 172513 524578 172547 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_3.VPWR
flabel nwell 172513 524578 172547 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_3.VPB
flabel pwell 172513 524034 172547 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_3.VNB
rlabel comment 172484 524051 172484 524051 4 dpga_flat_0.sr_0.FILLER_0_11_3.decap_12
flabel metal1 173617 524034 173651 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_15.VGND
flabel metal1 173617 524578 173651 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_15.VPWR
flabel nwell 173617 524578 173651 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_15.VPB
flabel pwell 173617 524034 173651 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_15.VNB
rlabel comment 173588 524051 173588 524051 4 dpga_flat_0.sr_0.FILLER_0_11_15.decap_12
flabel metal1 172237 524578 172271 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_11_Left_39.VPWR
flabel metal1 172237 524034 172271 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_11_Left_39.VGND
flabel nwell 172237 524578 172271 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_11_Left_39.VPB
flabel pwell 172237 524034 172271 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_11_Left_39.VNB
rlabel comment 172208 524051 172208 524051 4 dpga_flat_0.sr_0.PHY_EDGE_ROW_11_Left_39.decap_3
rlabel metal1 172208 524003 172484 524099 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_11_Left_39.VGND
rlabel metal1 172208 524547 172484 524643 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_11_Left_39.VPWR
flabel metal1 174721 524034 174755 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_27.VGND
flabel metal1 174721 524578 174755 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_27.VPWR
flabel nwell 174721 524578 174755 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_27.VPB
flabel pwell 174721 524034 174755 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_27.VNB
rlabel comment 174692 524051 174692 524051 4 dpga_flat_0.sr_0.FILLER_0_11_27.decap_12
flabel metal1 175825 524034 175859 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_39.VGND
flabel metal1 175825 524578 175859 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_39.VPWR
flabel nwell 175825 524578 175859 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_39.VPB
flabel pwell 175825 524034 175859 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_39.VNB
rlabel comment 175796 524051 175796 524051 4 dpga_flat_0.sr_0.FILLER_0_11_39.decap_12
flabel metal1 176929 524034 176963 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_51.VGND
flabel metal1 176929 524578 176963 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_51.VPWR
flabel nwell 176929 524578 176963 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_51.VPB
flabel pwell 176929 524034 176963 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_51.VNB
rlabel comment 176900 524051 176900 524051 4 dpga_flat_0.sr_0.FILLER_0_11_51.decap_4
rlabel metal1 176900 524003 177268 524099 1 dpga_flat_0.sr_0.FILLER_0_11_51.VGND
rlabel metal1 176900 524547 177268 524643 1 dpga_flat_0.sr_0.FILLER_0_11_51.VPWR
flabel metal1 177290 524578 177326 524608 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_55.VPWR
flabel metal1 177290 524038 177326 524067 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_55.VGND
flabel nwell 177299 524585 177319 524602 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_55.VPB
flabel pwell 177296 524040 177320 524062 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_55.VNB
rlabel comment 177268 524051 177268 524051 4 dpga_flat_0.sr_0.FILLER_0_11_55.fill_1
rlabel metal1 177268 524003 177360 524099 1 dpga_flat_0.sr_0.FILLER_0_11_55.VGND
rlabel metal1 177268 524547 177360 524643 1 dpga_flat_0.sr_0.FILLER_0_11_55.VPWR
flabel metal1 177481 524034 177515 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_57.VGND
flabel metal1 177481 524578 177515 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_57.VPWR
flabel nwell 177481 524578 177515 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_57.VPB
flabel pwell 177481 524034 177515 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_57.VNB
rlabel comment 177452 524051 177452 524051 4 dpga_flat_0.sr_0.FILLER_0_11_57.decap_12
flabel metal1 177382 524575 177435 524604 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_11_86.VPWR
flabel metal1 177381 524033 177432 524071 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_11_86.VGND
rlabel comment 177360 524051 177360 524051 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_11_86.tapvpwrvgnd_1
rlabel metal1 177360 524003 177452 524099 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_11_86.VGND
rlabel metal1 177360 524547 177452 524643 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_11_86.VPWR
flabel metal1 178585 524034 178619 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_69.VGND
flabel metal1 178585 524578 178619 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_69.VPWR
flabel nwell 178585 524578 178619 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_69.VPB
flabel pwell 178585 524034 178619 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_69.VNB
rlabel comment 178556 524051 178556 524051 4 dpga_flat_0.sr_0.FILLER_0_11_69.decap_12
flabel metal1 179689 524034 179723 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_81.VGND
flabel metal1 179689 524578 179723 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_81.VPWR
flabel nwell 179689 524578 179723 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_81.VPB
flabel pwell 179689 524034 179723 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_81.VNB
rlabel comment 179660 524051 179660 524051 4 dpga_flat_0.sr_0.FILLER_0_11_81.decap_12
flabel metal1 180793 524034 180827 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_93.VGND
flabel metal1 180793 524578 180827 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_93.VPWR
flabel nwell 180793 524578 180827 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_93.VPB
flabel pwell 180793 524034 180827 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_93.VNB
rlabel comment 180764 524051 180764 524051 4 dpga_flat_0.sr_0.FILLER_0_11_93.decap_12
flabel metal1 181897 524578 181931 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_105.VPWR
flabel metal1 181897 524034 181931 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_105.VGND
flabel nwell 181897 524578 181931 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_105.VPB
flabel pwell 181897 524034 181931 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_105.VNB
rlabel comment 181868 524051 181868 524051 4 dpga_flat_0.sr_0.FILLER_0_11_105.decap_6
rlabel metal1 181868 524003 182420 524099 1 dpga_flat_0.sr_0.FILLER_0_11_105.VGND
rlabel metal1 181868 524547 182420 524643 1 dpga_flat_0.sr_0.FILLER_0_11_105.VPWR
flabel metal1 182442 524578 182478 524608 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_111.VPWR
flabel metal1 182442 524038 182478 524067 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_111.VGND
flabel nwell 182451 524585 182471 524602 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_111.VPB
flabel pwell 182448 524040 182472 524062 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_111.VNB
rlabel comment 182420 524051 182420 524051 4 dpga_flat_0.sr_0.FILLER_0_11_111.fill_1
rlabel metal1 182420 524003 182512 524099 1 dpga_flat_0.sr_0.FILLER_0_11_111.VGND
rlabel metal1 182420 524547 182512 524643 1 dpga_flat_0.sr_0.FILLER_0_11_111.VPWR
flabel metal1 182633 524034 182667 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_113.VGND
flabel metal1 182633 524578 182667 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_113.VPWR
flabel nwell 182633 524578 182667 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_113.VPB
flabel pwell 182633 524034 182667 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_113.VNB
rlabel comment 182604 524051 182604 524051 4 dpga_flat_0.sr_0.FILLER_0_11_113.decap_12
flabel metal1 183737 524034 183771 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_125.VGND
flabel metal1 183737 524578 183771 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_125.VPWR
flabel nwell 183737 524578 183771 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_125.VPB
flabel pwell 183737 524034 183771 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_125.VNB
rlabel comment 183708 524051 183708 524051 4 dpga_flat_0.sr_0.FILLER_0_11_125.decap_12
flabel metal1 182534 524575 182587 524604 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_11_87.VPWR
flabel metal1 182533 524033 182584 524071 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_11_87.VGND
rlabel comment 182512 524051 182512 524051 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_11_87.tapvpwrvgnd_1
rlabel metal1 182512 524003 182604 524099 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_11_87.VGND
rlabel metal1 182512 524547 182604 524643 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_11_87.VPWR
flabel metal1 184841 524034 184875 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_137.VGND
flabel metal1 184841 524578 184875 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_137.VPWR
flabel nwell 184841 524578 184875 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_137.VPB
flabel pwell 184841 524034 184875 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_137.VNB
rlabel comment 184812 524051 184812 524051 4 dpga_flat_0.sr_0.FILLER_0_11_137.decap_12
flabel metal1 185945 524034 185979 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_149.VGND
flabel metal1 185945 524578 185979 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_149.VPWR
flabel nwell 185945 524578 185979 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_149.VPB
flabel pwell 185945 524034 185979 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_149.VNB
rlabel comment 185916 524051 185916 524051 4 dpga_flat_0.sr_0.FILLER_0_11_149.decap_12
flabel metal1 187040 524037 187093 524069 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_161.VGND
flabel metal1 187041 524581 187093 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_161.VPWR
flabel nwell 187048 524586 187082 524604 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_161.VPB
flabel pwell 187051 524041 187083 524063 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_161.VNB
rlabel comment 187020 524051 187020 524051 4 dpga_flat_0.sr_0.FILLER_0_11_161.fill_2
rlabel metal1 187020 524003 187204 524099 1 dpga_flat_0.sr_0.FILLER_0_11_161.VGND
rlabel metal1 187020 524547 187204 524643 1 dpga_flat_0.sr_0.FILLER_0_11_161.VPWR
flabel metal1 187417 524578 187451 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_11_Right_11.VPWR
flabel metal1 187417 524034 187451 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_11_Right_11.VGND
flabel nwell 187417 524578 187451 524612 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_11_Right_11.VPB
flabel pwell 187417 524034 187451 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_11_Right_11.VNB
rlabel comment 187480 524051 187480 524051 6 dpga_flat_0.sr_0.PHY_EDGE_ROW_11_Right_11.decap_3
rlabel metal1 187204 524003 187480 524099 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_11_Right_11.VGND
rlabel metal1 187204 524547 187480 524643 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_11_Right_11.VPWR
flabel metal1 172513 524034 172547 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_3.VGND
flabel metal1 172513 523490 172547 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_3.VPWR
flabel nwell 172513 523490 172547 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_3.VPB
flabel pwell 172513 524034 172547 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_3.VNB
rlabel comment 172484 524051 172484 524051 2 dpga_flat_0.sr_0.FILLER_0_12_3.decap_12
flabel metal1 173617 524034 173651 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_15.VGND
flabel metal1 173617 523490 173651 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_15.VPWR
flabel nwell 173617 523490 173651 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_15.VPB
flabel pwell 173617 524034 173651 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_15.VNB
rlabel comment 173588 524051 173588 524051 2 dpga_flat_0.sr_0.FILLER_0_12_15.decap_12
flabel metal1 172237 523490 172271 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_12_Left_40.VPWR
flabel metal1 172237 524034 172271 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_12_Left_40.VGND
flabel nwell 172237 523490 172271 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_12_Left_40.VPB
flabel pwell 172237 524034 172271 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_12_Left_40.VNB
rlabel comment 172208 524051 172208 524051 2 dpga_flat_0.sr_0.PHY_EDGE_ROW_12_Left_40.decap_3
rlabel metal1 172208 524003 172484 524099 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_12_Left_40.VGND
rlabel metal1 172208 523459 172484 523555 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_12_Left_40.VPWR
flabel metal1 174714 523494 174750 523524 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_27.VPWR
flabel metal1 174714 524035 174750 524064 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_27.VGND
flabel nwell 174723 523500 174743 523517 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_27.VPB
flabel pwell 174720 524040 174744 524062 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_27.VNB
rlabel comment 174692 524051 174692 524051 2 dpga_flat_0.sr_0.FILLER_0_12_27.fill_1
rlabel metal1 174692 524003 174784 524099 5 dpga_flat_0.sr_0.FILLER_0_12_27.VGND
rlabel metal1 174692 523459 174784 523555 5 dpga_flat_0.sr_0.FILLER_0_12_27.VPWR
flabel metal1 174905 524034 174939 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_29.VGND
flabel metal1 174905 523490 174939 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_29.VPWR
flabel nwell 174905 523490 174939 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_29.VPB
flabel pwell 174905 524034 174939 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_29.VNB
rlabel comment 174876 524051 174876 524051 2 dpga_flat_0.sr_0.FILLER_0_12_29.decap_12
flabel metal1 176009 524034 176043 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_41.VGND
flabel metal1 176009 523490 176043 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_41.VPWR
flabel nwell 176009 523490 176043 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_41.VPB
flabel pwell 176009 524034 176043 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_41.VNB
rlabel comment 175980 524051 175980 524051 2 dpga_flat_0.sr_0.FILLER_0_12_41.decap_12
flabel metal1 174806 523498 174859 523527 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_12_88.VPWR
flabel metal1 174805 524031 174856 524069 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_12_88.VGND
rlabel comment 174784 524051 174784 524051 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_12_88.tapvpwrvgnd_1
rlabel metal1 174784 524003 174876 524099 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_12_88.VGND
rlabel metal1 174784 523459 174876 523555 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_12_88.VPWR
flabel metal1 177113 524034 177147 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_53.VGND
flabel metal1 177113 523490 177147 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_53.VPWR
flabel nwell 177113 523490 177147 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_53.VPB
flabel pwell 177113 524034 177147 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_53.VNB
rlabel comment 177084 524051 177084 524051 2 dpga_flat_0.sr_0.FILLER_0_12_53.decap_12
flabel metal1 178217 524034 178251 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_65.VGND
flabel metal1 178217 523490 178251 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_65.VPWR
flabel nwell 178217 523490 178251 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_65.VPB
flabel pwell 178217 524034 178251 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_65.VNB
rlabel comment 178188 524051 178188 524051 2 dpga_flat_0.sr_0.FILLER_0_12_65.decap_12
flabel metal1 179321 523490 179355 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_77.VPWR
flabel metal1 179321 524034 179355 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_77.VGND
flabel nwell 179321 523490 179355 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_77.VPB
flabel pwell 179321 524034 179355 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_77.VNB
rlabel comment 179292 524051 179292 524051 2 dpga_flat_0.sr_0.FILLER_0_12_77.decap_6
rlabel metal1 179292 524003 179844 524099 5 dpga_flat_0.sr_0.FILLER_0_12_77.VGND
rlabel metal1 179292 523459 179844 523555 5 dpga_flat_0.sr_0.FILLER_0_12_77.VPWR
flabel metal1 179866 523494 179902 523524 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_83.VPWR
flabel metal1 179866 524035 179902 524064 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_83.VGND
flabel nwell 179875 523500 179895 523517 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_83.VPB
flabel pwell 179872 524040 179896 524062 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_83.VNB
rlabel comment 179844 524051 179844 524051 2 dpga_flat_0.sr_0.FILLER_0_12_83.fill_1
rlabel metal1 179844 524003 179936 524099 5 dpga_flat_0.sr_0.FILLER_0_12_83.VGND
rlabel metal1 179844 523459 179936 523555 5 dpga_flat_0.sr_0.FILLER_0_12_83.VPWR
flabel metal1 180057 524034 180091 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_85.VGND
flabel metal1 180057 523490 180091 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_85.VPWR
flabel nwell 180057 523490 180091 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_85.VPB
flabel pwell 180057 524034 180091 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_85.VNB
rlabel comment 180028 524051 180028 524051 2 dpga_flat_0.sr_0.FILLER_0_12_85.decap_12
flabel metal1 181161 524034 181195 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_97.VGND
flabel metal1 181161 523490 181195 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_97.VPWR
flabel nwell 181161 523490 181195 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_97.VPB
flabel pwell 181161 524034 181195 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_97.VNB
rlabel comment 181132 524051 181132 524051 2 dpga_flat_0.sr_0.FILLER_0_12_97.decap_12
flabel metal1 179958 523498 180011 523527 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_12_89.VPWR
flabel metal1 179957 524031 180008 524069 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_12_89.VGND
rlabel comment 179936 524051 179936 524051 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_12_89.tapvpwrvgnd_1
rlabel metal1 179936 524003 180028 524099 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_12_89.VGND
rlabel metal1 179936 523459 180028 523555 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_12_89.VPWR
flabel metal1 182265 524034 182299 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_109.VGND
flabel metal1 182265 523490 182299 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_109.VPWR
flabel nwell 182265 523490 182299 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_109.VPB
flabel pwell 182265 524034 182299 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_109.VNB
rlabel comment 182236 524051 182236 524051 2 dpga_flat_0.sr_0.FILLER_0_12_109.decap_12
flabel metal1 183369 524034 183403 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_121.VGND
flabel metal1 183369 523490 183403 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_121.VPWR
flabel nwell 183369 523490 183403 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_121.VPB
flabel pwell 183369 524034 183403 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_121.VNB
rlabel comment 183340 524051 183340 524051 2 dpga_flat_0.sr_0.FILLER_0_12_121.decap_12
flabel metal1 184473 523490 184507 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_133.VPWR
flabel metal1 184473 524034 184507 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_133.VGND
flabel nwell 184473 523490 184507 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_133.VPB
flabel pwell 184473 524034 184507 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_133.VNB
rlabel comment 184444 524051 184444 524051 2 dpga_flat_0.sr_0.FILLER_0_12_133.decap_6
rlabel metal1 184444 524003 184996 524099 5 dpga_flat_0.sr_0.FILLER_0_12_133.VGND
rlabel metal1 184444 523459 184996 523555 5 dpga_flat_0.sr_0.FILLER_0_12_133.VPWR
flabel metal1 185018 523494 185054 523524 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_139.VPWR
flabel metal1 185018 524035 185054 524064 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_139.VGND
flabel nwell 185027 523500 185047 523517 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_139.VPB
flabel pwell 185024 524040 185048 524062 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_139.VNB
rlabel comment 184996 524051 184996 524051 2 dpga_flat_0.sr_0.FILLER_0_12_139.fill_1
rlabel metal1 184996 524003 185088 524099 5 dpga_flat_0.sr_0.FILLER_0_12_139.VGND
rlabel metal1 184996 523459 185088 523555 5 dpga_flat_0.sr_0.FILLER_0_12_139.VPWR
flabel metal1 185209 524034 185243 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_141.VGND
flabel metal1 185209 523490 185243 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_141.VPWR
flabel nwell 185209 523490 185243 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_141.VPB
flabel pwell 185209 524034 185243 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_141.VNB
rlabel comment 185180 524051 185180 524051 2 dpga_flat_0.sr_0.FILLER_0_12_141.decap_12
flabel metal1 185110 523498 185163 523527 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_12_90.VPWR
flabel metal1 185109 524031 185160 524069 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_12_90.VGND
rlabel comment 185088 524051 185088 524051 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_12_90.tapvpwrvgnd_1
rlabel metal1 185088 524003 185180 524099 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_12_90.VGND
rlabel metal1 185088 523459 185180 523555 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_12_90.VPWR
flabel metal1 186313 523490 186347 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_153.VPWR
flabel metal1 186313 524034 186347 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_153.VGND
flabel nwell 186313 523490 186347 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_153.VPB
flabel pwell 186313 524034 186347 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_153.VNB
rlabel comment 186284 524051 186284 524051 2 dpga_flat_0.sr_0.FILLER_0_12_153.decap_8
rlabel metal1 186284 524003 187020 524099 5 dpga_flat_0.sr_0.FILLER_0_12_153.VGND
rlabel metal1 186284 523459 187020 523555 5 dpga_flat_0.sr_0.FILLER_0_12_153.VPWR
flabel metal1 187040 524033 187093 524065 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_161.VGND
flabel metal1 187041 523490 187093 523521 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_161.VPWR
flabel nwell 187048 523498 187082 523516 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_161.VPB
flabel pwell 187051 524039 187083 524061 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_161.VNB
rlabel comment 187020 524051 187020 524051 2 dpga_flat_0.sr_0.FILLER_0_12_161.fill_2
rlabel metal1 187020 524003 187204 524099 5 dpga_flat_0.sr_0.FILLER_0_12_161.VGND
rlabel metal1 187020 523459 187204 523555 5 dpga_flat_0.sr_0.FILLER_0_12_161.VPWR
flabel metal1 187417 523490 187451 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_12_Right_12.VPWR
flabel metal1 187417 524034 187451 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_12_Right_12.VGND
flabel nwell 187417 523490 187451 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_12_Right_12.VPB
flabel pwell 187417 524034 187451 524068 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_12_Right_12.VNB
rlabel comment 187480 524051 187480 524051 8 dpga_flat_0.sr_0.PHY_EDGE_ROW_12_Right_12.decap_3
rlabel metal1 187204 524003 187480 524099 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_12_Right_12.VGND
rlabel metal1 187204 523459 187480 523555 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_12_Right_12.VPWR
flabel metal1 172513 522946 172547 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_3.VGND
flabel metal1 172513 523490 172547 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_3.VPWR
flabel nwell 172513 523490 172547 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_3.VPB
flabel pwell 172513 522946 172547 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_3.VNB
rlabel comment 172484 522963 172484 522963 4 dpga_flat_0.sr_0.FILLER_0_13_3.decap_12
flabel metal1 173617 522946 173651 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_15.VGND
flabel metal1 173617 523490 173651 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_15.VPWR
flabel nwell 173617 523490 173651 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_15.VPB
flabel pwell 173617 522946 173651 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_15.VNB
rlabel comment 173588 522963 173588 522963 4 dpga_flat_0.sr_0.FILLER_0_13_15.decap_12
flabel metal1 172513 522946 172547 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_3.VGND
flabel metal1 172513 522402 172547 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_3.VPWR
flabel nwell 172513 522402 172547 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_3.VPB
flabel pwell 172513 522946 172547 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_3.VNB
rlabel comment 172484 522963 172484 522963 2 dpga_flat_0.sr_0.FILLER_0_14_3.decap_12
flabel metal1 173617 522946 173651 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_15.VGND
flabel metal1 173617 522402 173651 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_15.VPWR
flabel nwell 173617 522402 173651 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_15.VPB
flabel pwell 173617 522946 173651 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_15.VNB
rlabel comment 173588 522963 173588 522963 2 dpga_flat_0.sr_0.FILLER_0_14_15.decap_12
flabel metal1 172237 523490 172271 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_13_Left_41.VPWR
flabel metal1 172237 522946 172271 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_13_Left_41.VGND
flabel nwell 172237 523490 172271 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_13_Left_41.VPB
flabel pwell 172237 522946 172271 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_13_Left_41.VNB
rlabel comment 172208 522963 172208 522963 4 dpga_flat_0.sr_0.PHY_EDGE_ROW_13_Left_41.decap_3
rlabel metal1 172208 522915 172484 523011 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_13_Left_41.VGND
rlabel metal1 172208 523459 172484 523555 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_13_Left_41.VPWR
flabel metal1 172237 522402 172271 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_14_Left_42.VPWR
flabel metal1 172237 522946 172271 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_14_Left_42.VGND
flabel nwell 172237 522402 172271 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_14_Left_42.VPB
flabel pwell 172237 522946 172271 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_14_Left_42.VNB
rlabel comment 172208 522963 172208 522963 2 dpga_flat_0.sr_0.PHY_EDGE_ROW_14_Left_42.decap_3
rlabel metal1 172208 522915 172484 523011 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_14_Left_42.VGND
rlabel metal1 172208 522371 172484 522467 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_14_Left_42.VPWR
flabel metal1 174721 522946 174755 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_27.VGND
flabel metal1 174721 523490 174755 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_27.VPWR
flabel nwell 174721 523490 174755 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_27.VPB
flabel pwell 174721 522946 174755 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_27.VNB
rlabel comment 174692 522963 174692 522963 4 dpga_flat_0.sr_0.FILLER_0_13_27.decap_12
flabel metal1 175825 522946 175859 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_39.VGND
flabel metal1 175825 523490 175859 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_39.VPWR
flabel nwell 175825 523490 175859 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_39.VPB
flabel pwell 175825 522946 175859 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_39.VNB
rlabel comment 175796 522963 175796 522963 4 dpga_flat_0.sr_0.FILLER_0_13_39.decap_12
flabel metal1 174714 522406 174750 522436 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_27.VPWR
flabel metal1 174714 522947 174750 522976 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_27.VGND
flabel nwell 174723 522412 174743 522429 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_27.VPB
flabel pwell 174720 522952 174744 522974 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_27.VNB
rlabel comment 174692 522963 174692 522963 2 dpga_flat_0.sr_0.FILLER_0_14_27.fill_1
rlabel metal1 174692 522915 174784 523011 5 dpga_flat_0.sr_0.FILLER_0_14_27.VGND
rlabel metal1 174692 522371 174784 522467 5 dpga_flat_0.sr_0.FILLER_0_14_27.VPWR
flabel metal1 174905 522946 174939 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_29.VGND
flabel metal1 174905 522402 174939 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_29.VPWR
flabel nwell 174905 522402 174939 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_29.VPB
flabel pwell 174905 522946 174939 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_29.VNB
rlabel comment 174876 522963 174876 522963 2 dpga_flat_0.sr_0.FILLER_0_14_29.decap_12
flabel metal1 176009 522946 176043 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_41.VGND
flabel metal1 176009 522402 176043 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_41.VPWR
flabel nwell 176009 522402 176043 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_41.VPB
flabel pwell 176009 522946 176043 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_41.VNB
rlabel comment 175980 522963 175980 522963 2 dpga_flat_0.sr_0.FILLER_0_14_41.decap_12
flabel metal1 174806 522410 174859 522439 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_14_93.VPWR
flabel metal1 174805 522943 174856 522981 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_14_93.VGND
rlabel comment 174784 522963 174784 522963 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_14_93.tapvpwrvgnd_1
rlabel metal1 174784 522915 174876 523011 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_14_93.VGND
rlabel metal1 174784 522371 174876 522467 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_14_93.VPWR
flabel metal1 176929 522946 176963 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_51.VGND
flabel metal1 176929 523490 176963 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_51.VPWR
flabel nwell 176929 523490 176963 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_51.VPB
flabel pwell 176929 522946 176963 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_51.VNB
rlabel comment 176900 522963 176900 522963 4 dpga_flat_0.sr_0.FILLER_0_13_51.decap_4
rlabel metal1 176900 522915 177268 523011 1 dpga_flat_0.sr_0.FILLER_0_13_51.VGND
rlabel metal1 176900 523459 177268 523555 1 dpga_flat_0.sr_0.FILLER_0_13_51.VPWR
flabel metal1 177290 523490 177326 523520 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_55.VPWR
flabel metal1 177290 522950 177326 522979 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_55.VGND
flabel nwell 177299 523497 177319 523514 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_55.VPB
flabel pwell 177296 522952 177320 522974 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_55.VNB
rlabel comment 177268 522963 177268 522963 4 dpga_flat_0.sr_0.FILLER_0_13_55.fill_1
rlabel metal1 177268 522915 177360 523011 1 dpga_flat_0.sr_0.FILLER_0_13_55.VGND
rlabel metal1 177268 523459 177360 523555 1 dpga_flat_0.sr_0.FILLER_0_13_55.VPWR
flabel metal1 177481 522946 177515 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_57.VGND
flabel metal1 177481 523490 177515 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_57.VPWR
flabel nwell 177481 523490 177515 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_57.VPB
flabel pwell 177481 522946 177515 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_57.VNB
rlabel comment 177452 522963 177452 522963 4 dpga_flat_0.sr_0.FILLER_0_13_57.decap_12
flabel metal1 177113 522946 177147 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_53.VGND
flabel metal1 177113 522402 177147 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_53.VPWR
flabel nwell 177113 522402 177147 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_53.VPB
flabel pwell 177113 522946 177147 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_53.VNB
rlabel comment 177084 522963 177084 522963 2 dpga_flat_0.sr_0.FILLER_0_14_53.decap_12
flabel metal1 177382 523487 177435 523516 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_13_91.VPWR
flabel metal1 177381 522945 177432 522983 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_13_91.VGND
rlabel comment 177360 522963 177360 522963 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_13_91.tapvpwrvgnd_1
rlabel metal1 177360 522915 177452 523011 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_13_91.VGND
rlabel metal1 177360 523459 177452 523555 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_13_91.VPWR
flabel metal1 178585 522946 178619 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_69.VGND
flabel metal1 178585 523490 178619 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_69.VPWR
flabel nwell 178585 523490 178619 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_69.VPB
flabel pwell 178585 522946 178619 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_69.VNB
rlabel comment 178556 522963 178556 522963 4 dpga_flat_0.sr_0.FILLER_0_13_69.decap_12
flabel metal1 179689 522946 179723 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_81.VGND
flabel metal1 179689 523490 179723 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_81.VPWR
flabel nwell 179689 523490 179723 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_81.VPB
flabel pwell 179689 522946 179723 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_81.VNB
rlabel comment 179660 522963 179660 522963 4 dpga_flat_0.sr_0.FILLER_0_13_81.decap_12
flabel metal1 178217 522946 178251 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_65.VGND
flabel metal1 178217 522402 178251 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_65.VPWR
flabel nwell 178217 522402 178251 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_65.VPB
flabel pwell 178217 522946 178251 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_65.VNB
rlabel comment 178188 522963 178188 522963 2 dpga_flat_0.sr_0.FILLER_0_14_65.decap_12
flabel metal1 179321 522402 179355 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_77.VPWR
flabel metal1 179321 522946 179355 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_77.VGND
flabel nwell 179321 522402 179355 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_77.VPB
flabel pwell 179321 522946 179355 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_77.VNB
rlabel comment 179292 522963 179292 522963 2 dpga_flat_0.sr_0.FILLER_0_14_77.decap_6
rlabel metal1 179292 522915 179844 523011 5 dpga_flat_0.sr_0.FILLER_0_14_77.VGND
rlabel metal1 179292 522371 179844 522467 5 dpga_flat_0.sr_0.FILLER_0_14_77.VPWR
flabel metal1 179866 522406 179902 522436 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_83.VPWR
flabel metal1 179866 522947 179902 522976 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_83.VGND
flabel nwell 179875 522412 179895 522429 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_83.VPB
flabel pwell 179872 522952 179896 522974 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_83.VNB
rlabel comment 179844 522963 179844 522963 2 dpga_flat_0.sr_0.FILLER_0_14_83.fill_1
rlabel metal1 179844 522915 179936 523011 5 dpga_flat_0.sr_0.FILLER_0_14_83.VGND
rlabel metal1 179844 522371 179936 522467 5 dpga_flat_0.sr_0.FILLER_0_14_83.VPWR
flabel metal1 180793 522946 180827 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_93.VGND
flabel metal1 180793 523490 180827 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_93.VPWR
flabel nwell 180793 523490 180827 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_93.VPB
flabel pwell 180793 522946 180827 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_93.VNB
rlabel comment 180764 522963 180764 522963 4 dpga_flat_0.sr_0.FILLER_0_13_93.decap_12
flabel metal1 180057 522946 180091 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_85.VGND
flabel metal1 180057 522402 180091 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_85.VPWR
flabel nwell 180057 522402 180091 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_85.VPB
flabel pwell 180057 522946 180091 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_85.VNB
rlabel comment 180028 522963 180028 522963 2 dpga_flat_0.sr_0.FILLER_0_14_85.decap_12
flabel metal1 181161 522946 181195 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_97.VGND
flabel metal1 181161 522402 181195 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_97.VPWR
flabel nwell 181161 522402 181195 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_97.VPB
flabel pwell 181161 522946 181195 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_97.VNB
rlabel comment 181132 522963 181132 522963 2 dpga_flat_0.sr_0.FILLER_0_14_97.decap_12
flabel metal1 179958 522410 180011 522439 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_14_94.VPWR
flabel metal1 179957 522943 180008 522981 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_14_94.VGND
rlabel comment 179936 522963 179936 522963 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_14_94.tapvpwrvgnd_1
rlabel metal1 179936 522915 180028 523011 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_14_94.VGND
rlabel metal1 179936 522371 180028 522467 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_14_94.VPWR
flabel metal1 181897 523490 181931 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_105.VPWR
flabel metal1 181897 522946 181931 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_105.VGND
flabel nwell 181897 523490 181931 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_105.VPB
flabel pwell 181897 522946 181931 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_105.VNB
rlabel comment 181868 522963 181868 522963 4 dpga_flat_0.sr_0.FILLER_0_13_105.decap_6
rlabel metal1 181868 522915 182420 523011 1 dpga_flat_0.sr_0.FILLER_0_13_105.VGND
rlabel metal1 181868 523459 182420 523555 1 dpga_flat_0.sr_0.FILLER_0_13_105.VPWR
flabel metal1 182442 523490 182478 523520 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_111.VPWR
flabel metal1 182442 522950 182478 522979 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_111.VGND
flabel nwell 182451 523497 182471 523514 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_111.VPB
flabel pwell 182448 522952 182472 522974 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_111.VNB
rlabel comment 182420 522963 182420 522963 4 dpga_flat_0.sr_0.FILLER_0_13_111.fill_1
rlabel metal1 182420 522915 182512 523011 1 dpga_flat_0.sr_0.FILLER_0_13_111.VGND
rlabel metal1 182420 523459 182512 523555 1 dpga_flat_0.sr_0.FILLER_0_13_111.VPWR
flabel metal1 182633 522946 182667 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_113.VGND
flabel metal1 182633 523490 182667 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_113.VPWR
flabel nwell 182633 523490 182667 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_113.VPB
flabel pwell 182633 522946 182667 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_113.VNB
rlabel comment 182604 522963 182604 522963 4 dpga_flat_0.sr_0.FILLER_0_13_113.decap_12
flabel metal1 183737 522946 183771 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_125.VGND
flabel metal1 183737 523490 183771 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_125.VPWR
flabel nwell 183737 523490 183771 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_125.VPB
flabel pwell 183737 522946 183771 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_125.VNB
rlabel comment 183708 522963 183708 522963 4 dpga_flat_0.sr_0.FILLER_0_13_125.decap_12
flabel metal1 182265 522946 182299 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_109.VGND
flabel metal1 182265 522402 182299 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_109.VPWR
flabel nwell 182265 522402 182299 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_109.VPB
flabel pwell 182265 522946 182299 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_109.VNB
rlabel comment 182236 522963 182236 522963 2 dpga_flat_0.sr_0.FILLER_0_14_109.decap_12
flabel metal1 183369 522946 183403 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_121.VGND
flabel metal1 183369 522402 183403 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_121.VPWR
flabel nwell 183369 522402 183403 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_121.VPB
flabel pwell 183369 522946 183403 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_121.VNB
rlabel comment 183340 522963 183340 522963 2 dpga_flat_0.sr_0.FILLER_0_14_121.decap_12
flabel metal1 182534 523487 182587 523516 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_13_92.VPWR
flabel metal1 182533 522945 182584 522983 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_13_92.VGND
rlabel comment 182512 522963 182512 522963 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_13_92.tapvpwrvgnd_1
rlabel metal1 182512 522915 182604 523011 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_13_92.VGND
rlabel metal1 182512 523459 182604 523555 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_13_92.VPWR
flabel metal1 184841 522946 184875 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_137.VGND
flabel metal1 184841 523490 184875 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_137.VPWR
flabel nwell 184841 523490 184875 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_137.VPB
flabel pwell 184841 522946 184875 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_137.VNB
rlabel comment 184812 522963 184812 522963 4 dpga_flat_0.sr_0.FILLER_0_13_137.decap_12
flabel metal1 184473 522402 184507 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_133.VPWR
flabel metal1 184473 522946 184507 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_133.VGND
flabel nwell 184473 522402 184507 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_133.VPB
flabel pwell 184473 522946 184507 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_133.VNB
rlabel comment 184444 522963 184444 522963 2 dpga_flat_0.sr_0.FILLER_0_14_133.decap_6
rlabel metal1 184444 522915 184996 523011 5 dpga_flat_0.sr_0.FILLER_0_14_133.VGND
rlabel metal1 184444 522371 184996 522467 5 dpga_flat_0.sr_0.FILLER_0_14_133.VPWR
flabel metal1 185018 522406 185054 522436 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_139.VPWR
flabel metal1 185018 522947 185054 522976 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_139.VGND
flabel nwell 185027 522412 185047 522429 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_139.VPB
flabel pwell 185024 522952 185048 522974 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_139.VNB
rlabel comment 184996 522963 184996 522963 2 dpga_flat_0.sr_0.FILLER_0_14_139.fill_1
rlabel metal1 184996 522915 185088 523011 5 dpga_flat_0.sr_0.FILLER_0_14_139.VGND
rlabel metal1 184996 522371 185088 522467 5 dpga_flat_0.sr_0.FILLER_0_14_139.VPWR
flabel metal1 185209 522946 185243 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_141.VGND
flabel metal1 185209 522402 185243 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_141.VPWR
flabel nwell 185209 522402 185243 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_141.VPB
flabel pwell 185209 522946 185243 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_141.VNB
rlabel comment 185180 522963 185180 522963 2 dpga_flat_0.sr_0.FILLER_0_14_141.decap_12
flabel metal1 185110 522410 185163 522439 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_14_95.VPWR
flabel metal1 185109 522943 185160 522981 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_14_95.VGND
rlabel comment 185088 522963 185088 522963 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_14_95.tapvpwrvgnd_1
rlabel metal1 185088 522915 185180 523011 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_14_95.VGND
rlabel metal1 185088 522371 185180 522467 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_14_95.VPWR
flabel metal1 185945 522946 185979 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_149.VGND
flabel metal1 185945 523490 185979 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_149.VPWR
flabel nwell 185945 523490 185979 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_149.VPB
flabel pwell 185945 522946 185979 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_149.VNB
rlabel comment 185916 522963 185916 522963 4 dpga_flat_0.sr_0.FILLER_0_13_149.decap_12
flabel metal1 187040 522949 187093 522981 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_161.VGND
flabel metal1 187041 523493 187093 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_161.VPWR
flabel nwell 187048 523498 187082 523516 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_161.VPB
flabel pwell 187051 522953 187083 522975 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_161.VNB
rlabel comment 187020 522963 187020 522963 4 dpga_flat_0.sr_0.FILLER_0_13_161.fill_2
rlabel metal1 187020 522915 187204 523011 1 dpga_flat_0.sr_0.FILLER_0_13_161.VGND
rlabel metal1 187020 523459 187204 523555 1 dpga_flat_0.sr_0.FILLER_0_13_161.VPWR
flabel metal1 186313 522402 186347 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_153.VPWR
flabel metal1 186313 522946 186347 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_153.VGND
flabel nwell 186313 522402 186347 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_153.VPB
flabel pwell 186313 522946 186347 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_153.VNB
rlabel comment 186284 522963 186284 522963 2 dpga_flat_0.sr_0.FILLER_0_14_153.decap_8
rlabel metal1 186284 522915 187020 523011 5 dpga_flat_0.sr_0.FILLER_0_14_153.VGND
rlabel metal1 186284 522371 187020 522467 5 dpga_flat_0.sr_0.FILLER_0_14_153.VPWR
flabel metal1 187040 522945 187093 522977 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_161.VGND
flabel metal1 187041 522402 187093 522433 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_161.VPWR
flabel nwell 187048 522410 187082 522428 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_161.VPB
flabel pwell 187051 522951 187083 522973 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_161.VNB
rlabel comment 187020 522963 187020 522963 2 dpga_flat_0.sr_0.FILLER_0_14_161.fill_2
rlabel metal1 187020 522915 187204 523011 5 dpga_flat_0.sr_0.FILLER_0_14_161.VGND
rlabel metal1 187020 522371 187204 522467 5 dpga_flat_0.sr_0.FILLER_0_14_161.VPWR
flabel metal1 187417 523490 187451 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_13_Right_13.VPWR
flabel metal1 187417 522946 187451 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_13_Right_13.VGND
flabel nwell 187417 523490 187451 523524 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_13_Right_13.VPB
flabel pwell 187417 522946 187451 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_13_Right_13.VNB
rlabel comment 187480 522963 187480 522963 6 dpga_flat_0.sr_0.PHY_EDGE_ROW_13_Right_13.decap_3
rlabel metal1 187204 522915 187480 523011 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_13_Right_13.VGND
rlabel metal1 187204 523459 187480 523555 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_13_Right_13.VPWR
flabel metal1 187417 522402 187451 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_14_Right_14.VPWR
flabel metal1 187417 522946 187451 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_14_Right_14.VGND
flabel nwell 187417 522402 187451 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_14_Right_14.VPB
flabel pwell 187417 522946 187451 522980 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_14_Right_14.VNB
rlabel comment 187480 522963 187480 522963 8 dpga_flat_0.sr_0.PHY_EDGE_ROW_14_Right_14.decap_3
rlabel metal1 187204 522915 187480 523011 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_14_Right_14.VGND
rlabel metal1 187204 522371 187480 522467 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_14_Right_14.VPWR
flabel metal1 172513 521858 172547 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_3.VGND
flabel metal1 172513 522402 172547 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_3.VPWR
flabel nwell 172513 522402 172547 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_3.VPB
flabel pwell 172513 521858 172547 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_3.VNB
rlabel comment 172484 521875 172484 521875 4 dpga_flat_0.sr_0.FILLER_0_15_3.decap_12
flabel metal1 173617 521858 173651 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_15.VGND
flabel metal1 173617 522402 173651 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_15.VPWR
flabel nwell 173617 522402 173651 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_15.VPB
flabel pwell 173617 521858 173651 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_15.VNB
rlabel comment 173588 521875 173588 521875 4 dpga_flat_0.sr_0.FILLER_0_15_15.decap_12
flabel metal1 172237 522402 172271 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_15_Left_43.VPWR
flabel metal1 172237 521858 172271 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_15_Left_43.VGND
flabel nwell 172237 522402 172271 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_15_Left_43.VPB
flabel pwell 172237 521858 172271 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_15_Left_43.VNB
rlabel comment 172208 521875 172208 521875 4 dpga_flat_0.sr_0.PHY_EDGE_ROW_15_Left_43.decap_3
rlabel metal1 172208 521827 172484 521923 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_15_Left_43.VGND
rlabel metal1 172208 522371 172484 522467 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_15_Left_43.VPWR
flabel metal1 174721 521858 174755 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_27.VGND
flabel metal1 174721 522402 174755 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_27.VPWR
flabel nwell 174721 522402 174755 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_27.VPB
flabel pwell 174721 521858 174755 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_27.VNB
rlabel comment 174692 521875 174692 521875 4 dpga_flat_0.sr_0.FILLER_0_15_27.decap_12
flabel metal1 175825 521858 175859 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_39.VGND
flabel metal1 175825 522402 175859 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_39.VPWR
flabel nwell 175825 522402 175859 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_39.VPB
flabel pwell 175825 521858 175859 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_39.VNB
rlabel comment 175796 521875 175796 521875 4 dpga_flat_0.sr_0.FILLER_0_15_39.decap_12
flabel metal1 176929 521858 176963 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_51.VGND
flabel metal1 176929 522402 176963 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_51.VPWR
flabel nwell 176929 522402 176963 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_51.VPB
flabel pwell 176929 521858 176963 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_51.VNB
rlabel comment 176900 521875 176900 521875 4 dpga_flat_0.sr_0.FILLER_0_15_51.decap_4
rlabel metal1 176900 521827 177268 521923 1 dpga_flat_0.sr_0.FILLER_0_15_51.VGND
rlabel metal1 176900 522371 177268 522467 1 dpga_flat_0.sr_0.FILLER_0_15_51.VPWR
flabel metal1 177290 522402 177326 522432 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_55.VPWR
flabel metal1 177290 521862 177326 521891 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_55.VGND
flabel nwell 177299 522409 177319 522426 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_55.VPB
flabel pwell 177296 521864 177320 521886 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_55.VNB
rlabel comment 177268 521875 177268 521875 4 dpga_flat_0.sr_0.FILLER_0_15_55.fill_1
rlabel metal1 177268 521827 177360 521923 1 dpga_flat_0.sr_0.FILLER_0_15_55.VGND
rlabel metal1 177268 522371 177360 522467 1 dpga_flat_0.sr_0.FILLER_0_15_55.VPWR
flabel metal1 177481 521858 177515 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_57.VGND
flabel metal1 177481 522402 177515 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_57.VPWR
flabel nwell 177481 522402 177515 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_57.VPB
flabel pwell 177481 521858 177515 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_57.VNB
rlabel comment 177452 521875 177452 521875 4 dpga_flat_0.sr_0.FILLER_0_15_57.decap_12
flabel metal1 177382 522399 177435 522428 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_15_96.VPWR
flabel metal1 177381 521857 177432 521895 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_15_96.VGND
rlabel comment 177360 521875 177360 521875 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_15_96.tapvpwrvgnd_1
rlabel metal1 177360 521827 177452 521923 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_15_96.VGND
rlabel metal1 177360 522371 177452 522467 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_15_96.VPWR
flabel metal1 178585 521858 178619 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_69.VGND
flabel metal1 178585 522402 178619 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_69.VPWR
flabel nwell 178585 522402 178619 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_69.VPB
flabel pwell 178585 521858 178619 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_69.VNB
rlabel comment 178556 521875 178556 521875 4 dpga_flat_0.sr_0.FILLER_0_15_69.decap_12
flabel metal1 179689 521858 179723 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_81.VGND
flabel metal1 179689 522402 179723 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_81.VPWR
flabel nwell 179689 522402 179723 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_81.VPB
flabel pwell 179689 521858 179723 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_81.VNB
rlabel comment 179660 521875 179660 521875 4 dpga_flat_0.sr_0.FILLER_0_15_81.decap_12
flabel metal1 180793 521858 180827 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_93.VGND
flabel metal1 180793 522402 180827 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_93.VPWR
flabel nwell 180793 522402 180827 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_93.VPB
flabel pwell 180793 521858 180827 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_93.VNB
rlabel comment 180764 521875 180764 521875 4 dpga_flat_0.sr_0.FILLER_0_15_93.decap_12
flabel metal1 181897 522402 181931 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_105.VPWR
flabel metal1 181897 521858 181931 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_105.VGND
flabel nwell 181897 522402 181931 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_105.VPB
flabel pwell 181897 521858 181931 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_105.VNB
rlabel comment 181868 521875 181868 521875 4 dpga_flat_0.sr_0.FILLER_0_15_105.decap_6
rlabel metal1 181868 521827 182420 521923 1 dpga_flat_0.sr_0.FILLER_0_15_105.VGND
rlabel metal1 181868 522371 182420 522467 1 dpga_flat_0.sr_0.FILLER_0_15_105.VPWR
flabel metal1 182442 522402 182478 522432 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_111.VPWR
flabel metal1 182442 521862 182478 521891 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_111.VGND
flabel nwell 182451 522409 182471 522426 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_111.VPB
flabel pwell 182448 521864 182472 521886 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_111.VNB
rlabel comment 182420 521875 182420 521875 4 dpga_flat_0.sr_0.FILLER_0_15_111.fill_1
rlabel metal1 182420 521827 182512 521923 1 dpga_flat_0.sr_0.FILLER_0_15_111.VGND
rlabel metal1 182420 522371 182512 522467 1 dpga_flat_0.sr_0.FILLER_0_15_111.VPWR
flabel metal1 182633 521858 182667 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_113.VGND
flabel metal1 182633 522402 182667 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_113.VPWR
flabel nwell 182633 522402 182667 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_113.VPB
flabel pwell 182633 521858 182667 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_113.VNB
rlabel comment 182604 521875 182604 521875 4 dpga_flat_0.sr_0.FILLER_0_15_113.decap_12
flabel metal1 183737 521858 183771 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_125.VGND
flabel metal1 183737 522402 183771 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_125.VPWR
flabel nwell 183737 522402 183771 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_125.VPB
flabel pwell 183737 521858 183771 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_125.VNB
rlabel comment 183708 521875 183708 521875 4 dpga_flat_0.sr_0.FILLER_0_15_125.decap_12
flabel metal1 182534 522399 182587 522428 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_15_97.VPWR
flabel metal1 182533 521857 182584 521895 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_15_97.VGND
rlabel comment 182512 521875 182512 521875 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_15_97.tapvpwrvgnd_1
rlabel metal1 182512 521827 182604 521923 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_15_97.VGND
rlabel metal1 182512 522371 182604 522467 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_15_97.VPWR
flabel metal1 184841 521858 184875 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_137.VGND
flabel metal1 184841 522402 184875 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_137.VPWR
flabel nwell 184841 522402 184875 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_137.VPB
flabel pwell 184841 521858 184875 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_137.VNB
rlabel comment 184812 521875 184812 521875 4 dpga_flat_0.sr_0.FILLER_0_15_137.decap_12
flabel metal1 185945 521858 185979 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_149.VGND
flabel metal1 185945 522402 185979 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_149.VPWR
flabel nwell 185945 522402 185979 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_149.VPB
flabel pwell 185945 521858 185979 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_149.VNB
rlabel comment 185916 521875 185916 521875 4 dpga_flat_0.sr_0.FILLER_0_15_149.decap_12
flabel metal1 187040 521861 187093 521893 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_161.VGND
flabel metal1 187041 522405 187093 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_161.VPWR
flabel nwell 187048 522410 187082 522428 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_161.VPB
flabel pwell 187051 521865 187083 521887 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_161.VNB
rlabel comment 187020 521875 187020 521875 4 dpga_flat_0.sr_0.FILLER_0_15_161.fill_2
rlabel metal1 187020 521827 187204 521923 1 dpga_flat_0.sr_0.FILLER_0_15_161.VGND
rlabel metal1 187020 522371 187204 522467 1 dpga_flat_0.sr_0.FILLER_0_15_161.VPWR
flabel metal1 187417 522402 187451 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_15_Right_15.VPWR
flabel metal1 187417 521858 187451 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_15_Right_15.VGND
flabel nwell 187417 522402 187451 522436 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_15_Right_15.VPB
flabel pwell 187417 521858 187451 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_15_Right_15.VNB
rlabel comment 187480 521875 187480 521875 6 dpga_flat_0.sr_0.PHY_EDGE_ROW_15_Right_15.decap_3
rlabel metal1 187204 521827 187480 521923 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_15_Right_15.VGND
rlabel metal1 187204 522371 187480 522467 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_15_Right_15.VPWR
flabel metal1 172513 521858 172547 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_3.VGND
flabel metal1 172513 521314 172547 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_3.VPWR
flabel nwell 172513 521314 172547 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_3.VPB
flabel pwell 172513 521858 172547 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_3.VNB
rlabel comment 172484 521875 172484 521875 2 dpga_flat_0.sr_0.FILLER_0_16_3.decap_12
flabel metal1 173617 521858 173651 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_15.VGND
flabel metal1 173617 521314 173651 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_15.VPWR
flabel nwell 173617 521314 173651 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_15.VPB
flabel pwell 173617 521858 173651 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_15.VNB
rlabel comment 173588 521875 173588 521875 2 dpga_flat_0.sr_0.FILLER_0_16_15.decap_12
flabel metal1 172237 521314 172271 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_16_Left_44.VPWR
flabel metal1 172237 521858 172271 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_16_Left_44.VGND
flabel nwell 172237 521314 172271 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_16_Left_44.VPB
flabel pwell 172237 521858 172271 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_16_Left_44.VNB
rlabel comment 172208 521875 172208 521875 2 dpga_flat_0.sr_0.PHY_EDGE_ROW_16_Left_44.decap_3
rlabel metal1 172208 521827 172484 521923 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_16_Left_44.VGND
rlabel metal1 172208 521283 172484 521379 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_16_Left_44.VPWR
flabel metal1 174714 521318 174750 521348 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_27.VPWR
flabel metal1 174714 521859 174750 521888 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_27.VGND
flabel nwell 174723 521324 174743 521341 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_27.VPB
flabel pwell 174720 521864 174744 521886 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_27.VNB
rlabel comment 174692 521875 174692 521875 2 dpga_flat_0.sr_0.FILLER_0_16_27.fill_1
rlabel metal1 174692 521827 174784 521923 5 dpga_flat_0.sr_0.FILLER_0_16_27.VGND
rlabel metal1 174692 521283 174784 521379 5 dpga_flat_0.sr_0.FILLER_0_16_27.VPWR
flabel metal1 174905 521858 174939 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_29.VGND
flabel metal1 174905 521314 174939 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_29.VPWR
flabel nwell 174905 521314 174939 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_29.VPB
flabel pwell 174905 521858 174939 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_29.VNB
rlabel comment 174876 521875 174876 521875 2 dpga_flat_0.sr_0.FILLER_0_16_29.decap_12
flabel metal1 176009 521858 176043 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_41.VGND
flabel metal1 176009 521314 176043 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_41.VPWR
flabel nwell 176009 521314 176043 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_41.VPB
flabel pwell 176009 521858 176043 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_41.VNB
rlabel comment 175980 521875 175980 521875 2 dpga_flat_0.sr_0.FILLER_0_16_41.decap_12
flabel metal1 174806 521322 174859 521351 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_16_98.VPWR
flabel metal1 174805 521855 174856 521893 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_16_98.VGND
rlabel comment 174784 521875 174784 521875 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_16_98.tapvpwrvgnd_1
rlabel metal1 174784 521827 174876 521923 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_16_98.VGND
rlabel metal1 174784 521283 174876 521379 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_16_98.VPWR
flabel metal1 177113 521858 177147 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_53.VGND
flabel metal1 177113 521314 177147 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_53.VPWR
flabel nwell 177113 521314 177147 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_53.VPB
flabel pwell 177113 521858 177147 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_53.VNB
rlabel comment 177084 521875 177084 521875 2 dpga_flat_0.sr_0.FILLER_0_16_53.decap_12
flabel metal1 178217 521858 178251 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_65.VGND
flabel metal1 178217 521314 178251 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_65.VPWR
flabel nwell 178217 521314 178251 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_65.VPB
flabel pwell 178217 521858 178251 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_65.VNB
rlabel comment 178188 521875 178188 521875 2 dpga_flat_0.sr_0.FILLER_0_16_65.decap_12
flabel metal1 179321 521314 179355 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_77.VPWR
flabel metal1 179321 521858 179355 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_77.VGND
flabel nwell 179321 521314 179355 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_77.VPB
flabel pwell 179321 521858 179355 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_77.VNB
rlabel comment 179292 521875 179292 521875 2 dpga_flat_0.sr_0.FILLER_0_16_77.decap_6
rlabel metal1 179292 521827 179844 521923 5 dpga_flat_0.sr_0.FILLER_0_16_77.VGND
rlabel metal1 179292 521283 179844 521379 5 dpga_flat_0.sr_0.FILLER_0_16_77.VPWR
flabel metal1 179866 521318 179902 521348 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_83.VPWR
flabel metal1 179866 521859 179902 521888 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_83.VGND
flabel nwell 179875 521324 179895 521341 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_83.VPB
flabel pwell 179872 521864 179896 521886 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_83.VNB
rlabel comment 179844 521875 179844 521875 2 dpga_flat_0.sr_0.FILLER_0_16_83.fill_1
rlabel metal1 179844 521827 179936 521923 5 dpga_flat_0.sr_0.FILLER_0_16_83.VGND
rlabel metal1 179844 521283 179936 521379 5 dpga_flat_0.sr_0.FILLER_0_16_83.VPWR
flabel metal1 180057 521858 180091 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_85.VGND
flabel metal1 180057 521314 180091 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_85.VPWR
flabel nwell 180057 521314 180091 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_85.VPB
flabel pwell 180057 521858 180091 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_85.VNB
rlabel comment 180028 521875 180028 521875 2 dpga_flat_0.sr_0.FILLER_0_16_85.decap_12
flabel metal1 181161 521858 181195 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_97.VGND
flabel metal1 181161 521314 181195 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_97.VPWR
flabel nwell 181161 521314 181195 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_97.VPB
flabel pwell 181161 521858 181195 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_97.VNB
rlabel comment 181132 521875 181132 521875 2 dpga_flat_0.sr_0.FILLER_0_16_97.decap_12
flabel metal1 179958 521322 180011 521351 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_16_99.VPWR
flabel metal1 179957 521855 180008 521893 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_16_99.VGND
rlabel comment 179936 521875 179936 521875 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_16_99.tapvpwrvgnd_1
rlabel metal1 179936 521827 180028 521923 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_16_99.VGND
rlabel metal1 179936 521283 180028 521379 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_16_99.VPWR
flabel metal1 182265 521858 182299 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_109.VGND
flabel metal1 182265 521314 182299 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_109.VPWR
flabel nwell 182265 521314 182299 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_109.VPB
flabel pwell 182265 521858 182299 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_109.VNB
rlabel comment 182236 521875 182236 521875 2 dpga_flat_0.sr_0.FILLER_0_16_109.decap_12
flabel metal1 183369 521858 183403 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_121.VGND
flabel metal1 183369 521314 183403 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_121.VPWR
flabel nwell 183369 521314 183403 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_121.VPB
flabel pwell 183369 521858 183403 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_121.VNB
rlabel comment 183340 521875 183340 521875 2 dpga_flat_0.sr_0.FILLER_0_16_121.decap_12
flabel metal1 184473 521314 184507 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_133.VPWR
flabel metal1 184473 521858 184507 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_133.VGND
flabel nwell 184473 521314 184507 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_133.VPB
flabel pwell 184473 521858 184507 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_133.VNB
rlabel comment 184444 521875 184444 521875 2 dpga_flat_0.sr_0.FILLER_0_16_133.decap_6
rlabel metal1 184444 521827 184996 521923 5 dpga_flat_0.sr_0.FILLER_0_16_133.VGND
rlabel metal1 184444 521283 184996 521379 5 dpga_flat_0.sr_0.FILLER_0_16_133.VPWR
flabel metal1 185018 521318 185054 521348 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_139.VPWR
flabel metal1 185018 521859 185054 521888 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_139.VGND
flabel nwell 185027 521324 185047 521341 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_139.VPB
flabel pwell 185024 521864 185048 521886 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_139.VNB
rlabel comment 184996 521875 184996 521875 2 dpga_flat_0.sr_0.FILLER_0_16_139.fill_1
rlabel metal1 184996 521827 185088 521923 5 dpga_flat_0.sr_0.FILLER_0_16_139.VGND
rlabel metal1 184996 521283 185088 521379 5 dpga_flat_0.sr_0.FILLER_0_16_139.VPWR
flabel metal1 185209 521858 185243 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_141.VGND
flabel metal1 185209 521314 185243 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_141.VPWR
flabel nwell 185209 521314 185243 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_141.VPB
flabel pwell 185209 521858 185243 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_141.VNB
rlabel comment 185180 521875 185180 521875 2 dpga_flat_0.sr_0.FILLER_0_16_141.decap_12
flabel metal1 185110 521322 185163 521351 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_16_100.VPWR
flabel metal1 185109 521855 185160 521893 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_16_100.VGND
rlabel comment 185088 521875 185088 521875 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_16_100.tapvpwrvgnd_1
rlabel metal1 185088 521827 185180 521923 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_16_100.VGND
rlabel metal1 185088 521283 185180 521379 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_16_100.VPWR
flabel metal1 186313 521314 186347 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_153.VPWR
flabel metal1 186313 521858 186347 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_153.VGND
flabel nwell 186313 521314 186347 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_153.VPB
flabel pwell 186313 521858 186347 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_153.VNB
rlabel comment 186284 521875 186284 521875 2 dpga_flat_0.sr_0.FILLER_0_16_153.decap_8
rlabel metal1 186284 521827 187020 521923 5 dpga_flat_0.sr_0.FILLER_0_16_153.VGND
rlabel metal1 186284 521283 187020 521379 5 dpga_flat_0.sr_0.FILLER_0_16_153.VPWR
flabel metal1 187040 521857 187093 521889 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_161.VGND
flabel metal1 187041 521314 187093 521345 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_161.VPWR
flabel nwell 187048 521322 187082 521340 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_161.VPB
flabel pwell 187051 521863 187083 521885 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_161.VNB
rlabel comment 187020 521875 187020 521875 2 dpga_flat_0.sr_0.FILLER_0_16_161.fill_2
rlabel metal1 187020 521827 187204 521923 5 dpga_flat_0.sr_0.FILLER_0_16_161.VGND
rlabel metal1 187020 521283 187204 521379 5 dpga_flat_0.sr_0.FILLER_0_16_161.VPWR
flabel metal1 187417 521314 187451 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_16_Right_16.VPWR
flabel metal1 187417 521858 187451 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_16_Right_16.VGND
flabel nwell 187417 521314 187451 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_16_Right_16.VPB
flabel pwell 187417 521858 187451 521892 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_16_Right_16.VNB
rlabel comment 187480 521875 187480 521875 8 dpga_flat_0.sr_0.PHY_EDGE_ROW_16_Right_16.decap_3
rlabel metal1 187204 521827 187480 521923 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_16_Right_16.VGND
rlabel metal1 187204 521283 187480 521379 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_16_Right_16.VPWR
flabel metal1 172513 520770 172547 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_3.VGND
flabel metal1 172513 521314 172547 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_3.VPWR
flabel nwell 172513 521314 172547 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_3.VPB
flabel pwell 172513 520770 172547 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_3.VNB
rlabel comment 172484 520787 172484 520787 4 dpga_flat_0.sr_0.FILLER_0_17_3.decap_12
flabel metal1 173617 520770 173651 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_15.VGND
flabel metal1 173617 521314 173651 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_15.VPWR
flabel nwell 173617 521314 173651 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_15.VPB
flabel pwell 173617 520770 173651 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_15.VNB
rlabel comment 173588 520787 173588 520787 4 dpga_flat_0.sr_0.FILLER_0_17_15.decap_12
flabel metal1 172237 521314 172271 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_17_Left_45.VPWR
flabel metal1 172237 520770 172271 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_17_Left_45.VGND
flabel nwell 172237 521314 172271 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_17_Left_45.VPB
flabel pwell 172237 520770 172271 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_17_Left_45.VNB
rlabel comment 172208 520787 172208 520787 4 dpga_flat_0.sr_0.PHY_EDGE_ROW_17_Left_45.decap_3
rlabel metal1 172208 520739 172484 520835 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_17_Left_45.VGND
rlabel metal1 172208 521283 172484 521379 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_17_Left_45.VPWR
flabel metal1 174721 520770 174755 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_27.VGND
flabel metal1 174721 521314 174755 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_27.VPWR
flabel nwell 174721 521314 174755 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_27.VPB
flabel pwell 174721 520770 174755 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_27.VNB
rlabel comment 174692 520787 174692 520787 4 dpga_flat_0.sr_0.FILLER_0_17_27.decap_12
flabel metal1 175825 520770 175859 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_39.VGND
flabel metal1 175825 521314 175859 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_39.VPWR
flabel nwell 175825 521314 175859 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_39.VPB
flabel pwell 175825 520770 175859 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_39.VNB
rlabel comment 175796 520787 175796 520787 4 dpga_flat_0.sr_0.FILLER_0_17_39.decap_12
flabel metal1 176929 520770 176963 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_51.VGND
flabel metal1 176929 521314 176963 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_51.VPWR
flabel nwell 176929 521314 176963 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_51.VPB
flabel pwell 176929 520770 176963 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_51.VNB
rlabel comment 176900 520787 176900 520787 4 dpga_flat_0.sr_0.FILLER_0_17_51.decap_4
rlabel metal1 176900 520739 177268 520835 1 dpga_flat_0.sr_0.FILLER_0_17_51.VGND
rlabel metal1 176900 521283 177268 521379 1 dpga_flat_0.sr_0.FILLER_0_17_51.VPWR
flabel metal1 177290 521314 177326 521344 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_55.VPWR
flabel metal1 177290 520774 177326 520803 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_55.VGND
flabel nwell 177299 521321 177319 521338 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_55.VPB
flabel pwell 177296 520776 177320 520798 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_55.VNB
rlabel comment 177268 520787 177268 520787 4 dpga_flat_0.sr_0.FILLER_0_17_55.fill_1
rlabel metal1 177268 520739 177360 520835 1 dpga_flat_0.sr_0.FILLER_0_17_55.VGND
rlabel metal1 177268 521283 177360 521379 1 dpga_flat_0.sr_0.FILLER_0_17_55.VPWR
flabel metal1 177481 520770 177515 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_57.VGND
flabel metal1 177481 521314 177515 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_57.VPWR
flabel nwell 177481 521314 177515 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_57.VPB
flabel pwell 177481 520770 177515 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_57.VNB
rlabel comment 177452 520787 177452 520787 4 dpga_flat_0.sr_0.FILLER_0_17_57.decap_12
flabel metal1 177382 521311 177435 521340 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_17_101.VPWR
flabel metal1 177381 520769 177432 520807 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_17_101.VGND
rlabel comment 177360 520787 177360 520787 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_17_101.tapvpwrvgnd_1
rlabel metal1 177360 520739 177452 520835 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_17_101.VGND
rlabel metal1 177360 521283 177452 521379 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_17_101.VPWR
flabel metal1 178585 520770 178619 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_69.VGND
flabel metal1 178585 521314 178619 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_69.VPWR
flabel nwell 178585 521314 178619 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_69.VPB
flabel pwell 178585 520770 178619 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_69.VNB
rlabel comment 178556 520787 178556 520787 4 dpga_flat_0.sr_0.FILLER_0_17_69.decap_12
flabel metal1 179689 520770 179723 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_81.VGND
flabel metal1 179689 521314 179723 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_81.VPWR
flabel nwell 179689 521314 179723 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_81.VPB
flabel pwell 179689 520770 179723 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_81.VNB
rlabel comment 179660 520787 179660 520787 4 dpga_flat_0.sr_0.FILLER_0_17_81.decap_12
flabel metal1 180793 520770 180827 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_93.VGND
flabel metal1 180793 521314 180827 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_93.VPWR
flabel nwell 180793 521314 180827 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_93.VPB
flabel pwell 180793 520770 180827 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_93.VNB
rlabel comment 180764 520787 180764 520787 4 dpga_flat_0.sr_0.FILLER_0_17_93.decap_12
flabel metal1 181897 521314 181931 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_105.VPWR
flabel metal1 181897 520770 181931 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_105.VGND
flabel nwell 181897 521314 181931 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_105.VPB
flabel pwell 181897 520770 181931 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_105.VNB
rlabel comment 181868 520787 181868 520787 4 dpga_flat_0.sr_0.FILLER_0_17_105.decap_6
rlabel metal1 181868 520739 182420 520835 1 dpga_flat_0.sr_0.FILLER_0_17_105.VGND
rlabel metal1 181868 521283 182420 521379 1 dpga_flat_0.sr_0.FILLER_0_17_105.VPWR
flabel metal1 182442 521314 182478 521344 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_111.VPWR
flabel metal1 182442 520774 182478 520803 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_111.VGND
flabel nwell 182451 521321 182471 521338 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_111.VPB
flabel pwell 182448 520776 182472 520798 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_111.VNB
rlabel comment 182420 520787 182420 520787 4 dpga_flat_0.sr_0.FILLER_0_17_111.fill_1
rlabel metal1 182420 520739 182512 520835 1 dpga_flat_0.sr_0.FILLER_0_17_111.VGND
rlabel metal1 182420 521283 182512 521379 1 dpga_flat_0.sr_0.FILLER_0_17_111.VPWR
flabel metal1 182633 520770 182667 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_113.VGND
flabel metal1 182633 521314 182667 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_113.VPWR
flabel nwell 182633 521314 182667 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_113.VPB
flabel pwell 182633 520770 182667 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_113.VNB
rlabel comment 182604 520787 182604 520787 4 dpga_flat_0.sr_0.FILLER_0_17_113.decap_12
flabel metal1 183737 520770 183771 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_125.VGND
flabel metal1 183737 521314 183771 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_125.VPWR
flabel nwell 183737 521314 183771 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_125.VPB
flabel pwell 183737 520770 183771 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_125.VNB
rlabel comment 183708 520787 183708 520787 4 dpga_flat_0.sr_0.FILLER_0_17_125.decap_12
flabel metal1 182534 521311 182587 521340 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_17_102.VPWR
flabel metal1 182533 520769 182584 520807 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_17_102.VGND
rlabel comment 182512 520787 182512 520787 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_17_102.tapvpwrvgnd_1
rlabel metal1 182512 520739 182604 520835 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_17_102.VGND
rlabel metal1 182512 521283 182604 521379 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_17_102.VPWR
flabel metal1 184841 520770 184875 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_137.VGND
flabel metal1 184841 521314 184875 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_137.VPWR
flabel nwell 184841 521314 184875 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_137.VPB
flabel pwell 184841 520770 184875 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_137.VNB
rlabel comment 184812 520787 184812 520787 4 dpga_flat_0.sr_0.FILLER_0_17_137.decap_12
flabel metal1 185945 520770 185979 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_149.VGND
flabel metal1 185945 521314 185979 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_149.VPWR
flabel nwell 185945 521314 185979 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_149.VPB
flabel pwell 185945 520770 185979 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_149.VNB
rlabel comment 185916 520787 185916 520787 4 dpga_flat_0.sr_0.FILLER_0_17_149.decap_12
flabel metal1 187040 520773 187093 520805 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_161.VGND
flabel metal1 187041 521317 187093 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_161.VPWR
flabel nwell 187048 521322 187082 521340 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_161.VPB
flabel pwell 187051 520777 187083 520799 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_161.VNB
rlabel comment 187020 520787 187020 520787 4 dpga_flat_0.sr_0.FILLER_0_17_161.fill_2
rlabel metal1 187020 520739 187204 520835 1 dpga_flat_0.sr_0.FILLER_0_17_161.VGND
rlabel metal1 187020 521283 187204 521379 1 dpga_flat_0.sr_0.FILLER_0_17_161.VPWR
flabel metal1 187417 521314 187451 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_17_Right_17.VPWR
flabel metal1 187417 520770 187451 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_17_Right_17.VGND
flabel nwell 187417 521314 187451 521348 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_17_Right_17.VPB
flabel pwell 187417 520770 187451 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_17_Right_17.VNB
rlabel comment 187480 520787 187480 520787 6 dpga_flat_0.sr_0.PHY_EDGE_ROW_17_Right_17.decap_3
rlabel metal1 187204 520739 187480 520835 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_17_Right_17.VGND
rlabel metal1 187204 521283 187480 521379 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_17_Right_17.VPWR
flabel metal1 172513 520770 172547 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_3.VGND
flabel metal1 172513 520226 172547 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_3.VPWR
flabel nwell 172513 520226 172547 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_3.VPB
flabel pwell 172513 520770 172547 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_3.VNB
rlabel comment 172484 520787 172484 520787 2 dpga_flat_0.sr_0.FILLER_0_18_3.decap_12
flabel metal1 173617 520770 173651 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_15.VGND
flabel metal1 173617 520226 173651 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_15.VPWR
flabel nwell 173617 520226 173651 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_15.VPB
flabel pwell 173617 520770 173651 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_15.VNB
rlabel comment 173588 520787 173588 520787 2 dpga_flat_0.sr_0.FILLER_0_18_15.decap_12
flabel metal1 172237 520226 172271 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_18_Left_46.VPWR
flabel metal1 172237 520770 172271 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_18_Left_46.VGND
flabel nwell 172237 520226 172271 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_18_Left_46.VPB
flabel pwell 172237 520770 172271 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_18_Left_46.VNB
rlabel comment 172208 520787 172208 520787 2 dpga_flat_0.sr_0.PHY_EDGE_ROW_18_Left_46.decap_3
rlabel metal1 172208 520739 172484 520835 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_18_Left_46.VGND
rlabel metal1 172208 520195 172484 520291 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_18_Left_46.VPWR
flabel metal1 174714 520230 174750 520260 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_27.VPWR
flabel metal1 174714 520771 174750 520800 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_27.VGND
flabel nwell 174723 520236 174743 520253 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_27.VPB
flabel pwell 174720 520776 174744 520798 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_27.VNB
rlabel comment 174692 520787 174692 520787 2 dpga_flat_0.sr_0.FILLER_0_18_27.fill_1
rlabel metal1 174692 520739 174784 520835 5 dpga_flat_0.sr_0.FILLER_0_18_27.VGND
rlabel metal1 174692 520195 174784 520291 5 dpga_flat_0.sr_0.FILLER_0_18_27.VPWR
flabel metal1 174905 520770 174939 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_29.VGND
flabel metal1 174905 520226 174939 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_29.VPWR
flabel nwell 174905 520226 174939 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_29.VPB
flabel pwell 174905 520770 174939 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_29.VNB
rlabel comment 174876 520787 174876 520787 2 dpga_flat_0.sr_0.FILLER_0_18_29.decap_12
flabel metal1 176009 520770 176043 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_41.VGND
flabel metal1 176009 520226 176043 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_41.VPWR
flabel nwell 176009 520226 176043 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_41.VPB
flabel pwell 176009 520770 176043 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_41.VNB
rlabel comment 175980 520787 175980 520787 2 dpga_flat_0.sr_0.FILLER_0_18_41.decap_12
flabel metal1 174806 520234 174859 520263 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_18_103.VPWR
flabel metal1 174805 520767 174856 520805 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_18_103.VGND
rlabel comment 174784 520787 174784 520787 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_18_103.tapvpwrvgnd_1
rlabel metal1 174784 520739 174876 520835 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_18_103.VGND
rlabel metal1 174784 520195 174876 520291 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_18_103.VPWR
flabel metal1 177113 520770 177147 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_53.VGND
flabel metal1 177113 520226 177147 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_53.VPWR
flabel nwell 177113 520226 177147 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_53.VPB
flabel pwell 177113 520770 177147 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_53.VNB
rlabel comment 177084 520787 177084 520787 2 dpga_flat_0.sr_0.FILLER_0_18_53.decap_12
flabel metal1 178217 520770 178251 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_65.VGND
flabel metal1 178217 520226 178251 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_65.VPWR
flabel nwell 178217 520226 178251 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_65.VPB
flabel pwell 178217 520770 178251 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_65.VNB
rlabel comment 178188 520787 178188 520787 2 dpga_flat_0.sr_0.FILLER_0_18_65.decap_12
flabel metal1 179321 520226 179355 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_77.VPWR
flabel metal1 179321 520770 179355 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_77.VGND
flabel nwell 179321 520226 179355 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_77.VPB
flabel pwell 179321 520770 179355 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_77.VNB
rlabel comment 179292 520787 179292 520787 2 dpga_flat_0.sr_0.FILLER_0_18_77.decap_6
rlabel metal1 179292 520739 179844 520835 5 dpga_flat_0.sr_0.FILLER_0_18_77.VGND
rlabel metal1 179292 520195 179844 520291 5 dpga_flat_0.sr_0.FILLER_0_18_77.VPWR
flabel metal1 179866 520230 179902 520260 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_83.VPWR
flabel metal1 179866 520771 179902 520800 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_83.VGND
flabel nwell 179875 520236 179895 520253 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_83.VPB
flabel pwell 179872 520776 179896 520798 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_83.VNB
rlabel comment 179844 520787 179844 520787 2 dpga_flat_0.sr_0.FILLER_0_18_83.fill_1
rlabel metal1 179844 520739 179936 520835 5 dpga_flat_0.sr_0.FILLER_0_18_83.VGND
rlabel metal1 179844 520195 179936 520291 5 dpga_flat_0.sr_0.FILLER_0_18_83.VPWR
flabel metal1 180057 520770 180091 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_85.VGND
flabel metal1 180057 520226 180091 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_85.VPWR
flabel nwell 180057 520226 180091 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_85.VPB
flabel pwell 180057 520770 180091 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_85.VNB
rlabel comment 180028 520787 180028 520787 2 dpga_flat_0.sr_0.FILLER_0_18_85.decap_12
flabel metal1 181161 520770 181195 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_97.VGND
flabel metal1 181161 520226 181195 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_97.VPWR
flabel nwell 181161 520226 181195 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_97.VPB
flabel pwell 181161 520770 181195 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_97.VNB
rlabel comment 181132 520787 181132 520787 2 dpga_flat_0.sr_0.FILLER_0_18_97.decap_12
flabel metal1 179958 520234 180011 520263 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_18_104.VPWR
flabel metal1 179957 520767 180008 520805 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_18_104.VGND
rlabel comment 179936 520787 179936 520787 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_18_104.tapvpwrvgnd_1
rlabel metal1 179936 520739 180028 520835 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_18_104.VGND
rlabel metal1 179936 520195 180028 520291 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_18_104.VPWR
flabel metal1 182265 520770 182299 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_109.VGND
flabel metal1 182265 520226 182299 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_109.VPWR
flabel nwell 182265 520226 182299 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_109.VPB
flabel pwell 182265 520770 182299 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_109.VNB
rlabel comment 182236 520787 182236 520787 2 dpga_flat_0.sr_0.FILLER_0_18_109.decap_12
flabel metal1 183369 520770 183403 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_121.VGND
flabel metal1 183369 520226 183403 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_121.VPWR
flabel nwell 183369 520226 183403 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_121.VPB
flabel pwell 183369 520770 183403 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_121.VNB
rlabel comment 183340 520787 183340 520787 2 dpga_flat_0.sr_0.FILLER_0_18_121.decap_12
flabel metal1 184473 520226 184507 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_133.VPWR
flabel metal1 184473 520770 184507 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_133.VGND
flabel nwell 184473 520226 184507 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_133.VPB
flabel pwell 184473 520770 184507 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_133.VNB
rlabel comment 184444 520787 184444 520787 2 dpga_flat_0.sr_0.FILLER_0_18_133.decap_6
rlabel metal1 184444 520739 184996 520835 5 dpga_flat_0.sr_0.FILLER_0_18_133.VGND
rlabel metal1 184444 520195 184996 520291 5 dpga_flat_0.sr_0.FILLER_0_18_133.VPWR
flabel metal1 185018 520230 185054 520260 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_139.VPWR
flabel metal1 185018 520771 185054 520800 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_139.VGND
flabel nwell 185027 520236 185047 520253 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_139.VPB
flabel pwell 185024 520776 185048 520798 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_139.VNB
rlabel comment 184996 520787 184996 520787 2 dpga_flat_0.sr_0.FILLER_0_18_139.fill_1
rlabel metal1 184996 520739 185088 520835 5 dpga_flat_0.sr_0.FILLER_0_18_139.VGND
rlabel metal1 184996 520195 185088 520291 5 dpga_flat_0.sr_0.FILLER_0_18_139.VPWR
flabel metal1 185209 520770 185243 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_141.VGND
flabel metal1 185209 520226 185243 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_141.VPWR
flabel nwell 185209 520226 185243 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_141.VPB
flabel pwell 185209 520770 185243 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_141.VNB
rlabel comment 185180 520787 185180 520787 2 dpga_flat_0.sr_0.FILLER_0_18_141.decap_12
flabel metal1 185110 520234 185163 520263 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_18_105.VPWR
flabel metal1 185109 520767 185160 520805 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_18_105.VGND
rlabel comment 185088 520787 185088 520787 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_18_105.tapvpwrvgnd_1
rlabel metal1 185088 520739 185180 520835 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_18_105.VGND
rlabel metal1 185088 520195 185180 520291 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_18_105.VPWR
flabel metal1 186313 520226 186347 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_153.VPWR
flabel metal1 186313 520770 186347 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_153.VGND
flabel nwell 186313 520226 186347 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_153.VPB
flabel pwell 186313 520770 186347 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_153.VNB
rlabel comment 186284 520787 186284 520787 2 dpga_flat_0.sr_0.FILLER_0_18_153.decap_8
rlabel metal1 186284 520739 187020 520835 5 dpga_flat_0.sr_0.FILLER_0_18_153.VGND
rlabel metal1 186284 520195 187020 520291 5 dpga_flat_0.sr_0.FILLER_0_18_153.VPWR
flabel metal1 187040 520769 187093 520801 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_161.VGND
flabel metal1 187041 520226 187093 520257 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_161.VPWR
flabel nwell 187048 520234 187082 520252 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_161.VPB
flabel pwell 187051 520775 187083 520797 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_161.VNB
rlabel comment 187020 520787 187020 520787 2 dpga_flat_0.sr_0.FILLER_0_18_161.fill_2
rlabel metal1 187020 520739 187204 520835 5 dpga_flat_0.sr_0.FILLER_0_18_161.VGND
rlabel metal1 187020 520195 187204 520291 5 dpga_flat_0.sr_0.FILLER_0_18_161.VPWR
flabel metal1 187417 520226 187451 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_18_Right_18.VPWR
flabel metal1 187417 520770 187451 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_18_Right_18.VGND
flabel nwell 187417 520226 187451 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_18_Right_18.VPB
flabel pwell 187417 520770 187451 520804 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_18_Right_18.VNB
rlabel comment 187480 520787 187480 520787 8 dpga_flat_0.sr_0.PHY_EDGE_ROW_18_Right_18.decap_3
rlabel metal1 187204 520739 187480 520835 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_18_Right_18.VGND
rlabel metal1 187204 520195 187480 520291 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_18_Right_18.VPWR
flabel metal1 172513 519682 172547 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_3.VGND
flabel metal1 172513 520226 172547 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_3.VPWR
flabel nwell 172513 520226 172547 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_3.VPB
flabel pwell 172513 519682 172547 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_3.VNB
rlabel comment 172484 519699 172484 519699 4 dpga_flat_0.sr_0.FILLER_0_19_3.decap_12
flabel metal1 173617 519682 173651 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_15.VGND
flabel metal1 173617 520226 173651 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_15.VPWR
flabel nwell 173617 520226 173651 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_15.VPB
flabel pwell 173617 519682 173651 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_15.VNB
rlabel comment 173588 519699 173588 519699 4 dpga_flat_0.sr_0.FILLER_0_19_15.decap_12
flabel metal1 172513 519682 172547 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_3.VGND
flabel metal1 172513 519138 172547 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_3.VPWR
flabel nwell 172513 519138 172547 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_3.VPB
flabel pwell 172513 519682 172547 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_3.VNB
rlabel comment 172484 519699 172484 519699 2 dpga_flat_0.sr_0.FILLER_0_20_3.decap_12
flabel metal1 173617 519682 173651 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_15.VGND
flabel metal1 173617 519138 173651 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_15.VPWR
flabel nwell 173617 519138 173651 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_15.VPB
flabel pwell 173617 519682 173651 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_15.VNB
rlabel comment 173588 519699 173588 519699 2 dpga_flat_0.sr_0.FILLER_0_20_15.decap_12
flabel metal1 172237 520226 172271 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_19_Left_47.VPWR
flabel metal1 172237 519682 172271 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_19_Left_47.VGND
flabel nwell 172237 520226 172271 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_19_Left_47.VPB
flabel pwell 172237 519682 172271 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_19_Left_47.VNB
rlabel comment 172208 519699 172208 519699 4 dpga_flat_0.sr_0.PHY_EDGE_ROW_19_Left_47.decap_3
rlabel metal1 172208 519651 172484 519747 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_19_Left_47.VGND
rlabel metal1 172208 520195 172484 520291 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_19_Left_47.VPWR
flabel metal1 172237 519138 172271 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_20_Left_48.VPWR
flabel metal1 172237 519682 172271 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_20_Left_48.VGND
flabel nwell 172237 519138 172271 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_20_Left_48.VPB
flabel pwell 172237 519682 172271 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_20_Left_48.VNB
rlabel comment 172208 519699 172208 519699 2 dpga_flat_0.sr_0.PHY_EDGE_ROW_20_Left_48.decap_3
rlabel metal1 172208 519651 172484 519747 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_20_Left_48.VGND
rlabel metal1 172208 519107 172484 519203 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_20_Left_48.VPWR
flabel metal1 174721 519682 174755 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_27.VGND
flabel metal1 174721 520226 174755 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_27.VPWR
flabel nwell 174721 520226 174755 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_27.VPB
flabel pwell 174721 519682 174755 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_27.VNB
rlabel comment 174692 519699 174692 519699 4 dpga_flat_0.sr_0.FILLER_0_19_27.decap_12
flabel metal1 175825 519682 175859 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_39.VGND
flabel metal1 175825 520226 175859 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_39.VPWR
flabel nwell 175825 520226 175859 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_39.VPB
flabel pwell 175825 519682 175859 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_39.VNB
rlabel comment 175796 519699 175796 519699 4 dpga_flat_0.sr_0.FILLER_0_19_39.decap_12
flabel metal1 174714 519142 174750 519172 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_27.VPWR
flabel metal1 174714 519683 174750 519712 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_27.VGND
flabel nwell 174723 519148 174743 519165 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_27.VPB
flabel pwell 174720 519688 174744 519710 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_27.VNB
rlabel comment 174692 519699 174692 519699 2 dpga_flat_0.sr_0.FILLER_0_20_27.fill_1
rlabel metal1 174692 519651 174784 519747 5 dpga_flat_0.sr_0.FILLER_0_20_27.VGND
rlabel metal1 174692 519107 174784 519203 5 dpga_flat_0.sr_0.FILLER_0_20_27.VPWR
flabel metal1 174905 519682 174939 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_29.VGND
flabel metal1 174905 519138 174939 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_29.VPWR
flabel nwell 174905 519138 174939 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_29.VPB
flabel pwell 174905 519682 174939 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_29.VNB
rlabel comment 174876 519699 174876 519699 2 dpga_flat_0.sr_0.FILLER_0_20_29.decap_12
flabel metal1 176009 519682 176043 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_41.VGND
flabel metal1 176009 519138 176043 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_41.VPWR
flabel nwell 176009 519138 176043 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_41.VPB
flabel pwell 176009 519682 176043 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_41.VNB
rlabel comment 175980 519699 175980 519699 2 dpga_flat_0.sr_0.FILLER_0_20_41.decap_12
flabel metal1 174806 519146 174859 519175 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_20_108.VPWR
flabel metal1 174805 519679 174856 519717 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_20_108.VGND
rlabel comment 174784 519699 174784 519699 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_20_108.tapvpwrvgnd_1
rlabel metal1 174784 519651 174876 519747 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_20_108.VGND
rlabel metal1 174784 519107 174876 519203 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_20_108.VPWR
flabel metal1 176929 519682 176963 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_51.VGND
flabel metal1 176929 520226 176963 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_51.VPWR
flabel nwell 176929 520226 176963 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_51.VPB
flabel pwell 176929 519682 176963 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_51.VNB
rlabel comment 176900 519699 176900 519699 4 dpga_flat_0.sr_0.FILLER_0_19_51.decap_4
rlabel metal1 176900 519651 177268 519747 1 dpga_flat_0.sr_0.FILLER_0_19_51.VGND
rlabel metal1 176900 520195 177268 520291 1 dpga_flat_0.sr_0.FILLER_0_19_51.VPWR
flabel metal1 177290 520226 177326 520256 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_55.VPWR
flabel metal1 177290 519686 177326 519715 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_55.VGND
flabel nwell 177299 520233 177319 520250 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_55.VPB
flabel pwell 177296 519688 177320 519710 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_55.VNB
rlabel comment 177268 519699 177268 519699 4 dpga_flat_0.sr_0.FILLER_0_19_55.fill_1
rlabel metal1 177268 519651 177360 519747 1 dpga_flat_0.sr_0.FILLER_0_19_55.VGND
rlabel metal1 177268 520195 177360 520291 1 dpga_flat_0.sr_0.FILLER_0_19_55.VPWR
flabel metal1 177481 519682 177515 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_57.VGND
flabel metal1 177481 520226 177515 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_57.VPWR
flabel nwell 177481 520226 177515 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_57.VPB
flabel pwell 177481 519682 177515 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_57.VNB
rlabel comment 177452 519699 177452 519699 4 dpga_flat_0.sr_0.FILLER_0_19_57.decap_12
flabel metal1 177113 519682 177147 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_53.VGND
flabel metal1 177113 519138 177147 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_53.VPWR
flabel nwell 177113 519138 177147 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_53.VPB
flabel pwell 177113 519682 177147 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_53.VNB
rlabel comment 177084 519699 177084 519699 2 dpga_flat_0.sr_0.FILLER_0_20_53.decap_12
flabel metal1 177382 520223 177435 520252 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_19_106.VPWR
flabel metal1 177381 519681 177432 519719 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_19_106.VGND
rlabel comment 177360 519699 177360 519699 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_19_106.tapvpwrvgnd_1
rlabel metal1 177360 519651 177452 519747 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_19_106.VGND
rlabel metal1 177360 520195 177452 520291 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_19_106.VPWR
flabel metal1 178585 519682 178619 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_69.VGND
flabel metal1 178585 520226 178619 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_69.VPWR
flabel nwell 178585 520226 178619 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_69.VPB
flabel pwell 178585 519682 178619 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_69.VNB
rlabel comment 178556 519699 178556 519699 4 dpga_flat_0.sr_0.FILLER_0_19_69.decap_12
flabel metal1 179689 519682 179723 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_81.VGND
flabel metal1 179689 520226 179723 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_81.VPWR
flabel nwell 179689 520226 179723 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_81.VPB
flabel pwell 179689 519682 179723 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_81.VNB
rlabel comment 179660 519699 179660 519699 4 dpga_flat_0.sr_0.FILLER_0_19_81.decap_12
flabel metal1 178217 519682 178251 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_65.VGND
flabel metal1 178217 519138 178251 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_65.VPWR
flabel nwell 178217 519138 178251 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_65.VPB
flabel pwell 178217 519682 178251 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_65.VNB
rlabel comment 178188 519699 178188 519699 2 dpga_flat_0.sr_0.FILLER_0_20_65.decap_12
flabel metal1 179321 519138 179355 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_77.VPWR
flabel metal1 179321 519682 179355 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_77.VGND
flabel nwell 179321 519138 179355 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_77.VPB
flabel pwell 179321 519682 179355 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_77.VNB
rlabel comment 179292 519699 179292 519699 2 dpga_flat_0.sr_0.FILLER_0_20_77.decap_6
rlabel metal1 179292 519651 179844 519747 5 dpga_flat_0.sr_0.FILLER_0_20_77.VGND
rlabel metal1 179292 519107 179844 519203 5 dpga_flat_0.sr_0.FILLER_0_20_77.VPWR
flabel metal1 179866 519142 179902 519172 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_83.VPWR
flabel metal1 179866 519683 179902 519712 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_83.VGND
flabel nwell 179875 519148 179895 519165 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_83.VPB
flabel pwell 179872 519688 179896 519710 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_83.VNB
rlabel comment 179844 519699 179844 519699 2 dpga_flat_0.sr_0.FILLER_0_20_83.fill_1
rlabel metal1 179844 519651 179936 519747 5 dpga_flat_0.sr_0.FILLER_0_20_83.VGND
rlabel metal1 179844 519107 179936 519203 5 dpga_flat_0.sr_0.FILLER_0_20_83.VPWR
flabel metal1 180793 519682 180827 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_93.VGND
flabel metal1 180793 520226 180827 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_93.VPWR
flabel nwell 180793 520226 180827 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_93.VPB
flabel pwell 180793 519682 180827 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_93.VNB
rlabel comment 180764 519699 180764 519699 4 dpga_flat_0.sr_0.FILLER_0_19_93.decap_12
flabel metal1 180057 519682 180091 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_85.VGND
flabel metal1 180057 519138 180091 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_85.VPWR
flabel nwell 180057 519138 180091 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_85.VPB
flabel pwell 180057 519682 180091 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_85.VNB
rlabel comment 180028 519699 180028 519699 2 dpga_flat_0.sr_0.FILLER_0_20_85.decap_12
flabel metal1 181161 519682 181195 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_97.VGND
flabel metal1 181161 519138 181195 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_97.VPWR
flabel nwell 181161 519138 181195 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_97.VPB
flabel pwell 181161 519682 181195 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_97.VNB
rlabel comment 181132 519699 181132 519699 2 dpga_flat_0.sr_0.FILLER_0_20_97.decap_12
flabel metal1 179958 519146 180011 519175 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_20_109.VPWR
flabel metal1 179957 519679 180008 519717 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_20_109.VGND
rlabel comment 179936 519699 179936 519699 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_20_109.tapvpwrvgnd_1
rlabel metal1 179936 519651 180028 519747 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_20_109.VGND
rlabel metal1 179936 519107 180028 519203 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_20_109.VPWR
flabel metal1 181897 520226 181931 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_105.VPWR
flabel metal1 181897 519682 181931 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_105.VGND
flabel nwell 181897 520226 181931 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_105.VPB
flabel pwell 181897 519682 181931 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_105.VNB
rlabel comment 181868 519699 181868 519699 4 dpga_flat_0.sr_0.FILLER_0_19_105.decap_6
rlabel metal1 181868 519651 182420 519747 1 dpga_flat_0.sr_0.FILLER_0_19_105.VGND
rlabel metal1 181868 520195 182420 520291 1 dpga_flat_0.sr_0.FILLER_0_19_105.VPWR
flabel metal1 182442 520226 182478 520256 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_111.VPWR
flabel metal1 182442 519686 182478 519715 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_111.VGND
flabel nwell 182451 520233 182471 520250 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_111.VPB
flabel pwell 182448 519688 182472 519710 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_111.VNB
rlabel comment 182420 519699 182420 519699 4 dpga_flat_0.sr_0.FILLER_0_19_111.fill_1
rlabel metal1 182420 519651 182512 519747 1 dpga_flat_0.sr_0.FILLER_0_19_111.VGND
rlabel metal1 182420 520195 182512 520291 1 dpga_flat_0.sr_0.FILLER_0_19_111.VPWR
flabel metal1 182633 519682 182667 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_113.VGND
flabel metal1 182633 520226 182667 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_113.VPWR
flabel nwell 182633 520226 182667 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_113.VPB
flabel pwell 182633 519682 182667 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_113.VNB
rlabel comment 182604 519699 182604 519699 4 dpga_flat_0.sr_0.FILLER_0_19_113.decap_12
flabel metal1 183737 519682 183771 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_125.VGND
flabel metal1 183737 520226 183771 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_125.VPWR
flabel nwell 183737 520226 183771 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_125.VPB
flabel pwell 183737 519682 183771 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_125.VNB
rlabel comment 183708 519699 183708 519699 4 dpga_flat_0.sr_0.FILLER_0_19_125.decap_12
flabel metal1 182265 519682 182299 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_109.VGND
flabel metal1 182265 519138 182299 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_109.VPWR
flabel nwell 182265 519138 182299 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_109.VPB
flabel pwell 182265 519682 182299 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_109.VNB
rlabel comment 182236 519699 182236 519699 2 dpga_flat_0.sr_0.FILLER_0_20_109.decap_12
flabel metal1 183369 519682 183403 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_121.VGND
flabel metal1 183369 519138 183403 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_121.VPWR
flabel nwell 183369 519138 183403 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_121.VPB
flabel pwell 183369 519682 183403 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_121.VNB
rlabel comment 183340 519699 183340 519699 2 dpga_flat_0.sr_0.FILLER_0_20_121.decap_12
flabel metal1 182534 520223 182587 520252 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_19_107.VPWR
flabel metal1 182533 519681 182584 519719 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_19_107.VGND
rlabel comment 182512 519699 182512 519699 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_19_107.tapvpwrvgnd_1
rlabel metal1 182512 519651 182604 519747 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_19_107.VGND
rlabel metal1 182512 520195 182604 520291 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_19_107.VPWR
flabel metal1 184841 519682 184875 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_137.VGND
flabel metal1 184841 520226 184875 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_137.VPWR
flabel nwell 184841 520226 184875 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_137.VPB
flabel pwell 184841 519682 184875 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_137.VNB
rlabel comment 184812 519699 184812 519699 4 dpga_flat_0.sr_0.FILLER_0_19_137.decap_12
flabel metal1 184473 519138 184507 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_133.VPWR
flabel metal1 184473 519682 184507 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_133.VGND
flabel nwell 184473 519138 184507 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_133.VPB
flabel pwell 184473 519682 184507 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_133.VNB
rlabel comment 184444 519699 184444 519699 2 dpga_flat_0.sr_0.FILLER_0_20_133.decap_6
rlabel metal1 184444 519651 184996 519747 5 dpga_flat_0.sr_0.FILLER_0_20_133.VGND
rlabel metal1 184444 519107 184996 519203 5 dpga_flat_0.sr_0.FILLER_0_20_133.VPWR
flabel metal1 185018 519142 185054 519172 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_139.VPWR
flabel metal1 185018 519683 185054 519712 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_139.VGND
flabel nwell 185027 519148 185047 519165 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_139.VPB
flabel pwell 185024 519688 185048 519710 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_139.VNB
rlabel comment 184996 519699 184996 519699 2 dpga_flat_0.sr_0.FILLER_0_20_139.fill_1
rlabel metal1 184996 519651 185088 519747 5 dpga_flat_0.sr_0.FILLER_0_20_139.VGND
rlabel metal1 184996 519107 185088 519203 5 dpga_flat_0.sr_0.FILLER_0_20_139.VPWR
flabel metal1 185209 519682 185243 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_141.VGND
flabel metal1 185209 519138 185243 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_141.VPWR
flabel nwell 185209 519138 185243 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_141.VPB
flabel pwell 185209 519682 185243 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_141.VNB
rlabel comment 185180 519699 185180 519699 2 dpga_flat_0.sr_0.FILLER_0_20_141.decap_12
flabel metal1 185110 519146 185163 519175 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_20_110.VPWR
flabel metal1 185109 519679 185160 519717 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_20_110.VGND
rlabel comment 185088 519699 185088 519699 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_20_110.tapvpwrvgnd_1
rlabel metal1 185088 519651 185180 519747 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_20_110.VGND
rlabel metal1 185088 519107 185180 519203 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_20_110.VPWR
flabel metal1 185945 519682 185979 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_149.VGND
flabel metal1 185945 520226 185979 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_149.VPWR
flabel nwell 185945 520226 185979 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_149.VPB
flabel pwell 185945 519682 185979 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_149.VNB
rlabel comment 185916 519699 185916 519699 4 dpga_flat_0.sr_0.FILLER_0_19_149.decap_12
flabel metal1 187040 519685 187093 519717 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_161.VGND
flabel metal1 187041 520229 187093 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_161.VPWR
flabel nwell 187048 520234 187082 520252 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_161.VPB
flabel pwell 187051 519689 187083 519711 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_161.VNB
rlabel comment 187020 519699 187020 519699 4 dpga_flat_0.sr_0.FILLER_0_19_161.fill_2
rlabel metal1 187020 519651 187204 519747 1 dpga_flat_0.sr_0.FILLER_0_19_161.VGND
rlabel metal1 187020 520195 187204 520291 1 dpga_flat_0.sr_0.FILLER_0_19_161.VPWR
flabel metal1 186313 519138 186347 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_153.VPWR
flabel metal1 186313 519682 186347 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_153.VGND
flabel nwell 186313 519138 186347 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_153.VPB
flabel pwell 186313 519682 186347 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_153.VNB
rlabel comment 186284 519699 186284 519699 2 dpga_flat_0.sr_0.FILLER_0_20_153.decap_8
rlabel metal1 186284 519651 187020 519747 5 dpga_flat_0.sr_0.FILLER_0_20_153.VGND
rlabel metal1 186284 519107 187020 519203 5 dpga_flat_0.sr_0.FILLER_0_20_153.VPWR
flabel metal1 187040 519681 187093 519713 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_161.VGND
flabel metal1 187041 519138 187093 519169 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_161.VPWR
flabel nwell 187048 519146 187082 519164 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_161.VPB
flabel pwell 187051 519687 187083 519709 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_161.VNB
rlabel comment 187020 519699 187020 519699 2 dpga_flat_0.sr_0.FILLER_0_20_161.fill_2
rlabel metal1 187020 519651 187204 519747 5 dpga_flat_0.sr_0.FILLER_0_20_161.VGND
rlabel metal1 187020 519107 187204 519203 5 dpga_flat_0.sr_0.FILLER_0_20_161.VPWR
flabel metal1 187417 520226 187451 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_19_Right_19.VPWR
flabel metal1 187417 519682 187451 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_19_Right_19.VGND
flabel nwell 187417 520226 187451 520260 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_19_Right_19.VPB
flabel pwell 187417 519682 187451 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_19_Right_19.VNB
rlabel comment 187480 519699 187480 519699 6 dpga_flat_0.sr_0.PHY_EDGE_ROW_19_Right_19.decap_3
rlabel metal1 187204 519651 187480 519747 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_19_Right_19.VGND
rlabel metal1 187204 520195 187480 520291 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_19_Right_19.VPWR
flabel metal1 187417 519138 187451 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_20_Right_20.VPWR
flabel metal1 187417 519682 187451 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_20_Right_20.VGND
flabel nwell 187417 519138 187451 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_20_Right_20.VPB
flabel pwell 187417 519682 187451 519716 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_20_Right_20.VNB
rlabel comment 187480 519699 187480 519699 8 dpga_flat_0.sr_0.PHY_EDGE_ROW_20_Right_20.decap_3
rlabel metal1 187204 519651 187480 519747 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_20_Right_20.VGND
rlabel metal1 187204 519107 187480 519203 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_20_Right_20.VPWR
flabel metal1 172513 518594 172547 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_3.VGND
flabel metal1 172513 519138 172547 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_3.VPWR
flabel nwell 172513 519138 172547 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_3.VPB
flabel pwell 172513 518594 172547 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_3.VNB
rlabel comment 172484 518611 172484 518611 4 dpga_flat_0.sr_0.FILLER_0_21_3.decap_12
flabel metal1 173617 518594 173651 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_15.VGND
flabel metal1 173617 519138 173651 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_15.VPWR
flabel nwell 173617 519138 173651 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_15.VPB
flabel pwell 173617 518594 173651 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_15.VNB
rlabel comment 173588 518611 173588 518611 4 dpga_flat_0.sr_0.FILLER_0_21_15.decap_12
flabel metal1 172237 519138 172271 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_21_Left_49.VPWR
flabel metal1 172237 518594 172271 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_21_Left_49.VGND
flabel nwell 172237 519138 172271 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_21_Left_49.VPB
flabel pwell 172237 518594 172271 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_21_Left_49.VNB
rlabel comment 172208 518611 172208 518611 4 dpga_flat_0.sr_0.PHY_EDGE_ROW_21_Left_49.decap_3
rlabel metal1 172208 518563 172484 518659 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_21_Left_49.VGND
rlabel metal1 172208 519107 172484 519203 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_21_Left_49.VPWR
flabel metal1 174721 518594 174755 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_27.VGND
flabel metal1 174721 519138 174755 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_27.VPWR
flabel nwell 174721 519138 174755 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_27.VPB
flabel pwell 174721 518594 174755 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_27.VNB
rlabel comment 174692 518611 174692 518611 4 dpga_flat_0.sr_0.FILLER_0_21_27.decap_12
flabel metal1 175825 518594 175859 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_39.VGND
flabel metal1 175825 519138 175859 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_39.VPWR
flabel nwell 175825 519138 175859 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_39.VPB
flabel pwell 175825 518594 175859 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_39.VNB
rlabel comment 175796 518611 175796 518611 4 dpga_flat_0.sr_0.FILLER_0_21_39.decap_12
flabel metal1 176929 518594 176963 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_51.VGND
flabel metal1 176929 519138 176963 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_51.VPWR
flabel nwell 176929 519138 176963 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_51.VPB
flabel pwell 176929 518594 176963 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_51.VNB
rlabel comment 176900 518611 176900 518611 4 dpga_flat_0.sr_0.FILLER_0_21_51.decap_4
rlabel metal1 176900 518563 177268 518659 1 dpga_flat_0.sr_0.FILLER_0_21_51.VGND
rlabel metal1 176900 519107 177268 519203 1 dpga_flat_0.sr_0.FILLER_0_21_51.VPWR
flabel metal1 177290 519138 177326 519168 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_55.VPWR
flabel metal1 177290 518598 177326 518627 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_55.VGND
flabel nwell 177299 519145 177319 519162 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_55.VPB
flabel pwell 177296 518600 177320 518622 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_55.VNB
rlabel comment 177268 518611 177268 518611 4 dpga_flat_0.sr_0.FILLER_0_21_55.fill_1
rlabel metal1 177268 518563 177360 518659 1 dpga_flat_0.sr_0.FILLER_0_21_55.VGND
rlabel metal1 177268 519107 177360 519203 1 dpga_flat_0.sr_0.FILLER_0_21_55.VPWR
flabel metal1 177481 518594 177515 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_57.VGND
flabel metal1 177481 519138 177515 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_57.VPWR
flabel nwell 177481 519138 177515 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_57.VPB
flabel pwell 177481 518594 177515 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_57.VNB
rlabel comment 177452 518611 177452 518611 4 dpga_flat_0.sr_0.FILLER_0_21_57.decap_12
flabel metal1 177382 519135 177435 519164 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_21_111.VPWR
flabel metal1 177381 518593 177432 518631 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_21_111.VGND
rlabel comment 177360 518611 177360 518611 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_21_111.tapvpwrvgnd_1
rlabel metal1 177360 518563 177452 518659 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_21_111.VGND
rlabel metal1 177360 519107 177452 519203 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_21_111.VPWR
flabel metal1 178585 518594 178619 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_69.VGND
flabel metal1 178585 519138 178619 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_69.VPWR
flabel nwell 178585 519138 178619 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_69.VPB
flabel pwell 178585 518594 178619 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_69.VNB
rlabel comment 178556 518611 178556 518611 4 dpga_flat_0.sr_0.FILLER_0_21_69.decap_12
flabel metal1 179689 518594 179723 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_81.VGND
flabel metal1 179689 519138 179723 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_81.VPWR
flabel nwell 179689 519138 179723 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_81.VPB
flabel pwell 179689 518594 179723 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_81.VNB
rlabel comment 179660 518611 179660 518611 4 dpga_flat_0.sr_0.FILLER_0_21_81.decap_12
flabel metal1 180793 518594 180827 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_93.VGND
flabel metal1 180793 519138 180827 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_93.VPWR
flabel nwell 180793 519138 180827 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_93.VPB
flabel pwell 180793 518594 180827 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_93.VNB
rlabel comment 180764 518611 180764 518611 4 dpga_flat_0.sr_0.FILLER_0_21_93.decap_12
flabel metal1 181897 519138 181931 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_105.VPWR
flabel metal1 181897 518594 181931 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_105.VGND
flabel nwell 181897 519138 181931 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_105.VPB
flabel pwell 181897 518594 181931 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_105.VNB
rlabel comment 181868 518611 181868 518611 4 dpga_flat_0.sr_0.FILLER_0_21_105.decap_6
rlabel metal1 181868 518563 182420 518659 1 dpga_flat_0.sr_0.FILLER_0_21_105.VGND
rlabel metal1 181868 519107 182420 519203 1 dpga_flat_0.sr_0.FILLER_0_21_105.VPWR
flabel metal1 182442 519138 182478 519168 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_111.VPWR
flabel metal1 182442 518598 182478 518627 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_111.VGND
flabel nwell 182451 519145 182471 519162 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_111.VPB
flabel pwell 182448 518600 182472 518622 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_111.VNB
rlabel comment 182420 518611 182420 518611 4 dpga_flat_0.sr_0.FILLER_0_21_111.fill_1
rlabel metal1 182420 518563 182512 518659 1 dpga_flat_0.sr_0.FILLER_0_21_111.VGND
rlabel metal1 182420 519107 182512 519203 1 dpga_flat_0.sr_0.FILLER_0_21_111.VPWR
flabel metal1 182633 518594 182667 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_113.VGND
flabel metal1 182633 519138 182667 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_113.VPWR
flabel nwell 182633 519138 182667 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_113.VPB
flabel pwell 182633 518594 182667 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_113.VNB
rlabel comment 182604 518611 182604 518611 4 dpga_flat_0.sr_0.FILLER_0_21_113.decap_12
flabel metal1 183737 518594 183771 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_125.VGND
flabel metal1 183737 519138 183771 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_125.VPWR
flabel nwell 183737 519138 183771 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_125.VPB
flabel pwell 183737 518594 183771 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_125.VNB
rlabel comment 183708 518611 183708 518611 4 dpga_flat_0.sr_0.FILLER_0_21_125.decap_12
flabel metal1 182534 519135 182587 519164 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_21_112.VPWR
flabel metal1 182533 518593 182584 518631 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_21_112.VGND
rlabel comment 182512 518611 182512 518611 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_21_112.tapvpwrvgnd_1
rlabel metal1 182512 518563 182604 518659 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_21_112.VGND
rlabel metal1 182512 519107 182604 519203 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_21_112.VPWR
flabel metal1 184841 518594 184875 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_137.VGND
flabel metal1 184841 519138 184875 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_137.VPWR
flabel nwell 184841 519138 184875 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_137.VPB
flabel pwell 184841 518594 184875 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_137.VNB
rlabel comment 184812 518611 184812 518611 4 dpga_flat_0.sr_0.FILLER_0_21_137.decap_12
flabel metal1 185945 518594 185979 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_149.VGND
flabel metal1 185945 519138 185979 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_149.VPWR
flabel nwell 185945 519138 185979 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_149.VPB
flabel pwell 185945 518594 185979 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_149.VNB
rlabel comment 185916 518611 185916 518611 4 dpga_flat_0.sr_0.FILLER_0_21_149.decap_12
flabel metal1 187040 518597 187093 518629 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_161.VGND
flabel metal1 187041 519141 187093 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_161.VPWR
flabel nwell 187048 519146 187082 519164 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_161.VPB
flabel pwell 187051 518601 187083 518623 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_161.VNB
rlabel comment 187020 518611 187020 518611 4 dpga_flat_0.sr_0.FILLER_0_21_161.fill_2
rlabel metal1 187020 518563 187204 518659 1 dpga_flat_0.sr_0.FILLER_0_21_161.VGND
rlabel metal1 187020 519107 187204 519203 1 dpga_flat_0.sr_0.FILLER_0_21_161.VPWR
flabel metal1 187417 519138 187451 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_21_Right_21.VPWR
flabel metal1 187417 518594 187451 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_21_Right_21.VGND
flabel nwell 187417 519138 187451 519172 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_21_Right_21.VPB
flabel pwell 187417 518594 187451 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_21_Right_21.VNB
rlabel comment 187480 518611 187480 518611 6 dpga_flat_0.sr_0.PHY_EDGE_ROW_21_Right_21.decap_3
rlabel metal1 187204 518563 187480 518659 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_21_Right_21.VGND
rlabel metal1 187204 519107 187480 519203 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_21_Right_21.VPWR
flabel metal1 172513 518594 172547 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_3.VGND
flabel metal1 172513 518050 172547 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_3.VPWR
flabel nwell 172513 518050 172547 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_3.VPB
flabel pwell 172513 518594 172547 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_3.VNB
rlabel comment 172484 518611 172484 518611 2 dpga_flat_0.sr_0.FILLER_0_22_3.decap_12
flabel metal1 173617 518594 173651 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_15.VGND
flabel metal1 173617 518050 173651 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_15.VPWR
flabel nwell 173617 518050 173651 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_15.VPB
flabel pwell 173617 518594 173651 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_15.VNB
rlabel comment 173588 518611 173588 518611 2 dpga_flat_0.sr_0.FILLER_0_22_15.decap_12
flabel metal1 172237 518050 172271 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_22_Left_50.VPWR
flabel metal1 172237 518594 172271 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_22_Left_50.VGND
flabel nwell 172237 518050 172271 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_22_Left_50.VPB
flabel pwell 172237 518594 172271 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_22_Left_50.VNB
rlabel comment 172208 518611 172208 518611 2 dpga_flat_0.sr_0.PHY_EDGE_ROW_22_Left_50.decap_3
rlabel metal1 172208 518563 172484 518659 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_22_Left_50.VGND
rlabel metal1 172208 518019 172484 518115 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_22_Left_50.VPWR
flabel metal1 174714 518054 174750 518084 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_27.VPWR
flabel metal1 174714 518595 174750 518624 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_27.VGND
flabel nwell 174723 518060 174743 518077 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_27.VPB
flabel pwell 174720 518600 174744 518622 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_27.VNB
rlabel comment 174692 518611 174692 518611 2 dpga_flat_0.sr_0.FILLER_0_22_27.fill_1
rlabel metal1 174692 518563 174784 518659 5 dpga_flat_0.sr_0.FILLER_0_22_27.VGND
rlabel metal1 174692 518019 174784 518115 5 dpga_flat_0.sr_0.FILLER_0_22_27.VPWR
flabel metal1 174905 518594 174939 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_29.VGND
flabel metal1 174905 518050 174939 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_29.VPWR
flabel nwell 174905 518050 174939 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_29.VPB
flabel pwell 174905 518594 174939 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_29.VNB
rlabel comment 174876 518611 174876 518611 2 dpga_flat_0.sr_0.FILLER_0_22_29.decap_12
flabel metal1 176009 518594 176043 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_41.VGND
flabel metal1 176009 518050 176043 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_41.VPWR
flabel nwell 176009 518050 176043 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_41.VPB
flabel pwell 176009 518594 176043 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_41.VNB
rlabel comment 175980 518611 175980 518611 2 dpga_flat_0.sr_0.FILLER_0_22_41.decap_12
flabel metal1 174806 518058 174859 518087 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_22_113.VPWR
flabel metal1 174805 518591 174856 518629 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_22_113.VGND
rlabel comment 174784 518611 174784 518611 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_22_113.tapvpwrvgnd_1
rlabel metal1 174784 518563 174876 518659 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_22_113.VGND
rlabel metal1 174784 518019 174876 518115 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_22_113.VPWR
flabel metal1 177113 518594 177147 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_53.VGND
flabel metal1 177113 518050 177147 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_53.VPWR
flabel nwell 177113 518050 177147 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_53.VPB
flabel pwell 177113 518594 177147 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_53.VNB
rlabel comment 177084 518611 177084 518611 2 dpga_flat_0.sr_0.FILLER_0_22_53.decap_12
flabel metal1 178217 518594 178251 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_65.VGND
flabel metal1 178217 518050 178251 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_65.VPWR
flabel nwell 178217 518050 178251 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_65.VPB
flabel pwell 178217 518594 178251 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_65.VNB
rlabel comment 178188 518611 178188 518611 2 dpga_flat_0.sr_0.FILLER_0_22_65.decap_12
flabel metal1 179321 518050 179355 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_77.VPWR
flabel metal1 179321 518594 179355 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_77.VGND
flabel nwell 179321 518050 179355 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_77.VPB
flabel pwell 179321 518594 179355 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_77.VNB
rlabel comment 179292 518611 179292 518611 2 dpga_flat_0.sr_0.FILLER_0_22_77.decap_6
rlabel metal1 179292 518563 179844 518659 5 dpga_flat_0.sr_0.FILLER_0_22_77.VGND
rlabel metal1 179292 518019 179844 518115 5 dpga_flat_0.sr_0.FILLER_0_22_77.VPWR
flabel metal1 179866 518054 179902 518084 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_83.VPWR
flabel metal1 179866 518595 179902 518624 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_83.VGND
flabel nwell 179875 518060 179895 518077 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_83.VPB
flabel pwell 179872 518600 179896 518622 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_83.VNB
rlabel comment 179844 518611 179844 518611 2 dpga_flat_0.sr_0.FILLER_0_22_83.fill_1
rlabel metal1 179844 518563 179936 518659 5 dpga_flat_0.sr_0.FILLER_0_22_83.VGND
rlabel metal1 179844 518019 179936 518115 5 dpga_flat_0.sr_0.FILLER_0_22_83.VPWR
flabel metal1 180057 518594 180091 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_85.VGND
flabel metal1 180057 518050 180091 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_85.VPWR
flabel nwell 180057 518050 180091 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_85.VPB
flabel pwell 180057 518594 180091 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_85.VNB
rlabel comment 180028 518611 180028 518611 2 dpga_flat_0.sr_0.FILLER_0_22_85.decap_12
flabel metal1 181161 518594 181195 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_97.VGND
flabel metal1 181161 518050 181195 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_97.VPWR
flabel nwell 181161 518050 181195 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_97.VPB
flabel pwell 181161 518594 181195 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_97.VNB
rlabel comment 181132 518611 181132 518611 2 dpga_flat_0.sr_0.FILLER_0_22_97.decap_12
flabel metal1 179958 518058 180011 518087 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_22_114.VPWR
flabel metal1 179957 518591 180008 518629 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_22_114.VGND
rlabel comment 179936 518611 179936 518611 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_22_114.tapvpwrvgnd_1
rlabel metal1 179936 518563 180028 518659 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_22_114.VGND
rlabel metal1 179936 518019 180028 518115 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_22_114.VPWR
flabel metal1 182265 518594 182299 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_109.VGND
flabel metal1 182265 518050 182299 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_109.VPWR
flabel nwell 182265 518050 182299 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_109.VPB
flabel pwell 182265 518594 182299 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_109.VNB
rlabel comment 182236 518611 182236 518611 2 dpga_flat_0.sr_0.FILLER_0_22_109.decap_12
flabel metal1 183369 518594 183403 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_121.VGND
flabel metal1 183369 518050 183403 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_121.VPWR
flabel nwell 183369 518050 183403 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_121.VPB
flabel pwell 183369 518594 183403 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_121.VNB
rlabel comment 183340 518611 183340 518611 2 dpga_flat_0.sr_0.FILLER_0_22_121.decap_12
flabel metal1 184473 518050 184507 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_133.VPWR
flabel metal1 184473 518594 184507 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_133.VGND
flabel nwell 184473 518050 184507 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_133.VPB
flabel pwell 184473 518594 184507 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_133.VNB
rlabel comment 184444 518611 184444 518611 2 dpga_flat_0.sr_0.FILLER_0_22_133.decap_6
rlabel metal1 184444 518563 184996 518659 5 dpga_flat_0.sr_0.FILLER_0_22_133.VGND
rlabel metal1 184444 518019 184996 518115 5 dpga_flat_0.sr_0.FILLER_0_22_133.VPWR
flabel metal1 185018 518054 185054 518084 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_139.VPWR
flabel metal1 185018 518595 185054 518624 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_139.VGND
flabel nwell 185027 518060 185047 518077 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_139.VPB
flabel pwell 185024 518600 185048 518622 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_139.VNB
rlabel comment 184996 518611 184996 518611 2 dpga_flat_0.sr_0.FILLER_0_22_139.fill_1
rlabel metal1 184996 518563 185088 518659 5 dpga_flat_0.sr_0.FILLER_0_22_139.VGND
rlabel metal1 184996 518019 185088 518115 5 dpga_flat_0.sr_0.FILLER_0_22_139.VPWR
flabel metal1 185209 518594 185243 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_141.VGND
flabel metal1 185209 518050 185243 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_141.VPWR
flabel nwell 185209 518050 185243 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_141.VPB
flabel pwell 185209 518594 185243 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_141.VNB
rlabel comment 185180 518611 185180 518611 2 dpga_flat_0.sr_0.FILLER_0_22_141.decap_12
flabel metal1 185110 518058 185163 518087 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_22_115.VPWR
flabel metal1 185109 518591 185160 518629 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_22_115.VGND
rlabel comment 185088 518611 185088 518611 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_22_115.tapvpwrvgnd_1
rlabel metal1 185088 518563 185180 518659 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_22_115.VGND
rlabel metal1 185088 518019 185180 518115 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_22_115.VPWR
flabel metal1 186313 518050 186347 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_153.VPWR
flabel metal1 186313 518594 186347 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_153.VGND
flabel nwell 186313 518050 186347 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_153.VPB
flabel pwell 186313 518594 186347 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_153.VNB
rlabel comment 186284 518611 186284 518611 2 dpga_flat_0.sr_0.FILLER_0_22_153.decap_8
rlabel metal1 186284 518563 187020 518659 5 dpga_flat_0.sr_0.FILLER_0_22_153.VGND
rlabel metal1 186284 518019 187020 518115 5 dpga_flat_0.sr_0.FILLER_0_22_153.VPWR
flabel metal1 187040 518593 187093 518625 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_161.VGND
flabel metal1 187041 518050 187093 518081 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_161.VPWR
flabel nwell 187048 518058 187082 518076 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_161.VPB
flabel pwell 187051 518599 187083 518621 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_161.VNB
rlabel comment 187020 518611 187020 518611 2 dpga_flat_0.sr_0.FILLER_0_22_161.fill_2
rlabel metal1 187020 518563 187204 518659 5 dpga_flat_0.sr_0.FILLER_0_22_161.VGND
rlabel metal1 187020 518019 187204 518115 5 dpga_flat_0.sr_0.FILLER_0_22_161.VPWR
flabel metal1 187417 518050 187451 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_22_Right_22.VPWR
flabel metal1 187417 518594 187451 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_22_Right_22.VGND
flabel nwell 187417 518050 187451 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_22_Right_22.VPB
flabel pwell 187417 518594 187451 518628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_22_Right_22.VNB
rlabel comment 187480 518611 187480 518611 8 dpga_flat_0.sr_0.PHY_EDGE_ROW_22_Right_22.decap_3
rlabel metal1 187204 518563 187480 518659 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_22_Right_22.VGND
rlabel metal1 187204 518019 187480 518115 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_22_Right_22.VPWR
flabel metal1 172513 517506 172547 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_3.VGND
flabel metal1 172513 518050 172547 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_3.VPWR
flabel nwell 172513 518050 172547 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_3.VPB
flabel pwell 172513 517506 172547 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_3.VNB
rlabel comment 172484 517523 172484 517523 4 dpga_flat_0.sr_0.FILLER_0_23_3.decap_12
flabel metal1 173617 517506 173651 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_15.VGND
flabel metal1 173617 518050 173651 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_15.VPWR
flabel nwell 173617 518050 173651 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_15.VPB
flabel pwell 173617 517506 173651 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_15.VNB
rlabel comment 173588 517523 173588 517523 4 dpga_flat_0.sr_0.FILLER_0_23_15.decap_12
flabel metal1 172237 518050 172271 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_23_Left_51.VPWR
flabel metal1 172237 517506 172271 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_23_Left_51.VGND
flabel nwell 172237 518050 172271 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_23_Left_51.VPB
flabel pwell 172237 517506 172271 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_23_Left_51.VNB
rlabel comment 172208 517523 172208 517523 4 dpga_flat_0.sr_0.PHY_EDGE_ROW_23_Left_51.decap_3
rlabel metal1 172208 517475 172484 517571 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_23_Left_51.VGND
rlabel metal1 172208 518019 172484 518115 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_23_Left_51.VPWR
flabel metal1 174721 517506 174755 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_27.VGND
flabel metal1 174721 518050 174755 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_27.VPWR
flabel nwell 174721 518050 174755 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_27.VPB
flabel pwell 174721 517506 174755 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_27.VNB
rlabel comment 174692 517523 174692 517523 4 dpga_flat_0.sr_0.FILLER_0_23_27.decap_12
flabel metal1 175825 517506 175859 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_39.VGND
flabel metal1 175825 518050 175859 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_39.VPWR
flabel nwell 175825 518050 175859 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_39.VPB
flabel pwell 175825 517506 175859 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_39.VNB
rlabel comment 175796 517523 175796 517523 4 dpga_flat_0.sr_0.FILLER_0_23_39.decap_12
flabel metal1 176929 517506 176963 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_51.VGND
flabel metal1 176929 518050 176963 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_51.VPWR
flabel nwell 176929 518050 176963 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_51.VPB
flabel pwell 176929 517506 176963 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_51.VNB
rlabel comment 176900 517523 176900 517523 4 dpga_flat_0.sr_0.FILLER_0_23_51.decap_4
rlabel metal1 176900 517475 177268 517571 1 dpga_flat_0.sr_0.FILLER_0_23_51.VGND
rlabel metal1 176900 518019 177268 518115 1 dpga_flat_0.sr_0.FILLER_0_23_51.VPWR
flabel metal1 177290 518050 177326 518080 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_55.VPWR
flabel metal1 177290 517510 177326 517539 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_55.VGND
flabel nwell 177299 518057 177319 518074 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_55.VPB
flabel pwell 177296 517512 177320 517534 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_55.VNB
rlabel comment 177268 517523 177268 517523 4 dpga_flat_0.sr_0.FILLER_0_23_55.fill_1
rlabel metal1 177268 517475 177360 517571 1 dpga_flat_0.sr_0.FILLER_0_23_55.VGND
rlabel metal1 177268 518019 177360 518115 1 dpga_flat_0.sr_0.FILLER_0_23_55.VPWR
flabel metal1 177481 517506 177515 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_57.VGND
flabel metal1 177481 518050 177515 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_57.VPWR
flabel nwell 177481 518050 177515 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_57.VPB
flabel pwell 177481 517506 177515 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_57.VNB
rlabel comment 177452 517523 177452 517523 4 dpga_flat_0.sr_0.FILLER_0_23_57.decap_12
flabel metal1 177382 518047 177435 518076 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_23_116.VPWR
flabel metal1 177381 517505 177432 517543 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_23_116.VGND
rlabel comment 177360 517523 177360 517523 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_23_116.tapvpwrvgnd_1
rlabel metal1 177360 517475 177452 517571 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_23_116.VGND
rlabel metal1 177360 518019 177452 518115 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_23_116.VPWR
flabel metal1 178585 517506 178619 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_69.VGND
flabel metal1 178585 518050 178619 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_69.VPWR
flabel nwell 178585 518050 178619 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_69.VPB
flabel pwell 178585 517506 178619 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_69.VNB
rlabel comment 178556 517523 178556 517523 4 dpga_flat_0.sr_0.FILLER_0_23_69.decap_12
flabel metal1 179689 517506 179723 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_81.VGND
flabel metal1 179689 518050 179723 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_81.VPWR
flabel nwell 179689 518050 179723 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_81.VPB
flabel pwell 179689 517506 179723 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_81.VNB
rlabel comment 179660 517523 179660 517523 4 dpga_flat_0.sr_0.FILLER_0_23_81.decap_12
flabel metal1 180793 517506 180827 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_93.VGND
flabel metal1 180793 518050 180827 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_93.VPWR
flabel nwell 180793 518050 180827 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_93.VPB
flabel pwell 180793 517506 180827 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_93.VNB
rlabel comment 180764 517523 180764 517523 4 dpga_flat_0.sr_0.FILLER_0_23_93.decap_12
flabel metal1 181897 518050 181931 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_105.VPWR
flabel metal1 181897 517506 181931 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_105.VGND
flabel nwell 181897 518050 181931 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_105.VPB
flabel pwell 181897 517506 181931 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_105.VNB
rlabel comment 181868 517523 181868 517523 4 dpga_flat_0.sr_0.FILLER_0_23_105.decap_6
rlabel metal1 181868 517475 182420 517571 1 dpga_flat_0.sr_0.FILLER_0_23_105.VGND
rlabel metal1 181868 518019 182420 518115 1 dpga_flat_0.sr_0.FILLER_0_23_105.VPWR
flabel metal1 182442 518050 182478 518080 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_111.VPWR
flabel metal1 182442 517510 182478 517539 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_111.VGND
flabel nwell 182451 518057 182471 518074 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_111.VPB
flabel pwell 182448 517512 182472 517534 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_111.VNB
rlabel comment 182420 517523 182420 517523 4 dpga_flat_0.sr_0.FILLER_0_23_111.fill_1
rlabel metal1 182420 517475 182512 517571 1 dpga_flat_0.sr_0.FILLER_0_23_111.VGND
rlabel metal1 182420 518019 182512 518115 1 dpga_flat_0.sr_0.FILLER_0_23_111.VPWR
flabel metal1 182633 517506 182667 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_113.VGND
flabel metal1 182633 518050 182667 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_113.VPWR
flabel nwell 182633 518050 182667 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_113.VPB
flabel pwell 182633 517506 182667 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_113.VNB
rlabel comment 182604 517523 182604 517523 4 dpga_flat_0.sr_0.FILLER_0_23_113.decap_12
flabel metal1 183737 517506 183771 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_125.VGND
flabel metal1 183737 518050 183771 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_125.VPWR
flabel nwell 183737 518050 183771 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_125.VPB
flabel pwell 183737 517506 183771 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_125.VNB
rlabel comment 183708 517523 183708 517523 4 dpga_flat_0.sr_0.FILLER_0_23_125.decap_12
flabel metal1 182534 518047 182587 518076 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_23_117.VPWR
flabel metal1 182533 517505 182584 517543 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_23_117.VGND
rlabel comment 182512 517523 182512 517523 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_23_117.tapvpwrvgnd_1
rlabel metal1 182512 517475 182604 517571 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_23_117.VGND
rlabel metal1 182512 518019 182604 518115 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_23_117.VPWR
flabel metal1 184841 517506 184875 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_137.VGND
flabel metal1 184841 518050 184875 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_137.VPWR
flabel nwell 184841 518050 184875 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_137.VPB
flabel pwell 184841 517506 184875 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_137.VNB
rlabel comment 184812 517523 184812 517523 4 dpga_flat_0.sr_0.FILLER_0_23_137.decap_12
flabel metal1 185945 517506 185979 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_149.VGND
flabel metal1 185945 518050 185979 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_149.VPWR
flabel nwell 185945 518050 185979 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_149.VPB
flabel pwell 185945 517506 185979 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_149.VNB
rlabel comment 185916 517523 185916 517523 4 dpga_flat_0.sr_0.FILLER_0_23_149.decap_12
flabel metal1 187040 517509 187093 517541 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_161.VGND
flabel metal1 187041 518053 187093 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_161.VPWR
flabel nwell 187048 518058 187082 518076 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_161.VPB
flabel pwell 187051 517513 187083 517535 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_161.VNB
rlabel comment 187020 517523 187020 517523 4 dpga_flat_0.sr_0.FILLER_0_23_161.fill_2
rlabel metal1 187020 517475 187204 517571 1 dpga_flat_0.sr_0.FILLER_0_23_161.VGND
rlabel metal1 187020 518019 187204 518115 1 dpga_flat_0.sr_0.FILLER_0_23_161.VPWR
flabel metal1 187417 518050 187451 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_23_Right_23.VPWR
flabel metal1 187417 517506 187451 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_23_Right_23.VGND
flabel nwell 187417 518050 187451 518084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_23_Right_23.VPB
flabel pwell 187417 517506 187451 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_23_Right_23.VNB
rlabel comment 187480 517523 187480 517523 6 dpga_flat_0.sr_0.PHY_EDGE_ROW_23_Right_23.decap_3
rlabel metal1 187204 517475 187480 517571 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_23_Right_23.VGND
rlabel metal1 187204 518019 187480 518115 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_23_Right_23.VPWR
flabel metal1 172513 517506 172547 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_3.VGND
flabel metal1 172513 516962 172547 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_3.VPWR
flabel nwell 172513 516962 172547 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_3.VPB
flabel pwell 172513 517506 172547 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_3.VNB
rlabel comment 172484 517523 172484 517523 2 dpga_flat_0.sr_0.FILLER_0_24_3.decap_12
flabel metal1 173617 517506 173651 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_15.VGND
flabel metal1 173617 516962 173651 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_15.VPWR
flabel nwell 173617 516962 173651 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_15.VPB
flabel pwell 173617 517506 173651 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_15.VNB
rlabel comment 173588 517523 173588 517523 2 dpga_flat_0.sr_0.FILLER_0_24_15.decap_12
flabel metal1 172237 516962 172271 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_24_Left_52.VPWR
flabel metal1 172237 517506 172271 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_24_Left_52.VGND
flabel nwell 172237 516962 172271 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_24_Left_52.VPB
flabel pwell 172237 517506 172271 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_24_Left_52.VNB
rlabel comment 172208 517523 172208 517523 2 dpga_flat_0.sr_0.PHY_EDGE_ROW_24_Left_52.decap_3
rlabel metal1 172208 517475 172484 517571 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_24_Left_52.VGND
rlabel metal1 172208 516931 172484 517027 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_24_Left_52.VPWR
flabel metal1 174714 516966 174750 516996 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_27.VPWR
flabel metal1 174714 517507 174750 517536 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_27.VGND
flabel nwell 174723 516972 174743 516989 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_27.VPB
flabel pwell 174720 517512 174744 517534 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_27.VNB
rlabel comment 174692 517523 174692 517523 2 dpga_flat_0.sr_0.FILLER_0_24_27.fill_1
rlabel metal1 174692 517475 174784 517571 5 dpga_flat_0.sr_0.FILLER_0_24_27.VGND
rlabel metal1 174692 516931 174784 517027 5 dpga_flat_0.sr_0.FILLER_0_24_27.VPWR
flabel metal1 174905 517506 174939 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_29.VGND
flabel metal1 174905 516962 174939 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_29.VPWR
flabel nwell 174905 516962 174939 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_29.VPB
flabel pwell 174905 517506 174939 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_29.VNB
rlabel comment 174876 517523 174876 517523 2 dpga_flat_0.sr_0.FILLER_0_24_29.decap_12
flabel metal1 176009 517506 176043 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_41.VGND
flabel metal1 176009 516962 176043 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_41.VPWR
flabel nwell 176009 516962 176043 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_41.VPB
flabel pwell 176009 517506 176043 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_41.VNB
rlabel comment 175980 517523 175980 517523 2 dpga_flat_0.sr_0.FILLER_0_24_41.decap_12
flabel metal1 174806 516970 174859 516999 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_24_118.VPWR
flabel metal1 174805 517503 174856 517541 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_24_118.VGND
rlabel comment 174784 517523 174784 517523 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_24_118.tapvpwrvgnd_1
rlabel metal1 174784 517475 174876 517571 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_24_118.VGND
rlabel metal1 174784 516931 174876 517027 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_24_118.VPWR
flabel metal1 177113 517506 177147 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_53.VGND
flabel metal1 177113 516962 177147 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_53.VPWR
flabel nwell 177113 516962 177147 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_53.VPB
flabel pwell 177113 517506 177147 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_53.VNB
rlabel comment 177084 517523 177084 517523 2 dpga_flat_0.sr_0.FILLER_0_24_53.decap_12
flabel metal1 178217 517506 178251 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_65.VGND
flabel metal1 178217 516962 178251 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_65.VPWR
flabel nwell 178217 516962 178251 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_65.VPB
flabel pwell 178217 517506 178251 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_65.VNB
rlabel comment 178188 517523 178188 517523 2 dpga_flat_0.sr_0.FILLER_0_24_65.decap_12
flabel metal1 179321 516962 179355 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_77.VPWR
flabel metal1 179321 517506 179355 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_77.VGND
flabel nwell 179321 516962 179355 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_77.VPB
flabel pwell 179321 517506 179355 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_77.VNB
rlabel comment 179292 517523 179292 517523 2 dpga_flat_0.sr_0.FILLER_0_24_77.decap_6
rlabel metal1 179292 517475 179844 517571 5 dpga_flat_0.sr_0.FILLER_0_24_77.VGND
rlabel metal1 179292 516931 179844 517027 5 dpga_flat_0.sr_0.FILLER_0_24_77.VPWR
flabel metal1 179866 516966 179902 516996 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_83.VPWR
flabel metal1 179866 517507 179902 517536 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_83.VGND
flabel nwell 179875 516972 179895 516989 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_83.VPB
flabel pwell 179872 517512 179896 517534 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_83.VNB
rlabel comment 179844 517523 179844 517523 2 dpga_flat_0.sr_0.FILLER_0_24_83.fill_1
rlabel metal1 179844 517475 179936 517571 5 dpga_flat_0.sr_0.FILLER_0_24_83.VGND
rlabel metal1 179844 516931 179936 517027 5 dpga_flat_0.sr_0.FILLER_0_24_83.VPWR
flabel metal1 180057 517506 180091 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_85.VGND
flabel metal1 180057 516962 180091 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_85.VPWR
flabel nwell 180057 516962 180091 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_85.VPB
flabel pwell 180057 517506 180091 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_85.VNB
rlabel comment 180028 517523 180028 517523 2 dpga_flat_0.sr_0.FILLER_0_24_85.decap_12
flabel metal1 181161 517506 181195 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_97.VGND
flabel metal1 181161 516962 181195 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_97.VPWR
flabel nwell 181161 516962 181195 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_97.VPB
flabel pwell 181161 517506 181195 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_97.VNB
rlabel comment 181132 517523 181132 517523 2 dpga_flat_0.sr_0.FILLER_0_24_97.decap_12
flabel metal1 179958 516970 180011 516999 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_24_119.VPWR
flabel metal1 179957 517503 180008 517541 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_24_119.VGND
rlabel comment 179936 517523 179936 517523 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_24_119.tapvpwrvgnd_1
rlabel metal1 179936 517475 180028 517571 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_24_119.VGND
rlabel metal1 179936 516931 180028 517027 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_24_119.VPWR
flabel metal1 182265 517506 182299 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_109.VGND
flabel metal1 182265 516962 182299 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_109.VPWR
flabel nwell 182265 516962 182299 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_109.VPB
flabel pwell 182265 517506 182299 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_109.VNB
rlabel comment 182236 517523 182236 517523 2 dpga_flat_0.sr_0.FILLER_0_24_109.decap_12
flabel metal1 183369 517506 183403 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_121.VGND
flabel metal1 183369 516962 183403 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_121.VPWR
flabel nwell 183369 516962 183403 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_121.VPB
flabel pwell 183369 517506 183403 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_121.VNB
rlabel comment 183340 517523 183340 517523 2 dpga_flat_0.sr_0.FILLER_0_24_121.decap_12
flabel metal1 184473 516962 184507 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_133.VPWR
flabel metal1 184473 517506 184507 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_133.VGND
flabel nwell 184473 516962 184507 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_133.VPB
flabel pwell 184473 517506 184507 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_133.VNB
rlabel comment 184444 517523 184444 517523 2 dpga_flat_0.sr_0.FILLER_0_24_133.decap_6
rlabel metal1 184444 517475 184996 517571 5 dpga_flat_0.sr_0.FILLER_0_24_133.VGND
rlabel metal1 184444 516931 184996 517027 5 dpga_flat_0.sr_0.FILLER_0_24_133.VPWR
flabel metal1 185018 516966 185054 516996 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_139.VPWR
flabel metal1 185018 517507 185054 517536 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_139.VGND
flabel nwell 185027 516972 185047 516989 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_139.VPB
flabel pwell 185024 517512 185048 517534 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_139.VNB
rlabel comment 184996 517523 184996 517523 2 dpga_flat_0.sr_0.FILLER_0_24_139.fill_1
rlabel metal1 184996 517475 185088 517571 5 dpga_flat_0.sr_0.FILLER_0_24_139.VGND
rlabel metal1 184996 516931 185088 517027 5 dpga_flat_0.sr_0.FILLER_0_24_139.VPWR
flabel metal1 185209 517506 185243 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_141.VGND
flabel metal1 185209 516962 185243 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_141.VPWR
flabel nwell 185209 516962 185243 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_141.VPB
flabel pwell 185209 517506 185243 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_141.VNB
rlabel comment 185180 517523 185180 517523 2 dpga_flat_0.sr_0.FILLER_0_24_141.decap_12
flabel metal1 185110 516970 185163 516999 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_24_120.VPWR
flabel metal1 185109 517503 185160 517541 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_24_120.VGND
rlabel comment 185088 517523 185088 517523 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_24_120.tapvpwrvgnd_1
rlabel metal1 185088 517475 185180 517571 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_24_120.VGND
rlabel metal1 185088 516931 185180 517027 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_24_120.VPWR
flabel metal1 186313 516962 186347 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_153.VPWR
flabel metal1 186313 517506 186347 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_153.VGND
flabel nwell 186313 516962 186347 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_153.VPB
flabel pwell 186313 517506 186347 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_153.VNB
rlabel comment 186284 517523 186284 517523 2 dpga_flat_0.sr_0.FILLER_0_24_153.decap_8
rlabel metal1 186284 517475 187020 517571 5 dpga_flat_0.sr_0.FILLER_0_24_153.VGND
rlabel metal1 186284 516931 187020 517027 5 dpga_flat_0.sr_0.FILLER_0_24_153.VPWR
flabel metal1 187040 517505 187093 517537 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_161.VGND
flabel metal1 187041 516962 187093 516993 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_161.VPWR
flabel nwell 187048 516970 187082 516988 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_161.VPB
flabel pwell 187051 517511 187083 517533 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_161.VNB
rlabel comment 187020 517523 187020 517523 2 dpga_flat_0.sr_0.FILLER_0_24_161.fill_2
rlabel metal1 187020 517475 187204 517571 5 dpga_flat_0.sr_0.FILLER_0_24_161.VGND
rlabel metal1 187020 516931 187204 517027 5 dpga_flat_0.sr_0.FILLER_0_24_161.VPWR
flabel metal1 187417 516962 187451 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_24_Right_24.VPWR
flabel metal1 187417 517506 187451 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_24_Right_24.VGND
flabel nwell 187417 516962 187451 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_24_Right_24.VPB
flabel pwell 187417 517506 187451 517540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_24_Right_24.VNB
rlabel comment 187480 517523 187480 517523 8 dpga_flat_0.sr_0.PHY_EDGE_ROW_24_Right_24.decap_3
rlabel metal1 187204 517475 187480 517571 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_24_Right_24.VGND
rlabel metal1 187204 516931 187480 517027 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_24_Right_24.VPWR
flabel metal1 172513 516418 172547 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_3.VGND
flabel metal1 172513 516962 172547 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_3.VPWR
flabel nwell 172513 516962 172547 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_3.VPB
flabel pwell 172513 516418 172547 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_3.VNB
rlabel comment 172484 516435 172484 516435 4 dpga_flat_0.sr_0.FILLER_0_25_3.decap_12
flabel metal1 173617 516418 173651 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_15.VGND
flabel metal1 173617 516962 173651 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_15.VPWR
flabel nwell 173617 516962 173651 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_15.VPB
flabel pwell 173617 516418 173651 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_15.VNB
rlabel comment 173588 516435 173588 516435 4 dpga_flat_0.sr_0.FILLER_0_25_15.decap_12
flabel metal1 172237 516962 172271 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_25_Left_53.VPWR
flabel metal1 172237 516418 172271 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_25_Left_53.VGND
flabel nwell 172237 516962 172271 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_25_Left_53.VPB
flabel pwell 172237 516418 172271 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_25_Left_53.VNB
rlabel comment 172208 516435 172208 516435 4 dpga_flat_0.sr_0.PHY_EDGE_ROW_25_Left_53.decap_3
rlabel metal1 172208 516387 172484 516483 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_25_Left_53.VGND
rlabel metal1 172208 516931 172484 517027 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_25_Left_53.VPWR
flabel metal1 174721 516418 174755 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_27.VGND
flabel metal1 174721 516962 174755 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_27.VPWR
flabel nwell 174721 516962 174755 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_27.VPB
flabel pwell 174721 516418 174755 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_27.VNB
rlabel comment 174692 516435 174692 516435 4 dpga_flat_0.sr_0.FILLER_0_25_27.decap_12
flabel metal1 175825 516418 175859 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_39.VGND
flabel metal1 175825 516962 175859 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_39.VPWR
flabel nwell 175825 516962 175859 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_39.VPB
flabel pwell 175825 516418 175859 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_39.VNB
rlabel comment 175796 516435 175796 516435 4 dpga_flat_0.sr_0.FILLER_0_25_39.decap_12
flabel metal1 176929 516418 176963 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_51.VGND
flabel metal1 176929 516962 176963 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_51.VPWR
flabel nwell 176929 516962 176963 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_51.VPB
flabel pwell 176929 516418 176963 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_51.VNB
rlabel comment 176900 516435 176900 516435 4 dpga_flat_0.sr_0.FILLER_0_25_51.decap_4
rlabel metal1 176900 516387 177268 516483 1 dpga_flat_0.sr_0.FILLER_0_25_51.VGND
rlabel metal1 176900 516931 177268 517027 1 dpga_flat_0.sr_0.FILLER_0_25_51.VPWR
flabel metal1 177290 516962 177326 516992 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_55.VPWR
flabel metal1 177290 516422 177326 516451 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_55.VGND
flabel nwell 177299 516969 177319 516986 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_55.VPB
flabel pwell 177296 516424 177320 516446 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_55.VNB
rlabel comment 177268 516435 177268 516435 4 dpga_flat_0.sr_0.FILLER_0_25_55.fill_1
rlabel metal1 177268 516387 177360 516483 1 dpga_flat_0.sr_0.FILLER_0_25_55.VGND
rlabel metal1 177268 516931 177360 517027 1 dpga_flat_0.sr_0.FILLER_0_25_55.VPWR
flabel metal1 177481 516418 177515 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_57.VGND
flabel metal1 177481 516962 177515 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_57.VPWR
flabel nwell 177481 516962 177515 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_57.VPB
flabel pwell 177481 516418 177515 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_57.VNB
rlabel comment 177452 516435 177452 516435 4 dpga_flat_0.sr_0.FILLER_0_25_57.decap_12
flabel metal1 177382 516959 177435 516988 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_25_121.VPWR
flabel metal1 177381 516417 177432 516455 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_25_121.VGND
rlabel comment 177360 516435 177360 516435 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_25_121.tapvpwrvgnd_1
rlabel metal1 177360 516387 177452 516483 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_25_121.VGND
rlabel metal1 177360 516931 177452 517027 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_25_121.VPWR
flabel metal1 178585 516418 178619 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_69.VGND
flabel metal1 178585 516962 178619 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_69.VPWR
flabel nwell 178585 516962 178619 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_69.VPB
flabel pwell 178585 516418 178619 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_69.VNB
rlabel comment 178556 516435 178556 516435 4 dpga_flat_0.sr_0.FILLER_0_25_69.decap_12
flabel metal1 179689 516418 179723 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_81.VGND
flabel metal1 179689 516962 179723 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_81.VPWR
flabel nwell 179689 516962 179723 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_81.VPB
flabel pwell 179689 516418 179723 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_81.VNB
rlabel comment 179660 516435 179660 516435 4 dpga_flat_0.sr_0.FILLER_0_25_81.decap_12
flabel metal1 180793 516418 180827 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_93.VGND
flabel metal1 180793 516962 180827 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_93.VPWR
flabel nwell 180793 516962 180827 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_93.VPB
flabel pwell 180793 516418 180827 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_93.VNB
rlabel comment 180764 516435 180764 516435 4 dpga_flat_0.sr_0.FILLER_0_25_93.decap_12
flabel metal1 181897 516962 181931 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_105.VPWR
flabel metal1 181897 516418 181931 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_105.VGND
flabel nwell 181897 516962 181931 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_105.VPB
flabel pwell 181897 516418 181931 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_105.VNB
rlabel comment 181868 516435 181868 516435 4 dpga_flat_0.sr_0.FILLER_0_25_105.decap_6
rlabel metal1 181868 516387 182420 516483 1 dpga_flat_0.sr_0.FILLER_0_25_105.VGND
rlabel metal1 181868 516931 182420 517027 1 dpga_flat_0.sr_0.FILLER_0_25_105.VPWR
flabel metal1 182442 516962 182478 516992 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_111.VPWR
flabel metal1 182442 516422 182478 516451 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_111.VGND
flabel nwell 182451 516969 182471 516986 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_111.VPB
flabel pwell 182448 516424 182472 516446 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_111.VNB
rlabel comment 182420 516435 182420 516435 4 dpga_flat_0.sr_0.FILLER_0_25_111.fill_1
rlabel metal1 182420 516387 182512 516483 1 dpga_flat_0.sr_0.FILLER_0_25_111.VGND
rlabel metal1 182420 516931 182512 517027 1 dpga_flat_0.sr_0.FILLER_0_25_111.VPWR
flabel metal1 182633 516418 182667 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_113.VGND
flabel metal1 182633 516962 182667 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_113.VPWR
flabel nwell 182633 516962 182667 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_113.VPB
flabel pwell 182633 516418 182667 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_113.VNB
rlabel comment 182604 516435 182604 516435 4 dpga_flat_0.sr_0.FILLER_0_25_113.decap_12
flabel metal1 183737 516418 183771 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_125.VGND
flabel metal1 183737 516962 183771 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_125.VPWR
flabel nwell 183737 516962 183771 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_125.VPB
flabel pwell 183737 516418 183771 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_125.VNB
rlabel comment 183708 516435 183708 516435 4 dpga_flat_0.sr_0.FILLER_0_25_125.decap_12
flabel metal1 182534 516959 182587 516988 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_25_122.VPWR
flabel metal1 182533 516417 182584 516455 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_25_122.VGND
rlabel comment 182512 516435 182512 516435 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_25_122.tapvpwrvgnd_1
rlabel metal1 182512 516387 182604 516483 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_25_122.VGND
rlabel metal1 182512 516931 182604 517027 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_25_122.VPWR
flabel metal1 184841 516418 184875 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_137.VGND
flabel metal1 184841 516962 184875 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_137.VPWR
flabel nwell 184841 516962 184875 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_137.VPB
flabel pwell 184841 516418 184875 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_137.VNB
rlabel comment 184812 516435 184812 516435 4 dpga_flat_0.sr_0.FILLER_0_25_137.decap_12
flabel metal1 185945 516418 185979 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_149.VGND
flabel metal1 185945 516962 185979 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_149.VPWR
flabel nwell 185945 516962 185979 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_149.VPB
flabel pwell 185945 516418 185979 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_149.VNB
rlabel comment 185916 516435 185916 516435 4 dpga_flat_0.sr_0.FILLER_0_25_149.decap_12
flabel metal1 187040 516421 187093 516453 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_161.VGND
flabel metal1 187041 516965 187093 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_161.VPWR
flabel nwell 187048 516970 187082 516988 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_161.VPB
flabel pwell 187051 516425 187083 516447 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_161.VNB
rlabel comment 187020 516435 187020 516435 4 dpga_flat_0.sr_0.FILLER_0_25_161.fill_2
rlabel metal1 187020 516387 187204 516483 1 dpga_flat_0.sr_0.FILLER_0_25_161.VGND
rlabel metal1 187020 516931 187204 517027 1 dpga_flat_0.sr_0.FILLER_0_25_161.VPWR
flabel metal1 187417 516962 187451 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_25_Right_25.VPWR
flabel metal1 187417 516418 187451 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_25_Right_25.VGND
flabel nwell 187417 516962 187451 516996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_25_Right_25.VPB
flabel pwell 187417 516418 187451 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_25_Right_25.VNB
rlabel comment 187480 516435 187480 516435 6 dpga_flat_0.sr_0.PHY_EDGE_ROW_25_Right_25.decap_3
rlabel metal1 187204 516387 187480 516483 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_25_Right_25.VGND
rlabel metal1 187204 516931 187480 517027 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_25_Right_25.VPWR
flabel metal1 172513 516418 172547 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_3.VGND
flabel metal1 172513 515874 172547 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_3.VPWR
flabel nwell 172513 515874 172547 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_3.VPB
flabel pwell 172513 516418 172547 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_3.VNB
rlabel comment 172484 516435 172484 516435 2 dpga_flat_0.sr_0.FILLER_0_26_3.decap_12
flabel metal1 173617 516418 173651 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_15.VGND
flabel metal1 173617 515874 173651 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_15.VPWR
flabel nwell 173617 515874 173651 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_15.VPB
flabel pwell 173617 516418 173651 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_15.VNB
rlabel comment 173588 516435 173588 516435 2 dpga_flat_0.sr_0.FILLER_0_26_15.decap_12
flabel metal1 172513 515874 172547 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_3.VPWR
flabel metal1 172513 515330 172547 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_3.VGND
flabel nwell 172513 515874 172547 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_3.VPB
flabel pwell 172513 515330 172547 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_3.VNB
rlabel comment 172484 515347 172484 515347 4 dpga_flat_0.sr_0.FILLER_0_27_3.decap_8
rlabel metal1 172484 515299 173220 515395 1 dpga_flat_0.sr_0.FILLER_0_27_3.VGND
rlabel metal1 172484 515843 173220 515939 1 dpga_flat_0.sr_0.FILLER_0_27_3.VPWR
flabel metal1 173240 515333 173293 515365 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_11.VGND
flabel metal1 173241 515877 173293 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_11.VPWR
flabel nwell 173248 515882 173282 515900 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_11.VPB
flabel pwell 173251 515337 173283 515359 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_11.VNB
rlabel comment 173220 515347 173220 515347 4 dpga_flat_0.sr_0.FILLER_0_27_11.fill_2
rlabel metal1 173220 515299 173404 515395 1 dpga_flat_0.sr_0.FILLER_0_27_11.VGND
rlabel metal1 173220 515843 173404 515939 1 dpga_flat_0.sr_0.FILLER_0_27_11.VPWR
flabel metal1 173985 515874 174019 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_19.VPWR
flabel metal1 173985 515330 174019 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_19.VGND
flabel nwell 173985 515874 174019 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_19.VPB
flabel pwell 173985 515330 174019 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_19.VNB
rlabel comment 173956 515347 173956 515347 4 dpga_flat_0.sr_0.FILLER_0_27_19.decap_8
rlabel metal1 173956 515299 174692 515395 1 dpga_flat_0.sr_0.FILLER_0_27_19.VGND
rlabel metal1 173956 515843 174692 515939 1 dpga_flat_0.sr_0.FILLER_0_27_19.VPWR
flabel metal1 172237 515874 172271 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_26_Left_54.VPWR
flabel metal1 172237 516418 172271 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_26_Left_54.VGND
flabel nwell 172237 515874 172271 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_26_Left_54.VPB
flabel pwell 172237 516418 172271 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_26_Left_54.VNB
rlabel comment 172208 516435 172208 516435 2 dpga_flat_0.sr_0.PHY_EDGE_ROW_26_Left_54.decap_3
rlabel metal1 172208 516387 172484 516483 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_26_Left_54.VGND
rlabel metal1 172208 515843 172484 515939 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_26_Left_54.VPWR
flabel metal1 172237 515874 172271 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_27_Left_55.VPWR
flabel metal1 172237 515330 172271 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_27_Left_55.VGND
flabel nwell 172237 515874 172271 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_27_Left_55.VPB
flabel pwell 172237 515330 172271 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_27_Left_55.VNB
rlabel comment 172208 515347 172208 515347 4 dpga_flat_0.sr_0.PHY_EDGE_ROW_27_Left_55.decap_3
rlabel metal1 172208 515299 172484 515395 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_27_Left_55.VGND
rlabel metal1 172208 515843 172484 515939 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_27_Left_55.VPWR
flabel locali 173801 515636 173835 515670 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input3.X
flabel locali 173525 515500 173559 515534 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input3.A
flabel locali 173893 515500 173927 515534 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input3.X
flabel locali 173525 515568 173559 515602 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input3.A
flabel locali 173893 515568 173927 515602 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input3.X
flabel metal1 173433 515330 173467 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input3.VGND
flabel metal1 173433 515874 173467 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input3.VPWR
flabel nwell 173433 515874 173467 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input3.VPB
flabel pwell 173433 515330 173467 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input3.VNB
rlabel comment 173404 515347 173404 515347 4 dpga_flat_0.sr_0.input3.clkbuf_4
rlabel metal1 173404 515299 173956 515395 1 dpga_flat_0.sr_0.input3.VGND
rlabel metal1 173404 515843 173956 515939 1 dpga_flat_0.sr_0.input3.VPWR
flabel metal1 174714 515878 174750 515908 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_27.VPWR
flabel metal1 174714 516419 174750 516448 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_27.VGND
flabel nwell 174723 515884 174743 515901 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_27.VPB
flabel pwell 174720 516424 174744 516446 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_27.VNB
rlabel comment 174692 516435 174692 516435 2 dpga_flat_0.sr_0.FILLER_0_26_27.fill_1
rlabel metal1 174692 516387 174784 516483 5 dpga_flat_0.sr_0.FILLER_0_26_27.VGND
rlabel metal1 174692 515843 174784 515939 5 dpga_flat_0.sr_0.FILLER_0_26_27.VPWR
flabel metal1 174905 516418 174939 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_29.VGND
flabel metal1 174905 515874 174939 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_29.VPWR
flabel nwell 174905 515874 174939 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_29.VPB
flabel pwell 174905 516418 174939 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_29.VNB
rlabel comment 174876 516435 174876 516435 2 dpga_flat_0.sr_0.FILLER_0_26_29.decap_12
flabel metal1 176009 516418 176043 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_41.VGND
flabel metal1 176009 515874 176043 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_41.VPWR
flabel nwell 176009 515874 176043 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_41.VPB
flabel pwell 176009 516418 176043 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_41.VNB
rlabel comment 175980 516435 175980 516435 2 dpga_flat_0.sr_0.FILLER_0_26_41.decap_12
flabel metal1 174714 515874 174750 515904 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_27.VPWR
flabel metal1 174714 515334 174750 515363 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_27.VGND
flabel nwell 174723 515881 174743 515898 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_27.VPB
flabel pwell 174720 515336 174744 515358 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_27.VNB
rlabel comment 174692 515347 174692 515347 4 dpga_flat_0.sr_0.FILLER_0_27_27.fill_1
rlabel metal1 174692 515299 174784 515395 1 dpga_flat_0.sr_0.FILLER_0_27_27.VGND
rlabel metal1 174692 515843 174784 515939 1 dpga_flat_0.sr_0.FILLER_0_27_27.VPWR
flabel metal1 174905 515330 174939 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_29.VGND
flabel metal1 174905 515874 174939 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_29.VPWR
flabel nwell 174905 515874 174939 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_29.VPB
flabel pwell 174905 515330 174939 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_29.VNB
rlabel comment 174876 515347 174876 515347 4 dpga_flat_0.sr_0.FILLER_0_27_29.decap_12
flabel metal1 176009 515330 176043 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_41.VGND
flabel metal1 176009 515874 176043 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_41.VPWR
flabel nwell 176009 515874 176043 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_41.VPB
flabel pwell 176009 515330 176043 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_41.VNB
rlabel comment 175980 515347 175980 515347 4 dpga_flat_0.sr_0.FILLER_0_27_41.decap_12
flabel metal1 174806 515882 174859 515911 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_26_123.VPWR
flabel metal1 174805 516415 174856 516453 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_26_123.VGND
rlabel comment 174784 516435 174784 516435 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_26_123.tapvpwrvgnd_1
rlabel metal1 174784 516387 174876 516483 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_26_123.VGND
rlabel metal1 174784 515843 174876 515939 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_26_123.VPWR
flabel metal1 174806 515871 174859 515900 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_126.VPWR
flabel metal1 174805 515329 174856 515367 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_126.VGND
rlabel comment 174784 515347 174784 515347 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_126.tapvpwrvgnd_1
rlabel metal1 174784 515299 174876 515395 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_126.VGND
rlabel metal1 174784 515843 174876 515939 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_126.VPWR
flabel metal1 177113 516418 177147 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_53.VGND
flabel metal1 177113 515874 177147 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_53.VPWR
flabel nwell 177113 515874 177147 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_53.VPB
flabel pwell 177113 516418 177147 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_53.VNB
rlabel comment 177084 516435 177084 516435 2 dpga_flat_0.sr_0.FILLER_0_26_53.decap_12
flabel metal1 177113 515874 177147 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_53.VPWR
flabel metal1 177113 515330 177147 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_53.VGND
flabel nwell 177113 515874 177147 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_53.VPB
flabel pwell 177113 515330 177147 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_53.VNB
rlabel comment 177084 515347 177084 515347 4 dpga_flat_0.sr_0.FILLER_0_27_53.decap_3
rlabel metal1 177084 515299 177360 515395 1 dpga_flat_0.sr_0.FILLER_0_27_53.VGND
rlabel metal1 177084 515843 177360 515939 1 dpga_flat_0.sr_0.FILLER_0_27_53.VPWR
flabel metal1 177481 515330 177515 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_57.VGND
flabel metal1 177481 515874 177515 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_57.VPWR
flabel nwell 177481 515874 177515 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_57.VPB
flabel pwell 177481 515330 177515 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_57.VNB
rlabel comment 177452 515347 177452 515347 4 dpga_flat_0.sr_0.FILLER_0_27_57.decap_12
flabel metal1 177382 515871 177435 515900 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_127.VPWR
flabel metal1 177381 515329 177432 515367 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_127.VGND
rlabel comment 177360 515347 177360 515347 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_127.tapvpwrvgnd_1
rlabel metal1 177360 515299 177452 515395 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_127.VGND
rlabel metal1 177360 515843 177452 515939 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_127.VPWR
flabel metal1 178217 516418 178251 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_65.VGND
flabel metal1 178217 515874 178251 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_65.VPWR
flabel nwell 178217 515874 178251 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_65.VPB
flabel pwell 178217 516418 178251 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_65.VNB
rlabel comment 178188 516435 178188 516435 2 dpga_flat_0.sr_0.FILLER_0_26_65.decap_12
flabel metal1 179321 515874 179355 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_77.VPWR
flabel metal1 179321 516418 179355 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_77.VGND
flabel nwell 179321 515874 179355 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_77.VPB
flabel pwell 179321 516418 179355 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_77.VNB
rlabel comment 179292 516435 179292 516435 2 dpga_flat_0.sr_0.FILLER_0_26_77.decap_6
rlabel metal1 179292 516387 179844 516483 5 dpga_flat_0.sr_0.FILLER_0_26_77.VGND
rlabel metal1 179292 515843 179844 515939 5 dpga_flat_0.sr_0.FILLER_0_26_77.VPWR
flabel metal1 179866 515878 179902 515908 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_83.VPWR
flabel metal1 179866 516419 179902 516448 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_83.VGND
flabel nwell 179875 515884 179895 515901 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_83.VPB
flabel pwell 179872 516424 179896 516446 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_83.VNB
rlabel comment 179844 516435 179844 516435 2 dpga_flat_0.sr_0.FILLER_0_26_83.fill_1
rlabel metal1 179844 516387 179936 516483 5 dpga_flat_0.sr_0.FILLER_0_26_83.VGND
rlabel metal1 179844 515843 179936 515939 5 dpga_flat_0.sr_0.FILLER_0_26_83.VPWR
flabel metal1 178585 515330 178619 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_69.VGND
flabel metal1 178585 515874 178619 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_69.VPWR
flabel nwell 178585 515874 178619 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_69.VPB
flabel pwell 178585 515330 178619 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_69.VNB
rlabel comment 178556 515347 178556 515347 4 dpga_flat_0.sr_0.FILLER_0_27_69.decap_12
flabel metal1 179689 515874 179723 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_81.VPWR
flabel metal1 179689 515330 179723 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_81.VGND
flabel nwell 179689 515874 179723 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_81.VPB
flabel pwell 179689 515330 179723 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_81.VNB
rlabel comment 179660 515347 179660 515347 4 dpga_flat_0.sr_0.FILLER_0_27_81.decap_3
rlabel metal1 179660 515299 179936 515395 1 dpga_flat_0.sr_0.FILLER_0_27_81.VGND
rlabel metal1 179660 515843 179936 515939 1 dpga_flat_0.sr_0.FILLER_0_27_81.VPWR
flabel metal1 180057 516418 180091 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_85.VGND
flabel metal1 180057 515874 180091 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_85.VPWR
flabel nwell 180057 515874 180091 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_85.VPB
flabel pwell 180057 516418 180091 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_85.VNB
rlabel comment 180028 516435 180028 516435 2 dpga_flat_0.sr_0.FILLER_0_26_85.decap_12
flabel metal1 181161 516418 181195 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_97.VGND
flabel metal1 181161 515874 181195 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_97.VPWR
flabel nwell 181161 515874 181195 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_97.VPB
flabel pwell 181161 516418 181195 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_97.VNB
rlabel comment 181132 516435 181132 516435 2 dpga_flat_0.sr_0.FILLER_0_26_97.decap_12
flabel metal1 180057 515330 180091 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_85.VGND
flabel metal1 180057 515874 180091 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_85.VPWR
flabel nwell 180057 515874 180091 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_85.VPB
flabel pwell 180057 515330 180091 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_85.VNB
rlabel comment 180028 515347 180028 515347 4 dpga_flat_0.sr_0.FILLER_0_27_85.decap_12
flabel metal1 181161 515874 181195 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_97.VPWR
flabel metal1 181161 515330 181195 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_97.VGND
flabel nwell 181161 515874 181195 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_97.VPB
flabel pwell 181161 515330 181195 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_97.VNB
rlabel comment 181132 515347 181132 515347 4 dpga_flat_0.sr_0.FILLER_0_27_97.decap_8
rlabel metal1 181132 515299 181868 515395 1 dpga_flat_0.sr_0.FILLER_0_27_97.VGND
rlabel metal1 181132 515843 181868 515939 1 dpga_flat_0.sr_0.FILLER_0_27_97.VPWR
flabel metal1 179958 515882 180011 515911 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_26_124.VPWR
flabel metal1 179957 516415 180008 516453 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_26_124.VGND
rlabel comment 179936 516435 179936 516435 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_26_124.tapvpwrvgnd_1
rlabel metal1 179936 516387 180028 516483 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_26_124.VGND
rlabel metal1 179936 515843 180028 515939 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_26_124.VPWR
flabel metal1 179958 515871 180011 515900 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_128.VPWR
flabel metal1 179957 515329 180008 515367 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_128.VGND
rlabel comment 179936 515347 179936 515347 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_128.tapvpwrvgnd_1
rlabel metal1 179936 515299 180028 515395 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_128.VGND
rlabel metal1 179936 515843 180028 515939 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_128.VPWR
flabel metal1 182265 516418 182299 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_109.VGND
flabel metal1 182265 515874 182299 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_109.VPWR
flabel nwell 182265 515874 182299 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_109.VPB
flabel pwell 182265 516418 182299 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_109.VNB
rlabel comment 182236 516435 182236 516435 2 dpga_flat_0.sr_0.FILLER_0_26_109.decap_12
flabel metal1 183369 516418 183403 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_121.VGND
flabel metal1 183369 515874 183403 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_121.VPWR
flabel nwell 183369 515874 183403 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_121.VPB
flabel pwell 183369 516418 183403 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_121.VNB
rlabel comment 183340 516435 183340 516435 2 dpga_flat_0.sr_0.FILLER_0_26_121.decap_12
flabel metal1 181888 515333 181941 515365 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_105.VGND
flabel metal1 181889 515877 181941 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_105.VPWR
flabel nwell 181896 515882 181930 515900 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_105.VPB
flabel pwell 181899 515337 181931 515359 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_105.VNB
rlabel comment 181868 515347 181868 515347 4 dpga_flat_0.sr_0.FILLER_0_27_105.fill_2
rlabel metal1 181868 515299 182052 515395 1 dpga_flat_0.sr_0.FILLER_0_27_105.VGND
rlabel metal1 181868 515843 182052 515939 1 dpga_flat_0.sr_0.FILLER_0_27_105.VPWR
flabel metal1 182348 515333 182401 515365 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_110.VGND
flabel metal1 182349 515877 182401 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_110.VPWR
flabel nwell 182356 515882 182390 515900 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_110.VPB
flabel pwell 182359 515337 182391 515359 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_110.VNB
rlabel comment 182328 515347 182328 515347 4 dpga_flat_0.sr_0.FILLER_0_27_110.fill_2
rlabel metal1 182328 515299 182512 515395 1 dpga_flat_0.sr_0.FILLER_0_27_110.VGND
rlabel metal1 182328 515843 182512 515939 1 dpga_flat_0.sr_0.FILLER_0_27_110.VPWR
flabel metal1 182633 515330 182667 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_113.VGND
flabel metal1 182633 515874 182667 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_113.VPWR
flabel nwell 182633 515874 182667 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_113.VPB
flabel pwell 182633 515330 182667 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_113.VNB
rlabel comment 182604 515347 182604 515347 4 dpga_flat_0.sr_0.FILLER_0_27_113.decap_12
flabel metal1 183737 515330 183771 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_125.VGND
flabel metal1 183737 515874 183771 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_125.VPWR
flabel nwell 183737 515874 183771 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_125.VPB
flabel pwell 183737 515330 183771 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_125.VNB
rlabel comment 183708 515347 183708 515347 4 dpga_flat_0.sr_0.FILLER_0_27_125.decap_12
flabel metal1 182534 515871 182587 515900 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_129.VPWR
flabel metal1 182533 515329 182584 515367 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_129.VGND
rlabel comment 182512 515347 182512 515347 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_129.tapvpwrvgnd_1
rlabel metal1 182512 515299 182604 515395 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_129.VGND
rlabel metal1 182512 515843 182604 515939 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_129.VPWR
flabel metal1 182263 515330 182297 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input2.VGND
flabel metal1 182265 515874 182299 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input2.VPWR
flabel locali 182265 515874 182299 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input2.VPWR
flabel locali 182263 515330 182297 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input2.VGND
flabel locali 182083 515432 182117 515466 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input2.X
flabel locali 182083 515704 182117 515738 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input2.X
flabel locali 182083 515772 182117 515806 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input2.X
flabel locali 182265 515568 182299 515602 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input2.A
flabel nwell 182265 515874 182299 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input2.VPB
flabel pwell 182263 515330 182297 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input2.VNB
rlabel comment 182328 515347 182328 515347 6 dpga_flat_0.sr_0.input2.buf_1
rlabel metal1 182052 515299 182328 515395 1 dpga_flat_0.sr_0.input2.VGND
rlabel metal1 182052 515843 182328 515939 1 dpga_flat_0.sr_0.input2.VPWR
flabel metal1 184473 515874 184507 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_133.VPWR
flabel metal1 184473 516418 184507 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_133.VGND
flabel nwell 184473 515874 184507 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_133.VPB
flabel pwell 184473 516418 184507 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_133.VNB
rlabel comment 184444 516435 184444 516435 2 dpga_flat_0.sr_0.FILLER_0_26_133.decap_6
rlabel metal1 184444 516387 184996 516483 5 dpga_flat_0.sr_0.FILLER_0_26_133.VGND
rlabel metal1 184444 515843 184996 515939 5 dpga_flat_0.sr_0.FILLER_0_26_133.VPWR
flabel metal1 185018 515878 185054 515908 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_139.VPWR
flabel metal1 185018 516419 185054 516448 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_139.VGND
flabel nwell 185027 515884 185047 515901 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_139.VPB
flabel pwell 185024 516424 185048 516446 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_139.VNB
rlabel comment 184996 516435 184996 516435 2 dpga_flat_0.sr_0.FILLER_0_26_139.fill_1
rlabel metal1 184996 516387 185088 516483 5 dpga_flat_0.sr_0.FILLER_0_26_139.VGND
rlabel metal1 184996 515843 185088 515939 5 dpga_flat_0.sr_0.FILLER_0_26_139.VPWR
flabel metal1 185209 516418 185243 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_141.VGND
flabel metal1 185209 515874 185243 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_141.VPWR
flabel nwell 185209 515874 185243 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_141.VPB
flabel pwell 185209 516418 185243 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_141.VNB
rlabel comment 185180 516435 185180 516435 2 dpga_flat_0.sr_0.FILLER_0_26_141.decap_12
flabel metal1 184841 515874 184875 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_137.VPWR
flabel metal1 184841 515330 184875 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_137.VGND
flabel nwell 184841 515874 184875 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_137.VPB
flabel pwell 184841 515330 184875 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_137.VNB
rlabel comment 184812 515347 184812 515347 4 dpga_flat_0.sr_0.FILLER_0_27_137.decap_3
rlabel metal1 184812 515299 185088 515395 1 dpga_flat_0.sr_0.FILLER_0_27_137.VGND
rlabel metal1 184812 515843 185088 515939 1 dpga_flat_0.sr_0.FILLER_0_27_137.VPWR
flabel metal1 185209 515330 185243 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_141.VGND
flabel metal1 185209 515874 185243 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_141.VPWR
flabel nwell 185209 515874 185243 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_141.VPB
flabel pwell 185209 515330 185243 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_141.VNB
rlabel comment 185180 515347 185180 515347 4 dpga_flat_0.sr_0.FILLER_0_27_141.decap_12
flabel metal1 185110 515882 185163 515911 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_26_125.VPWR
flabel metal1 185109 516415 185160 516453 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_26_125.VGND
rlabel comment 185088 516435 185088 516435 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_26_125.tapvpwrvgnd_1
rlabel metal1 185088 516387 185180 516483 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_26_125.VGND
rlabel metal1 185088 515843 185180 515939 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_26_125.VPWR
flabel metal1 185110 515871 185163 515900 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_130.VPWR
flabel metal1 185109 515329 185160 515367 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_130.VGND
rlabel comment 185088 515347 185088 515347 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_130.tapvpwrvgnd_1
rlabel metal1 185088 515299 185180 515395 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_130.VGND
rlabel metal1 185088 515843 185180 515939 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_130.VPWR
flabel metal1 186313 515874 186347 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_153.VPWR
flabel metal1 186313 516418 186347 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_153.VGND
flabel nwell 186313 515874 186347 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_153.VPB
flabel pwell 186313 516418 186347 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_153.VNB
rlabel comment 186284 516435 186284 516435 2 dpga_flat_0.sr_0.FILLER_0_26_153.decap_8
rlabel metal1 186284 516387 187020 516483 5 dpga_flat_0.sr_0.FILLER_0_26_153.VGND
rlabel metal1 186284 515843 187020 515939 5 dpga_flat_0.sr_0.FILLER_0_26_153.VPWR
flabel metal1 187040 516417 187093 516449 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_161.VGND
flabel metal1 187041 515874 187093 515905 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_161.VPWR
flabel nwell 187048 515882 187082 515900 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_161.VPB
flabel pwell 187051 516423 187083 516445 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_161.VNB
rlabel comment 187020 516435 187020 516435 2 dpga_flat_0.sr_0.FILLER_0_26_161.fill_2
rlabel metal1 187020 516387 187204 516483 5 dpga_flat_0.sr_0.FILLER_0_26_161.VGND
rlabel metal1 187020 515843 187204 515939 5 dpga_flat_0.sr_0.FILLER_0_26_161.VPWR
flabel metal1 186306 515874 186342 515904 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_153.VPWR
flabel metal1 186306 515334 186342 515363 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_153.VGND
flabel nwell 186315 515881 186335 515898 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_153.VPB
flabel pwell 186312 515336 186336 515358 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_153.VNB
rlabel comment 186284 515347 186284 515347 4 dpga_flat_0.sr_0.FILLER_0_27_153.fill_1
rlabel metal1 186284 515299 186376 515395 1 dpga_flat_0.sr_0.FILLER_0_27_153.VGND
rlabel metal1 186284 515843 186376 515939 1 dpga_flat_0.sr_0.FILLER_0_27_153.VPWR
flabel metal1 186957 515874 186991 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_160.VPWR
flabel metal1 186957 515330 186991 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_160.VGND
flabel nwell 186957 515874 186991 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_160.VPB
flabel pwell 186957 515330 186991 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_160.VNB
rlabel comment 186928 515347 186928 515347 4 dpga_flat_0.sr_0.FILLER_0_27_160.decap_3
rlabel metal1 186928 515299 187204 515395 1 dpga_flat_0.sr_0.FILLER_0_27_160.VGND
rlabel metal1 186928 515843 187204 515939 1 dpga_flat_0.sr_0.FILLER_0_27_160.VPWR
flabel metal1 187417 515874 187451 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_26_Right_26.VPWR
flabel metal1 187417 516418 187451 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_26_Right_26.VGND
flabel nwell 187417 515874 187451 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_26_Right_26.VPB
flabel pwell 187417 516418 187451 516452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_26_Right_26.VNB
rlabel comment 187480 516435 187480 516435 8 dpga_flat_0.sr_0.PHY_EDGE_ROW_26_Right_26.decap_3
rlabel metal1 187204 516387 187480 516483 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_26_Right_26.VGND
rlabel metal1 187204 515843 187480 515939 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_26_Right_26.VPWR
flabel metal1 187417 515874 187451 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_27_Right_27.VPWR
flabel metal1 187417 515330 187451 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_27_Right_27.VGND
flabel nwell 187417 515874 187451 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_27_Right_27.VPB
flabel pwell 187417 515330 187451 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_27_Right_27.VNB
rlabel comment 187480 515347 187480 515347 6 dpga_flat_0.sr_0.PHY_EDGE_ROW_27_Right_27.decap_3
rlabel metal1 187204 515299 187480 515395 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_27_Right_27.VGND
rlabel metal1 187204 515843 187480 515939 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_27_Right_27.VPWR
flabel locali 186773 515636 186807 515670 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input1.X
flabel locali 186497 515500 186531 515534 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input1.A
flabel locali 186865 515500 186899 515534 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input1.X
flabel locali 186497 515568 186531 515602 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input1.A
flabel locali 186865 515568 186899 515602 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input1.X
flabel metal1 186405 515330 186439 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input1.VGND
flabel metal1 186405 515874 186439 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input1.VPWR
flabel nwell 186405 515874 186439 515908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input1.VPB
flabel pwell 186405 515330 186439 515364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input1.VNB
rlabel comment 186376 515347 186376 515347 4 dpga_flat_0.sr_0.input1.clkbuf_4
rlabel metal1 186376 515299 186928 515395 1 dpga_flat_0.sr_0.input1.VGND
rlabel metal1 186376 515843 186928 515939 1 dpga_flat_0.sr_0.input1.VPWR
flabel metal1 156998 536765 157198 536955 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.out
flabel metal1 192228 540065 192428 540255 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.gnd
flabel metal1 192228 539115 192428 539315 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.vd
flabel metal1 163528 542565 163728 542755 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.inp
flabel metal1 178178 542525 178378 542715 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.inn
flabel metal1 163028 533315 163228 533505 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.ib
flabel metal1 167518 533305 167718 533505 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.c0
flabel metal1 171048 533305 171248 533505 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.c1
flabel metal1 174678 533305 174878 533505 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.c2
flabel metal1 178218 533305 178418 533505 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.c3
flabel metal1 181728 533305 181928 533505 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.c4
flabel metal1 184968 533305 185168 533505 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.c5
flabel metal1 188198 533305 188398 533505 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.c6
flabel metal1 191478 533305 191678 533505 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.c7
flabel metal1 163028 538675 163228 538875 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.ota_0.vs
flabel metal1 163018 536995 163218 537195 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.ota_0.inn
flabel metal1 163018 537835 163218 538035 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.ota_0.inp
flabel metal1 163028 536565 163228 536765 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.ota_0.ib
flabel metal1 160178 535385 160378 535585 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.ota_0.vd
flabel metal1 157198 536755 157398 536955 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.ota_0.out
flabel metal1 161448 538045 161488 538065 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.ota_0.d
flabel metal1 162188 538045 162188 538065 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.ota_0.c
flabel metal2 161648 536825 161668 536845 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.ota_0.b
flabel metal1 167518 535215 167718 535415 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.c0
flabel metal1 171048 535215 171248 535415 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.c1
flabel metal1 174678 535215 174878 535415 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.c2
flabel metal1 178218 535215 178418 535415 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.c3
flabel metal1 181728 535215 181928 535415 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.c4
flabel metal1 184968 535215 185168 535415 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.c5
flabel metal1 188198 535215 188398 535415 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.c6
flabel metal1 191478 535215 191678 535415 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.c7
flabel metal1 178178 542065 178378 542265 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.n0
flabel metal1 163528 536005 163728 536205 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.n8
flabel metal1 192028 540055 192228 540255 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.gnd
flabel metal1 192028 539115 192228 539315 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.vd
flabel metal1 170478 539115 170678 539315 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_7.vd
flabel metal1 168078 539555 168278 539755 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_7.b
flabel metal1 170478 540055 170678 540255 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_7.vgnd
flabel metal1 170478 540695 170678 540895 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_7.ctrl
flabel metal1 168078 540835 168278 541035 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_7.a
flabel metal1 169938 538485 169958 538495 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_7.nctrl
flabel metal1 174178 539115 174378 539315 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_6.vd
flabel metal1 171778 539555 171978 539755 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_6.b
flabel metal1 174178 540055 174378 540255 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_6.vgnd
flabel metal1 174178 540695 174378 540895 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_6.ctrl
flabel metal1 171778 540835 171978 541035 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_6.a
flabel metal1 173638 538485 173658 538495 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_6.nctrl
flabel metal1 177678 539115 177878 539315 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_5.vd
flabel metal1 175278 539555 175478 539755 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_5.b
flabel metal1 177678 540055 177878 540255 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_5.vgnd
flabel metal1 177678 540695 177878 540895 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_5.ctrl
flabel metal1 175278 540835 175478 541035 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_5.a
flabel metal1 177138 538485 177158 538495 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_5.nctrl
flabel metal1 166678 539115 166878 539315 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_4.vd
flabel metal1 164278 539555 164478 539755 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_4.b
flabel metal1 166678 540055 166878 540255 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_4.vgnd
flabel metal1 166678 540695 166878 540895 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_4.ctrl
flabel metal1 164278 540835 164478 541035 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_4.a
flabel metal1 166138 538485 166158 538495 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_4.nctrl
flabel metal1 181278 539115 181478 539315 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_3.vd
flabel metal1 178878 539555 179078 539755 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_3.b
flabel metal1 181278 540055 181478 540255 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_3.vgnd
flabel metal1 181278 540695 181478 540895 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_3.ctrl
flabel metal1 178878 540835 179078 541035 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_3.a
flabel metal1 180738 538485 180758 538495 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_3.nctrl
flabel metal1 184578 539115 184778 539315 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_2.vd
flabel metal1 182178 539555 182378 539755 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_2.b
flabel metal1 184578 540055 184778 540255 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_2.vgnd
flabel metal1 184578 540695 184778 540895 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_2.ctrl
flabel metal1 182178 540835 182378 541035 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_2.a
flabel metal1 184038 538485 184058 538495 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_2.nctrl
flabel metal1 191178 539115 191378 539315 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_1.vd
flabel metal1 188778 539555 188978 539755 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_1.b
flabel metal1 191178 540055 191378 540255 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_1.vgnd
flabel metal1 191178 540695 191378 540895 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_1.ctrl
flabel metal1 188778 540835 188978 541035 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_1.a
flabel metal1 190638 538485 190658 538495 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_1.nctrl
flabel metal1 187878 539115 188078 539315 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_0.vd
flabel metal1 185478 539555 185678 539755 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_0.b
flabel metal1 187878 540055 188078 540255 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_0.vgnd
flabel metal1 187878 540695 188078 540895 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_0.ctrl
flabel metal1 185478 540835 185678 541035 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_0.a
flabel metal1 187338 538485 187358 538495 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_0.nctrl
flabel metal1 193000 540000 195000 542000 0 FreeSans 1600 0 0 0 gnd_ota
port 70 nsew
flabel metal1 193000 537320 195000 539320 0 FreeSans 1600 0 0 0 vd_ota
port 68 nsew
<< end >>

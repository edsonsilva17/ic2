magic
tech sky130A
magscale 1 2
timestamp 1699055702
use cafeina_top_level  cafeina_top_level_0
timestamp 1699054617
transform 1 0 0 0 1 9
box 217294 450753 583581 703284
use gme_cefet_top_level  gme_cefet_top_level_0
timestamp 1699054617
transform 1 0 78 0 1 -9
box 326 15091 583606 406686
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>

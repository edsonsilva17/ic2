magic
tech sky130A
magscale 1 2
timestamp 1699054617
<< nwell >>
rect 106133 277914 107804 279258
rect 106272 276894 107744 277360
rect 106670 274677 109883 275970
rect 109052 270485 109897 272638
rect 114419 272669 115786 280999
rect 112237 270724 115567 271722
rect 120201 279136 121769 280849
rect 122142 280643 123674 280644
rect 120201 273034 121764 279136
rect 122133 278930 123674 280643
rect 122218 277151 124406 278518
rect 122242 276273 124028 276887
rect 122247 275515 124993 276007
rect 120201 268958 123590 273034
rect 120201 268942 121884 268958
<< pwell >>
rect 105948 281071 106173 281091
rect 111020 281073 119185 281205
rect 105948 279515 110339 281071
rect 105948 274645 106086 279515
rect 110027 279211 110213 279515
rect 111020 279451 111226 281073
rect 111498 279451 112650 280904
rect 112944 280716 114379 281073
rect 112944 280120 114096 280716
rect 112974 280086 114096 280120
rect 112974 279451 114126 280086
rect 111020 279309 114292 279451
rect 109591 276574 110249 279211
rect 111020 277785 111226 279309
rect 111498 277785 112650 279309
rect 112944 279268 114292 279309
rect 112944 279050 114379 279268
rect 112944 278454 114096 279050
rect 112974 278420 114096 278454
rect 112974 277785 114126 278420
rect 111020 277643 114292 277785
rect 109591 276517 110250 276574
rect 110119 274645 110250 276517
rect 105948 274501 110250 274645
rect 111020 276119 111226 277643
rect 111498 276119 112650 277643
rect 112944 277602 114292 277643
rect 112944 277384 114379 277602
rect 112944 276788 114096 277384
rect 112974 276754 114096 276788
rect 112974 276119 114126 276754
rect 111020 275977 114292 276119
rect 111020 274453 111226 275977
rect 111498 274453 112650 275977
rect 112944 275936 114292 275977
rect 112944 275718 114379 275936
rect 112944 275122 114096 275718
rect 112974 275088 114096 275122
rect 112974 274453 114126 275088
rect 111020 274311 114292 274453
rect 106255 272760 110285 272977
rect 106255 270360 106485 272760
rect 106689 272273 108829 272393
rect 106689 271997 106815 272273
rect 107375 271997 108163 272273
rect 106689 271781 108163 271997
rect 106689 270827 106815 271781
rect 107375 271573 108163 271781
rect 107147 270827 108399 271573
rect 108703 270827 108829 272273
rect 106689 270707 108829 270827
rect 110055 270360 110285 272760
rect 111020 272787 111226 274311
rect 111498 272787 112650 274311
rect 112944 274270 114292 274311
rect 112944 274052 114379 274270
rect 112944 273456 114096 274052
rect 112974 273422 114096 273456
rect 112974 272792 114126 273422
rect 112974 272787 114292 272792
rect 111020 272645 114292 272787
rect 115826 280716 117261 281073
rect 116109 280120 117261 280716
rect 116109 280086 117231 280120
rect 116079 279451 117231 280086
rect 117555 279451 118707 280904
rect 118979 279451 119185 281073
rect 115913 279309 119185 279451
rect 115913 279268 117261 279309
rect 115826 279050 117261 279268
rect 116109 278454 117261 279050
rect 116109 278420 117231 278454
rect 116079 277785 117231 278420
rect 117555 277785 118707 279309
rect 118979 277785 119185 279309
rect 115913 277643 119185 277785
rect 115913 277602 117261 277643
rect 115826 277384 117261 277602
rect 116109 276788 117261 277384
rect 116109 276754 117231 276788
rect 116079 276119 117231 276754
rect 117555 276119 118707 277643
rect 118979 276119 119185 277643
rect 115913 275977 119185 276119
rect 115913 275936 117261 275977
rect 115826 275718 117261 275936
rect 116109 275122 117261 275718
rect 116109 275088 117231 275122
rect 116079 274453 117231 275088
rect 117555 274453 118707 275977
rect 118979 274453 119185 275977
rect 115913 274311 119185 274453
rect 115913 274270 117261 274311
rect 115826 274052 117261 274270
rect 116109 273456 117261 274052
rect 116109 273422 117231 273456
rect 116079 272792 117231 273422
rect 115913 272787 117231 272792
rect 117555 272787 118707 274311
rect 118979 272787 119185 274311
rect 114117 272577 114292 272645
rect 115913 272645 119185 272787
rect 119912 280986 125198 281191
rect 115913 272577 116088 272645
rect 106255 270143 110285 270360
rect 111913 272275 112095 272299
rect 114117 272275 116088 272577
rect 118995 272275 119177 272299
rect 111913 272099 119177 272275
rect 111913 268852 112095 272099
rect 115797 270798 119177 272099
rect 112476 269098 118804 270250
rect 118995 268852 119177 270798
rect 111913 268676 119177 268852
rect 119912 268887 120130 280986
rect 122001 276238 122170 278669
rect 122001 276071 124347 276238
rect 122001 275481 122170 276071
rect 122766 274608 124138 275062
rect 125021 274608 125197 280986
rect 122766 274588 125197 274608
rect 122034 274462 125197 274588
rect 122034 274358 124840 274462
rect 122036 273519 124840 274358
rect 125021 272803 125197 274462
rect 123952 269167 125197 272803
rect 125021 268887 125197 269167
rect 119912 268682 125225 268887
rect 111913 268625 112095 268676
rect 118995 268625 119177 268676
<< nmos >>
rect 106981 271807 107191 271971
<< pmos >>
rect 106951 274935 107129 275713
rect 107451 274935 107629 275713
rect 107951 274935 108129 275713
rect 108451 274935 108629 275713
rect 108951 274935 109129 275713
rect 109451 274935 109629 275713
rect 122414 277792 123290 278266
rect 122466 275711 122866 275811
rect 123102 275711 123502 275811
rect 123738 275711 124138 275811
rect 124374 275711 124774 275811
<< pmoslvt >>
rect 106368 278757 107582 279011
rect 106368 278157 107582 278411
rect 106491 277090 107525 277164
rect 109440 270706 109510 272426
rect 114657 280403 114857 280803
rect 114657 279957 114857 280117
rect 114657 279549 114857 279709
rect 115348 280403 115548 280803
rect 115348 279957 115548 280117
rect 115348 279549 115548 279709
rect 114657 278737 114857 279137
rect 114657 278291 114857 278451
rect 114657 277883 114857 278043
rect 115348 278737 115548 279137
rect 115348 278291 115548 278451
rect 115348 277883 115548 278043
rect 114657 277071 114857 277471
rect 114657 276625 114857 276785
rect 114657 276217 114857 276377
rect 115348 277071 115548 277471
rect 115348 276625 115548 276785
rect 115348 276217 115548 276377
rect 114657 275405 114857 275805
rect 114657 274959 114857 275119
rect 114657 274551 114857 274711
rect 115348 275405 115548 275805
rect 115348 274959 115548 275119
rect 115348 274551 115548 274711
rect 114657 273739 114857 274139
rect 114657 273293 114857 273453
rect 114657 272885 114857 273045
rect 115348 273739 115548 274139
rect 115348 273293 115548 273453
rect 115348 272885 115548 273045
rect 112578 271106 112738 271306
rect 112978 271106 113138 271306
rect 113378 271106 113538 271306
rect 113778 271106 113938 271306
rect 114637 271077 114797 271277
rect 115037 271077 115197 271277
rect 120429 280537 120829 280637
rect 121129 280537 121529 280637
rect 120429 279753 120829 280253
rect 121129 279753 121529 280253
rect 120429 278969 120829 279469
rect 121129 278969 121529 279469
rect 122356 279923 122756 280423
rect 123056 279923 123456 280423
rect 122356 279139 122756 279639
rect 123056 279139 123456 279639
rect 120429 278185 120829 278685
rect 121129 278185 121529 278685
rect 120429 277401 120829 277901
rect 121129 277401 121529 277901
rect 120429 276617 120829 277117
rect 121129 276617 121529 277117
rect 120429 275833 120829 276333
rect 121129 275833 121529 276333
rect 120429 275049 120829 275549
rect 121129 275049 121529 275549
rect 122416 277400 123216 277500
rect 123656 277394 124210 278080
rect 122438 276492 123832 276668
rect 120429 274265 120829 274765
rect 121129 274265 121529 274765
rect 120429 273481 120829 273981
rect 121129 273481 121529 273981
rect 120429 272697 120829 273197
rect 121129 272697 121529 273197
rect 120429 271913 120829 272413
rect 121129 271913 121529 272413
rect 120429 271129 120829 271629
rect 121129 271129 121529 271629
rect 120429 270345 120829 270845
rect 121129 270345 121529 270845
rect 120429 269561 120829 270061
rect 121129 269561 121529 270061
rect 120429 269177 120829 269277
rect 121129 269177 121529 269277
rect 122125 272713 122525 272813
rect 122825 272713 123225 272813
rect 122125 271929 122525 272429
rect 122825 271929 123225 272429
rect 122125 271145 122525 271645
rect 122825 271145 123225 271645
rect 122125 270361 122525 270861
rect 122825 270361 123225 270861
rect 122125 269577 122525 270077
rect 122825 269577 123225 270077
rect 122125 269193 122525 269293
rect 122825 269193 123225 269293
<< nmoslvt >>
rect 106357 279793 106489 280813
rect 106757 279793 106889 280813
rect 107157 279793 107289 280813
rect 107557 279793 107689 280813
rect 107957 279793 108089 280813
rect 108357 279793 108489 280813
rect 108757 279793 108889 280813
rect 109157 279793 109289 280813
rect 109557 279793 109689 280813
rect 109957 279793 110089 280813
rect 109777 277973 110063 279011
rect 109777 276717 110063 277755
rect 107459 271735 108079 272079
rect 107173 271311 108373 271489
rect 107173 270941 108373 271119
rect 111524 280660 112624 280820
rect 112970 280628 114070 280828
rect 111524 280300 112624 280460
rect 112970 280204 114070 280404
rect 111524 279940 112624 280100
rect 113000 279922 114100 280002
rect 111524 279580 112624 279740
rect 113000 279624 114100 279704
rect 116135 280628 117235 280828
rect 117581 280660 118681 280820
rect 116135 280204 117235 280404
rect 117581 280300 118681 280460
rect 116105 279922 117205 280002
rect 117581 279940 118681 280100
rect 116105 279624 117205 279704
rect 117581 279580 118681 279740
rect 111524 278994 112624 279154
rect 112970 278962 114070 279162
rect 111524 278634 112624 278794
rect 112970 278538 114070 278738
rect 111524 278274 112624 278434
rect 113000 278256 114100 278336
rect 111524 277914 112624 278074
rect 113000 277958 114100 278038
rect 116135 278962 117235 279162
rect 117581 278994 118681 279154
rect 116135 278538 117235 278738
rect 117581 278634 118681 278794
rect 116105 278256 117205 278336
rect 117581 278274 118681 278434
rect 116105 277958 117205 278038
rect 117581 277914 118681 278074
rect 111524 277328 112624 277488
rect 112970 277296 114070 277496
rect 111524 276968 112624 277128
rect 112970 276872 114070 277072
rect 111524 276608 112624 276768
rect 113000 276590 114100 276670
rect 111524 276248 112624 276408
rect 113000 276292 114100 276372
rect 116135 277296 117235 277496
rect 117581 277328 118681 277488
rect 116135 276872 117235 277072
rect 117581 276968 118681 277128
rect 116105 276590 117205 276670
rect 117581 276608 118681 276768
rect 116105 276292 117205 276372
rect 117581 276248 118681 276408
rect 111524 275662 112624 275822
rect 112970 275630 114070 275830
rect 111524 275302 112624 275462
rect 112970 275206 114070 275406
rect 111524 274942 112624 275102
rect 113000 274924 114100 275004
rect 111524 274582 112624 274742
rect 113000 274626 114100 274706
rect 116135 275630 117235 275830
rect 117581 275662 118681 275822
rect 116135 275206 117235 275406
rect 117581 275302 118681 275462
rect 116105 274924 117205 275004
rect 117581 274942 118681 275102
rect 116105 274626 117205 274706
rect 117581 274582 118681 274742
rect 111524 273996 112624 274156
rect 112970 273964 114070 274164
rect 111524 273636 112624 273796
rect 112970 273540 114070 273740
rect 111524 273276 112624 273436
rect 113000 273258 114100 273338
rect 111524 272916 112624 273076
rect 113000 272960 114100 273040
rect 116135 273964 117235 274164
rect 117581 273996 118681 274156
rect 116135 273540 117235 273740
rect 117581 273636 118681 273796
rect 116105 273258 117205 273338
rect 117581 273276 118681 273436
rect 116105 272960 117205 273040
rect 117581 272916 118681 273076
rect 115881 270824 116041 271924
rect 116281 270824 116441 271924
rect 116681 270824 116841 271924
rect 117081 270824 117241 271924
rect 117481 270824 117641 271924
rect 117881 270824 118041 271924
rect 118281 270824 118441 271924
rect 118681 270824 118841 271924
rect 112560 269124 112720 270224
rect 112960 269124 113120 270224
rect 113360 269124 113520 270224
rect 113760 269124 113920 270224
rect 114160 269124 114320 270224
rect 114560 269124 114720 270224
rect 114960 269124 115120 270224
rect 115360 269124 115520 270224
rect 115760 269124 115920 270224
rect 116160 269124 116320 270224
rect 116560 269124 116720 270224
rect 116960 269124 117120 270224
rect 117360 269124 117520 270224
rect 117760 269124 117920 270224
rect 118160 269124 118320 270224
rect 118560 269124 118720 270224
rect 122952 274662 123952 274862
rect 122277 273778 122477 274278
rect 122693 273778 122893 274278
rect 123109 273778 123309 274278
rect 123525 273778 123725 274278
rect 123941 273778 124141 274278
rect 124357 273778 124557 274278
rect 124192 272320 124692 272520
rect 124192 271904 124692 272104
rect 124192 271488 124692 271688
rect 124192 271072 124692 271272
rect 124192 270656 124692 270856
rect 124192 270240 124692 270440
rect 124192 269824 124692 270024
rect 124192 269408 124692 269608
<< ndiff >>
rect 106299 280796 106357 280813
rect 106299 280762 106311 280796
rect 106345 280762 106357 280796
rect 106299 280728 106357 280762
rect 106299 280694 106311 280728
rect 106345 280694 106357 280728
rect 106299 280660 106357 280694
rect 106299 280626 106311 280660
rect 106345 280626 106357 280660
rect 106299 280592 106357 280626
rect 106299 280558 106311 280592
rect 106345 280558 106357 280592
rect 106299 280524 106357 280558
rect 106299 280490 106311 280524
rect 106345 280490 106357 280524
rect 106299 280456 106357 280490
rect 106299 280422 106311 280456
rect 106345 280422 106357 280456
rect 106299 280388 106357 280422
rect 106299 280354 106311 280388
rect 106345 280354 106357 280388
rect 106299 280320 106357 280354
rect 106299 280286 106311 280320
rect 106345 280286 106357 280320
rect 106299 280252 106357 280286
rect 106299 280218 106311 280252
rect 106345 280218 106357 280252
rect 106299 280184 106357 280218
rect 106299 280150 106311 280184
rect 106345 280150 106357 280184
rect 106299 280116 106357 280150
rect 106299 280082 106311 280116
rect 106345 280082 106357 280116
rect 106299 280048 106357 280082
rect 106299 280014 106311 280048
rect 106345 280014 106357 280048
rect 106299 279980 106357 280014
rect 106299 279946 106311 279980
rect 106345 279946 106357 279980
rect 106299 279912 106357 279946
rect 106299 279878 106311 279912
rect 106345 279878 106357 279912
rect 106299 279844 106357 279878
rect 106299 279810 106311 279844
rect 106345 279810 106357 279844
rect 106299 279793 106357 279810
rect 106489 280796 106547 280813
rect 106489 280762 106501 280796
rect 106535 280762 106547 280796
rect 106489 280728 106547 280762
rect 106489 280694 106501 280728
rect 106535 280694 106547 280728
rect 106489 280660 106547 280694
rect 106489 280626 106501 280660
rect 106535 280626 106547 280660
rect 106489 280592 106547 280626
rect 106489 280558 106501 280592
rect 106535 280558 106547 280592
rect 106489 280524 106547 280558
rect 106489 280490 106501 280524
rect 106535 280490 106547 280524
rect 106489 280456 106547 280490
rect 106489 280422 106501 280456
rect 106535 280422 106547 280456
rect 106489 280388 106547 280422
rect 106489 280354 106501 280388
rect 106535 280354 106547 280388
rect 106489 280320 106547 280354
rect 106489 280286 106501 280320
rect 106535 280286 106547 280320
rect 106489 280252 106547 280286
rect 106489 280218 106501 280252
rect 106535 280218 106547 280252
rect 106489 280184 106547 280218
rect 106489 280150 106501 280184
rect 106535 280150 106547 280184
rect 106489 280116 106547 280150
rect 106489 280082 106501 280116
rect 106535 280082 106547 280116
rect 106489 280048 106547 280082
rect 106489 280014 106501 280048
rect 106535 280014 106547 280048
rect 106489 279980 106547 280014
rect 106489 279946 106501 279980
rect 106535 279946 106547 279980
rect 106489 279912 106547 279946
rect 106489 279878 106501 279912
rect 106535 279878 106547 279912
rect 106489 279844 106547 279878
rect 106489 279810 106501 279844
rect 106535 279810 106547 279844
rect 106489 279793 106547 279810
rect 106699 280796 106757 280813
rect 106699 280762 106711 280796
rect 106745 280762 106757 280796
rect 106699 280728 106757 280762
rect 106699 280694 106711 280728
rect 106745 280694 106757 280728
rect 106699 280660 106757 280694
rect 106699 280626 106711 280660
rect 106745 280626 106757 280660
rect 106699 280592 106757 280626
rect 106699 280558 106711 280592
rect 106745 280558 106757 280592
rect 106699 280524 106757 280558
rect 106699 280490 106711 280524
rect 106745 280490 106757 280524
rect 106699 280456 106757 280490
rect 106699 280422 106711 280456
rect 106745 280422 106757 280456
rect 106699 280388 106757 280422
rect 106699 280354 106711 280388
rect 106745 280354 106757 280388
rect 106699 280320 106757 280354
rect 106699 280286 106711 280320
rect 106745 280286 106757 280320
rect 106699 280252 106757 280286
rect 106699 280218 106711 280252
rect 106745 280218 106757 280252
rect 106699 280184 106757 280218
rect 106699 280150 106711 280184
rect 106745 280150 106757 280184
rect 106699 280116 106757 280150
rect 106699 280082 106711 280116
rect 106745 280082 106757 280116
rect 106699 280048 106757 280082
rect 106699 280014 106711 280048
rect 106745 280014 106757 280048
rect 106699 279980 106757 280014
rect 106699 279946 106711 279980
rect 106745 279946 106757 279980
rect 106699 279912 106757 279946
rect 106699 279878 106711 279912
rect 106745 279878 106757 279912
rect 106699 279844 106757 279878
rect 106699 279810 106711 279844
rect 106745 279810 106757 279844
rect 106699 279793 106757 279810
rect 106889 280796 106947 280813
rect 106889 280762 106901 280796
rect 106935 280762 106947 280796
rect 106889 280728 106947 280762
rect 106889 280694 106901 280728
rect 106935 280694 106947 280728
rect 106889 280660 106947 280694
rect 106889 280626 106901 280660
rect 106935 280626 106947 280660
rect 106889 280592 106947 280626
rect 106889 280558 106901 280592
rect 106935 280558 106947 280592
rect 106889 280524 106947 280558
rect 106889 280490 106901 280524
rect 106935 280490 106947 280524
rect 106889 280456 106947 280490
rect 106889 280422 106901 280456
rect 106935 280422 106947 280456
rect 106889 280388 106947 280422
rect 106889 280354 106901 280388
rect 106935 280354 106947 280388
rect 106889 280320 106947 280354
rect 106889 280286 106901 280320
rect 106935 280286 106947 280320
rect 106889 280252 106947 280286
rect 106889 280218 106901 280252
rect 106935 280218 106947 280252
rect 106889 280184 106947 280218
rect 106889 280150 106901 280184
rect 106935 280150 106947 280184
rect 106889 280116 106947 280150
rect 106889 280082 106901 280116
rect 106935 280082 106947 280116
rect 106889 280048 106947 280082
rect 106889 280014 106901 280048
rect 106935 280014 106947 280048
rect 106889 279980 106947 280014
rect 106889 279946 106901 279980
rect 106935 279946 106947 279980
rect 106889 279912 106947 279946
rect 106889 279878 106901 279912
rect 106935 279878 106947 279912
rect 106889 279844 106947 279878
rect 106889 279810 106901 279844
rect 106935 279810 106947 279844
rect 106889 279793 106947 279810
rect 107099 280796 107157 280813
rect 107099 280762 107111 280796
rect 107145 280762 107157 280796
rect 107099 280728 107157 280762
rect 107099 280694 107111 280728
rect 107145 280694 107157 280728
rect 107099 280660 107157 280694
rect 107099 280626 107111 280660
rect 107145 280626 107157 280660
rect 107099 280592 107157 280626
rect 107099 280558 107111 280592
rect 107145 280558 107157 280592
rect 107099 280524 107157 280558
rect 107099 280490 107111 280524
rect 107145 280490 107157 280524
rect 107099 280456 107157 280490
rect 107099 280422 107111 280456
rect 107145 280422 107157 280456
rect 107099 280388 107157 280422
rect 107099 280354 107111 280388
rect 107145 280354 107157 280388
rect 107099 280320 107157 280354
rect 107099 280286 107111 280320
rect 107145 280286 107157 280320
rect 107099 280252 107157 280286
rect 107099 280218 107111 280252
rect 107145 280218 107157 280252
rect 107099 280184 107157 280218
rect 107099 280150 107111 280184
rect 107145 280150 107157 280184
rect 107099 280116 107157 280150
rect 107099 280082 107111 280116
rect 107145 280082 107157 280116
rect 107099 280048 107157 280082
rect 107099 280014 107111 280048
rect 107145 280014 107157 280048
rect 107099 279980 107157 280014
rect 107099 279946 107111 279980
rect 107145 279946 107157 279980
rect 107099 279912 107157 279946
rect 107099 279878 107111 279912
rect 107145 279878 107157 279912
rect 107099 279844 107157 279878
rect 107099 279810 107111 279844
rect 107145 279810 107157 279844
rect 107099 279793 107157 279810
rect 107289 280796 107347 280813
rect 107289 280762 107301 280796
rect 107335 280762 107347 280796
rect 107289 280728 107347 280762
rect 107289 280694 107301 280728
rect 107335 280694 107347 280728
rect 107289 280660 107347 280694
rect 107289 280626 107301 280660
rect 107335 280626 107347 280660
rect 107289 280592 107347 280626
rect 107289 280558 107301 280592
rect 107335 280558 107347 280592
rect 107289 280524 107347 280558
rect 107289 280490 107301 280524
rect 107335 280490 107347 280524
rect 107289 280456 107347 280490
rect 107289 280422 107301 280456
rect 107335 280422 107347 280456
rect 107289 280388 107347 280422
rect 107289 280354 107301 280388
rect 107335 280354 107347 280388
rect 107289 280320 107347 280354
rect 107289 280286 107301 280320
rect 107335 280286 107347 280320
rect 107289 280252 107347 280286
rect 107289 280218 107301 280252
rect 107335 280218 107347 280252
rect 107289 280184 107347 280218
rect 107289 280150 107301 280184
rect 107335 280150 107347 280184
rect 107289 280116 107347 280150
rect 107289 280082 107301 280116
rect 107335 280082 107347 280116
rect 107289 280048 107347 280082
rect 107289 280014 107301 280048
rect 107335 280014 107347 280048
rect 107289 279980 107347 280014
rect 107289 279946 107301 279980
rect 107335 279946 107347 279980
rect 107289 279912 107347 279946
rect 107289 279878 107301 279912
rect 107335 279878 107347 279912
rect 107289 279844 107347 279878
rect 107289 279810 107301 279844
rect 107335 279810 107347 279844
rect 107289 279793 107347 279810
rect 107499 280796 107557 280813
rect 107499 280762 107511 280796
rect 107545 280762 107557 280796
rect 107499 280728 107557 280762
rect 107499 280694 107511 280728
rect 107545 280694 107557 280728
rect 107499 280660 107557 280694
rect 107499 280626 107511 280660
rect 107545 280626 107557 280660
rect 107499 280592 107557 280626
rect 107499 280558 107511 280592
rect 107545 280558 107557 280592
rect 107499 280524 107557 280558
rect 107499 280490 107511 280524
rect 107545 280490 107557 280524
rect 107499 280456 107557 280490
rect 107499 280422 107511 280456
rect 107545 280422 107557 280456
rect 107499 280388 107557 280422
rect 107499 280354 107511 280388
rect 107545 280354 107557 280388
rect 107499 280320 107557 280354
rect 107499 280286 107511 280320
rect 107545 280286 107557 280320
rect 107499 280252 107557 280286
rect 107499 280218 107511 280252
rect 107545 280218 107557 280252
rect 107499 280184 107557 280218
rect 107499 280150 107511 280184
rect 107545 280150 107557 280184
rect 107499 280116 107557 280150
rect 107499 280082 107511 280116
rect 107545 280082 107557 280116
rect 107499 280048 107557 280082
rect 107499 280014 107511 280048
rect 107545 280014 107557 280048
rect 107499 279980 107557 280014
rect 107499 279946 107511 279980
rect 107545 279946 107557 279980
rect 107499 279912 107557 279946
rect 107499 279878 107511 279912
rect 107545 279878 107557 279912
rect 107499 279844 107557 279878
rect 107499 279810 107511 279844
rect 107545 279810 107557 279844
rect 107499 279793 107557 279810
rect 107689 280796 107747 280813
rect 107689 280762 107701 280796
rect 107735 280762 107747 280796
rect 107689 280728 107747 280762
rect 107689 280694 107701 280728
rect 107735 280694 107747 280728
rect 107689 280660 107747 280694
rect 107689 280626 107701 280660
rect 107735 280626 107747 280660
rect 107689 280592 107747 280626
rect 107689 280558 107701 280592
rect 107735 280558 107747 280592
rect 107689 280524 107747 280558
rect 107689 280490 107701 280524
rect 107735 280490 107747 280524
rect 107689 280456 107747 280490
rect 107689 280422 107701 280456
rect 107735 280422 107747 280456
rect 107689 280388 107747 280422
rect 107689 280354 107701 280388
rect 107735 280354 107747 280388
rect 107689 280320 107747 280354
rect 107689 280286 107701 280320
rect 107735 280286 107747 280320
rect 107689 280252 107747 280286
rect 107689 280218 107701 280252
rect 107735 280218 107747 280252
rect 107689 280184 107747 280218
rect 107689 280150 107701 280184
rect 107735 280150 107747 280184
rect 107689 280116 107747 280150
rect 107689 280082 107701 280116
rect 107735 280082 107747 280116
rect 107689 280048 107747 280082
rect 107689 280014 107701 280048
rect 107735 280014 107747 280048
rect 107689 279980 107747 280014
rect 107689 279946 107701 279980
rect 107735 279946 107747 279980
rect 107689 279912 107747 279946
rect 107689 279878 107701 279912
rect 107735 279878 107747 279912
rect 107689 279844 107747 279878
rect 107689 279810 107701 279844
rect 107735 279810 107747 279844
rect 107689 279793 107747 279810
rect 107899 280796 107957 280813
rect 107899 280762 107911 280796
rect 107945 280762 107957 280796
rect 107899 280728 107957 280762
rect 107899 280694 107911 280728
rect 107945 280694 107957 280728
rect 107899 280660 107957 280694
rect 107899 280626 107911 280660
rect 107945 280626 107957 280660
rect 107899 280592 107957 280626
rect 107899 280558 107911 280592
rect 107945 280558 107957 280592
rect 107899 280524 107957 280558
rect 107899 280490 107911 280524
rect 107945 280490 107957 280524
rect 107899 280456 107957 280490
rect 107899 280422 107911 280456
rect 107945 280422 107957 280456
rect 107899 280388 107957 280422
rect 107899 280354 107911 280388
rect 107945 280354 107957 280388
rect 107899 280320 107957 280354
rect 107899 280286 107911 280320
rect 107945 280286 107957 280320
rect 107899 280252 107957 280286
rect 107899 280218 107911 280252
rect 107945 280218 107957 280252
rect 107899 280184 107957 280218
rect 107899 280150 107911 280184
rect 107945 280150 107957 280184
rect 107899 280116 107957 280150
rect 107899 280082 107911 280116
rect 107945 280082 107957 280116
rect 107899 280048 107957 280082
rect 107899 280014 107911 280048
rect 107945 280014 107957 280048
rect 107899 279980 107957 280014
rect 107899 279946 107911 279980
rect 107945 279946 107957 279980
rect 107899 279912 107957 279946
rect 107899 279878 107911 279912
rect 107945 279878 107957 279912
rect 107899 279844 107957 279878
rect 107899 279810 107911 279844
rect 107945 279810 107957 279844
rect 107899 279793 107957 279810
rect 108089 280796 108147 280813
rect 108089 280762 108101 280796
rect 108135 280762 108147 280796
rect 108089 280728 108147 280762
rect 108089 280694 108101 280728
rect 108135 280694 108147 280728
rect 108089 280660 108147 280694
rect 108089 280626 108101 280660
rect 108135 280626 108147 280660
rect 108089 280592 108147 280626
rect 108089 280558 108101 280592
rect 108135 280558 108147 280592
rect 108089 280524 108147 280558
rect 108089 280490 108101 280524
rect 108135 280490 108147 280524
rect 108089 280456 108147 280490
rect 108089 280422 108101 280456
rect 108135 280422 108147 280456
rect 108089 280388 108147 280422
rect 108089 280354 108101 280388
rect 108135 280354 108147 280388
rect 108089 280320 108147 280354
rect 108089 280286 108101 280320
rect 108135 280286 108147 280320
rect 108089 280252 108147 280286
rect 108089 280218 108101 280252
rect 108135 280218 108147 280252
rect 108089 280184 108147 280218
rect 108089 280150 108101 280184
rect 108135 280150 108147 280184
rect 108089 280116 108147 280150
rect 108089 280082 108101 280116
rect 108135 280082 108147 280116
rect 108089 280048 108147 280082
rect 108089 280014 108101 280048
rect 108135 280014 108147 280048
rect 108089 279980 108147 280014
rect 108089 279946 108101 279980
rect 108135 279946 108147 279980
rect 108089 279912 108147 279946
rect 108089 279878 108101 279912
rect 108135 279878 108147 279912
rect 108089 279844 108147 279878
rect 108089 279810 108101 279844
rect 108135 279810 108147 279844
rect 108089 279793 108147 279810
rect 108299 280796 108357 280813
rect 108299 280762 108311 280796
rect 108345 280762 108357 280796
rect 108299 280728 108357 280762
rect 108299 280694 108311 280728
rect 108345 280694 108357 280728
rect 108299 280660 108357 280694
rect 108299 280626 108311 280660
rect 108345 280626 108357 280660
rect 108299 280592 108357 280626
rect 108299 280558 108311 280592
rect 108345 280558 108357 280592
rect 108299 280524 108357 280558
rect 108299 280490 108311 280524
rect 108345 280490 108357 280524
rect 108299 280456 108357 280490
rect 108299 280422 108311 280456
rect 108345 280422 108357 280456
rect 108299 280388 108357 280422
rect 108299 280354 108311 280388
rect 108345 280354 108357 280388
rect 108299 280320 108357 280354
rect 108299 280286 108311 280320
rect 108345 280286 108357 280320
rect 108299 280252 108357 280286
rect 108299 280218 108311 280252
rect 108345 280218 108357 280252
rect 108299 280184 108357 280218
rect 108299 280150 108311 280184
rect 108345 280150 108357 280184
rect 108299 280116 108357 280150
rect 108299 280082 108311 280116
rect 108345 280082 108357 280116
rect 108299 280048 108357 280082
rect 108299 280014 108311 280048
rect 108345 280014 108357 280048
rect 108299 279980 108357 280014
rect 108299 279946 108311 279980
rect 108345 279946 108357 279980
rect 108299 279912 108357 279946
rect 108299 279878 108311 279912
rect 108345 279878 108357 279912
rect 108299 279844 108357 279878
rect 108299 279810 108311 279844
rect 108345 279810 108357 279844
rect 108299 279793 108357 279810
rect 108489 280796 108547 280813
rect 108489 280762 108501 280796
rect 108535 280762 108547 280796
rect 108489 280728 108547 280762
rect 108489 280694 108501 280728
rect 108535 280694 108547 280728
rect 108489 280660 108547 280694
rect 108489 280626 108501 280660
rect 108535 280626 108547 280660
rect 108489 280592 108547 280626
rect 108489 280558 108501 280592
rect 108535 280558 108547 280592
rect 108489 280524 108547 280558
rect 108489 280490 108501 280524
rect 108535 280490 108547 280524
rect 108489 280456 108547 280490
rect 108489 280422 108501 280456
rect 108535 280422 108547 280456
rect 108489 280388 108547 280422
rect 108489 280354 108501 280388
rect 108535 280354 108547 280388
rect 108489 280320 108547 280354
rect 108489 280286 108501 280320
rect 108535 280286 108547 280320
rect 108489 280252 108547 280286
rect 108489 280218 108501 280252
rect 108535 280218 108547 280252
rect 108489 280184 108547 280218
rect 108489 280150 108501 280184
rect 108535 280150 108547 280184
rect 108489 280116 108547 280150
rect 108489 280082 108501 280116
rect 108535 280082 108547 280116
rect 108489 280048 108547 280082
rect 108489 280014 108501 280048
rect 108535 280014 108547 280048
rect 108489 279980 108547 280014
rect 108489 279946 108501 279980
rect 108535 279946 108547 279980
rect 108489 279912 108547 279946
rect 108489 279878 108501 279912
rect 108535 279878 108547 279912
rect 108489 279844 108547 279878
rect 108489 279810 108501 279844
rect 108535 279810 108547 279844
rect 108489 279793 108547 279810
rect 108699 280796 108757 280813
rect 108699 280762 108711 280796
rect 108745 280762 108757 280796
rect 108699 280728 108757 280762
rect 108699 280694 108711 280728
rect 108745 280694 108757 280728
rect 108699 280660 108757 280694
rect 108699 280626 108711 280660
rect 108745 280626 108757 280660
rect 108699 280592 108757 280626
rect 108699 280558 108711 280592
rect 108745 280558 108757 280592
rect 108699 280524 108757 280558
rect 108699 280490 108711 280524
rect 108745 280490 108757 280524
rect 108699 280456 108757 280490
rect 108699 280422 108711 280456
rect 108745 280422 108757 280456
rect 108699 280388 108757 280422
rect 108699 280354 108711 280388
rect 108745 280354 108757 280388
rect 108699 280320 108757 280354
rect 108699 280286 108711 280320
rect 108745 280286 108757 280320
rect 108699 280252 108757 280286
rect 108699 280218 108711 280252
rect 108745 280218 108757 280252
rect 108699 280184 108757 280218
rect 108699 280150 108711 280184
rect 108745 280150 108757 280184
rect 108699 280116 108757 280150
rect 108699 280082 108711 280116
rect 108745 280082 108757 280116
rect 108699 280048 108757 280082
rect 108699 280014 108711 280048
rect 108745 280014 108757 280048
rect 108699 279980 108757 280014
rect 108699 279946 108711 279980
rect 108745 279946 108757 279980
rect 108699 279912 108757 279946
rect 108699 279878 108711 279912
rect 108745 279878 108757 279912
rect 108699 279844 108757 279878
rect 108699 279810 108711 279844
rect 108745 279810 108757 279844
rect 108699 279793 108757 279810
rect 108889 280796 108947 280813
rect 108889 280762 108901 280796
rect 108935 280762 108947 280796
rect 108889 280728 108947 280762
rect 108889 280694 108901 280728
rect 108935 280694 108947 280728
rect 108889 280660 108947 280694
rect 108889 280626 108901 280660
rect 108935 280626 108947 280660
rect 108889 280592 108947 280626
rect 108889 280558 108901 280592
rect 108935 280558 108947 280592
rect 108889 280524 108947 280558
rect 108889 280490 108901 280524
rect 108935 280490 108947 280524
rect 108889 280456 108947 280490
rect 108889 280422 108901 280456
rect 108935 280422 108947 280456
rect 108889 280388 108947 280422
rect 108889 280354 108901 280388
rect 108935 280354 108947 280388
rect 108889 280320 108947 280354
rect 108889 280286 108901 280320
rect 108935 280286 108947 280320
rect 108889 280252 108947 280286
rect 108889 280218 108901 280252
rect 108935 280218 108947 280252
rect 108889 280184 108947 280218
rect 108889 280150 108901 280184
rect 108935 280150 108947 280184
rect 108889 280116 108947 280150
rect 108889 280082 108901 280116
rect 108935 280082 108947 280116
rect 108889 280048 108947 280082
rect 108889 280014 108901 280048
rect 108935 280014 108947 280048
rect 108889 279980 108947 280014
rect 108889 279946 108901 279980
rect 108935 279946 108947 279980
rect 108889 279912 108947 279946
rect 108889 279878 108901 279912
rect 108935 279878 108947 279912
rect 108889 279844 108947 279878
rect 108889 279810 108901 279844
rect 108935 279810 108947 279844
rect 108889 279793 108947 279810
rect 109099 280796 109157 280813
rect 109099 280762 109111 280796
rect 109145 280762 109157 280796
rect 109099 280728 109157 280762
rect 109099 280694 109111 280728
rect 109145 280694 109157 280728
rect 109099 280660 109157 280694
rect 109099 280626 109111 280660
rect 109145 280626 109157 280660
rect 109099 280592 109157 280626
rect 109099 280558 109111 280592
rect 109145 280558 109157 280592
rect 109099 280524 109157 280558
rect 109099 280490 109111 280524
rect 109145 280490 109157 280524
rect 109099 280456 109157 280490
rect 109099 280422 109111 280456
rect 109145 280422 109157 280456
rect 109099 280388 109157 280422
rect 109099 280354 109111 280388
rect 109145 280354 109157 280388
rect 109099 280320 109157 280354
rect 109099 280286 109111 280320
rect 109145 280286 109157 280320
rect 109099 280252 109157 280286
rect 109099 280218 109111 280252
rect 109145 280218 109157 280252
rect 109099 280184 109157 280218
rect 109099 280150 109111 280184
rect 109145 280150 109157 280184
rect 109099 280116 109157 280150
rect 109099 280082 109111 280116
rect 109145 280082 109157 280116
rect 109099 280048 109157 280082
rect 109099 280014 109111 280048
rect 109145 280014 109157 280048
rect 109099 279980 109157 280014
rect 109099 279946 109111 279980
rect 109145 279946 109157 279980
rect 109099 279912 109157 279946
rect 109099 279878 109111 279912
rect 109145 279878 109157 279912
rect 109099 279844 109157 279878
rect 109099 279810 109111 279844
rect 109145 279810 109157 279844
rect 109099 279793 109157 279810
rect 109289 280796 109347 280813
rect 109289 280762 109301 280796
rect 109335 280762 109347 280796
rect 109289 280728 109347 280762
rect 109289 280694 109301 280728
rect 109335 280694 109347 280728
rect 109289 280660 109347 280694
rect 109289 280626 109301 280660
rect 109335 280626 109347 280660
rect 109289 280592 109347 280626
rect 109289 280558 109301 280592
rect 109335 280558 109347 280592
rect 109289 280524 109347 280558
rect 109289 280490 109301 280524
rect 109335 280490 109347 280524
rect 109289 280456 109347 280490
rect 109289 280422 109301 280456
rect 109335 280422 109347 280456
rect 109289 280388 109347 280422
rect 109289 280354 109301 280388
rect 109335 280354 109347 280388
rect 109289 280320 109347 280354
rect 109289 280286 109301 280320
rect 109335 280286 109347 280320
rect 109289 280252 109347 280286
rect 109289 280218 109301 280252
rect 109335 280218 109347 280252
rect 109289 280184 109347 280218
rect 109289 280150 109301 280184
rect 109335 280150 109347 280184
rect 109289 280116 109347 280150
rect 109289 280082 109301 280116
rect 109335 280082 109347 280116
rect 109289 280048 109347 280082
rect 109289 280014 109301 280048
rect 109335 280014 109347 280048
rect 109289 279980 109347 280014
rect 109289 279946 109301 279980
rect 109335 279946 109347 279980
rect 109289 279912 109347 279946
rect 109289 279878 109301 279912
rect 109335 279878 109347 279912
rect 109289 279844 109347 279878
rect 109289 279810 109301 279844
rect 109335 279810 109347 279844
rect 109289 279793 109347 279810
rect 109499 280796 109557 280813
rect 109499 280762 109511 280796
rect 109545 280762 109557 280796
rect 109499 280728 109557 280762
rect 109499 280694 109511 280728
rect 109545 280694 109557 280728
rect 109499 280660 109557 280694
rect 109499 280626 109511 280660
rect 109545 280626 109557 280660
rect 109499 280592 109557 280626
rect 109499 280558 109511 280592
rect 109545 280558 109557 280592
rect 109499 280524 109557 280558
rect 109499 280490 109511 280524
rect 109545 280490 109557 280524
rect 109499 280456 109557 280490
rect 109499 280422 109511 280456
rect 109545 280422 109557 280456
rect 109499 280388 109557 280422
rect 109499 280354 109511 280388
rect 109545 280354 109557 280388
rect 109499 280320 109557 280354
rect 109499 280286 109511 280320
rect 109545 280286 109557 280320
rect 109499 280252 109557 280286
rect 109499 280218 109511 280252
rect 109545 280218 109557 280252
rect 109499 280184 109557 280218
rect 109499 280150 109511 280184
rect 109545 280150 109557 280184
rect 109499 280116 109557 280150
rect 109499 280082 109511 280116
rect 109545 280082 109557 280116
rect 109499 280048 109557 280082
rect 109499 280014 109511 280048
rect 109545 280014 109557 280048
rect 109499 279980 109557 280014
rect 109499 279946 109511 279980
rect 109545 279946 109557 279980
rect 109499 279912 109557 279946
rect 109499 279878 109511 279912
rect 109545 279878 109557 279912
rect 109499 279844 109557 279878
rect 109499 279810 109511 279844
rect 109545 279810 109557 279844
rect 109499 279793 109557 279810
rect 109689 280796 109747 280813
rect 109689 280762 109701 280796
rect 109735 280762 109747 280796
rect 109689 280728 109747 280762
rect 109689 280694 109701 280728
rect 109735 280694 109747 280728
rect 109689 280660 109747 280694
rect 109689 280626 109701 280660
rect 109735 280626 109747 280660
rect 109689 280592 109747 280626
rect 109689 280558 109701 280592
rect 109735 280558 109747 280592
rect 109689 280524 109747 280558
rect 109689 280490 109701 280524
rect 109735 280490 109747 280524
rect 109689 280456 109747 280490
rect 109689 280422 109701 280456
rect 109735 280422 109747 280456
rect 109689 280388 109747 280422
rect 109689 280354 109701 280388
rect 109735 280354 109747 280388
rect 109689 280320 109747 280354
rect 109689 280286 109701 280320
rect 109735 280286 109747 280320
rect 109689 280252 109747 280286
rect 109689 280218 109701 280252
rect 109735 280218 109747 280252
rect 109689 280184 109747 280218
rect 109689 280150 109701 280184
rect 109735 280150 109747 280184
rect 109689 280116 109747 280150
rect 109689 280082 109701 280116
rect 109735 280082 109747 280116
rect 109689 280048 109747 280082
rect 109689 280014 109701 280048
rect 109735 280014 109747 280048
rect 109689 279980 109747 280014
rect 109689 279946 109701 279980
rect 109735 279946 109747 279980
rect 109689 279912 109747 279946
rect 109689 279878 109701 279912
rect 109735 279878 109747 279912
rect 109689 279844 109747 279878
rect 109689 279810 109701 279844
rect 109735 279810 109747 279844
rect 109689 279793 109747 279810
rect 109899 280796 109957 280813
rect 109899 280762 109911 280796
rect 109945 280762 109957 280796
rect 109899 280728 109957 280762
rect 109899 280694 109911 280728
rect 109945 280694 109957 280728
rect 109899 280660 109957 280694
rect 109899 280626 109911 280660
rect 109945 280626 109957 280660
rect 109899 280592 109957 280626
rect 109899 280558 109911 280592
rect 109945 280558 109957 280592
rect 109899 280524 109957 280558
rect 109899 280490 109911 280524
rect 109945 280490 109957 280524
rect 109899 280456 109957 280490
rect 109899 280422 109911 280456
rect 109945 280422 109957 280456
rect 109899 280388 109957 280422
rect 109899 280354 109911 280388
rect 109945 280354 109957 280388
rect 109899 280320 109957 280354
rect 109899 280286 109911 280320
rect 109945 280286 109957 280320
rect 109899 280252 109957 280286
rect 109899 280218 109911 280252
rect 109945 280218 109957 280252
rect 109899 280184 109957 280218
rect 109899 280150 109911 280184
rect 109945 280150 109957 280184
rect 109899 280116 109957 280150
rect 109899 280082 109911 280116
rect 109945 280082 109957 280116
rect 109899 280048 109957 280082
rect 109899 280014 109911 280048
rect 109945 280014 109957 280048
rect 109899 279980 109957 280014
rect 109899 279946 109911 279980
rect 109945 279946 109957 279980
rect 109899 279912 109957 279946
rect 109899 279878 109911 279912
rect 109945 279878 109957 279912
rect 109899 279844 109957 279878
rect 109899 279810 109911 279844
rect 109945 279810 109957 279844
rect 109899 279793 109957 279810
rect 110089 280796 110147 280813
rect 110089 280762 110101 280796
rect 110135 280762 110147 280796
rect 110089 280728 110147 280762
rect 110089 280694 110101 280728
rect 110135 280694 110147 280728
rect 110089 280660 110147 280694
rect 110089 280626 110101 280660
rect 110135 280626 110147 280660
rect 110089 280592 110147 280626
rect 110089 280558 110101 280592
rect 110135 280558 110147 280592
rect 110089 280524 110147 280558
rect 110089 280490 110101 280524
rect 110135 280490 110147 280524
rect 110089 280456 110147 280490
rect 110089 280422 110101 280456
rect 110135 280422 110147 280456
rect 110089 280388 110147 280422
rect 110089 280354 110101 280388
rect 110135 280354 110147 280388
rect 110089 280320 110147 280354
rect 110089 280286 110101 280320
rect 110135 280286 110147 280320
rect 110089 280252 110147 280286
rect 110089 280218 110101 280252
rect 110135 280218 110147 280252
rect 110089 280184 110147 280218
rect 110089 280150 110101 280184
rect 110135 280150 110147 280184
rect 110089 280116 110147 280150
rect 110089 280082 110101 280116
rect 110135 280082 110147 280116
rect 110089 280048 110147 280082
rect 110089 280014 110101 280048
rect 110135 280014 110147 280048
rect 110089 279980 110147 280014
rect 110089 279946 110101 279980
rect 110135 279946 110147 279980
rect 110089 279912 110147 279946
rect 110089 279878 110101 279912
rect 110135 279878 110147 279912
rect 110089 279844 110147 279878
rect 110089 279810 110101 279844
rect 110135 279810 110147 279844
rect 110089 279793 110147 279810
rect 109719 278985 109777 279011
rect 109719 278951 109731 278985
rect 109765 278951 109777 278985
rect 109719 278917 109777 278951
rect 109719 278883 109731 278917
rect 109765 278883 109777 278917
rect 109719 278849 109777 278883
rect 109719 278815 109731 278849
rect 109765 278815 109777 278849
rect 109719 278781 109777 278815
rect 109719 278747 109731 278781
rect 109765 278747 109777 278781
rect 109719 278713 109777 278747
rect 109719 278679 109731 278713
rect 109765 278679 109777 278713
rect 109719 278645 109777 278679
rect 109719 278611 109731 278645
rect 109765 278611 109777 278645
rect 109719 278577 109777 278611
rect 109719 278543 109731 278577
rect 109765 278543 109777 278577
rect 109719 278509 109777 278543
rect 109719 278475 109731 278509
rect 109765 278475 109777 278509
rect 109719 278441 109777 278475
rect 109719 278407 109731 278441
rect 109765 278407 109777 278441
rect 109719 278373 109777 278407
rect 109719 278339 109731 278373
rect 109765 278339 109777 278373
rect 109719 278305 109777 278339
rect 109719 278271 109731 278305
rect 109765 278271 109777 278305
rect 109719 278237 109777 278271
rect 109719 278203 109731 278237
rect 109765 278203 109777 278237
rect 109719 278169 109777 278203
rect 109719 278135 109731 278169
rect 109765 278135 109777 278169
rect 109719 278101 109777 278135
rect 109719 278067 109731 278101
rect 109765 278067 109777 278101
rect 109719 278033 109777 278067
rect 109719 277999 109731 278033
rect 109765 277999 109777 278033
rect 109719 277973 109777 277999
rect 110063 278985 110121 279011
rect 110063 278951 110075 278985
rect 110109 278951 110121 278985
rect 110063 278917 110121 278951
rect 110063 278883 110075 278917
rect 110109 278883 110121 278917
rect 110063 278849 110121 278883
rect 110063 278815 110075 278849
rect 110109 278815 110121 278849
rect 110063 278781 110121 278815
rect 110063 278747 110075 278781
rect 110109 278747 110121 278781
rect 110063 278713 110121 278747
rect 110063 278679 110075 278713
rect 110109 278679 110121 278713
rect 110063 278645 110121 278679
rect 110063 278611 110075 278645
rect 110109 278611 110121 278645
rect 110063 278577 110121 278611
rect 110063 278543 110075 278577
rect 110109 278543 110121 278577
rect 110063 278509 110121 278543
rect 110063 278475 110075 278509
rect 110109 278475 110121 278509
rect 110063 278441 110121 278475
rect 110063 278407 110075 278441
rect 110109 278407 110121 278441
rect 110063 278373 110121 278407
rect 110063 278339 110075 278373
rect 110109 278339 110121 278373
rect 110063 278305 110121 278339
rect 110063 278271 110075 278305
rect 110109 278271 110121 278305
rect 110063 278237 110121 278271
rect 110063 278203 110075 278237
rect 110109 278203 110121 278237
rect 110063 278169 110121 278203
rect 110063 278135 110075 278169
rect 110109 278135 110121 278169
rect 110063 278101 110121 278135
rect 110063 278067 110075 278101
rect 110109 278067 110121 278101
rect 110063 278033 110121 278067
rect 110063 277999 110075 278033
rect 110109 277999 110121 278033
rect 110063 277973 110121 277999
rect 109719 277729 109777 277755
rect 109719 277695 109731 277729
rect 109765 277695 109777 277729
rect 109719 277661 109777 277695
rect 109719 277627 109731 277661
rect 109765 277627 109777 277661
rect 109719 277593 109777 277627
rect 109719 277559 109731 277593
rect 109765 277559 109777 277593
rect 109719 277525 109777 277559
rect 109719 277491 109731 277525
rect 109765 277491 109777 277525
rect 109719 277457 109777 277491
rect 109719 277423 109731 277457
rect 109765 277423 109777 277457
rect 109719 277389 109777 277423
rect 109719 277355 109731 277389
rect 109765 277355 109777 277389
rect 109719 277321 109777 277355
rect 109719 277287 109731 277321
rect 109765 277287 109777 277321
rect 109719 277253 109777 277287
rect 109719 277219 109731 277253
rect 109765 277219 109777 277253
rect 109719 277185 109777 277219
rect 109719 277151 109731 277185
rect 109765 277151 109777 277185
rect 109719 277117 109777 277151
rect 109719 277083 109731 277117
rect 109765 277083 109777 277117
rect 109719 277049 109777 277083
rect 109719 277015 109731 277049
rect 109765 277015 109777 277049
rect 109719 276981 109777 277015
rect 109719 276947 109731 276981
rect 109765 276947 109777 276981
rect 109719 276913 109777 276947
rect 109719 276879 109731 276913
rect 109765 276879 109777 276913
rect 109719 276845 109777 276879
rect 109719 276811 109731 276845
rect 109765 276811 109777 276845
rect 109719 276777 109777 276811
rect 109719 276743 109731 276777
rect 109765 276743 109777 276777
rect 109719 276717 109777 276743
rect 110063 277729 110121 277755
rect 110063 277695 110075 277729
rect 110109 277695 110121 277729
rect 110063 277661 110121 277695
rect 110063 277627 110075 277661
rect 110109 277627 110121 277661
rect 110063 277593 110121 277627
rect 110063 277559 110075 277593
rect 110109 277559 110121 277593
rect 110063 277525 110121 277559
rect 110063 277491 110075 277525
rect 110109 277491 110121 277525
rect 110063 277457 110121 277491
rect 110063 277423 110075 277457
rect 110109 277423 110121 277457
rect 110063 277389 110121 277423
rect 110063 277355 110075 277389
rect 110109 277355 110121 277389
rect 110063 277321 110121 277355
rect 110063 277287 110075 277321
rect 110109 277287 110121 277321
rect 110063 277253 110121 277287
rect 110063 277219 110075 277253
rect 110109 277219 110121 277253
rect 110063 277185 110121 277219
rect 110063 277151 110075 277185
rect 110109 277151 110121 277185
rect 110063 277117 110121 277151
rect 110063 277083 110075 277117
rect 110109 277083 110121 277117
rect 110063 277049 110121 277083
rect 110063 277015 110075 277049
rect 110109 277015 110121 277049
rect 110063 276981 110121 277015
rect 110063 276947 110075 276981
rect 110109 276947 110121 276981
rect 110063 276913 110121 276947
rect 110063 276879 110075 276913
rect 110109 276879 110121 276913
rect 110063 276845 110121 276879
rect 110063 276811 110075 276845
rect 110109 276811 110121 276845
rect 110063 276777 110121 276811
rect 110063 276743 110075 276777
rect 110109 276743 110121 276777
rect 110063 276717 110121 276743
rect 107401 272060 107459 272079
rect 107401 272026 107413 272060
rect 107447 272026 107459 272060
rect 107401 271992 107459 272026
rect 106923 271940 106981 271971
rect 106923 271906 106935 271940
rect 106969 271906 106981 271940
rect 106923 271872 106981 271906
rect 106923 271838 106935 271872
rect 106969 271838 106981 271872
rect 106923 271807 106981 271838
rect 107191 271940 107249 271971
rect 107191 271906 107203 271940
rect 107237 271906 107249 271940
rect 107191 271872 107249 271906
rect 107191 271838 107203 271872
rect 107237 271838 107249 271872
rect 107191 271807 107249 271838
rect 107401 271958 107413 271992
rect 107447 271958 107459 271992
rect 107401 271924 107459 271958
rect 107401 271890 107413 271924
rect 107447 271890 107459 271924
rect 107401 271856 107459 271890
rect 107401 271822 107413 271856
rect 107447 271822 107459 271856
rect 107401 271788 107459 271822
rect 107401 271754 107413 271788
rect 107447 271754 107459 271788
rect 107401 271735 107459 271754
rect 108079 272060 108137 272079
rect 108079 272026 108091 272060
rect 108125 272026 108137 272060
rect 108079 271992 108137 272026
rect 108079 271958 108091 271992
rect 108125 271958 108137 271992
rect 108079 271924 108137 271958
rect 108079 271890 108091 271924
rect 108125 271890 108137 271924
rect 108079 271856 108137 271890
rect 108079 271822 108091 271856
rect 108125 271822 108137 271856
rect 108079 271788 108137 271822
rect 108079 271754 108091 271788
rect 108125 271754 108137 271788
rect 108079 271735 108137 271754
rect 107173 271535 108373 271547
rect 107173 271501 107212 271535
rect 107246 271501 107280 271535
rect 107314 271501 107348 271535
rect 107382 271501 107416 271535
rect 107450 271501 107484 271535
rect 107518 271501 107552 271535
rect 107586 271501 107620 271535
rect 107654 271501 107688 271535
rect 107722 271501 107756 271535
rect 107790 271501 107824 271535
rect 107858 271501 107892 271535
rect 107926 271501 107960 271535
rect 107994 271501 108028 271535
rect 108062 271501 108096 271535
rect 108130 271501 108164 271535
rect 108198 271501 108232 271535
rect 108266 271501 108300 271535
rect 108334 271501 108373 271535
rect 107173 271489 108373 271501
rect 107173 271299 108373 271311
rect 107173 271265 107212 271299
rect 107246 271265 107280 271299
rect 107314 271265 107348 271299
rect 107382 271265 107416 271299
rect 107450 271265 107484 271299
rect 107518 271265 107552 271299
rect 107586 271265 107620 271299
rect 107654 271265 107688 271299
rect 107722 271265 107756 271299
rect 107790 271265 107824 271299
rect 107858 271265 107892 271299
rect 107926 271265 107960 271299
rect 107994 271265 108028 271299
rect 108062 271265 108096 271299
rect 108130 271265 108164 271299
rect 108198 271265 108232 271299
rect 108266 271265 108300 271299
rect 108334 271265 108373 271299
rect 107173 271253 108373 271265
rect 107173 271165 108373 271177
rect 107173 271131 107212 271165
rect 107246 271131 107280 271165
rect 107314 271131 107348 271165
rect 107382 271131 107416 271165
rect 107450 271131 107484 271165
rect 107518 271131 107552 271165
rect 107586 271131 107620 271165
rect 107654 271131 107688 271165
rect 107722 271131 107756 271165
rect 107790 271131 107824 271165
rect 107858 271131 107892 271165
rect 107926 271131 107960 271165
rect 107994 271131 108028 271165
rect 108062 271131 108096 271165
rect 108130 271131 108164 271165
rect 108198 271131 108232 271165
rect 108266 271131 108300 271165
rect 108334 271131 108373 271165
rect 107173 271119 108373 271131
rect 107173 270929 108373 270941
rect 107173 270895 107212 270929
rect 107246 270895 107280 270929
rect 107314 270895 107348 270929
rect 107382 270895 107416 270929
rect 107450 270895 107484 270929
rect 107518 270895 107552 270929
rect 107586 270895 107620 270929
rect 107654 270895 107688 270929
rect 107722 270895 107756 270929
rect 107790 270895 107824 270929
rect 107858 270895 107892 270929
rect 107926 270895 107960 270929
rect 107994 270895 108028 270929
rect 108062 270895 108096 270929
rect 108130 270895 108164 270929
rect 108198 270895 108232 270929
rect 108266 270895 108300 270929
rect 108334 270895 108373 270929
rect 107173 270883 108373 270895
rect 111524 280866 112624 280878
rect 111524 280832 111547 280866
rect 111581 280832 111615 280866
rect 111649 280832 111683 280866
rect 111717 280832 111751 280866
rect 111785 280832 111819 280866
rect 111853 280832 111887 280866
rect 111921 280832 111955 280866
rect 111989 280832 112023 280866
rect 112057 280832 112091 280866
rect 112125 280832 112159 280866
rect 112193 280832 112227 280866
rect 112261 280832 112295 280866
rect 112329 280832 112363 280866
rect 112397 280832 112431 280866
rect 112465 280832 112499 280866
rect 112533 280832 112567 280866
rect 112601 280832 112624 280866
rect 111524 280820 112624 280832
rect 112970 280874 114070 280886
rect 112970 280840 112993 280874
rect 113027 280840 113061 280874
rect 113095 280840 113129 280874
rect 113163 280840 113197 280874
rect 113231 280840 113265 280874
rect 113299 280840 113333 280874
rect 113367 280840 113401 280874
rect 113435 280840 113469 280874
rect 113503 280840 113537 280874
rect 113571 280840 113605 280874
rect 113639 280840 113673 280874
rect 113707 280840 113741 280874
rect 113775 280840 113809 280874
rect 113843 280840 113877 280874
rect 113911 280840 113945 280874
rect 113979 280840 114013 280874
rect 114047 280840 114070 280874
rect 112970 280828 114070 280840
rect 111524 280648 112624 280660
rect 111524 280614 111547 280648
rect 111581 280614 111615 280648
rect 111649 280614 111683 280648
rect 111717 280614 111751 280648
rect 111785 280614 111819 280648
rect 111853 280614 111887 280648
rect 111921 280614 111955 280648
rect 111989 280614 112023 280648
rect 112057 280614 112091 280648
rect 112125 280614 112159 280648
rect 112193 280614 112227 280648
rect 112261 280614 112295 280648
rect 112329 280614 112363 280648
rect 112397 280614 112431 280648
rect 112465 280614 112499 280648
rect 112533 280614 112567 280648
rect 112601 280614 112624 280648
rect 111524 280602 112624 280614
rect 112970 280616 114070 280628
rect 112970 280582 112993 280616
rect 113027 280582 113061 280616
rect 113095 280582 113129 280616
rect 113163 280582 113197 280616
rect 113231 280582 113265 280616
rect 113299 280582 113333 280616
rect 113367 280582 113401 280616
rect 113435 280582 113469 280616
rect 113503 280582 113537 280616
rect 113571 280582 113605 280616
rect 113639 280582 113673 280616
rect 113707 280582 113741 280616
rect 113775 280582 113809 280616
rect 113843 280582 113877 280616
rect 113911 280582 113945 280616
rect 113979 280582 114013 280616
rect 114047 280582 114070 280616
rect 112970 280570 114070 280582
rect 111524 280506 112624 280518
rect 111524 280472 111547 280506
rect 111581 280472 111615 280506
rect 111649 280472 111683 280506
rect 111717 280472 111751 280506
rect 111785 280472 111819 280506
rect 111853 280472 111887 280506
rect 111921 280472 111955 280506
rect 111989 280472 112023 280506
rect 112057 280472 112091 280506
rect 112125 280472 112159 280506
rect 112193 280472 112227 280506
rect 112261 280472 112295 280506
rect 112329 280472 112363 280506
rect 112397 280472 112431 280506
rect 112465 280472 112499 280506
rect 112533 280472 112567 280506
rect 112601 280472 112624 280506
rect 111524 280460 112624 280472
rect 112970 280450 114070 280462
rect 112970 280416 112993 280450
rect 113027 280416 113061 280450
rect 113095 280416 113129 280450
rect 113163 280416 113197 280450
rect 113231 280416 113265 280450
rect 113299 280416 113333 280450
rect 113367 280416 113401 280450
rect 113435 280416 113469 280450
rect 113503 280416 113537 280450
rect 113571 280416 113605 280450
rect 113639 280416 113673 280450
rect 113707 280416 113741 280450
rect 113775 280416 113809 280450
rect 113843 280416 113877 280450
rect 113911 280416 113945 280450
rect 113979 280416 114013 280450
rect 114047 280416 114070 280450
rect 112970 280404 114070 280416
rect 111524 280288 112624 280300
rect 111524 280254 111547 280288
rect 111581 280254 111615 280288
rect 111649 280254 111683 280288
rect 111717 280254 111751 280288
rect 111785 280254 111819 280288
rect 111853 280254 111887 280288
rect 111921 280254 111955 280288
rect 111989 280254 112023 280288
rect 112057 280254 112091 280288
rect 112125 280254 112159 280288
rect 112193 280254 112227 280288
rect 112261 280254 112295 280288
rect 112329 280254 112363 280288
rect 112397 280254 112431 280288
rect 112465 280254 112499 280288
rect 112533 280254 112567 280288
rect 112601 280254 112624 280288
rect 111524 280242 112624 280254
rect 112970 280192 114070 280204
rect 112970 280158 112993 280192
rect 113027 280158 113061 280192
rect 113095 280158 113129 280192
rect 113163 280158 113197 280192
rect 113231 280158 113265 280192
rect 113299 280158 113333 280192
rect 113367 280158 113401 280192
rect 113435 280158 113469 280192
rect 113503 280158 113537 280192
rect 113571 280158 113605 280192
rect 113639 280158 113673 280192
rect 113707 280158 113741 280192
rect 113775 280158 113809 280192
rect 113843 280158 113877 280192
rect 113911 280158 113945 280192
rect 113979 280158 114013 280192
rect 114047 280158 114070 280192
rect 111524 280146 112624 280158
rect 112970 280146 114070 280158
rect 111524 280112 111547 280146
rect 111581 280112 111615 280146
rect 111649 280112 111683 280146
rect 111717 280112 111751 280146
rect 111785 280112 111819 280146
rect 111853 280112 111887 280146
rect 111921 280112 111955 280146
rect 111989 280112 112023 280146
rect 112057 280112 112091 280146
rect 112125 280112 112159 280146
rect 112193 280112 112227 280146
rect 112261 280112 112295 280146
rect 112329 280112 112363 280146
rect 112397 280112 112431 280146
rect 112465 280112 112499 280146
rect 112533 280112 112567 280146
rect 112601 280112 112624 280146
rect 111524 280100 112624 280112
rect 113000 280048 114100 280060
rect 113000 280014 113023 280048
rect 113057 280014 113091 280048
rect 113125 280014 113159 280048
rect 113193 280014 113227 280048
rect 113261 280014 113295 280048
rect 113329 280014 113363 280048
rect 113397 280014 113431 280048
rect 113465 280014 113499 280048
rect 113533 280014 113567 280048
rect 113601 280014 113635 280048
rect 113669 280014 113703 280048
rect 113737 280014 113771 280048
rect 113805 280014 113839 280048
rect 113873 280014 113907 280048
rect 113941 280014 113975 280048
rect 114009 280014 114043 280048
rect 114077 280014 114100 280048
rect 113000 280002 114100 280014
rect 111524 279928 112624 279940
rect 111524 279894 111547 279928
rect 111581 279894 111615 279928
rect 111649 279894 111683 279928
rect 111717 279894 111751 279928
rect 111785 279894 111819 279928
rect 111853 279894 111887 279928
rect 111921 279894 111955 279928
rect 111989 279894 112023 279928
rect 112057 279894 112091 279928
rect 112125 279894 112159 279928
rect 112193 279894 112227 279928
rect 112261 279894 112295 279928
rect 112329 279894 112363 279928
rect 112397 279894 112431 279928
rect 112465 279894 112499 279928
rect 112533 279894 112567 279928
rect 112601 279894 112624 279928
rect 111524 279882 112624 279894
rect 113000 279910 114100 279922
rect 113000 279876 113023 279910
rect 113057 279876 113091 279910
rect 113125 279876 113159 279910
rect 113193 279876 113227 279910
rect 113261 279876 113295 279910
rect 113329 279876 113363 279910
rect 113397 279876 113431 279910
rect 113465 279876 113499 279910
rect 113533 279876 113567 279910
rect 113601 279876 113635 279910
rect 113669 279876 113703 279910
rect 113737 279876 113771 279910
rect 113805 279876 113839 279910
rect 113873 279876 113907 279910
rect 113941 279876 113975 279910
rect 114009 279876 114043 279910
rect 114077 279876 114100 279910
rect 113000 279864 114100 279876
rect 111524 279786 112624 279798
rect 111524 279752 111547 279786
rect 111581 279752 111615 279786
rect 111649 279752 111683 279786
rect 111717 279752 111751 279786
rect 111785 279752 111819 279786
rect 111853 279752 111887 279786
rect 111921 279752 111955 279786
rect 111989 279752 112023 279786
rect 112057 279752 112091 279786
rect 112125 279752 112159 279786
rect 112193 279752 112227 279786
rect 112261 279752 112295 279786
rect 112329 279752 112363 279786
rect 112397 279752 112431 279786
rect 112465 279752 112499 279786
rect 112533 279752 112567 279786
rect 112601 279752 112624 279786
rect 111524 279740 112624 279752
rect 113000 279750 114100 279762
rect 113000 279716 113023 279750
rect 113057 279716 113091 279750
rect 113125 279716 113159 279750
rect 113193 279716 113227 279750
rect 113261 279716 113295 279750
rect 113329 279716 113363 279750
rect 113397 279716 113431 279750
rect 113465 279716 113499 279750
rect 113533 279716 113567 279750
rect 113601 279716 113635 279750
rect 113669 279716 113703 279750
rect 113737 279716 113771 279750
rect 113805 279716 113839 279750
rect 113873 279716 113907 279750
rect 113941 279716 113975 279750
rect 114009 279716 114043 279750
rect 114077 279716 114100 279750
rect 113000 279704 114100 279716
rect 113000 279612 114100 279624
rect 111524 279568 112624 279580
rect 111524 279534 111547 279568
rect 111581 279534 111615 279568
rect 111649 279534 111683 279568
rect 111717 279534 111751 279568
rect 111785 279534 111819 279568
rect 111853 279534 111887 279568
rect 111921 279534 111955 279568
rect 111989 279534 112023 279568
rect 112057 279534 112091 279568
rect 112125 279534 112159 279568
rect 112193 279534 112227 279568
rect 112261 279534 112295 279568
rect 112329 279534 112363 279568
rect 112397 279534 112431 279568
rect 112465 279534 112499 279568
rect 112533 279534 112567 279568
rect 112601 279534 112624 279568
rect 113000 279578 113023 279612
rect 113057 279578 113091 279612
rect 113125 279578 113159 279612
rect 113193 279578 113227 279612
rect 113261 279578 113295 279612
rect 113329 279578 113363 279612
rect 113397 279578 113431 279612
rect 113465 279578 113499 279612
rect 113533 279578 113567 279612
rect 113601 279578 113635 279612
rect 113669 279578 113703 279612
rect 113737 279578 113771 279612
rect 113805 279578 113839 279612
rect 113873 279578 113907 279612
rect 113941 279578 113975 279612
rect 114009 279578 114043 279612
rect 114077 279578 114100 279612
rect 113000 279566 114100 279578
rect 111524 279522 112624 279534
rect 116135 280874 117235 280886
rect 116135 280840 116158 280874
rect 116192 280840 116226 280874
rect 116260 280840 116294 280874
rect 116328 280840 116362 280874
rect 116396 280840 116430 280874
rect 116464 280840 116498 280874
rect 116532 280840 116566 280874
rect 116600 280840 116634 280874
rect 116668 280840 116702 280874
rect 116736 280840 116770 280874
rect 116804 280840 116838 280874
rect 116872 280840 116906 280874
rect 116940 280840 116974 280874
rect 117008 280840 117042 280874
rect 117076 280840 117110 280874
rect 117144 280840 117178 280874
rect 117212 280840 117235 280874
rect 116135 280828 117235 280840
rect 117581 280866 118681 280878
rect 117581 280832 117604 280866
rect 117638 280832 117672 280866
rect 117706 280832 117740 280866
rect 117774 280832 117808 280866
rect 117842 280832 117876 280866
rect 117910 280832 117944 280866
rect 117978 280832 118012 280866
rect 118046 280832 118080 280866
rect 118114 280832 118148 280866
rect 118182 280832 118216 280866
rect 118250 280832 118284 280866
rect 118318 280832 118352 280866
rect 118386 280832 118420 280866
rect 118454 280832 118488 280866
rect 118522 280832 118556 280866
rect 118590 280832 118624 280866
rect 118658 280832 118681 280866
rect 117581 280820 118681 280832
rect 117581 280648 118681 280660
rect 116135 280616 117235 280628
rect 116135 280582 116158 280616
rect 116192 280582 116226 280616
rect 116260 280582 116294 280616
rect 116328 280582 116362 280616
rect 116396 280582 116430 280616
rect 116464 280582 116498 280616
rect 116532 280582 116566 280616
rect 116600 280582 116634 280616
rect 116668 280582 116702 280616
rect 116736 280582 116770 280616
rect 116804 280582 116838 280616
rect 116872 280582 116906 280616
rect 116940 280582 116974 280616
rect 117008 280582 117042 280616
rect 117076 280582 117110 280616
rect 117144 280582 117178 280616
rect 117212 280582 117235 280616
rect 117581 280614 117604 280648
rect 117638 280614 117672 280648
rect 117706 280614 117740 280648
rect 117774 280614 117808 280648
rect 117842 280614 117876 280648
rect 117910 280614 117944 280648
rect 117978 280614 118012 280648
rect 118046 280614 118080 280648
rect 118114 280614 118148 280648
rect 118182 280614 118216 280648
rect 118250 280614 118284 280648
rect 118318 280614 118352 280648
rect 118386 280614 118420 280648
rect 118454 280614 118488 280648
rect 118522 280614 118556 280648
rect 118590 280614 118624 280648
rect 118658 280614 118681 280648
rect 117581 280602 118681 280614
rect 116135 280570 117235 280582
rect 117581 280506 118681 280518
rect 117581 280472 117604 280506
rect 117638 280472 117672 280506
rect 117706 280472 117740 280506
rect 117774 280472 117808 280506
rect 117842 280472 117876 280506
rect 117910 280472 117944 280506
rect 117978 280472 118012 280506
rect 118046 280472 118080 280506
rect 118114 280472 118148 280506
rect 118182 280472 118216 280506
rect 118250 280472 118284 280506
rect 118318 280472 118352 280506
rect 118386 280472 118420 280506
rect 118454 280472 118488 280506
rect 118522 280472 118556 280506
rect 118590 280472 118624 280506
rect 118658 280472 118681 280506
rect 116135 280450 117235 280462
rect 117581 280460 118681 280472
rect 116135 280416 116158 280450
rect 116192 280416 116226 280450
rect 116260 280416 116294 280450
rect 116328 280416 116362 280450
rect 116396 280416 116430 280450
rect 116464 280416 116498 280450
rect 116532 280416 116566 280450
rect 116600 280416 116634 280450
rect 116668 280416 116702 280450
rect 116736 280416 116770 280450
rect 116804 280416 116838 280450
rect 116872 280416 116906 280450
rect 116940 280416 116974 280450
rect 117008 280416 117042 280450
rect 117076 280416 117110 280450
rect 117144 280416 117178 280450
rect 117212 280416 117235 280450
rect 116135 280404 117235 280416
rect 117581 280288 118681 280300
rect 117581 280254 117604 280288
rect 117638 280254 117672 280288
rect 117706 280254 117740 280288
rect 117774 280254 117808 280288
rect 117842 280254 117876 280288
rect 117910 280254 117944 280288
rect 117978 280254 118012 280288
rect 118046 280254 118080 280288
rect 118114 280254 118148 280288
rect 118182 280254 118216 280288
rect 118250 280254 118284 280288
rect 118318 280254 118352 280288
rect 118386 280254 118420 280288
rect 118454 280254 118488 280288
rect 118522 280254 118556 280288
rect 118590 280254 118624 280288
rect 118658 280254 118681 280288
rect 117581 280242 118681 280254
rect 116135 280192 117235 280204
rect 116135 280158 116158 280192
rect 116192 280158 116226 280192
rect 116260 280158 116294 280192
rect 116328 280158 116362 280192
rect 116396 280158 116430 280192
rect 116464 280158 116498 280192
rect 116532 280158 116566 280192
rect 116600 280158 116634 280192
rect 116668 280158 116702 280192
rect 116736 280158 116770 280192
rect 116804 280158 116838 280192
rect 116872 280158 116906 280192
rect 116940 280158 116974 280192
rect 117008 280158 117042 280192
rect 117076 280158 117110 280192
rect 117144 280158 117178 280192
rect 117212 280158 117235 280192
rect 116135 280146 117235 280158
rect 117581 280146 118681 280158
rect 117581 280112 117604 280146
rect 117638 280112 117672 280146
rect 117706 280112 117740 280146
rect 117774 280112 117808 280146
rect 117842 280112 117876 280146
rect 117910 280112 117944 280146
rect 117978 280112 118012 280146
rect 118046 280112 118080 280146
rect 118114 280112 118148 280146
rect 118182 280112 118216 280146
rect 118250 280112 118284 280146
rect 118318 280112 118352 280146
rect 118386 280112 118420 280146
rect 118454 280112 118488 280146
rect 118522 280112 118556 280146
rect 118590 280112 118624 280146
rect 118658 280112 118681 280146
rect 117581 280100 118681 280112
rect 116105 280048 117205 280060
rect 116105 280014 116128 280048
rect 116162 280014 116196 280048
rect 116230 280014 116264 280048
rect 116298 280014 116332 280048
rect 116366 280014 116400 280048
rect 116434 280014 116468 280048
rect 116502 280014 116536 280048
rect 116570 280014 116604 280048
rect 116638 280014 116672 280048
rect 116706 280014 116740 280048
rect 116774 280014 116808 280048
rect 116842 280014 116876 280048
rect 116910 280014 116944 280048
rect 116978 280014 117012 280048
rect 117046 280014 117080 280048
rect 117114 280014 117148 280048
rect 117182 280014 117205 280048
rect 116105 280002 117205 280014
rect 117581 279928 118681 279940
rect 116105 279910 117205 279922
rect 116105 279876 116128 279910
rect 116162 279876 116196 279910
rect 116230 279876 116264 279910
rect 116298 279876 116332 279910
rect 116366 279876 116400 279910
rect 116434 279876 116468 279910
rect 116502 279876 116536 279910
rect 116570 279876 116604 279910
rect 116638 279876 116672 279910
rect 116706 279876 116740 279910
rect 116774 279876 116808 279910
rect 116842 279876 116876 279910
rect 116910 279876 116944 279910
rect 116978 279876 117012 279910
rect 117046 279876 117080 279910
rect 117114 279876 117148 279910
rect 117182 279876 117205 279910
rect 117581 279894 117604 279928
rect 117638 279894 117672 279928
rect 117706 279894 117740 279928
rect 117774 279894 117808 279928
rect 117842 279894 117876 279928
rect 117910 279894 117944 279928
rect 117978 279894 118012 279928
rect 118046 279894 118080 279928
rect 118114 279894 118148 279928
rect 118182 279894 118216 279928
rect 118250 279894 118284 279928
rect 118318 279894 118352 279928
rect 118386 279894 118420 279928
rect 118454 279894 118488 279928
rect 118522 279894 118556 279928
rect 118590 279894 118624 279928
rect 118658 279894 118681 279928
rect 117581 279882 118681 279894
rect 116105 279864 117205 279876
rect 117581 279786 118681 279798
rect 116105 279750 117205 279762
rect 116105 279716 116128 279750
rect 116162 279716 116196 279750
rect 116230 279716 116264 279750
rect 116298 279716 116332 279750
rect 116366 279716 116400 279750
rect 116434 279716 116468 279750
rect 116502 279716 116536 279750
rect 116570 279716 116604 279750
rect 116638 279716 116672 279750
rect 116706 279716 116740 279750
rect 116774 279716 116808 279750
rect 116842 279716 116876 279750
rect 116910 279716 116944 279750
rect 116978 279716 117012 279750
rect 117046 279716 117080 279750
rect 117114 279716 117148 279750
rect 117182 279716 117205 279750
rect 117581 279752 117604 279786
rect 117638 279752 117672 279786
rect 117706 279752 117740 279786
rect 117774 279752 117808 279786
rect 117842 279752 117876 279786
rect 117910 279752 117944 279786
rect 117978 279752 118012 279786
rect 118046 279752 118080 279786
rect 118114 279752 118148 279786
rect 118182 279752 118216 279786
rect 118250 279752 118284 279786
rect 118318 279752 118352 279786
rect 118386 279752 118420 279786
rect 118454 279752 118488 279786
rect 118522 279752 118556 279786
rect 118590 279752 118624 279786
rect 118658 279752 118681 279786
rect 117581 279740 118681 279752
rect 116105 279704 117205 279716
rect 116105 279612 117205 279624
rect 116105 279578 116128 279612
rect 116162 279578 116196 279612
rect 116230 279578 116264 279612
rect 116298 279578 116332 279612
rect 116366 279578 116400 279612
rect 116434 279578 116468 279612
rect 116502 279578 116536 279612
rect 116570 279578 116604 279612
rect 116638 279578 116672 279612
rect 116706 279578 116740 279612
rect 116774 279578 116808 279612
rect 116842 279578 116876 279612
rect 116910 279578 116944 279612
rect 116978 279578 117012 279612
rect 117046 279578 117080 279612
rect 117114 279578 117148 279612
rect 117182 279578 117205 279612
rect 116105 279566 117205 279578
rect 117581 279568 118681 279580
rect 117581 279534 117604 279568
rect 117638 279534 117672 279568
rect 117706 279534 117740 279568
rect 117774 279534 117808 279568
rect 117842 279534 117876 279568
rect 117910 279534 117944 279568
rect 117978 279534 118012 279568
rect 118046 279534 118080 279568
rect 118114 279534 118148 279568
rect 118182 279534 118216 279568
rect 118250 279534 118284 279568
rect 118318 279534 118352 279568
rect 118386 279534 118420 279568
rect 118454 279534 118488 279568
rect 118522 279534 118556 279568
rect 118590 279534 118624 279568
rect 118658 279534 118681 279568
rect 117581 279522 118681 279534
rect 111524 279200 112624 279212
rect 111524 279166 111547 279200
rect 111581 279166 111615 279200
rect 111649 279166 111683 279200
rect 111717 279166 111751 279200
rect 111785 279166 111819 279200
rect 111853 279166 111887 279200
rect 111921 279166 111955 279200
rect 111989 279166 112023 279200
rect 112057 279166 112091 279200
rect 112125 279166 112159 279200
rect 112193 279166 112227 279200
rect 112261 279166 112295 279200
rect 112329 279166 112363 279200
rect 112397 279166 112431 279200
rect 112465 279166 112499 279200
rect 112533 279166 112567 279200
rect 112601 279166 112624 279200
rect 111524 279154 112624 279166
rect 112970 279208 114070 279220
rect 112970 279174 112993 279208
rect 113027 279174 113061 279208
rect 113095 279174 113129 279208
rect 113163 279174 113197 279208
rect 113231 279174 113265 279208
rect 113299 279174 113333 279208
rect 113367 279174 113401 279208
rect 113435 279174 113469 279208
rect 113503 279174 113537 279208
rect 113571 279174 113605 279208
rect 113639 279174 113673 279208
rect 113707 279174 113741 279208
rect 113775 279174 113809 279208
rect 113843 279174 113877 279208
rect 113911 279174 113945 279208
rect 113979 279174 114013 279208
rect 114047 279174 114070 279208
rect 112970 279162 114070 279174
rect 111524 278982 112624 278994
rect 111524 278948 111547 278982
rect 111581 278948 111615 278982
rect 111649 278948 111683 278982
rect 111717 278948 111751 278982
rect 111785 278948 111819 278982
rect 111853 278948 111887 278982
rect 111921 278948 111955 278982
rect 111989 278948 112023 278982
rect 112057 278948 112091 278982
rect 112125 278948 112159 278982
rect 112193 278948 112227 278982
rect 112261 278948 112295 278982
rect 112329 278948 112363 278982
rect 112397 278948 112431 278982
rect 112465 278948 112499 278982
rect 112533 278948 112567 278982
rect 112601 278948 112624 278982
rect 111524 278936 112624 278948
rect 112970 278950 114070 278962
rect 112970 278916 112993 278950
rect 113027 278916 113061 278950
rect 113095 278916 113129 278950
rect 113163 278916 113197 278950
rect 113231 278916 113265 278950
rect 113299 278916 113333 278950
rect 113367 278916 113401 278950
rect 113435 278916 113469 278950
rect 113503 278916 113537 278950
rect 113571 278916 113605 278950
rect 113639 278916 113673 278950
rect 113707 278916 113741 278950
rect 113775 278916 113809 278950
rect 113843 278916 113877 278950
rect 113911 278916 113945 278950
rect 113979 278916 114013 278950
rect 114047 278916 114070 278950
rect 112970 278904 114070 278916
rect 111524 278840 112624 278852
rect 111524 278806 111547 278840
rect 111581 278806 111615 278840
rect 111649 278806 111683 278840
rect 111717 278806 111751 278840
rect 111785 278806 111819 278840
rect 111853 278806 111887 278840
rect 111921 278806 111955 278840
rect 111989 278806 112023 278840
rect 112057 278806 112091 278840
rect 112125 278806 112159 278840
rect 112193 278806 112227 278840
rect 112261 278806 112295 278840
rect 112329 278806 112363 278840
rect 112397 278806 112431 278840
rect 112465 278806 112499 278840
rect 112533 278806 112567 278840
rect 112601 278806 112624 278840
rect 111524 278794 112624 278806
rect 112970 278784 114070 278796
rect 112970 278750 112993 278784
rect 113027 278750 113061 278784
rect 113095 278750 113129 278784
rect 113163 278750 113197 278784
rect 113231 278750 113265 278784
rect 113299 278750 113333 278784
rect 113367 278750 113401 278784
rect 113435 278750 113469 278784
rect 113503 278750 113537 278784
rect 113571 278750 113605 278784
rect 113639 278750 113673 278784
rect 113707 278750 113741 278784
rect 113775 278750 113809 278784
rect 113843 278750 113877 278784
rect 113911 278750 113945 278784
rect 113979 278750 114013 278784
rect 114047 278750 114070 278784
rect 112970 278738 114070 278750
rect 111524 278622 112624 278634
rect 111524 278588 111547 278622
rect 111581 278588 111615 278622
rect 111649 278588 111683 278622
rect 111717 278588 111751 278622
rect 111785 278588 111819 278622
rect 111853 278588 111887 278622
rect 111921 278588 111955 278622
rect 111989 278588 112023 278622
rect 112057 278588 112091 278622
rect 112125 278588 112159 278622
rect 112193 278588 112227 278622
rect 112261 278588 112295 278622
rect 112329 278588 112363 278622
rect 112397 278588 112431 278622
rect 112465 278588 112499 278622
rect 112533 278588 112567 278622
rect 112601 278588 112624 278622
rect 111524 278576 112624 278588
rect 112970 278526 114070 278538
rect 112970 278492 112993 278526
rect 113027 278492 113061 278526
rect 113095 278492 113129 278526
rect 113163 278492 113197 278526
rect 113231 278492 113265 278526
rect 113299 278492 113333 278526
rect 113367 278492 113401 278526
rect 113435 278492 113469 278526
rect 113503 278492 113537 278526
rect 113571 278492 113605 278526
rect 113639 278492 113673 278526
rect 113707 278492 113741 278526
rect 113775 278492 113809 278526
rect 113843 278492 113877 278526
rect 113911 278492 113945 278526
rect 113979 278492 114013 278526
rect 114047 278492 114070 278526
rect 111524 278480 112624 278492
rect 112970 278480 114070 278492
rect 111524 278446 111547 278480
rect 111581 278446 111615 278480
rect 111649 278446 111683 278480
rect 111717 278446 111751 278480
rect 111785 278446 111819 278480
rect 111853 278446 111887 278480
rect 111921 278446 111955 278480
rect 111989 278446 112023 278480
rect 112057 278446 112091 278480
rect 112125 278446 112159 278480
rect 112193 278446 112227 278480
rect 112261 278446 112295 278480
rect 112329 278446 112363 278480
rect 112397 278446 112431 278480
rect 112465 278446 112499 278480
rect 112533 278446 112567 278480
rect 112601 278446 112624 278480
rect 111524 278434 112624 278446
rect 113000 278382 114100 278394
rect 113000 278348 113023 278382
rect 113057 278348 113091 278382
rect 113125 278348 113159 278382
rect 113193 278348 113227 278382
rect 113261 278348 113295 278382
rect 113329 278348 113363 278382
rect 113397 278348 113431 278382
rect 113465 278348 113499 278382
rect 113533 278348 113567 278382
rect 113601 278348 113635 278382
rect 113669 278348 113703 278382
rect 113737 278348 113771 278382
rect 113805 278348 113839 278382
rect 113873 278348 113907 278382
rect 113941 278348 113975 278382
rect 114009 278348 114043 278382
rect 114077 278348 114100 278382
rect 113000 278336 114100 278348
rect 111524 278262 112624 278274
rect 111524 278228 111547 278262
rect 111581 278228 111615 278262
rect 111649 278228 111683 278262
rect 111717 278228 111751 278262
rect 111785 278228 111819 278262
rect 111853 278228 111887 278262
rect 111921 278228 111955 278262
rect 111989 278228 112023 278262
rect 112057 278228 112091 278262
rect 112125 278228 112159 278262
rect 112193 278228 112227 278262
rect 112261 278228 112295 278262
rect 112329 278228 112363 278262
rect 112397 278228 112431 278262
rect 112465 278228 112499 278262
rect 112533 278228 112567 278262
rect 112601 278228 112624 278262
rect 111524 278216 112624 278228
rect 113000 278244 114100 278256
rect 113000 278210 113023 278244
rect 113057 278210 113091 278244
rect 113125 278210 113159 278244
rect 113193 278210 113227 278244
rect 113261 278210 113295 278244
rect 113329 278210 113363 278244
rect 113397 278210 113431 278244
rect 113465 278210 113499 278244
rect 113533 278210 113567 278244
rect 113601 278210 113635 278244
rect 113669 278210 113703 278244
rect 113737 278210 113771 278244
rect 113805 278210 113839 278244
rect 113873 278210 113907 278244
rect 113941 278210 113975 278244
rect 114009 278210 114043 278244
rect 114077 278210 114100 278244
rect 113000 278198 114100 278210
rect 111524 278120 112624 278132
rect 111524 278086 111547 278120
rect 111581 278086 111615 278120
rect 111649 278086 111683 278120
rect 111717 278086 111751 278120
rect 111785 278086 111819 278120
rect 111853 278086 111887 278120
rect 111921 278086 111955 278120
rect 111989 278086 112023 278120
rect 112057 278086 112091 278120
rect 112125 278086 112159 278120
rect 112193 278086 112227 278120
rect 112261 278086 112295 278120
rect 112329 278086 112363 278120
rect 112397 278086 112431 278120
rect 112465 278086 112499 278120
rect 112533 278086 112567 278120
rect 112601 278086 112624 278120
rect 111524 278074 112624 278086
rect 113000 278084 114100 278096
rect 113000 278050 113023 278084
rect 113057 278050 113091 278084
rect 113125 278050 113159 278084
rect 113193 278050 113227 278084
rect 113261 278050 113295 278084
rect 113329 278050 113363 278084
rect 113397 278050 113431 278084
rect 113465 278050 113499 278084
rect 113533 278050 113567 278084
rect 113601 278050 113635 278084
rect 113669 278050 113703 278084
rect 113737 278050 113771 278084
rect 113805 278050 113839 278084
rect 113873 278050 113907 278084
rect 113941 278050 113975 278084
rect 114009 278050 114043 278084
rect 114077 278050 114100 278084
rect 113000 278038 114100 278050
rect 113000 277946 114100 277958
rect 111524 277902 112624 277914
rect 111524 277868 111547 277902
rect 111581 277868 111615 277902
rect 111649 277868 111683 277902
rect 111717 277868 111751 277902
rect 111785 277868 111819 277902
rect 111853 277868 111887 277902
rect 111921 277868 111955 277902
rect 111989 277868 112023 277902
rect 112057 277868 112091 277902
rect 112125 277868 112159 277902
rect 112193 277868 112227 277902
rect 112261 277868 112295 277902
rect 112329 277868 112363 277902
rect 112397 277868 112431 277902
rect 112465 277868 112499 277902
rect 112533 277868 112567 277902
rect 112601 277868 112624 277902
rect 113000 277912 113023 277946
rect 113057 277912 113091 277946
rect 113125 277912 113159 277946
rect 113193 277912 113227 277946
rect 113261 277912 113295 277946
rect 113329 277912 113363 277946
rect 113397 277912 113431 277946
rect 113465 277912 113499 277946
rect 113533 277912 113567 277946
rect 113601 277912 113635 277946
rect 113669 277912 113703 277946
rect 113737 277912 113771 277946
rect 113805 277912 113839 277946
rect 113873 277912 113907 277946
rect 113941 277912 113975 277946
rect 114009 277912 114043 277946
rect 114077 277912 114100 277946
rect 113000 277900 114100 277912
rect 111524 277856 112624 277868
rect 116135 279208 117235 279220
rect 116135 279174 116158 279208
rect 116192 279174 116226 279208
rect 116260 279174 116294 279208
rect 116328 279174 116362 279208
rect 116396 279174 116430 279208
rect 116464 279174 116498 279208
rect 116532 279174 116566 279208
rect 116600 279174 116634 279208
rect 116668 279174 116702 279208
rect 116736 279174 116770 279208
rect 116804 279174 116838 279208
rect 116872 279174 116906 279208
rect 116940 279174 116974 279208
rect 117008 279174 117042 279208
rect 117076 279174 117110 279208
rect 117144 279174 117178 279208
rect 117212 279174 117235 279208
rect 116135 279162 117235 279174
rect 117581 279200 118681 279212
rect 117581 279166 117604 279200
rect 117638 279166 117672 279200
rect 117706 279166 117740 279200
rect 117774 279166 117808 279200
rect 117842 279166 117876 279200
rect 117910 279166 117944 279200
rect 117978 279166 118012 279200
rect 118046 279166 118080 279200
rect 118114 279166 118148 279200
rect 118182 279166 118216 279200
rect 118250 279166 118284 279200
rect 118318 279166 118352 279200
rect 118386 279166 118420 279200
rect 118454 279166 118488 279200
rect 118522 279166 118556 279200
rect 118590 279166 118624 279200
rect 118658 279166 118681 279200
rect 117581 279154 118681 279166
rect 117581 278982 118681 278994
rect 116135 278950 117235 278962
rect 116135 278916 116158 278950
rect 116192 278916 116226 278950
rect 116260 278916 116294 278950
rect 116328 278916 116362 278950
rect 116396 278916 116430 278950
rect 116464 278916 116498 278950
rect 116532 278916 116566 278950
rect 116600 278916 116634 278950
rect 116668 278916 116702 278950
rect 116736 278916 116770 278950
rect 116804 278916 116838 278950
rect 116872 278916 116906 278950
rect 116940 278916 116974 278950
rect 117008 278916 117042 278950
rect 117076 278916 117110 278950
rect 117144 278916 117178 278950
rect 117212 278916 117235 278950
rect 117581 278948 117604 278982
rect 117638 278948 117672 278982
rect 117706 278948 117740 278982
rect 117774 278948 117808 278982
rect 117842 278948 117876 278982
rect 117910 278948 117944 278982
rect 117978 278948 118012 278982
rect 118046 278948 118080 278982
rect 118114 278948 118148 278982
rect 118182 278948 118216 278982
rect 118250 278948 118284 278982
rect 118318 278948 118352 278982
rect 118386 278948 118420 278982
rect 118454 278948 118488 278982
rect 118522 278948 118556 278982
rect 118590 278948 118624 278982
rect 118658 278948 118681 278982
rect 117581 278936 118681 278948
rect 116135 278904 117235 278916
rect 117581 278840 118681 278852
rect 117581 278806 117604 278840
rect 117638 278806 117672 278840
rect 117706 278806 117740 278840
rect 117774 278806 117808 278840
rect 117842 278806 117876 278840
rect 117910 278806 117944 278840
rect 117978 278806 118012 278840
rect 118046 278806 118080 278840
rect 118114 278806 118148 278840
rect 118182 278806 118216 278840
rect 118250 278806 118284 278840
rect 118318 278806 118352 278840
rect 118386 278806 118420 278840
rect 118454 278806 118488 278840
rect 118522 278806 118556 278840
rect 118590 278806 118624 278840
rect 118658 278806 118681 278840
rect 116135 278784 117235 278796
rect 117581 278794 118681 278806
rect 116135 278750 116158 278784
rect 116192 278750 116226 278784
rect 116260 278750 116294 278784
rect 116328 278750 116362 278784
rect 116396 278750 116430 278784
rect 116464 278750 116498 278784
rect 116532 278750 116566 278784
rect 116600 278750 116634 278784
rect 116668 278750 116702 278784
rect 116736 278750 116770 278784
rect 116804 278750 116838 278784
rect 116872 278750 116906 278784
rect 116940 278750 116974 278784
rect 117008 278750 117042 278784
rect 117076 278750 117110 278784
rect 117144 278750 117178 278784
rect 117212 278750 117235 278784
rect 116135 278738 117235 278750
rect 117581 278622 118681 278634
rect 117581 278588 117604 278622
rect 117638 278588 117672 278622
rect 117706 278588 117740 278622
rect 117774 278588 117808 278622
rect 117842 278588 117876 278622
rect 117910 278588 117944 278622
rect 117978 278588 118012 278622
rect 118046 278588 118080 278622
rect 118114 278588 118148 278622
rect 118182 278588 118216 278622
rect 118250 278588 118284 278622
rect 118318 278588 118352 278622
rect 118386 278588 118420 278622
rect 118454 278588 118488 278622
rect 118522 278588 118556 278622
rect 118590 278588 118624 278622
rect 118658 278588 118681 278622
rect 117581 278576 118681 278588
rect 116135 278526 117235 278538
rect 116135 278492 116158 278526
rect 116192 278492 116226 278526
rect 116260 278492 116294 278526
rect 116328 278492 116362 278526
rect 116396 278492 116430 278526
rect 116464 278492 116498 278526
rect 116532 278492 116566 278526
rect 116600 278492 116634 278526
rect 116668 278492 116702 278526
rect 116736 278492 116770 278526
rect 116804 278492 116838 278526
rect 116872 278492 116906 278526
rect 116940 278492 116974 278526
rect 117008 278492 117042 278526
rect 117076 278492 117110 278526
rect 117144 278492 117178 278526
rect 117212 278492 117235 278526
rect 116135 278480 117235 278492
rect 117581 278480 118681 278492
rect 117581 278446 117604 278480
rect 117638 278446 117672 278480
rect 117706 278446 117740 278480
rect 117774 278446 117808 278480
rect 117842 278446 117876 278480
rect 117910 278446 117944 278480
rect 117978 278446 118012 278480
rect 118046 278446 118080 278480
rect 118114 278446 118148 278480
rect 118182 278446 118216 278480
rect 118250 278446 118284 278480
rect 118318 278446 118352 278480
rect 118386 278446 118420 278480
rect 118454 278446 118488 278480
rect 118522 278446 118556 278480
rect 118590 278446 118624 278480
rect 118658 278446 118681 278480
rect 117581 278434 118681 278446
rect 116105 278382 117205 278394
rect 116105 278348 116128 278382
rect 116162 278348 116196 278382
rect 116230 278348 116264 278382
rect 116298 278348 116332 278382
rect 116366 278348 116400 278382
rect 116434 278348 116468 278382
rect 116502 278348 116536 278382
rect 116570 278348 116604 278382
rect 116638 278348 116672 278382
rect 116706 278348 116740 278382
rect 116774 278348 116808 278382
rect 116842 278348 116876 278382
rect 116910 278348 116944 278382
rect 116978 278348 117012 278382
rect 117046 278348 117080 278382
rect 117114 278348 117148 278382
rect 117182 278348 117205 278382
rect 116105 278336 117205 278348
rect 117581 278262 118681 278274
rect 116105 278244 117205 278256
rect 116105 278210 116128 278244
rect 116162 278210 116196 278244
rect 116230 278210 116264 278244
rect 116298 278210 116332 278244
rect 116366 278210 116400 278244
rect 116434 278210 116468 278244
rect 116502 278210 116536 278244
rect 116570 278210 116604 278244
rect 116638 278210 116672 278244
rect 116706 278210 116740 278244
rect 116774 278210 116808 278244
rect 116842 278210 116876 278244
rect 116910 278210 116944 278244
rect 116978 278210 117012 278244
rect 117046 278210 117080 278244
rect 117114 278210 117148 278244
rect 117182 278210 117205 278244
rect 117581 278228 117604 278262
rect 117638 278228 117672 278262
rect 117706 278228 117740 278262
rect 117774 278228 117808 278262
rect 117842 278228 117876 278262
rect 117910 278228 117944 278262
rect 117978 278228 118012 278262
rect 118046 278228 118080 278262
rect 118114 278228 118148 278262
rect 118182 278228 118216 278262
rect 118250 278228 118284 278262
rect 118318 278228 118352 278262
rect 118386 278228 118420 278262
rect 118454 278228 118488 278262
rect 118522 278228 118556 278262
rect 118590 278228 118624 278262
rect 118658 278228 118681 278262
rect 117581 278216 118681 278228
rect 116105 278198 117205 278210
rect 117581 278120 118681 278132
rect 116105 278084 117205 278096
rect 116105 278050 116128 278084
rect 116162 278050 116196 278084
rect 116230 278050 116264 278084
rect 116298 278050 116332 278084
rect 116366 278050 116400 278084
rect 116434 278050 116468 278084
rect 116502 278050 116536 278084
rect 116570 278050 116604 278084
rect 116638 278050 116672 278084
rect 116706 278050 116740 278084
rect 116774 278050 116808 278084
rect 116842 278050 116876 278084
rect 116910 278050 116944 278084
rect 116978 278050 117012 278084
rect 117046 278050 117080 278084
rect 117114 278050 117148 278084
rect 117182 278050 117205 278084
rect 117581 278086 117604 278120
rect 117638 278086 117672 278120
rect 117706 278086 117740 278120
rect 117774 278086 117808 278120
rect 117842 278086 117876 278120
rect 117910 278086 117944 278120
rect 117978 278086 118012 278120
rect 118046 278086 118080 278120
rect 118114 278086 118148 278120
rect 118182 278086 118216 278120
rect 118250 278086 118284 278120
rect 118318 278086 118352 278120
rect 118386 278086 118420 278120
rect 118454 278086 118488 278120
rect 118522 278086 118556 278120
rect 118590 278086 118624 278120
rect 118658 278086 118681 278120
rect 117581 278074 118681 278086
rect 116105 278038 117205 278050
rect 116105 277946 117205 277958
rect 116105 277912 116128 277946
rect 116162 277912 116196 277946
rect 116230 277912 116264 277946
rect 116298 277912 116332 277946
rect 116366 277912 116400 277946
rect 116434 277912 116468 277946
rect 116502 277912 116536 277946
rect 116570 277912 116604 277946
rect 116638 277912 116672 277946
rect 116706 277912 116740 277946
rect 116774 277912 116808 277946
rect 116842 277912 116876 277946
rect 116910 277912 116944 277946
rect 116978 277912 117012 277946
rect 117046 277912 117080 277946
rect 117114 277912 117148 277946
rect 117182 277912 117205 277946
rect 116105 277900 117205 277912
rect 117581 277902 118681 277914
rect 117581 277868 117604 277902
rect 117638 277868 117672 277902
rect 117706 277868 117740 277902
rect 117774 277868 117808 277902
rect 117842 277868 117876 277902
rect 117910 277868 117944 277902
rect 117978 277868 118012 277902
rect 118046 277868 118080 277902
rect 118114 277868 118148 277902
rect 118182 277868 118216 277902
rect 118250 277868 118284 277902
rect 118318 277868 118352 277902
rect 118386 277868 118420 277902
rect 118454 277868 118488 277902
rect 118522 277868 118556 277902
rect 118590 277868 118624 277902
rect 118658 277868 118681 277902
rect 117581 277856 118681 277868
rect 111524 277534 112624 277546
rect 111524 277500 111547 277534
rect 111581 277500 111615 277534
rect 111649 277500 111683 277534
rect 111717 277500 111751 277534
rect 111785 277500 111819 277534
rect 111853 277500 111887 277534
rect 111921 277500 111955 277534
rect 111989 277500 112023 277534
rect 112057 277500 112091 277534
rect 112125 277500 112159 277534
rect 112193 277500 112227 277534
rect 112261 277500 112295 277534
rect 112329 277500 112363 277534
rect 112397 277500 112431 277534
rect 112465 277500 112499 277534
rect 112533 277500 112567 277534
rect 112601 277500 112624 277534
rect 111524 277488 112624 277500
rect 112970 277542 114070 277554
rect 112970 277508 112993 277542
rect 113027 277508 113061 277542
rect 113095 277508 113129 277542
rect 113163 277508 113197 277542
rect 113231 277508 113265 277542
rect 113299 277508 113333 277542
rect 113367 277508 113401 277542
rect 113435 277508 113469 277542
rect 113503 277508 113537 277542
rect 113571 277508 113605 277542
rect 113639 277508 113673 277542
rect 113707 277508 113741 277542
rect 113775 277508 113809 277542
rect 113843 277508 113877 277542
rect 113911 277508 113945 277542
rect 113979 277508 114013 277542
rect 114047 277508 114070 277542
rect 112970 277496 114070 277508
rect 111524 277316 112624 277328
rect 111524 277282 111547 277316
rect 111581 277282 111615 277316
rect 111649 277282 111683 277316
rect 111717 277282 111751 277316
rect 111785 277282 111819 277316
rect 111853 277282 111887 277316
rect 111921 277282 111955 277316
rect 111989 277282 112023 277316
rect 112057 277282 112091 277316
rect 112125 277282 112159 277316
rect 112193 277282 112227 277316
rect 112261 277282 112295 277316
rect 112329 277282 112363 277316
rect 112397 277282 112431 277316
rect 112465 277282 112499 277316
rect 112533 277282 112567 277316
rect 112601 277282 112624 277316
rect 111524 277270 112624 277282
rect 112970 277284 114070 277296
rect 112970 277250 112993 277284
rect 113027 277250 113061 277284
rect 113095 277250 113129 277284
rect 113163 277250 113197 277284
rect 113231 277250 113265 277284
rect 113299 277250 113333 277284
rect 113367 277250 113401 277284
rect 113435 277250 113469 277284
rect 113503 277250 113537 277284
rect 113571 277250 113605 277284
rect 113639 277250 113673 277284
rect 113707 277250 113741 277284
rect 113775 277250 113809 277284
rect 113843 277250 113877 277284
rect 113911 277250 113945 277284
rect 113979 277250 114013 277284
rect 114047 277250 114070 277284
rect 112970 277238 114070 277250
rect 111524 277174 112624 277186
rect 111524 277140 111547 277174
rect 111581 277140 111615 277174
rect 111649 277140 111683 277174
rect 111717 277140 111751 277174
rect 111785 277140 111819 277174
rect 111853 277140 111887 277174
rect 111921 277140 111955 277174
rect 111989 277140 112023 277174
rect 112057 277140 112091 277174
rect 112125 277140 112159 277174
rect 112193 277140 112227 277174
rect 112261 277140 112295 277174
rect 112329 277140 112363 277174
rect 112397 277140 112431 277174
rect 112465 277140 112499 277174
rect 112533 277140 112567 277174
rect 112601 277140 112624 277174
rect 111524 277128 112624 277140
rect 112970 277118 114070 277130
rect 112970 277084 112993 277118
rect 113027 277084 113061 277118
rect 113095 277084 113129 277118
rect 113163 277084 113197 277118
rect 113231 277084 113265 277118
rect 113299 277084 113333 277118
rect 113367 277084 113401 277118
rect 113435 277084 113469 277118
rect 113503 277084 113537 277118
rect 113571 277084 113605 277118
rect 113639 277084 113673 277118
rect 113707 277084 113741 277118
rect 113775 277084 113809 277118
rect 113843 277084 113877 277118
rect 113911 277084 113945 277118
rect 113979 277084 114013 277118
rect 114047 277084 114070 277118
rect 112970 277072 114070 277084
rect 111524 276956 112624 276968
rect 111524 276922 111547 276956
rect 111581 276922 111615 276956
rect 111649 276922 111683 276956
rect 111717 276922 111751 276956
rect 111785 276922 111819 276956
rect 111853 276922 111887 276956
rect 111921 276922 111955 276956
rect 111989 276922 112023 276956
rect 112057 276922 112091 276956
rect 112125 276922 112159 276956
rect 112193 276922 112227 276956
rect 112261 276922 112295 276956
rect 112329 276922 112363 276956
rect 112397 276922 112431 276956
rect 112465 276922 112499 276956
rect 112533 276922 112567 276956
rect 112601 276922 112624 276956
rect 111524 276910 112624 276922
rect 112970 276860 114070 276872
rect 112970 276826 112993 276860
rect 113027 276826 113061 276860
rect 113095 276826 113129 276860
rect 113163 276826 113197 276860
rect 113231 276826 113265 276860
rect 113299 276826 113333 276860
rect 113367 276826 113401 276860
rect 113435 276826 113469 276860
rect 113503 276826 113537 276860
rect 113571 276826 113605 276860
rect 113639 276826 113673 276860
rect 113707 276826 113741 276860
rect 113775 276826 113809 276860
rect 113843 276826 113877 276860
rect 113911 276826 113945 276860
rect 113979 276826 114013 276860
rect 114047 276826 114070 276860
rect 111524 276814 112624 276826
rect 112970 276814 114070 276826
rect 111524 276780 111547 276814
rect 111581 276780 111615 276814
rect 111649 276780 111683 276814
rect 111717 276780 111751 276814
rect 111785 276780 111819 276814
rect 111853 276780 111887 276814
rect 111921 276780 111955 276814
rect 111989 276780 112023 276814
rect 112057 276780 112091 276814
rect 112125 276780 112159 276814
rect 112193 276780 112227 276814
rect 112261 276780 112295 276814
rect 112329 276780 112363 276814
rect 112397 276780 112431 276814
rect 112465 276780 112499 276814
rect 112533 276780 112567 276814
rect 112601 276780 112624 276814
rect 111524 276768 112624 276780
rect 113000 276716 114100 276728
rect 113000 276682 113023 276716
rect 113057 276682 113091 276716
rect 113125 276682 113159 276716
rect 113193 276682 113227 276716
rect 113261 276682 113295 276716
rect 113329 276682 113363 276716
rect 113397 276682 113431 276716
rect 113465 276682 113499 276716
rect 113533 276682 113567 276716
rect 113601 276682 113635 276716
rect 113669 276682 113703 276716
rect 113737 276682 113771 276716
rect 113805 276682 113839 276716
rect 113873 276682 113907 276716
rect 113941 276682 113975 276716
rect 114009 276682 114043 276716
rect 114077 276682 114100 276716
rect 113000 276670 114100 276682
rect 111524 276596 112624 276608
rect 111524 276562 111547 276596
rect 111581 276562 111615 276596
rect 111649 276562 111683 276596
rect 111717 276562 111751 276596
rect 111785 276562 111819 276596
rect 111853 276562 111887 276596
rect 111921 276562 111955 276596
rect 111989 276562 112023 276596
rect 112057 276562 112091 276596
rect 112125 276562 112159 276596
rect 112193 276562 112227 276596
rect 112261 276562 112295 276596
rect 112329 276562 112363 276596
rect 112397 276562 112431 276596
rect 112465 276562 112499 276596
rect 112533 276562 112567 276596
rect 112601 276562 112624 276596
rect 111524 276550 112624 276562
rect 113000 276578 114100 276590
rect 113000 276544 113023 276578
rect 113057 276544 113091 276578
rect 113125 276544 113159 276578
rect 113193 276544 113227 276578
rect 113261 276544 113295 276578
rect 113329 276544 113363 276578
rect 113397 276544 113431 276578
rect 113465 276544 113499 276578
rect 113533 276544 113567 276578
rect 113601 276544 113635 276578
rect 113669 276544 113703 276578
rect 113737 276544 113771 276578
rect 113805 276544 113839 276578
rect 113873 276544 113907 276578
rect 113941 276544 113975 276578
rect 114009 276544 114043 276578
rect 114077 276544 114100 276578
rect 113000 276532 114100 276544
rect 111524 276454 112624 276466
rect 111524 276420 111547 276454
rect 111581 276420 111615 276454
rect 111649 276420 111683 276454
rect 111717 276420 111751 276454
rect 111785 276420 111819 276454
rect 111853 276420 111887 276454
rect 111921 276420 111955 276454
rect 111989 276420 112023 276454
rect 112057 276420 112091 276454
rect 112125 276420 112159 276454
rect 112193 276420 112227 276454
rect 112261 276420 112295 276454
rect 112329 276420 112363 276454
rect 112397 276420 112431 276454
rect 112465 276420 112499 276454
rect 112533 276420 112567 276454
rect 112601 276420 112624 276454
rect 111524 276408 112624 276420
rect 113000 276418 114100 276430
rect 113000 276384 113023 276418
rect 113057 276384 113091 276418
rect 113125 276384 113159 276418
rect 113193 276384 113227 276418
rect 113261 276384 113295 276418
rect 113329 276384 113363 276418
rect 113397 276384 113431 276418
rect 113465 276384 113499 276418
rect 113533 276384 113567 276418
rect 113601 276384 113635 276418
rect 113669 276384 113703 276418
rect 113737 276384 113771 276418
rect 113805 276384 113839 276418
rect 113873 276384 113907 276418
rect 113941 276384 113975 276418
rect 114009 276384 114043 276418
rect 114077 276384 114100 276418
rect 113000 276372 114100 276384
rect 113000 276280 114100 276292
rect 111524 276236 112624 276248
rect 111524 276202 111547 276236
rect 111581 276202 111615 276236
rect 111649 276202 111683 276236
rect 111717 276202 111751 276236
rect 111785 276202 111819 276236
rect 111853 276202 111887 276236
rect 111921 276202 111955 276236
rect 111989 276202 112023 276236
rect 112057 276202 112091 276236
rect 112125 276202 112159 276236
rect 112193 276202 112227 276236
rect 112261 276202 112295 276236
rect 112329 276202 112363 276236
rect 112397 276202 112431 276236
rect 112465 276202 112499 276236
rect 112533 276202 112567 276236
rect 112601 276202 112624 276236
rect 113000 276246 113023 276280
rect 113057 276246 113091 276280
rect 113125 276246 113159 276280
rect 113193 276246 113227 276280
rect 113261 276246 113295 276280
rect 113329 276246 113363 276280
rect 113397 276246 113431 276280
rect 113465 276246 113499 276280
rect 113533 276246 113567 276280
rect 113601 276246 113635 276280
rect 113669 276246 113703 276280
rect 113737 276246 113771 276280
rect 113805 276246 113839 276280
rect 113873 276246 113907 276280
rect 113941 276246 113975 276280
rect 114009 276246 114043 276280
rect 114077 276246 114100 276280
rect 113000 276234 114100 276246
rect 111524 276190 112624 276202
rect 116135 277542 117235 277554
rect 116135 277508 116158 277542
rect 116192 277508 116226 277542
rect 116260 277508 116294 277542
rect 116328 277508 116362 277542
rect 116396 277508 116430 277542
rect 116464 277508 116498 277542
rect 116532 277508 116566 277542
rect 116600 277508 116634 277542
rect 116668 277508 116702 277542
rect 116736 277508 116770 277542
rect 116804 277508 116838 277542
rect 116872 277508 116906 277542
rect 116940 277508 116974 277542
rect 117008 277508 117042 277542
rect 117076 277508 117110 277542
rect 117144 277508 117178 277542
rect 117212 277508 117235 277542
rect 116135 277496 117235 277508
rect 117581 277534 118681 277546
rect 117581 277500 117604 277534
rect 117638 277500 117672 277534
rect 117706 277500 117740 277534
rect 117774 277500 117808 277534
rect 117842 277500 117876 277534
rect 117910 277500 117944 277534
rect 117978 277500 118012 277534
rect 118046 277500 118080 277534
rect 118114 277500 118148 277534
rect 118182 277500 118216 277534
rect 118250 277500 118284 277534
rect 118318 277500 118352 277534
rect 118386 277500 118420 277534
rect 118454 277500 118488 277534
rect 118522 277500 118556 277534
rect 118590 277500 118624 277534
rect 118658 277500 118681 277534
rect 117581 277488 118681 277500
rect 117581 277316 118681 277328
rect 116135 277284 117235 277296
rect 116135 277250 116158 277284
rect 116192 277250 116226 277284
rect 116260 277250 116294 277284
rect 116328 277250 116362 277284
rect 116396 277250 116430 277284
rect 116464 277250 116498 277284
rect 116532 277250 116566 277284
rect 116600 277250 116634 277284
rect 116668 277250 116702 277284
rect 116736 277250 116770 277284
rect 116804 277250 116838 277284
rect 116872 277250 116906 277284
rect 116940 277250 116974 277284
rect 117008 277250 117042 277284
rect 117076 277250 117110 277284
rect 117144 277250 117178 277284
rect 117212 277250 117235 277284
rect 117581 277282 117604 277316
rect 117638 277282 117672 277316
rect 117706 277282 117740 277316
rect 117774 277282 117808 277316
rect 117842 277282 117876 277316
rect 117910 277282 117944 277316
rect 117978 277282 118012 277316
rect 118046 277282 118080 277316
rect 118114 277282 118148 277316
rect 118182 277282 118216 277316
rect 118250 277282 118284 277316
rect 118318 277282 118352 277316
rect 118386 277282 118420 277316
rect 118454 277282 118488 277316
rect 118522 277282 118556 277316
rect 118590 277282 118624 277316
rect 118658 277282 118681 277316
rect 117581 277270 118681 277282
rect 116135 277238 117235 277250
rect 117581 277174 118681 277186
rect 117581 277140 117604 277174
rect 117638 277140 117672 277174
rect 117706 277140 117740 277174
rect 117774 277140 117808 277174
rect 117842 277140 117876 277174
rect 117910 277140 117944 277174
rect 117978 277140 118012 277174
rect 118046 277140 118080 277174
rect 118114 277140 118148 277174
rect 118182 277140 118216 277174
rect 118250 277140 118284 277174
rect 118318 277140 118352 277174
rect 118386 277140 118420 277174
rect 118454 277140 118488 277174
rect 118522 277140 118556 277174
rect 118590 277140 118624 277174
rect 118658 277140 118681 277174
rect 116135 277118 117235 277130
rect 117581 277128 118681 277140
rect 116135 277084 116158 277118
rect 116192 277084 116226 277118
rect 116260 277084 116294 277118
rect 116328 277084 116362 277118
rect 116396 277084 116430 277118
rect 116464 277084 116498 277118
rect 116532 277084 116566 277118
rect 116600 277084 116634 277118
rect 116668 277084 116702 277118
rect 116736 277084 116770 277118
rect 116804 277084 116838 277118
rect 116872 277084 116906 277118
rect 116940 277084 116974 277118
rect 117008 277084 117042 277118
rect 117076 277084 117110 277118
rect 117144 277084 117178 277118
rect 117212 277084 117235 277118
rect 116135 277072 117235 277084
rect 117581 276956 118681 276968
rect 117581 276922 117604 276956
rect 117638 276922 117672 276956
rect 117706 276922 117740 276956
rect 117774 276922 117808 276956
rect 117842 276922 117876 276956
rect 117910 276922 117944 276956
rect 117978 276922 118012 276956
rect 118046 276922 118080 276956
rect 118114 276922 118148 276956
rect 118182 276922 118216 276956
rect 118250 276922 118284 276956
rect 118318 276922 118352 276956
rect 118386 276922 118420 276956
rect 118454 276922 118488 276956
rect 118522 276922 118556 276956
rect 118590 276922 118624 276956
rect 118658 276922 118681 276956
rect 117581 276910 118681 276922
rect 116135 276860 117235 276872
rect 116135 276826 116158 276860
rect 116192 276826 116226 276860
rect 116260 276826 116294 276860
rect 116328 276826 116362 276860
rect 116396 276826 116430 276860
rect 116464 276826 116498 276860
rect 116532 276826 116566 276860
rect 116600 276826 116634 276860
rect 116668 276826 116702 276860
rect 116736 276826 116770 276860
rect 116804 276826 116838 276860
rect 116872 276826 116906 276860
rect 116940 276826 116974 276860
rect 117008 276826 117042 276860
rect 117076 276826 117110 276860
rect 117144 276826 117178 276860
rect 117212 276826 117235 276860
rect 116135 276814 117235 276826
rect 117581 276814 118681 276826
rect 117581 276780 117604 276814
rect 117638 276780 117672 276814
rect 117706 276780 117740 276814
rect 117774 276780 117808 276814
rect 117842 276780 117876 276814
rect 117910 276780 117944 276814
rect 117978 276780 118012 276814
rect 118046 276780 118080 276814
rect 118114 276780 118148 276814
rect 118182 276780 118216 276814
rect 118250 276780 118284 276814
rect 118318 276780 118352 276814
rect 118386 276780 118420 276814
rect 118454 276780 118488 276814
rect 118522 276780 118556 276814
rect 118590 276780 118624 276814
rect 118658 276780 118681 276814
rect 117581 276768 118681 276780
rect 116105 276716 117205 276728
rect 116105 276682 116128 276716
rect 116162 276682 116196 276716
rect 116230 276682 116264 276716
rect 116298 276682 116332 276716
rect 116366 276682 116400 276716
rect 116434 276682 116468 276716
rect 116502 276682 116536 276716
rect 116570 276682 116604 276716
rect 116638 276682 116672 276716
rect 116706 276682 116740 276716
rect 116774 276682 116808 276716
rect 116842 276682 116876 276716
rect 116910 276682 116944 276716
rect 116978 276682 117012 276716
rect 117046 276682 117080 276716
rect 117114 276682 117148 276716
rect 117182 276682 117205 276716
rect 116105 276670 117205 276682
rect 117581 276596 118681 276608
rect 116105 276578 117205 276590
rect 116105 276544 116128 276578
rect 116162 276544 116196 276578
rect 116230 276544 116264 276578
rect 116298 276544 116332 276578
rect 116366 276544 116400 276578
rect 116434 276544 116468 276578
rect 116502 276544 116536 276578
rect 116570 276544 116604 276578
rect 116638 276544 116672 276578
rect 116706 276544 116740 276578
rect 116774 276544 116808 276578
rect 116842 276544 116876 276578
rect 116910 276544 116944 276578
rect 116978 276544 117012 276578
rect 117046 276544 117080 276578
rect 117114 276544 117148 276578
rect 117182 276544 117205 276578
rect 117581 276562 117604 276596
rect 117638 276562 117672 276596
rect 117706 276562 117740 276596
rect 117774 276562 117808 276596
rect 117842 276562 117876 276596
rect 117910 276562 117944 276596
rect 117978 276562 118012 276596
rect 118046 276562 118080 276596
rect 118114 276562 118148 276596
rect 118182 276562 118216 276596
rect 118250 276562 118284 276596
rect 118318 276562 118352 276596
rect 118386 276562 118420 276596
rect 118454 276562 118488 276596
rect 118522 276562 118556 276596
rect 118590 276562 118624 276596
rect 118658 276562 118681 276596
rect 117581 276550 118681 276562
rect 116105 276532 117205 276544
rect 117581 276454 118681 276466
rect 116105 276418 117205 276430
rect 116105 276384 116128 276418
rect 116162 276384 116196 276418
rect 116230 276384 116264 276418
rect 116298 276384 116332 276418
rect 116366 276384 116400 276418
rect 116434 276384 116468 276418
rect 116502 276384 116536 276418
rect 116570 276384 116604 276418
rect 116638 276384 116672 276418
rect 116706 276384 116740 276418
rect 116774 276384 116808 276418
rect 116842 276384 116876 276418
rect 116910 276384 116944 276418
rect 116978 276384 117012 276418
rect 117046 276384 117080 276418
rect 117114 276384 117148 276418
rect 117182 276384 117205 276418
rect 117581 276420 117604 276454
rect 117638 276420 117672 276454
rect 117706 276420 117740 276454
rect 117774 276420 117808 276454
rect 117842 276420 117876 276454
rect 117910 276420 117944 276454
rect 117978 276420 118012 276454
rect 118046 276420 118080 276454
rect 118114 276420 118148 276454
rect 118182 276420 118216 276454
rect 118250 276420 118284 276454
rect 118318 276420 118352 276454
rect 118386 276420 118420 276454
rect 118454 276420 118488 276454
rect 118522 276420 118556 276454
rect 118590 276420 118624 276454
rect 118658 276420 118681 276454
rect 117581 276408 118681 276420
rect 116105 276372 117205 276384
rect 116105 276280 117205 276292
rect 116105 276246 116128 276280
rect 116162 276246 116196 276280
rect 116230 276246 116264 276280
rect 116298 276246 116332 276280
rect 116366 276246 116400 276280
rect 116434 276246 116468 276280
rect 116502 276246 116536 276280
rect 116570 276246 116604 276280
rect 116638 276246 116672 276280
rect 116706 276246 116740 276280
rect 116774 276246 116808 276280
rect 116842 276246 116876 276280
rect 116910 276246 116944 276280
rect 116978 276246 117012 276280
rect 117046 276246 117080 276280
rect 117114 276246 117148 276280
rect 117182 276246 117205 276280
rect 116105 276234 117205 276246
rect 117581 276236 118681 276248
rect 117581 276202 117604 276236
rect 117638 276202 117672 276236
rect 117706 276202 117740 276236
rect 117774 276202 117808 276236
rect 117842 276202 117876 276236
rect 117910 276202 117944 276236
rect 117978 276202 118012 276236
rect 118046 276202 118080 276236
rect 118114 276202 118148 276236
rect 118182 276202 118216 276236
rect 118250 276202 118284 276236
rect 118318 276202 118352 276236
rect 118386 276202 118420 276236
rect 118454 276202 118488 276236
rect 118522 276202 118556 276236
rect 118590 276202 118624 276236
rect 118658 276202 118681 276236
rect 117581 276190 118681 276202
rect 111524 275868 112624 275880
rect 111524 275834 111547 275868
rect 111581 275834 111615 275868
rect 111649 275834 111683 275868
rect 111717 275834 111751 275868
rect 111785 275834 111819 275868
rect 111853 275834 111887 275868
rect 111921 275834 111955 275868
rect 111989 275834 112023 275868
rect 112057 275834 112091 275868
rect 112125 275834 112159 275868
rect 112193 275834 112227 275868
rect 112261 275834 112295 275868
rect 112329 275834 112363 275868
rect 112397 275834 112431 275868
rect 112465 275834 112499 275868
rect 112533 275834 112567 275868
rect 112601 275834 112624 275868
rect 111524 275822 112624 275834
rect 112970 275876 114070 275888
rect 112970 275842 112993 275876
rect 113027 275842 113061 275876
rect 113095 275842 113129 275876
rect 113163 275842 113197 275876
rect 113231 275842 113265 275876
rect 113299 275842 113333 275876
rect 113367 275842 113401 275876
rect 113435 275842 113469 275876
rect 113503 275842 113537 275876
rect 113571 275842 113605 275876
rect 113639 275842 113673 275876
rect 113707 275842 113741 275876
rect 113775 275842 113809 275876
rect 113843 275842 113877 275876
rect 113911 275842 113945 275876
rect 113979 275842 114013 275876
rect 114047 275842 114070 275876
rect 112970 275830 114070 275842
rect 111524 275650 112624 275662
rect 111524 275616 111547 275650
rect 111581 275616 111615 275650
rect 111649 275616 111683 275650
rect 111717 275616 111751 275650
rect 111785 275616 111819 275650
rect 111853 275616 111887 275650
rect 111921 275616 111955 275650
rect 111989 275616 112023 275650
rect 112057 275616 112091 275650
rect 112125 275616 112159 275650
rect 112193 275616 112227 275650
rect 112261 275616 112295 275650
rect 112329 275616 112363 275650
rect 112397 275616 112431 275650
rect 112465 275616 112499 275650
rect 112533 275616 112567 275650
rect 112601 275616 112624 275650
rect 111524 275604 112624 275616
rect 112970 275618 114070 275630
rect 112970 275584 112993 275618
rect 113027 275584 113061 275618
rect 113095 275584 113129 275618
rect 113163 275584 113197 275618
rect 113231 275584 113265 275618
rect 113299 275584 113333 275618
rect 113367 275584 113401 275618
rect 113435 275584 113469 275618
rect 113503 275584 113537 275618
rect 113571 275584 113605 275618
rect 113639 275584 113673 275618
rect 113707 275584 113741 275618
rect 113775 275584 113809 275618
rect 113843 275584 113877 275618
rect 113911 275584 113945 275618
rect 113979 275584 114013 275618
rect 114047 275584 114070 275618
rect 112970 275572 114070 275584
rect 111524 275508 112624 275520
rect 111524 275474 111547 275508
rect 111581 275474 111615 275508
rect 111649 275474 111683 275508
rect 111717 275474 111751 275508
rect 111785 275474 111819 275508
rect 111853 275474 111887 275508
rect 111921 275474 111955 275508
rect 111989 275474 112023 275508
rect 112057 275474 112091 275508
rect 112125 275474 112159 275508
rect 112193 275474 112227 275508
rect 112261 275474 112295 275508
rect 112329 275474 112363 275508
rect 112397 275474 112431 275508
rect 112465 275474 112499 275508
rect 112533 275474 112567 275508
rect 112601 275474 112624 275508
rect 111524 275462 112624 275474
rect 112970 275452 114070 275464
rect 112970 275418 112993 275452
rect 113027 275418 113061 275452
rect 113095 275418 113129 275452
rect 113163 275418 113197 275452
rect 113231 275418 113265 275452
rect 113299 275418 113333 275452
rect 113367 275418 113401 275452
rect 113435 275418 113469 275452
rect 113503 275418 113537 275452
rect 113571 275418 113605 275452
rect 113639 275418 113673 275452
rect 113707 275418 113741 275452
rect 113775 275418 113809 275452
rect 113843 275418 113877 275452
rect 113911 275418 113945 275452
rect 113979 275418 114013 275452
rect 114047 275418 114070 275452
rect 112970 275406 114070 275418
rect 111524 275290 112624 275302
rect 111524 275256 111547 275290
rect 111581 275256 111615 275290
rect 111649 275256 111683 275290
rect 111717 275256 111751 275290
rect 111785 275256 111819 275290
rect 111853 275256 111887 275290
rect 111921 275256 111955 275290
rect 111989 275256 112023 275290
rect 112057 275256 112091 275290
rect 112125 275256 112159 275290
rect 112193 275256 112227 275290
rect 112261 275256 112295 275290
rect 112329 275256 112363 275290
rect 112397 275256 112431 275290
rect 112465 275256 112499 275290
rect 112533 275256 112567 275290
rect 112601 275256 112624 275290
rect 111524 275244 112624 275256
rect 112970 275194 114070 275206
rect 112970 275160 112993 275194
rect 113027 275160 113061 275194
rect 113095 275160 113129 275194
rect 113163 275160 113197 275194
rect 113231 275160 113265 275194
rect 113299 275160 113333 275194
rect 113367 275160 113401 275194
rect 113435 275160 113469 275194
rect 113503 275160 113537 275194
rect 113571 275160 113605 275194
rect 113639 275160 113673 275194
rect 113707 275160 113741 275194
rect 113775 275160 113809 275194
rect 113843 275160 113877 275194
rect 113911 275160 113945 275194
rect 113979 275160 114013 275194
rect 114047 275160 114070 275194
rect 111524 275148 112624 275160
rect 112970 275148 114070 275160
rect 111524 275114 111547 275148
rect 111581 275114 111615 275148
rect 111649 275114 111683 275148
rect 111717 275114 111751 275148
rect 111785 275114 111819 275148
rect 111853 275114 111887 275148
rect 111921 275114 111955 275148
rect 111989 275114 112023 275148
rect 112057 275114 112091 275148
rect 112125 275114 112159 275148
rect 112193 275114 112227 275148
rect 112261 275114 112295 275148
rect 112329 275114 112363 275148
rect 112397 275114 112431 275148
rect 112465 275114 112499 275148
rect 112533 275114 112567 275148
rect 112601 275114 112624 275148
rect 111524 275102 112624 275114
rect 113000 275050 114100 275062
rect 113000 275016 113023 275050
rect 113057 275016 113091 275050
rect 113125 275016 113159 275050
rect 113193 275016 113227 275050
rect 113261 275016 113295 275050
rect 113329 275016 113363 275050
rect 113397 275016 113431 275050
rect 113465 275016 113499 275050
rect 113533 275016 113567 275050
rect 113601 275016 113635 275050
rect 113669 275016 113703 275050
rect 113737 275016 113771 275050
rect 113805 275016 113839 275050
rect 113873 275016 113907 275050
rect 113941 275016 113975 275050
rect 114009 275016 114043 275050
rect 114077 275016 114100 275050
rect 113000 275004 114100 275016
rect 111524 274930 112624 274942
rect 111524 274896 111547 274930
rect 111581 274896 111615 274930
rect 111649 274896 111683 274930
rect 111717 274896 111751 274930
rect 111785 274896 111819 274930
rect 111853 274896 111887 274930
rect 111921 274896 111955 274930
rect 111989 274896 112023 274930
rect 112057 274896 112091 274930
rect 112125 274896 112159 274930
rect 112193 274896 112227 274930
rect 112261 274896 112295 274930
rect 112329 274896 112363 274930
rect 112397 274896 112431 274930
rect 112465 274896 112499 274930
rect 112533 274896 112567 274930
rect 112601 274896 112624 274930
rect 111524 274884 112624 274896
rect 113000 274912 114100 274924
rect 113000 274878 113023 274912
rect 113057 274878 113091 274912
rect 113125 274878 113159 274912
rect 113193 274878 113227 274912
rect 113261 274878 113295 274912
rect 113329 274878 113363 274912
rect 113397 274878 113431 274912
rect 113465 274878 113499 274912
rect 113533 274878 113567 274912
rect 113601 274878 113635 274912
rect 113669 274878 113703 274912
rect 113737 274878 113771 274912
rect 113805 274878 113839 274912
rect 113873 274878 113907 274912
rect 113941 274878 113975 274912
rect 114009 274878 114043 274912
rect 114077 274878 114100 274912
rect 113000 274866 114100 274878
rect 111524 274788 112624 274800
rect 111524 274754 111547 274788
rect 111581 274754 111615 274788
rect 111649 274754 111683 274788
rect 111717 274754 111751 274788
rect 111785 274754 111819 274788
rect 111853 274754 111887 274788
rect 111921 274754 111955 274788
rect 111989 274754 112023 274788
rect 112057 274754 112091 274788
rect 112125 274754 112159 274788
rect 112193 274754 112227 274788
rect 112261 274754 112295 274788
rect 112329 274754 112363 274788
rect 112397 274754 112431 274788
rect 112465 274754 112499 274788
rect 112533 274754 112567 274788
rect 112601 274754 112624 274788
rect 111524 274742 112624 274754
rect 113000 274752 114100 274764
rect 113000 274718 113023 274752
rect 113057 274718 113091 274752
rect 113125 274718 113159 274752
rect 113193 274718 113227 274752
rect 113261 274718 113295 274752
rect 113329 274718 113363 274752
rect 113397 274718 113431 274752
rect 113465 274718 113499 274752
rect 113533 274718 113567 274752
rect 113601 274718 113635 274752
rect 113669 274718 113703 274752
rect 113737 274718 113771 274752
rect 113805 274718 113839 274752
rect 113873 274718 113907 274752
rect 113941 274718 113975 274752
rect 114009 274718 114043 274752
rect 114077 274718 114100 274752
rect 113000 274706 114100 274718
rect 113000 274614 114100 274626
rect 111524 274570 112624 274582
rect 111524 274536 111547 274570
rect 111581 274536 111615 274570
rect 111649 274536 111683 274570
rect 111717 274536 111751 274570
rect 111785 274536 111819 274570
rect 111853 274536 111887 274570
rect 111921 274536 111955 274570
rect 111989 274536 112023 274570
rect 112057 274536 112091 274570
rect 112125 274536 112159 274570
rect 112193 274536 112227 274570
rect 112261 274536 112295 274570
rect 112329 274536 112363 274570
rect 112397 274536 112431 274570
rect 112465 274536 112499 274570
rect 112533 274536 112567 274570
rect 112601 274536 112624 274570
rect 113000 274580 113023 274614
rect 113057 274580 113091 274614
rect 113125 274580 113159 274614
rect 113193 274580 113227 274614
rect 113261 274580 113295 274614
rect 113329 274580 113363 274614
rect 113397 274580 113431 274614
rect 113465 274580 113499 274614
rect 113533 274580 113567 274614
rect 113601 274580 113635 274614
rect 113669 274580 113703 274614
rect 113737 274580 113771 274614
rect 113805 274580 113839 274614
rect 113873 274580 113907 274614
rect 113941 274580 113975 274614
rect 114009 274580 114043 274614
rect 114077 274580 114100 274614
rect 113000 274568 114100 274580
rect 111524 274524 112624 274536
rect 116135 275876 117235 275888
rect 116135 275842 116158 275876
rect 116192 275842 116226 275876
rect 116260 275842 116294 275876
rect 116328 275842 116362 275876
rect 116396 275842 116430 275876
rect 116464 275842 116498 275876
rect 116532 275842 116566 275876
rect 116600 275842 116634 275876
rect 116668 275842 116702 275876
rect 116736 275842 116770 275876
rect 116804 275842 116838 275876
rect 116872 275842 116906 275876
rect 116940 275842 116974 275876
rect 117008 275842 117042 275876
rect 117076 275842 117110 275876
rect 117144 275842 117178 275876
rect 117212 275842 117235 275876
rect 116135 275830 117235 275842
rect 117581 275868 118681 275880
rect 117581 275834 117604 275868
rect 117638 275834 117672 275868
rect 117706 275834 117740 275868
rect 117774 275834 117808 275868
rect 117842 275834 117876 275868
rect 117910 275834 117944 275868
rect 117978 275834 118012 275868
rect 118046 275834 118080 275868
rect 118114 275834 118148 275868
rect 118182 275834 118216 275868
rect 118250 275834 118284 275868
rect 118318 275834 118352 275868
rect 118386 275834 118420 275868
rect 118454 275834 118488 275868
rect 118522 275834 118556 275868
rect 118590 275834 118624 275868
rect 118658 275834 118681 275868
rect 117581 275822 118681 275834
rect 117581 275650 118681 275662
rect 116135 275618 117235 275630
rect 116135 275584 116158 275618
rect 116192 275584 116226 275618
rect 116260 275584 116294 275618
rect 116328 275584 116362 275618
rect 116396 275584 116430 275618
rect 116464 275584 116498 275618
rect 116532 275584 116566 275618
rect 116600 275584 116634 275618
rect 116668 275584 116702 275618
rect 116736 275584 116770 275618
rect 116804 275584 116838 275618
rect 116872 275584 116906 275618
rect 116940 275584 116974 275618
rect 117008 275584 117042 275618
rect 117076 275584 117110 275618
rect 117144 275584 117178 275618
rect 117212 275584 117235 275618
rect 117581 275616 117604 275650
rect 117638 275616 117672 275650
rect 117706 275616 117740 275650
rect 117774 275616 117808 275650
rect 117842 275616 117876 275650
rect 117910 275616 117944 275650
rect 117978 275616 118012 275650
rect 118046 275616 118080 275650
rect 118114 275616 118148 275650
rect 118182 275616 118216 275650
rect 118250 275616 118284 275650
rect 118318 275616 118352 275650
rect 118386 275616 118420 275650
rect 118454 275616 118488 275650
rect 118522 275616 118556 275650
rect 118590 275616 118624 275650
rect 118658 275616 118681 275650
rect 117581 275604 118681 275616
rect 116135 275572 117235 275584
rect 117581 275508 118681 275520
rect 117581 275474 117604 275508
rect 117638 275474 117672 275508
rect 117706 275474 117740 275508
rect 117774 275474 117808 275508
rect 117842 275474 117876 275508
rect 117910 275474 117944 275508
rect 117978 275474 118012 275508
rect 118046 275474 118080 275508
rect 118114 275474 118148 275508
rect 118182 275474 118216 275508
rect 118250 275474 118284 275508
rect 118318 275474 118352 275508
rect 118386 275474 118420 275508
rect 118454 275474 118488 275508
rect 118522 275474 118556 275508
rect 118590 275474 118624 275508
rect 118658 275474 118681 275508
rect 116135 275452 117235 275464
rect 117581 275462 118681 275474
rect 116135 275418 116158 275452
rect 116192 275418 116226 275452
rect 116260 275418 116294 275452
rect 116328 275418 116362 275452
rect 116396 275418 116430 275452
rect 116464 275418 116498 275452
rect 116532 275418 116566 275452
rect 116600 275418 116634 275452
rect 116668 275418 116702 275452
rect 116736 275418 116770 275452
rect 116804 275418 116838 275452
rect 116872 275418 116906 275452
rect 116940 275418 116974 275452
rect 117008 275418 117042 275452
rect 117076 275418 117110 275452
rect 117144 275418 117178 275452
rect 117212 275418 117235 275452
rect 116135 275406 117235 275418
rect 117581 275290 118681 275302
rect 117581 275256 117604 275290
rect 117638 275256 117672 275290
rect 117706 275256 117740 275290
rect 117774 275256 117808 275290
rect 117842 275256 117876 275290
rect 117910 275256 117944 275290
rect 117978 275256 118012 275290
rect 118046 275256 118080 275290
rect 118114 275256 118148 275290
rect 118182 275256 118216 275290
rect 118250 275256 118284 275290
rect 118318 275256 118352 275290
rect 118386 275256 118420 275290
rect 118454 275256 118488 275290
rect 118522 275256 118556 275290
rect 118590 275256 118624 275290
rect 118658 275256 118681 275290
rect 117581 275244 118681 275256
rect 116135 275194 117235 275206
rect 116135 275160 116158 275194
rect 116192 275160 116226 275194
rect 116260 275160 116294 275194
rect 116328 275160 116362 275194
rect 116396 275160 116430 275194
rect 116464 275160 116498 275194
rect 116532 275160 116566 275194
rect 116600 275160 116634 275194
rect 116668 275160 116702 275194
rect 116736 275160 116770 275194
rect 116804 275160 116838 275194
rect 116872 275160 116906 275194
rect 116940 275160 116974 275194
rect 117008 275160 117042 275194
rect 117076 275160 117110 275194
rect 117144 275160 117178 275194
rect 117212 275160 117235 275194
rect 116135 275148 117235 275160
rect 117581 275148 118681 275160
rect 117581 275114 117604 275148
rect 117638 275114 117672 275148
rect 117706 275114 117740 275148
rect 117774 275114 117808 275148
rect 117842 275114 117876 275148
rect 117910 275114 117944 275148
rect 117978 275114 118012 275148
rect 118046 275114 118080 275148
rect 118114 275114 118148 275148
rect 118182 275114 118216 275148
rect 118250 275114 118284 275148
rect 118318 275114 118352 275148
rect 118386 275114 118420 275148
rect 118454 275114 118488 275148
rect 118522 275114 118556 275148
rect 118590 275114 118624 275148
rect 118658 275114 118681 275148
rect 117581 275102 118681 275114
rect 116105 275050 117205 275062
rect 116105 275016 116128 275050
rect 116162 275016 116196 275050
rect 116230 275016 116264 275050
rect 116298 275016 116332 275050
rect 116366 275016 116400 275050
rect 116434 275016 116468 275050
rect 116502 275016 116536 275050
rect 116570 275016 116604 275050
rect 116638 275016 116672 275050
rect 116706 275016 116740 275050
rect 116774 275016 116808 275050
rect 116842 275016 116876 275050
rect 116910 275016 116944 275050
rect 116978 275016 117012 275050
rect 117046 275016 117080 275050
rect 117114 275016 117148 275050
rect 117182 275016 117205 275050
rect 116105 275004 117205 275016
rect 117581 274930 118681 274942
rect 116105 274912 117205 274924
rect 116105 274878 116128 274912
rect 116162 274878 116196 274912
rect 116230 274878 116264 274912
rect 116298 274878 116332 274912
rect 116366 274878 116400 274912
rect 116434 274878 116468 274912
rect 116502 274878 116536 274912
rect 116570 274878 116604 274912
rect 116638 274878 116672 274912
rect 116706 274878 116740 274912
rect 116774 274878 116808 274912
rect 116842 274878 116876 274912
rect 116910 274878 116944 274912
rect 116978 274878 117012 274912
rect 117046 274878 117080 274912
rect 117114 274878 117148 274912
rect 117182 274878 117205 274912
rect 117581 274896 117604 274930
rect 117638 274896 117672 274930
rect 117706 274896 117740 274930
rect 117774 274896 117808 274930
rect 117842 274896 117876 274930
rect 117910 274896 117944 274930
rect 117978 274896 118012 274930
rect 118046 274896 118080 274930
rect 118114 274896 118148 274930
rect 118182 274896 118216 274930
rect 118250 274896 118284 274930
rect 118318 274896 118352 274930
rect 118386 274896 118420 274930
rect 118454 274896 118488 274930
rect 118522 274896 118556 274930
rect 118590 274896 118624 274930
rect 118658 274896 118681 274930
rect 117581 274884 118681 274896
rect 116105 274866 117205 274878
rect 117581 274788 118681 274800
rect 116105 274752 117205 274764
rect 116105 274718 116128 274752
rect 116162 274718 116196 274752
rect 116230 274718 116264 274752
rect 116298 274718 116332 274752
rect 116366 274718 116400 274752
rect 116434 274718 116468 274752
rect 116502 274718 116536 274752
rect 116570 274718 116604 274752
rect 116638 274718 116672 274752
rect 116706 274718 116740 274752
rect 116774 274718 116808 274752
rect 116842 274718 116876 274752
rect 116910 274718 116944 274752
rect 116978 274718 117012 274752
rect 117046 274718 117080 274752
rect 117114 274718 117148 274752
rect 117182 274718 117205 274752
rect 117581 274754 117604 274788
rect 117638 274754 117672 274788
rect 117706 274754 117740 274788
rect 117774 274754 117808 274788
rect 117842 274754 117876 274788
rect 117910 274754 117944 274788
rect 117978 274754 118012 274788
rect 118046 274754 118080 274788
rect 118114 274754 118148 274788
rect 118182 274754 118216 274788
rect 118250 274754 118284 274788
rect 118318 274754 118352 274788
rect 118386 274754 118420 274788
rect 118454 274754 118488 274788
rect 118522 274754 118556 274788
rect 118590 274754 118624 274788
rect 118658 274754 118681 274788
rect 117581 274742 118681 274754
rect 116105 274706 117205 274718
rect 116105 274614 117205 274626
rect 116105 274580 116128 274614
rect 116162 274580 116196 274614
rect 116230 274580 116264 274614
rect 116298 274580 116332 274614
rect 116366 274580 116400 274614
rect 116434 274580 116468 274614
rect 116502 274580 116536 274614
rect 116570 274580 116604 274614
rect 116638 274580 116672 274614
rect 116706 274580 116740 274614
rect 116774 274580 116808 274614
rect 116842 274580 116876 274614
rect 116910 274580 116944 274614
rect 116978 274580 117012 274614
rect 117046 274580 117080 274614
rect 117114 274580 117148 274614
rect 117182 274580 117205 274614
rect 116105 274568 117205 274580
rect 117581 274570 118681 274582
rect 117581 274536 117604 274570
rect 117638 274536 117672 274570
rect 117706 274536 117740 274570
rect 117774 274536 117808 274570
rect 117842 274536 117876 274570
rect 117910 274536 117944 274570
rect 117978 274536 118012 274570
rect 118046 274536 118080 274570
rect 118114 274536 118148 274570
rect 118182 274536 118216 274570
rect 118250 274536 118284 274570
rect 118318 274536 118352 274570
rect 118386 274536 118420 274570
rect 118454 274536 118488 274570
rect 118522 274536 118556 274570
rect 118590 274536 118624 274570
rect 118658 274536 118681 274570
rect 117581 274524 118681 274536
rect 111524 274202 112624 274214
rect 111524 274168 111547 274202
rect 111581 274168 111615 274202
rect 111649 274168 111683 274202
rect 111717 274168 111751 274202
rect 111785 274168 111819 274202
rect 111853 274168 111887 274202
rect 111921 274168 111955 274202
rect 111989 274168 112023 274202
rect 112057 274168 112091 274202
rect 112125 274168 112159 274202
rect 112193 274168 112227 274202
rect 112261 274168 112295 274202
rect 112329 274168 112363 274202
rect 112397 274168 112431 274202
rect 112465 274168 112499 274202
rect 112533 274168 112567 274202
rect 112601 274168 112624 274202
rect 111524 274156 112624 274168
rect 112970 274210 114070 274222
rect 112970 274176 112993 274210
rect 113027 274176 113061 274210
rect 113095 274176 113129 274210
rect 113163 274176 113197 274210
rect 113231 274176 113265 274210
rect 113299 274176 113333 274210
rect 113367 274176 113401 274210
rect 113435 274176 113469 274210
rect 113503 274176 113537 274210
rect 113571 274176 113605 274210
rect 113639 274176 113673 274210
rect 113707 274176 113741 274210
rect 113775 274176 113809 274210
rect 113843 274176 113877 274210
rect 113911 274176 113945 274210
rect 113979 274176 114013 274210
rect 114047 274176 114070 274210
rect 112970 274164 114070 274176
rect 111524 273984 112624 273996
rect 111524 273950 111547 273984
rect 111581 273950 111615 273984
rect 111649 273950 111683 273984
rect 111717 273950 111751 273984
rect 111785 273950 111819 273984
rect 111853 273950 111887 273984
rect 111921 273950 111955 273984
rect 111989 273950 112023 273984
rect 112057 273950 112091 273984
rect 112125 273950 112159 273984
rect 112193 273950 112227 273984
rect 112261 273950 112295 273984
rect 112329 273950 112363 273984
rect 112397 273950 112431 273984
rect 112465 273950 112499 273984
rect 112533 273950 112567 273984
rect 112601 273950 112624 273984
rect 111524 273938 112624 273950
rect 112970 273952 114070 273964
rect 112970 273918 112993 273952
rect 113027 273918 113061 273952
rect 113095 273918 113129 273952
rect 113163 273918 113197 273952
rect 113231 273918 113265 273952
rect 113299 273918 113333 273952
rect 113367 273918 113401 273952
rect 113435 273918 113469 273952
rect 113503 273918 113537 273952
rect 113571 273918 113605 273952
rect 113639 273918 113673 273952
rect 113707 273918 113741 273952
rect 113775 273918 113809 273952
rect 113843 273918 113877 273952
rect 113911 273918 113945 273952
rect 113979 273918 114013 273952
rect 114047 273918 114070 273952
rect 112970 273906 114070 273918
rect 111524 273842 112624 273854
rect 111524 273808 111547 273842
rect 111581 273808 111615 273842
rect 111649 273808 111683 273842
rect 111717 273808 111751 273842
rect 111785 273808 111819 273842
rect 111853 273808 111887 273842
rect 111921 273808 111955 273842
rect 111989 273808 112023 273842
rect 112057 273808 112091 273842
rect 112125 273808 112159 273842
rect 112193 273808 112227 273842
rect 112261 273808 112295 273842
rect 112329 273808 112363 273842
rect 112397 273808 112431 273842
rect 112465 273808 112499 273842
rect 112533 273808 112567 273842
rect 112601 273808 112624 273842
rect 111524 273796 112624 273808
rect 112970 273786 114070 273798
rect 112970 273752 112993 273786
rect 113027 273752 113061 273786
rect 113095 273752 113129 273786
rect 113163 273752 113197 273786
rect 113231 273752 113265 273786
rect 113299 273752 113333 273786
rect 113367 273752 113401 273786
rect 113435 273752 113469 273786
rect 113503 273752 113537 273786
rect 113571 273752 113605 273786
rect 113639 273752 113673 273786
rect 113707 273752 113741 273786
rect 113775 273752 113809 273786
rect 113843 273752 113877 273786
rect 113911 273752 113945 273786
rect 113979 273752 114013 273786
rect 114047 273752 114070 273786
rect 112970 273740 114070 273752
rect 111524 273624 112624 273636
rect 111524 273590 111547 273624
rect 111581 273590 111615 273624
rect 111649 273590 111683 273624
rect 111717 273590 111751 273624
rect 111785 273590 111819 273624
rect 111853 273590 111887 273624
rect 111921 273590 111955 273624
rect 111989 273590 112023 273624
rect 112057 273590 112091 273624
rect 112125 273590 112159 273624
rect 112193 273590 112227 273624
rect 112261 273590 112295 273624
rect 112329 273590 112363 273624
rect 112397 273590 112431 273624
rect 112465 273590 112499 273624
rect 112533 273590 112567 273624
rect 112601 273590 112624 273624
rect 111524 273578 112624 273590
rect 112970 273528 114070 273540
rect 112970 273494 112993 273528
rect 113027 273494 113061 273528
rect 113095 273494 113129 273528
rect 113163 273494 113197 273528
rect 113231 273494 113265 273528
rect 113299 273494 113333 273528
rect 113367 273494 113401 273528
rect 113435 273494 113469 273528
rect 113503 273494 113537 273528
rect 113571 273494 113605 273528
rect 113639 273494 113673 273528
rect 113707 273494 113741 273528
rect 113775 273494 113809 273528
rect 113843 273494 113877 273528
rect 113911 273494 113945 273528
rect 113979 273494 114013 273528
rect 114047 273494 114070 273528
rect 111524 273482 112624 273494
rect 112970 273482 114070 273494
rect 111524 273448 111547 273482
rect 111581 273448 111615 273482
rect 111649 273448 111683 273482
rect 111717 273448 111751 273482
rect 111785 273448 111819 273482
rect 111853 273448 111887 273482
rect 111921 273448 111955 273482
rect 111989 273448 112023 273482
rect 112057 273448 112091 273482
rect 112125 273448 112159 273482
rect 112193 273448 112227 273482
rect 112261 273448 112295 273482
rect 112329 273448 112363 273482
rect 112397 273448 112431 273482
rect 112465 273448 112499 273482
rect 112533 273448 112567 273482
rect 112601 273448 112624 273482
rect 111524 273436 112624 273448
rect 113000 273384 114100 273396
rect 113000 273350 113023 273384
rect 113057 273350 113091 273384
rect 113125 273350 113159 273384
rect 113193 273350 113227 273384
rect 113261 273350 113295 273384
rect 113329 273350 113363 273384
rect 113397 273350 113431 273384
rect 113465 273350 113499 273384
rect 113533 273350 113567 273384
rect 113601 273350 113635 273384
rect 113669 273350 113703 273384
rect 113737 273350 113771 273384
rect 113805 273350 113839 273384
rect 113873 273350 113907 273384
rect 113941 273350 113975 273384
rect 114009 273350 114043 273384
rect 114077 273350 114100 273384
rect 113000 273338 114100 273350
rect 111524 273264 112624 273276
rect 111524 273230 111547 273264
rect 111581 273230 111615 273264
rect 111649 273230 111683 273264
rect 111717 273230 111751 273264
rect 111785 273230 111819 273264
rect 111853 273230 111887 273264
rect 111921 273230 111955 273264
rect 111989 273230 112023 273264
rect 112057 273230 112091 273264
rect 112125 273230 112159 273264
rect 112193 273230 112227 273264
rect 112261 273230 112295 273264
rect 112329 273230 112363 273264
rect 112397 273230 112431 273264
rect 112465 273230 112499 273264
rect 112533 273230 112567 273264
rect 112601 273230 112624 273264
rect 111524 273218 112624 273230
rect 113000 273246 114100 273258
rect 113000 273212 113023 273246
rect 113057 273212 113091 273246
rect 113125 273212 113159 273246
rect 113193 273212 113227 273246
rect 113261 273212 113295 273246
rect 113329 273212 113363 273246
rect 113397 273212 113431 273246
rect 113465 273212 113499 273246
rect 113533 273212 113567 273246
rect 113601 273212 113635 273246
rect 113669 273212 113703 273246
rect 113737 273212 113771 273246
rect 113805 273212 113839 273246
rect 113873 273212 113907 273246
rect 113941 273212 113975 273246
rect 114009 273212 114043 273246
rect 114077 273212 114100 273246
rect 113000 273200 114100 273212
rect 111524 273122 112624 273134
rect 111524 273088 111547 273122
rect 111581 273088 111615 273122
rect 111649 273088 111683 273122
rect 111717 273088 111751 273122
rect 111785 273088 111819 273122
rect 111853 273088 111887 273122
rect 111921 273088 111955 273122
rect 111989 273088 112023 273122
rect 112057 273088 112091 273122
rect 112125 273088 112159 273122
rect 112193 273088 112227 273122
rect 112261 273088 112295 273122
rect 112329 273088 112363 273122
rect 112397 273088 112431 273122
rect 112465 273088 112499 273122
rect 112533 273088 112567 273122
rect 112601 273088 112624 273122
rect 111524 273076 112624 273088
rect 113000 273086 114100 273098
rect 113000 273052 113023 273086
rect 113057 273052 113091 273086
rect 113125 273052 113159 273086
rect 113193 273052 113227 273086
rect 113261 273052 113295 273086
rect 113329 273052 113363 273086
rect 113397 273052 113431 273086
rect 113465 273052 113499 273086
rect 113533 273052 113567 273086
rect 113601 273052 113635 273086
rect 113669 273052 113703 273086
rect 113737 273052 113771 273086
rect 113805 273052 113839 273086
rect 113873 273052 113907 273086
rect 113941 273052 113975 273086
rect 114009 273052 114043 273086
rect 114077 273052 114100 273086
rect 113000 273040 114100 273052
rect 113000 272948 114100 272960
rect 111524 272904 112624 272916
rect 111524 272870 111547 272904
rect 111581 272870 111615 272904
rect 111649 272870 111683 272904
rect 111717 272870 111751 272904
rect 111785 272870 111819 272904
rect 111853 272870 111887 272904
rect 111921 272870 111955 272904
rect 111989 272870 112023 272904
rect 112057 272870 112091 272904
rect 112125 272870 112159 272904
rect 112193 272870 112227 272904
rect 112261 272870 112295 272904
rect 112329 272870 112363 272904
rect 112397 272870 112431 272904
rect 112465 272870 112499 272904
rect 112533 272870 112567 272904
rect 112601 272870 112624 272904
rect 113000 272914 113023 272948
rect 113057 272914 113091 272948
rect 113125 272914 113159 272948
rect 113193 272914 113227 272948
rect 113261 272914 113295 272948
rect 113329 272914 113363 272948
rect 113397 272914 113431 272948
rect 113465 272914 113499 272948
rect 113533 272914 113567 272948
rect 113601 272914 113635 272948
rect 113669 272914 113703 272948
rect 113737 272914 113771 272948
rect 113805 272914 113839 272948
rect 113873 272914 113907 272948
rect 113941 272914 113975 272948
rect 114009 272914 114043 272948
rect 114077 272914 114100 272948
rect 113000 272902 114100 272914
rect 111524 272858 112624 272870
rect 116135 274210 117235 274222
rect 116135 274176 116158 274210
rect 116192 274176 116226 274210
rect 116260 274176 116294 274210
rect 116328 274176 116362 274210
rect 116396 274176 116430 274210
rect 116464 274176 116498 274210
rect 116532 274176 116566 274210
rect 116600 274176 116634 274210
rect 116668 274176 116702 274210
rect 116736 274176 116770 274210
rect 116804 274176 116838 274210
rect 116872 274176 116906 274210
rect 116940 274176 116974 274210
rect 117008 274176 117042 274210
rect 117076 274176 117110 274210
rect 117144 274176 117178 274210
rect 117212 274176 117235 274210
rect 116135 274164 117235 274176
rect 117581 274202 118681 274214
rect 117581 274168 117604 274202
rect 117638 274168 117672 274202
rect 117706 274168 117740 274202
rect 117774 274168 117808 274202
rect 117842 274168 117876 274202
rect 117910 274168 117944 274202
rect 117978 274168 118012 274202
rect 118046 274168 118080 274202
rect 118114 274168 118148 274202
rect 118182 274168 118216 274202
rect 118250 274168 118284 274202
rect 118318 274168 118352 274202
rect 118386 274168 118420 274202
rect 118454 274168 118488 274202
rect 118522 274168 118556 274202
rect 118590 274168 118624 274202
rect 118658 274168 118681 274202
rect 117581 274156 118681 274168
rect 117581 273984 118681 273996
rect 116135 273952 117235 273964
rect 116135 273918 116158 273952
rect 116192 273918 116226 273952
rect 116260 273918 116294 273952
rect 116328 273918 116362 273952
rect 116396 273918 116430 273952
rect 116464 273918 116498 273952
rect 116532 273918 116566 273952
rect 116600 273918 116634 273952
rect 116668 273918 116702 273952
rect 116736 273918 116770 273952
rect 116804 273918 116838 273952
rect 116872 273918 116906 273952
rect 116940 273918 116974 273952
rect 117008 273918 117042 273952
rect 117076 273918 117110 273952
rect 117144 273918 117178 273952
rect 117212 273918 117235 273952
rect 117581 273950 117604 273984
rect 117638 273950 117672 273984
rect 117706 273950 117740 273984
rect 117774 273950 117808 273984
rect 117842 273950 117876 273984
rect 117910 273950 117944 273984
rect 117978 273950 118012 273984
rect 118046 273950 118080 273984
rect 118114 273950 118148 273984
rect 118182 273950 118216 273984
rect 118250 273950 118284 273984
rect 118318 273950 118352 273984
rect 118386 273950 118420 273984
rect 118454 273950 118488 273984
rect 118522 273950 118556 273984
rect 118590 273950 118624 273984
rect 118658 273950 118681 273984
rect 117581 273938 118681 273950
rect 116135 273906 117235 273918
rect 117581 273842 118681 273854
rect 117581 273808 117604 273842
rect 117638 273808 117672 273842
rect 117706 273808 117740 273842
rect 117774 273808 117808 273842
rect 117842 273808 117876 273842
rect 117910 273808 117944 273842
rect 117978 273808 118012 273842
rect 118046 273808 118080 273842
rect 118114 273808 118148 273842
rect 118182 273808 118216 273842
rect 118250 273808 118284 273842
rect 118318 273808 118352 273842
rect 118386 273808 118420 273842
rect 118454 273808 118488 273842
rect 118522 273808 118556 273842
rect 118590 273808 118624 273842
rect 118658 273808 118681 273842
rect 116135 273786 117235 273798
rect 117581 273796 118681 273808
rect 116135 273752 116158 273786
rect 116192 273752 116226 273786
rect 116260 273752 116294 273786
rect 116328 273752 116362 273786
rect 116396 273752 116430 273786
rect 116464 273752 116498 273786
rect 116532 273752 116566 273786
rect 116600 273752 116634 273786
rect 116668 273752 116702 273786
rect 116736 273752 116770 273786
rect 116804 273752 116838 273786
rect 116872 273752 116906 273786
rect 116940 273752 116974 273786
rect 117008 273752 117042 273786
rect 117076 273752 117110 273786
rect 117144 273752 117178 273786
rect 117212 273752 117235 273786
rect 116135 273740 117235 273752
rect 117581 273624 118681 273636
rect 117581 273590 117604 273624
rect 117638 273590 117672 273624
rect 117706 273590 117740 273624
rect 117774 273590 117808 273624
rect 117842 273590 117876 273624
rect 117910 273590 117944 273624
rect 117978 273590 118012 273624
rect 118046 273590 118080 273624
rect 118114 273590 118148 273624
rect 118182 273590 118216 273624
rect 118250 273590 118284 273624
rect 118318 273590 118352 273624
rect 118386 273590 118420 273624
rect 118454 273590 118488 273624
rect 118522 273590 118556 273624
rect 118590 273590 118624 273624
rect 118658 273590 118681 273624
rect 117581 273578 118681 273590
rect 116135 273528 117235 273540
rect 116135 273494 116158 273528
rect 116192 273494 116226 273528
rect 116260 273494 116294 273528
rect 116328 273494 116362 273528
rect 116396 273494 116430 273528
rect 116464 273494 116498 273528
rect 116532 273494 116566 273528
rect 116600 273494 116634 273528
rect 116668 273494 116702 273528
rect 116736 273494 116770 273528
rect 116804 273494 116838 273528
rect 116872 273494 116906 273528
rect 116940 273494 116974 273528
rect 117008 273494 117042 273528
rect 117076 273494 117110 273528
rect 117144 273494 117178 273528
rect 117212 273494 117235 273528
rect 116135 273482 117235 273494
rect 117581 273482 118681 273494
rect 117581 273448 117604 273482
rect 117638 273448 117672 273482
rect 117706 273448 117740 273482
rect 117774 273448 117808 273482
rect 117842 273448 117876 273482
rect 117910 273448 117944 273482
rect 117978 273448 118012 273482
rect 118046 273448 118080 273482
rect 118114 273448 118148 273482
rect 118182 273448 118216 273482
rect 118250 273448 118284 273482
rect 118318 273448 118352 273482
rect 118386 273448 118420 273482
rect 118454 273448 118488 273482
rect 118522 273448 118556 273482
rect 118590 273448 118624 273482
rect 118658 273448 118681 273482
rect 117581 273436 118681 273448
rect 116105 273384 117205 273396
rect 116105 273350 116128 273384
rect 116162 273350 116196 273384
rect 116230 273350 116264 273384
rect 116298 273350 116332 273384
rect 116366 273350 116400 273384
rect 116434 273350 116468 273384
rect 116502 273350 116536 273384
rect 116570 273350 116604 273384
rect 116638 273350 116672 273384
rect 116706 273350 116740 273384
rect 116774 273350 116808 273384
rect 116842 273350 116876 273384
rect 116910 273350 116944 273384
rect 116978 273350 117012 273384
rect 117046 273350 117080 273384
rect 117114 273350 117148 273384
rect 117182 273350 117205 273384
rect 116105 273338 117205 273350
rect 117581 273264 118681 273276
rect 116105 273246 117205 273258
rect 116105 273212 116128 273246
rect 116162 273212 116196 273246
rect 116230 273212 116264 273246
rect 116298 273212 116332 273246
rect 116366 273212 116400 273246
rect 116434 273212 116468 273246
rect 116502 273212 116536 273246
rect 116570 273212 116604 273246
rect 116638 273212 116672 273246
rect 116706 273212 116740 273246
rect 116774 273212 116808 273246
rect 116842 273212 116876 273246
rect 116910 273212 116944 273246
rect 116978 273212 117012 273246
rect 117046 273212 117080 273246
rect 117114 273212 117148 273246
rect 117182 273212 117205 273246
rect 117581 273230 117604 273264
rect 117638 273230 117672 273264
rect 117706 273230 117740 273264
rect 117774 273230 117808 273264
rect 117842 273230 117876 273264
rect 117910 273230 117944 273264
rect 117978 273230 118012 273264
rect 118046 273230 118080 273264
rect 118114 273230 118148 273264
rect 118182 273230 118216 273264
rect 118250 273230 118284 273264
rect 118318 273230 118352 273264
rect 118386 273230 118420 273264
rect 118454 273230 118488 273264
rect 118522 273230 118556 273264
rect 118590 273230 118624 273264
rect 118658 273230 118681 273264
rect 117581 273218 118681 273230
rect 116105 273200 117205 273212
rect 117581 273122 118681 273134
rect 116105 273086 117205 273098
rect 116105 273052 116128 273086
rect 116162 273052 116196 273086
rect 116230 273052 116264 273086
rect 116298 273052 116332 273086
rect 116366 273052 116400 273086
rect 116434 273052 116468 273086
rect 116502 273052 116536 273086
rect 116570 273052 116604 273086
rect 116638 273052 116672 273086
rect 116706 273052 116740 273086
rect 116774 273052 116808 273086
rect 116842 273052 116876 273086
rect 116910 273052 116944 273086
rect 116978 273052 117012 273086
rect 117046 273052 117080 273086
rect 117114 273052 117148 273086
rect 117182 273052 117205 273086
rect 117581 273088 117604 273122
rect 117638 273088 117672 273122
rect 117706 273088 117740 273122
rect 117774 273088 117808 273122
rect 117842 273088 117876 273122
rect 117910 273088 117944 273122
rect 117978 273088 118012 273122
rect 118046 273088 118080 273122
rect 118114 273088 118148 273122
rect 118182 273088 118216 273122
rect 118250 273088 118284 273122
rect 118318 273088 118352 273122
rect 118386 273088 118420 273122
rect 118454 273088 118488 273122
rect 118522 273088 118556 273122
rect 118590 273088 118624 273122
rect 118658 273088 118681 273122
rect 117581 273076 118681 273088
rect 116105 273040 117205 273052
rect 116105 272948 117205 272960
rect 116105 272914 116128 272948
rect 116162 272914 116196 272948
rect 116230 272914 116264 272948
rect 116298 272914 116332 272948
rect 116366 272914 116400 272948
rect 116434 272914 116468 272948
rect 116502 272914 116536 272948
rect 116570 272914 116604 272948
rect 116638 272914 116672 272948
rect 116706 272914 116740 272948
rect 116774 272914 116808 272948
rect 116842 272914 116876 272948
rect 116910 272914 116944 272948
rect 116978 272914 117012 272948
rect 117046 272914 117080 272948
rect 117114 272914 117148 272948
rect 117182 272914 117205 272948
rect 116105 272902 117205 272914
rect 117581 272904 118681 272916
rect 117581 272870 117604 272904
rect 117638 272870 117672 272904
rect 117706 272870 117740 272904
rect 117774 272870 117808 272904
rect 117842 272870 117876 272904
rect 117910 272870 117944 272904
rect 117978 272870 118012 272904
rect 118046 272870 118080 272904
rect 118114 272870 118148 272904
rect 118182 272870 118216 272904
rect 118250 272870 118284 272904
rect 118318 272870 118352 272904
rect 118386 272870 118420 272904
rect 118454 272870 118488 272904
rect 118522 272870 118556 272904
rect 118590 272870 118624 272904
rect 118658 272870 118681 272904
rect 117581 272858 118681 272870
rect 115823 271901 115881 271924
rect 115823 271867 115835 271901
rect 115869 271867 115881 271901
rect 115823 271833 115881 271867
rect 115823 271799 115835 271833
rect 115869 271799 115881 271833
rect 115823 271765 115881 271799
rect 115823 271731 115835 271765
rect 115869 271731 115881 271765
rect 115823 271697 115881 271731
rect 115823 271663 115835 271697
rect 115869 271663 115881 271697
rect 115823 271629 115881 271663
rect 115823 271595 115835 271629
rect 115869 271595 115881 271629
rect 115823 271561 115881 271595
rect 115823 271527 115835 271561
rect 115869 271527 115881 271561
rect 115823 271493 115881 271527
rect 115823 271459 115835 271493
rect 115869 271459 115881 271493
rect 115823 271425 115881 271459
rect 115823 271391 115835 271425
rect 115869 271391 115881 271425
rect 115823 271357 115881 271391
rect 115823 271323 115835 271357
rect 115869 271323 115881 271357
rect 115823 271289 115881 271323
rect 115823 271255 115835 271289
rect 115869 271255 115881 271289
rect 115823 271221 115881 271255
rect 115823 271187 115835 271221
rect 115869 271187 115881 271221
rect 115823 271153 115881 271187
rect 115823 271119 115835 271153
rect 115869 271119 115881 271153
rect 115823 271085 115881 271119
rect 115823 271051 115835 271085
rect 115869 271051 115881 271085
rect 115823 271017 115881 271051
rect 115823 270983 115835 271017
rect 115869 270983 115881 271017
rect 115823 270949 115881 270983
rect 115823 270915 115835 270949
rect 115869 270915 115881 270949
rect 115823 270881 115881 270915
rect 115823 270847 115835 270881
rect 115869 270847 115881 270881
rect 115823 270824 115881 270847
rect 116041 271901 116099 271924
rect 116041 271867 116053 271901
rect 116087 271867 116099 271901
rect 116041 271833 116099 271867
rect 116041 271799 116053 271833
rect 116087 271799 116099 271833
rect 116041 271765 116099 271799
rect 116041 271731 116053 271765
rect 116087 271731 116099 271765
rect 116041 271697 116099 271731
rect 116041 271663 116053 271697
rect 116087 271663 116099 271697
rect 116041 271629 116099 271663
rect 116041 271595 116053 271629
rect 116087 271595 116099 271629
rect 116041 271561 116099 271595
rect 116041 271527 116053 271561
rect 116087 271527 116099 271561
rect 116041 271493 116099 271527
rect 116041 271459 116053 271493
rect 116087 271459 116099 271493
rect 116041 271425 116099 271459
rect 116041 271391 116053 271425
rect 116087 271391 116099 271425
rect 116041 271357 116099 271391
rect 116041 271323 116053 271357
rect 116087 271323 116099 271357
rect 116041 271289 116099 271323
rect 116041 271255 116053 271289
rect 116087 271255 116099 271289
rect 116041 271221 116099 271255
rect 116041 271187 116053 271221
rect 116087 271187 116099 271221
rect 116041 271153 116099 271187
rect 116041 271119 116053 271153
rect 116087 271119 116099 271153
rect 116041 271085 116099 271119
rect 116041 271051 116053 271085
rect 116087 271051 116099 271085
rect 116041 271017 116099 271051
rect 116041 270983 116053 271017
rect 116087 270983 116099 271017
rect 116041 270949 116099 270983
rect 116041 270915 116053 270949
rect 116087 270915 116099 270949
rect 116041 270881 116099 270915
rect 116041 270847 116053 270881
rect 116087 270847 116099 270881
rect 116041 270824 116099 270847
rect 116223 271901 116281 271924
rect 116223 271867 116235 271901
rect 116269 271867 116281 271901
rect 116223 271833 116281 271867
rect 116223 271799 116235 271833
rect 116269 271799 116281 271833
rect 116223 271765 116281 271799
rect 116223 271731 116235 271765
rect 116269 271731 116281 271765
rect 116223 271697 116281 271731
rect 116223 271663 116235 271697
rect 116269 271663 116281 271697
rect 116223 271629 116281 271663
rect 116223 271595 116235 271629
rect 116269 271595 116281 271629
rect 116223 271561 116281 271595
rect 116223 271527 116235 271561
rect 116269 271527 116281 271561
rect 116223 271493 116281 271527
rect 116223 271459 116235 271493
rect 116269 271459 116281 271493
rect 116223 271425 116281 271459
rect 116223 271391 116235 271425
rect 116269 271391 116281 271425
rect 116223 271357 116281 271391
rect 116223 271323 116235 271357
rect 116269 271323 116281 271357
rect 116223 271289 116281 271323
rect 116223 271255 116235 271289
rect 116269 271255 116281 271289
rect 116223 271221 116281 271255
rect 116223 271187 116235 271221
rect 116269 271187 116281 271221
rect 116223 271153 116281 271187
rect 116223 271119 116235 271153
rect 116269 271119 116281 271153
rect 116223 271085 116281 271119
rect 116223 271051 116235 271085
rect 116269 271051 116281 271085
rect 116223 271017 116281 271051
rect 116223 270983 116235 271017
rect 116269 270983 116281 271017
rect 116223 270949 116281 270983
rect 116223 270915 116235 270949
rect 116269 270915 116281 270949
rect 116223 270881 116281 270915
rect 116223 270847 116235 270881
rect 116269 270847 116281 270881
rect 116223 270824 116281 270847
rect 116441 271901 116499 271924
rect 116441 271867 116453 271901
rect 116487 271867 116499 271901
rect 116441 271833 116499 271867
rect 116441 271799 116453 271833
rect 116487 271799 116499 271833
rect 116441 271765 116499 271799
rect 116441 271731 116453 271765
rect 116487 271731 116499 271765
rect 116441 271697 116499 271731
rect 116441 271663 116453 271697
rect 116487 271663 116499 271697
rect 116441 271629 116499 271663
rect 116441 271595 116453 271629
rect 116487 271595 116499 271629
rect 116441 271561 116499 271595
rect 116441 271527 116453 271561
rect 116487 271527 116499 271561
rect 116441 271493 116499 271527
rect 116441 271459 116453 271493
rect 116487 271459 116499 271493
rect 116441 271425 116499 271459
rect 116441 271391 116453 271425
rect 116487 271391 116499 271425
rect 116441 271357 116499 271391
rect 116441 271323 116453 271357
rect 116487 271323 116499 271357
rect 116441 271289 116499 271323
rect 116441 271255 116453 271289
rect 116487 271255 116499 271289
rect 116441 271221 116499 271255
rect 116441 271187 116453 271221
rect 116487 271187 116499 271221
rect 116441 271153 116499 271187
rect 116441 271119 116453 271153
rect 116487 271119 116499 271153
rect 116441 271085 116499 271119
rect 116441 271051 116453 271085
rect 116487 271051 116499 271085
rect 116441 271017 116499 271051
rect 116441 270983 116453 271017
rect 116487 270983 116499 271017
rect 116441 270949 116499 270983
rect 116441 270915 116453 270949
rect 116487 270915 116499 270949
rect 116441 270881 116499 270915
rect 116441 270847 116453 270881
rect 116487 270847 116499 270881
rect 116441 270824 116499 270847
rect 116623 271901 116681 271924
rect 116623 271867 116635 271901
rect 116669 271867 116681 271901
rect 116623 271833 116681 271867
rect 116623 271799 116635 271833
rect 116669 271799 116681 271833
rect 116623 271765 116681 271799
rect 116623 271731 116635 271765
rect 116669 271731 116681 271765
rect 116623 271697 116681 271731
rect 116623 271663 116635 271697
rect 116669 271663 116681 271697
rect 116623 271629 116681 271663
rect 116623 271595 116635 271629
rect 116669 271595 116681 271629
rect 116623 271561 116681 271595
rect 116623 271527 116635 271561
rect 116669 271527 116681 271561
rect 116623 271493 116681 271527
rect 116623 271459 116635 271493
rect 116669 271459 116681 271493
rect 116623 271425 116681 271459
rect 116623 271391 116635 271425
rect 116669 271391 116681 271425
rect 116623 271357 116681 271391
rect 116623 271323 116635 271357
rect 116669 271323 116681 271357
rect 116623 271289 116681 271323
rect 116623 271255 116635 271289
rect 116669 271255 116681 271289
rect 116623 271221 116681 271255
rect 116623 271187 116635 271221
rect 116669 271187 116681 271221
rect 116623 271153 116681 271187
rect 116623 271119 116635 271153
rect 116669 271119 116681 271153
rect 116623 271085 116681 271119
rect 116623 271051 116635 271085
rect 116669 271051 116681 271085
rect 116623 271017 116681 271051
rect 116623 270983 116635 271017
rect 116669 270983 116681 271017
rect 116623 270949 116681 270983
rect 116623 270915 116635 270949
rect 116669 270915 116681 270949
rect 116623 270881 116681 270915
rect 116623 270847 116635 270881
rect 116669 270847 116681 270881
rect 116623 270824 116681 270847
rect 116841 271901 116899 271924
rect 116841 271867 116853 271901
rect 116887 271867 116899 271901
rect 116841 271833 116899 271867
rect 116841 271799 116853 271833
rect 116887 271799 116899 271833
rect 116841 271765 116899 271799
rect 116841 271731 116853 271765
rect 116887 271731 116899 271765
rect 116841 271697 116899 271731
rect 116841 271663 116853 271697
rect 116887 271663 116899 271697
rect 116841 271629 116899 271663
rect 116841 271595 116853 271629
rect 116887 271595 116899 271629
rect 116841 271561 116899 271595
rect 116841 271527 116853 271561
rect 116887 271527 116899 271561
rect 116841 271493 116899 271527
rect 116841 271459 116853 271493
rect 116887 271459 116899 271493
rect 116841 271425 116899 271459
rect 116841 271391 116853 271425
rect 116887 271391 116899 271425
rect 116841 271357 116899 271391
rect 116841 271323 116853 271357
rect 116887 271323 116899 271357
rect 116841 271289 116899 271323
rect 116841 271255 116853 271289
rect 116887 271255 116899 271289
rect 116841 271221 116899 271255
rect 116841 271187 116853 271221
rect 116887 271187 116899 271221
rect 116841 271153 116899 271187
rect 116841 271119 116853 271153
rect 116887 271119 116899 271153
rect 116841 271085 116899 271119
rect 116841 271051 116853 271085
rect 116887 271051 116899 271085
rect 116841 271017 116899 271051
rect 116841 270983 116853 271017
rect 116887 270983 116899 271017
rect 116841 270949 116899 270983
rect 116841 270915 116853 270949
rect 116887 270915 116899 270949
rect 116841 270881 116899 270915
rect 116841 270847 116853 270881
rect 116887 270847 116899 270881
rect 116841 270824 116899 270847
rect 117023 271901 117081 271924
rect 117023 271867 117035 271901
rect 117069 271867 117081 271901
rect 117023 271833 117081 271867
rect 117023 271799 117035 271833
rect 117069 271799 117081 271833
rect 117023 271765 117081 271799
rect 117023 271731 117035 271765
rect 117069 271731 117081 271765
rect 117023 271697 117081 271731
rect 117023 271663 117035 271697
rect 117069 271663 117081 271697
rect 117023 271629 117081 271663
rect 117023 271595 117035 271629
rect 117069 271595 117081 271629
rect 117023 271561 117081 271595
rect 117023 271527 117035 271561
rect 117069 271527 117081 271561
rect 117023 271493 117081 271527
rect 117023 271459 117035 271493
rect 117069 271459 117081 271493
rect 117023 271425 117081 271459
rect 117023 271391 117035 271425
rect 117069 271391 117081 271425
rect 117023 271357 117081 271391
rect 117023 271323 117035 271357
rect 117069 271323 117081 271357
rect 117023 271289 117081 271323
rect 117023 271255 117035 271289
rect 117069 271255 117081 271289
rect 117023 271221 117081 271255
rect 117023 271187 117035 271221
rect 117069 271187 117081 271221
rect 117023 271153 117081 271187
rect 117023 271119 117035 271153
rect 117069 271119 117081 271153
rect 117023 271085 117081 271119
rect 117023 271051 117035 271085
rect 117069 271051 117081 271085
rect 117023 271017 117081 271051
rect 117023 270983 117035 271017
rect 117069 270983 117081 271017
rect 117023 270949 117081 270983
rect 117023 270915 117035 270949
rect 117069 270915 117081 270949
rect 117023 270881 117081 270915
rect 117023 270847 117035 270881
rect 117069 270847 117081 270881
rect 117023 270824 117081 270847
rect 117241 271901 117299 271924
rect 117241 271867 117253 271901
rect 117287 271867 117299 271901
rect 117241 271833 117299 271867
rect 117241 271799 117253 271833
rect 117287 271799 117299 271833
rect 117241 271765 117299 271799
rect 117241 271731 117253 271765
rect 117287 271731 117299 271765
rect 117241 271697 117299 271731
rect 117241 271663 117253 271697
rect 117287 271663 117299 271697
rect 117241 271629 117299 271663
rect 117241 271595 117253 271629
rect 117287 271595 117299 271629
rect 117241 271561 117299 271595
rect 117241 271527 117253 271561
rect 117287 271527 117299 271561
rect 117241 271493 117299 271527
rect 117241 271459 117253 271493
rect 117287 271459 117299 271493
rect 117241 271425 117299 271459
rect 117241 271391 117253 271425
rect 117287 271391 117299 271425
rect 117241 271357 117299 271391
rect 117241 271323 117253 271357
rect 117287 271323 117299 271357
rect 117241 271289 117299 271323
rect 117241 271255 117253 271289
rect 117287 271255 117299 271289
rect 117241 271221 117299 271255
rect 117241 271187 117253 271221
rect 117287 271187 117299 271221
rect 117241 271153 117299 271187
rect 117241 271119 117253 271153
rect 117287 271119 117299 271153
rect 117241 271085 117299 271119
rect 117241 271051 117253 271085
rect 117287 271051 117299 271085
rect 117241 271017 117299 271051
rect 117241 270983 117253 271017
rect 117287 270983 117299 271017
rect 117241 270949 117299 270983
rect 117241 270915 117253 270949
rect 117287 270915 117299 270949
rect 117241 270881 117299 270915
rect 117241 270847 117253 270881
rect 117287 270847 117299 270881
rect 117241 270824 117299 270847
rect 117423 271901 117481 271924
rect 117423 271867 117435 271901
rect 117469 271867 117481 271901
rect 117423 271833 117481 271867
rect 117423 271799 117435 271833
rect 117469 271799 117481 271833
rect 117423 271765 117481 271799
rect 117423 271731 117435 271765
rect 117469 271731 117481 271765
rect 117423 271697 117481 271731
rect 117423 271663 117435 271697
rect 117469 271663 117481 271697
rect 117423 271629 117481 271663
rect 117423 271595 117435 271629
rect 117469 271595 117481 271629
rect 117423 271561 117481 271595
rect 117423 271527 117435 271561
rect 117469 271527 117481 271561
rect 117423 271493 117481 271527
rect 117423 271459 117435 271493
rect 117469 271459 117481 271493
rect 117423 271425 117481 271459
rect 117423 271391 117435 271425
rect 117469 271391 117481 271425
rect 117423 271357 117481 271391
rect 117423 271323 117435 271357
rect 117469 271323 117481 271357
rect 117423 271289 117481 271323
rect 117423 271255 117435 271289
rect 117469 271255 117481 271289
rect 117423 271221 117481 271255
rect 117423 271187 117435 271221
rect 117469 271187 117481 271221
rect 117423 271153 117481 271187
rect 117423 271119 117435 271153
rect 117469 271119 117481 271153
rect 117423 271085 117481 271119
rect 117423 271051 117435 271085
rect 117469 271051 117481 271085
rect 117423 271017 117481 271051
rect 117423 270983 117435 271017
rect 117469 270983 117481 271017
rect 117423 270949 117481 270983
rect 117423 270915 117435 270949
rect 117469 270915 117481 270949
rect 117423 270881 117481 270915
rect 117423 270847 117435 270881
rect 117469 270847 117481 270881
rect 117423 270824 117481 270847
rect 117641 271901 117699 271924
rect 117641 271867 117653 271901
rect 117687 271867 117699 271901
rect 117641 271833 117699 271867
rect 117641 271799 117653 271833
rect 117687 271799 117699 271833
rect 117641 271765 117699 271799
rect 117641 271731 117653 271765
rect 117687 271731 117699 271765
rect 117641 271697 117699 271731
rect 117641 271663 117653 271697
rect 117687 271663 117699 271697
rect 117641 271629 117699 271663
rect 117641 271595 117653 271629
rect 117687 271595 117699 271629
rect 117641 271561 117699 271595
rect 117641 271527 117653 271561
rect 117687 271527 117699 271561
rect 117641 271493 117699 271527
rect 117641 271459 117653 271493
rect 117687 271459 117699 271493
rect 117641 271425 117699 271459
rect 117641 271391 117653 271425
rect 117687 271391 117699 271425
rect 117641 271357 117699 271391
rect 117641 271323 117653 271357
rect 117687 271323 117699 271357
rect 117641 271289 117699 271323
rect 117641 271255 117653 271289
rect 117687 271255 117699 271289
rect 117641 271221 117699 271255
rect 117641 271187 117653 271221
rect 117687 271187 117699 271221
rect 117641 271153 117699 271187
rect 117641 271119 117653 271153
rect 117687 271119 117699 271153
rect 117641 271085 117699 271119
rect 117641 271051 117653 271085
rect 117687 271051 117699 271085
rect 117641 271017 117699 271051
rect 117641 270983 117653 271017
rect 117687 270983 117699 271017
rect 117641 270949 117699 270983
rect 117641 270915 117653 270949
rect 117687 270915 117699 270949
rect 117641 270881 117699 270915
rect 117641 270847 117653 270881
rect 117687 270847 117699 270881
rect 117641 270824 117699 270847
rect 117823 271901 117881 271924
rect 117823 271867 117835 271901
rect 117869 271867 117881 271901
rect 117823 271833 117881 271867
rect 117823 271799 117835 271833
rect 117869 271799 117881 271833
rect 117823 271765 117881 271799
rect 117823 271731 117835 271765
rect 117869 271731 117881 271765
rect 117823 271697 117881 271731
rect 117823 271663 117835 271697
rect 117869 271663 117881 271697
rect 117823 271629 117881 271663
rect 117823 271595 117835 271629
rect 117869 271595 117881 271629
rect 117823 271561 117881 271595
rect 117823 271527 117835 271561
rect 117869 271527 117881 271561
rect 117823 271493 117881 271527
rect 117823 271459 117835 271493
rect 117869 271459 117881 271493
rect 117823 271425 117881 271459
rect 117823 271391 117835 271425
rect 117869 271391 117881 271425
rect 117823 271357 117881 271391
rect 117823 271323 117835 271357
rect 117869 271323 117881 271357
rect 117823 271289 117881 271323
rect 117823 271255 117835 271289
rect 117869 271255 117881 271289
rect 117823 271221 117881 271255
rect 117823 271187 117835 271221
rect 117869 271187 117881 271221
rect 117823 271153 117881 271187
rect 117823 271119 117835 271153
rect 117869 271119 117881 271153
rect 117823 271085 117881 271119
rect 117823 271051 117835 271085
rect 117869 271051 117881 271085
rect 117823 271017 117881 271051
rect 117823 270983 117835 271017
rect 117869 270983 117881 271017
rect 117823 270949 117881 270983
rect 117823 270915 117835 270949
rect 117869 270915 117881 270949
rect 117823 270881 117881 270915
rect 117823 270847 117835 270881
rect 117869 270847 117881 270881
rect 117823 270824 117881 270847
rect 118041 271901 118099 271924
rect 118041 271867 118053 271901
rect 118087 271867 118099 271901
rect 118041 271833 118099 271867
rect 118041 271799 118053 271833
rect 118087 271799 118099 271833
rect 118041 271765 118099 271799
rect 118041 271731 118053 271765
rect 118087 271731 118099 271765
rect 118041 271697 118099 271731
rect 118041 271663 118053 271697
rect 118087 271663 118099 271697
rect 118041 271629 118099 271663
rect 118041 271595 118053 271629
rect 118087 271595 118099 271629
rect 118041 271561 118099 271595
rect 118041 271527 118053 271561
rect 118087 271527 118099 271561
rect 118041 271493 118099 271527
rect 118041 271459 118053 271493
rect 118087 271459 118099 271493
rect 118041 271425 118099 271459
rect 118041 271391 118053 271425
rect 118087 271391 118099 271425
rect 118041 271357 118099 271391
rect 118041 271323 118053 271357
rect 118087 271323 118099 271357
rect 118041 271289 118099 271323
rect 118041 271255 118053 271289
rect 118087 271255 118099 271289
rect 118041 271221 118099 271255
rect 118041 271187 118053 271221
rect 118087 271187 118099 271221
rect 118041 271153 118099 271187
rect 118041 271119 118053 271153
rect 118087 271119 118099 271153
rect 118041 271085 118099 271119
rect 118041 271051 118053 271085
rect 118087 271051 118099 271085
rect 118041 271017 118099 271051
rect 118041 270983 118053 271017
rect 118087 270983 118099 271017
rect 118041 270949 118099 270983
rect 118041 270915 118053 270949
rect 118087 270915 118099 270949
rect 118041 270881 118099 270915
rect 118041 270847 118053 270881
rect 118087 270847 118099 270881
rect 118041 270824 118099 270847
rect 118223 271901 118281 271924
rect 118223 271867 118235 271901
rect 118269 271867 118281 271901
rect 118223 271833 118281 271867
rect 118223 271799 118235 271833
rect 118269 271799 118281 271833
rect 118223 271765 118281 271799
rect 118223 271731 118235 271765
rect 118269 271731 118281 271765
rect 118223 271697 118281 271731
rect 118223 271663 118235 271697
rect 118269 271663 118281 271697
rect 118223 271629 118281 271663
rect 118223 271595 118235 271629
rect 118269 271595 118281 271629
rect 118223 271561 118281 271595
rect 118223 271527 118235 271561
rect 118269 271527 118281 271561
rect 118223 271493 118281 271527
rect 118223 271459 118235 271493
rect 118269 271459 118281 271493
rect 118223 271425 118281 271459
rect 118223 271391 118235 271425
rect 118269 271391 118281 271425
rect 118223 271357 118281 271391
rect 118223 271323 118235 271357
rect 118269 271323 118281 271357
rect 118223 271289 118281 271323
rect 118223 271255 118235 271289
rect 118269 271255 118281 271289
rect 118223 271221 118281 271255
rect 118223 271187 118235 271221
rect 118269 271187 118281 271221
rect 118223 271153 118281 271187
rect 118223 271119 118235 271153
rect 118269 271119 118281 271153
rect 118223 271085 118281 271119
rect 118223 271051 118235 271085
rect 118269 271051 118281 271085
rect 118223 271017 118281 271051
rect 118223 270983 118235 271017
rect 118269 270983 118281 271017
rect 118223 270949 118281 270983
rect 118223 270915 118235 270949
rect 118269 270915 118281 270949
rect 118223 270881 118281 270915
rect 118223 270847 118235 270881
rect 118269 270847 118281 270881
rect 118223 270824 118281 270847
rect 118441 271901 118499 271924
rect 118441 271867 118453 271901
rect 118487 271867 118499 271901
rect 118441 271833 118499 271867
rect 118441 271799 118453 271833
rect 118487 271799 118499 271833
rect 118441 271765 118499 271799
rect 118441 271731 118453 271765
rect 118487 271731 118499 271765
rect 118441 271697 118499 271731
rect 118441 271663 118453 271697
rect 118487 271663 118499 271697
rect 118441 271629 118499 271663
rect 118441 271595 118453 271629
rect 118487 271595 118499 271629
rect 118441 271561 118499 271595
rect 118441 271527 118453 271561
rect 118487 271527 118499 271561
rect 118441 271493 118499 271527
rect 118441 271459 118453 271493
rect 118487 271459 118499 271493
rect 118441 271425 118499 271459
rect 118441 271391 118453 271425
rect 118487 271391 118499 271425
rect 118441 271357 118499 271391
rect 118441 271323 118453 271357
rect 118487 271323 118499 271357
rect 118441 271289 118499 271323
rect 118441 271255 118453 271289
rect 118487 271255 118499 271289
rect 118441 271221 118499 271255
rect 118441 271187 118453 271221
rect 118487 271187 118499 271221
rect 118441 271153 118499 271187
rect 118441 271119 118453 271153
rect 118487 271119 118499 271153
rect 118441 271085 118499 271119
rect 118441 271051 118453 271085
rect 118487 271051 118499 271085
rect 118441 271017 118499 271051
rect 118441 270983 118453 271017
rect 118487 270983 118499 271017
rect 118441 270949 118499 270983
rect 118441 270915 118453 270949
rect 118487 270915 118499 270949
rect 118441 270881 118499 270915
rect 118441 270847 118453 270881
rect 118487 270847 118499 270881
rect 118441 270824 118499 270847
rect 118623 271901 118681 271924
rect 118623 271867 118635 271901
rect 118669 271867 118681 271901
rect 118623 271833 118681 271867
rect 118623 271799 118635 271833
rect 118669 271799 118681 271833
rect 118623 271765 118681 271799
rect 118623 271731 118635 271765
rect 118669 271731 118681 271765
rect 118623 271697 118681 271731
rect 118623 271663 118635 271697
rect 118669 271663 118681 271697
rect 118623 271629 118681 271663
rect 118623 271595 118635 271629
rect 118669 271595 118681 271629
rect 118623 271561 118681 271595
rect 118623 271527 118635 271561
rect 118669 271527 118681 271561
rect 118623 271493 118681 271527
rect 118623 271459 118635 271493
rect 118669 271459 118681 271493
rect 118623 271425 118681 271459
rect 118623 271391 118635 271425
rect 118669 271391 118681 271425
rect 118623 271357 118681 271391
rect 118623 271323 118635 271357
rect 118669 271323 118681 271357
rect 118623 271289 118681 271323
rect 118623 271255 118635 271289
rect 118669 271255 118681 271289
rect 118623 271221 118681 271255
rect 118623 271187 118635 271221
rect 118669 271187 118681 271221
rect 118623 271153 118681 271187
rect 118623 271119 118635 271153
rect 118669 271119 118681 271153
rect 118623 271085 118681 271119
rect 118623 271051 118635 271085
rect 118669 271051 118681 271085
rect 118623 271017 118681 271051
rect 118623 270983 118635 271017
rect 118669 270983 118681 271017
rect 118623 270949 118681 270983
rect 118623 270915 118635 270949
rect 118669 270915 118681 270949
rect 118623 270881 118681 270915
rect 118623 270847 118635 270881
rect 118669 270847 118681 270881
rect 118623 270824 118681 270847
rect 118841 271901 118899 271924
rect 118841 271867 118853 271901
rect 118887 271867 118899 271901
rect 118841 271833 118899 271867
rect 118841 271799 118853 271833
rect 118887 271799 118899 271833
rect 118841 271765 118899 271799
rect 118841 271731 118853 271765
rect 118887 271731 118899 271765
rect 118841 271697 118899 271731
rect 118841 271663 118853 271697
rect 118887 271663 118899 271697
rect 118841 271629 118899 271663
rect 118841 271595 118853 271629
rect 118887 271595 118899 271629
rect 118841 271561 118899 271595
rect 118841 271527 118853 271561
rect 118887 271527 118899 271561
rect 118841 271493 118899 271527
rect 118841 271459 118853 271493
rect 118887 271459 118899 271493
rect 118841 271425 118899 271459
rect 118841 271391 118853 271425
rect 118887 271391 118899 271425
rect 118841 271357 118899 271391
rect 118841 271323 118853 271357
rect 118887 271323 118899 271357
rect 118841 271289 118899 271323
rect 118841 271255 118853 271289
rect 118887 271255 118899 271289
rect 118841 271221 118899 271255
rect 118841 271187 118853 271221
rect 118887 271187 118899 271221
rect 118841 271153 118899 271187
rect 118841 271119 118853 271153
rect 118887 271119 118899 271153
rect 118841 271085 118899 271119
rect 118841 271051 118853 271085
rect 118887 271051 118899 271085
rect 118841 271017 118899 271051
rect 118841 270983 118853 271017
rect 118887 270983 118899 271017
rect 118841 270949 118899 270983
rect 118841 270915 118853 270949
rect 118887 270915 118899 270949
rect 118841 270881 118899 270915
rect 118841 270847 118853 270881
rect 118887 270847 118899 270881
rect 118841 270824 118899 270847
rect 112502 270201 112560 270224
rect 112502 270167 112514 270201
rect 112548 270167 112560 270201
rect 112502 270133 112560 270167
rect 112502 270099 112514 270133
rect 112548 270099 112560 270133
rect 112502 270065 112560 270099
rect 112502 270031 112514 270065
rect 112548 270031 112560 270065
rect 112502 269997 112560 270031
rect 112502 269963 112514 269997
rect 112548 269963 112560 269997
rect 112502 269929 112560 269963
rect 112502 269895 112514 269929
rect 112548 269895 112560 269929
rect 112502 269861 112560 269895
rect 112502 269827 112514 269861
rect 112548 269827 112560 269861
rect 112502 269793 112560 269827
rect 112502 269759 112514 269793
rect 112548 269759 112560 269793
rect 112502 269725 112560 269759
rect 112502 269691 112514 269725
rect 112548 269691 112560 269725
rect 112502 269657 112560 269691
rect 112502 269623 112514 269657
rect 112548 269623 112560 269657
rect 112502 269589 112560 269623
rect 112502 269555 112514 269589
rect 112548 269555 112560 269589
rect 112502 269521 112560 269555
rect 112502 269487 112514 269521
rect 112548 269487 112560 269521
rect 112502 269453 112560 269487
rect 112502 269419 112514 269453
rect 112548 269419 112560 269453
rect 112502 269385 112560 269419
rect 112502 269351 112514 269385
rect 112548 269351 112560 269385
rect 112502 269317 112560 269351
rect 112502 269283 112514 269317
rect 112548 269283 112560 269317
rect 112502 269249 112560 269283
rect 112502 269215 112514 269249
rect 112548 269215 112560 269249
rect 112502 269181 112560 269215
rect 112502 269147 112514 269181
rect 112548 269147 112560 269181
rect 112502 269124 112560 269147
rect 112720 270201 112778 270224
rect 112720 270167 112732 270201
rect 112766 270167 112778 270201
rect 112720 270133 112778 270167
rect 112720 270099 112732 270133
rect 112766 270099 112778 270133
rect 112720 270065 112778 270099
rect 112720 270031 112732 270065
rect 112766 270031 112778 270065
rect 112720 269997 112778 270031
rect 112720 269963 112732 269997
rect 112766 269963 112778 269997
rect 112720 269929 112778 269963
rect 112720 269895 112732 269929
rect 112766 269895 112778 269929
rect 112720 269861 112778 269895
rect 112720 269827 112732 269861
rect 112766 269827 112778 269861
rect 112720 269793 112778 269827
rect 112720 269759 112732 269793
rect 112766 269759 112778 269793
rect 112720 269725 112778 269759
rect 112720 269691 112732 269725
rect 112766 269691 112778 269725
rect 112720 269657 112778 269691
rect 112720 269623 112732 269657
rect 112766 269623 112778 269657
rect 112720 269589 112778 269623
rect 112720 269555 112732 269589
rect 112766 269555 112778 269589
rect 112720 269521 112778 269555
rect 112720 269487 112732 269521
rect 112766 269487 112778 269521
rect 112720 269453 112778 269487
rect 112720 269419 112732 269453
rect 112766 269419 112778 269453
rect 112720 269385 112778 269419
rect 112720 269351 112732 269385
rect 112766 269351 112778 269385
rect 112720 269317 112778 269351
rect 112720 269283 112732 269317
rect 112766 269283 112778 269317
rect 112720 269249 112778 269283
rect 112720 269215 112732 269249
rect 112766 269215 112778 269249
rect 112720 269181 112778 269215
rect 112720 269147 112732 269181
rect 112766 269147 112778 269181
rect 112720 269124 112778 269147
rect 112902 270201 112960 270224
rect 112902 270167 112914 270201
rect 112948 270167 112960 270201
rect 112902 270133 112960 270167
rect 112902 270099 112914 270133
rect 112948 270099 112960 270133
rect 112902 270065 112960 270099
rect 112902 270031 112914 270065
rect 112948 270031 112960 270065
rect 112902 269997 112960 270031
rect 112902 269963 112914 269997
rect 112948 269963 112960 269997
rect 112902 269929 112960 269963
rect 112902 269895 112914 269929
rect 112948 269895 112960 269929
rect 112902 269861 112960 269895
rect 112902 269827 112914 269861
rect 112948 269827 112960 269861
rect 112902 269793 112960 269827
rect 112902 269759 112914 269793
rect 112948 269759 112960 269793
rect 112902 269725 112960 269759
rect 112902 269691 112914 269725
rect 112948 269691 112960 269725
rect 112902 269657 112960 269691
rect 112902 269623 112914 269657
rect 112948 269623 112960 269657
rect 112902 269589 112960 269623
rect 112902 269555 112914 269589
rect 112948 269555 112960 269589
rect 112902 269521 112960 269555
rect 112902 269487 112914 269521
rect 112948 269487 112960 269521
rect 112902 269453 112960 269487
rect 112902 269419 112914 269453
rect 112948 269419 112960 269453
rect 112902 269385 112960 269419
rect 112902 269351 112914 269385
rect 112948 269351 112960 269385
rect 112902 269317 112960 269351
rect 112902 269283 112914 269317
rect 112948 269283 112960 269317
rect 112902 269249 112960 269283
rect 112902 269215 112914 269249
rect 112948 269215 112960 269249
rect 112902 269181 112960 269215
rect 112902 269147 112914 269181
rect 112948 269147 112960 269181
rect 112902 269124 112960 269147
rect 113120 270201 113178 270224
rect 113120 270167 113132 270201
rect 113166 270167 113178 270201
rect 113120 270133 113178 270167
rect 113120 270099 113132 270133
rect 113166 270099 113178 270133
rect 113120 270065 113178 270099
rect 113120 270031 113132 270065
rect 113166 270031 113178 270065
rect 113120 269997 113178 270031
rect 113120 269963 113132 269997
rect 113166 269963 113178 269997
rect 113120 269929 113178 269963
rect 113120 269895 113132 269929
rect 113166 269895 113178 269929
rect 113120 269861 113178 269895
rect 113120 269827 113132 269861
rect 113166 269827 113178 269861
rect 113120 269793 113178 269827
rect 113120 269759 113132 269793
rect 113166 269759 113178 269793
rect 113120 269725 113178 269759
rect 113120 269691 113132 269725
rect 113166 269691 113178 269725
rect 113120 269657 113178 269691
rect 113120 269623 113132 269657
rect 113166 269623 113178 269657
rect 113120 269589 113178 269623
rect 113120 269555 113132 269589
rect 113166 269555 113178 269589
rect 113120 269521 113178 269555
rect 113120 269487 113132 269521
rect 113166 269487 113178 269521
rect 113120 269453 113178 269487
rect 113120 269419 113132 269453
rect 113166 269419 113178 269453
rect 113120 269385 113178 269419
rect 113120 269351 113132 269385
rect 113166 269351 113178 269385
rect 113120 269317 113178 269351
rect 113120 269283 113132 269317
rect 113166 269283 113178 269317
rect 113120 269249 113178 269283
rect 113120 269215 113132 269249
rect 113166 269215 113178 269249
rect 113120 269181 113178 269215
rect 113120 269147 113132 269181
rect 113166 269147 113178 269181
rect 113120 269124 113178 269147
rect 113302 270201 113360 270224
rect 113302 270167 113314 270201
rect 113348 270167 113360 270201
rect 113302 270133 113360 270167
rect 113302 270099 113314 270133
rect 113348 270099 113360 270133
rect 113302 270065 113360 270099
rect 113302 270031 113314 270065
rect 113348 270031 113360 270065
rect 113302 269997 113360 270031
rect 113302 269963 113314 269997
rect 113348 269963 113360 269997
rect 113302 269929 113360 269963
rect 113302 269895 113314 269929
rect 113348 269895 113360 269929
rect 113302 269861 113360 269895
rect 113302 269827 113314 269861
rect 113348 269827 113360 269861
rect 113302 269793 113360 269827
rect 113302 269759 113314 269793
rect 113348 269759 113360 269793
rect 113302 269725 113360 269759
rect 113302 269691 113314 269725
rect 113348 269691 113360 269725
rect 113302 269657 113360 269691
rect 113302 269623 113314 269657
rect 113348 269623 113360 269657
rect 113302 269589 113360 269623
rect 113302 269555 113314 269589
rect 113348 269555 113360 269589
rect 113302 269521 113360 269555
rect 113302 269487 113314 269521
rect 113348 269487 113360 269521
rect 113302 269453 113360 269487
rect 113302 269419 113314 269453
rect 113348 269419 113360 269453
rect 113302 269385 113360 269419
rect 113302 269351 113314 269385
rect 113348 269351 113360 269385
rect 113302 269317 113360 269351
rect 113302 269283 113314 269317
rect 113348 269283 113360 269317
rect 113302 269249 113360 269283
rect 113302 269215 113314 269249
rect 113348 269215 113360 269249
rect 113302 269181 113360 269215
rect 113302 269147 113314 269181
rect 113348 269147 113360 269181
rect 113302 269124 113360 269147
rect 113520 270201 113578 270224
rect 113520 270167 113532 270201
rect 113566 270167 113578 270201
rect 113520 270133 113578 270167
rect 113520 270099 113532 270133
rect 113566 270099 113578 270133
rect 113520 270065 113578 270099
rect 113520 270031 113532 270065
rect 113566 270031 113578 270065
rect 113520 269997 113578 270031
rect 113520 269963 113532 269997
rect 113566 269963 113578 269997
rect 113520 269929 113578 269963
rect 113520 269895 113532 269929
rect 113566 269895 113578 269929
rect 113520 269861 113578 269895
rect 113520 269827 113532 269861
rect 113566 269827 113578 269861
rect 113520 269793 113578 269827
rect 113520 269759 113532 269793
rect 113566 269759 113578 269793
rect 113520 269725 113578 269759
rect 113520 269691 113532 269725
rect 113566 269691 113578 269725
rect 113520 269657 113578 269691
rect 113520 269623 113532 269657
rect 113566 269623 113578 269657
rect 113520 269589 113578 269623
rect 113520 269555 113532 269589
rect 113566 269555 113578 269589
rect 113520 269521 113578 269555
rect 113520 269487 113532 269521
rect 113566 269487 113578 269521
rect 113520 269453 113578 269487
rect 113520 269419 113532 269453
rect 113566 269419 113578 269453
rect 113520 269385 113578 269419
rect 113520 269351 113532 269385
rect 113566 269351 113578 269385
rect 113520 269317 113578 269351
rect 113520 269283 113532 269317
rect 113566 269283 113578 269317
rect 113520 269249 113578 269283
rect 113520 269215 113532 269249
rect 113566 269215 113578 269249
rect 113520 269181 113578 269215
rect 113520 269147 113532 269181
rect 113566 269147 113578 269181
rect 113520 269124 113578 269147
rect 113702 270201 113760 270224
rect 113702 270167 113714 270201
rect 113748 270167 113760 270201
rect 113702 270133 113760 270167
rect 113702 270099 113714 270133
rect 113748 270099 113760 270133
rect 113702 270065 113760 270099
rect 113702 270031 113714 270065
rect 113748 270031 113760 270065
rect 113702 269997 113760 270031
rect 113702 269963 113714 269997
rect 113748 269963 113760 269997
rect 113702 269929 113760 269963
rect 113702 269895 113714 269929
rect 113748 269895 113760 269929
rect 113702 269861 113760 269895
rect 113702 269827 113714 269861
rect 113748 269827 113760 269861
rect 113702 269793 113760 269827
rect 113702 269759 113714 269793
rect 113748 269759 113760 269793
rect 113702 269725 113760 269759
rect 113702 269691 113714 269725
rect 113748 269691 113760 269725
rect 113702 269657 113760 269691
rect 113702 269623 113714 269657
rect 113748 269623 113760 269657
rect 113702 269589 113760 269623
rect 113702 269555 113714 269589
rect 113748 269555 113760 269589
rect 113702 269521 113760 269555
rect 113702 269487 113714 269521
rect 113748 269487 113760 269521
rect 113702 269453 113760 269487
rect 113702 269419 113714 269453
rect 113748 269419 113760 269453
rect 113702 269385 113760 269419
rect 113702 269351 113714 269385
rect 113748 269351 113760 269385
rect 113702 269317 113760 269351
rect 113702 269283 113714 269317
rect 113748 269283 113760 269317
rect 113702 269249 113760 269283
rect 113702 269215 113714 269249
rect 113748 269215 113760 269249
rect 113702 269181 113760 269215
rect 113702 269147 113714 269181
rect 113748 269147 113760 269181
rect 113702 269124 113760 269147
rect 113920 270201 113978 270224
rect 113920 270167 113932 270201
rect 113966 270167 113978 270201
rect 113920 270133 113978 270167
rect 113920 270099 113932 270133
rect 113966 270099 113978 270133
rect 113920 270065 113978 270099
rect 113920 270031 113932 270065
rect 113966 270031 113978 270065
rect 113920 269997 113978 270031
rect 113920 269963 113932 269997
rect 113966 269963 113978 269997
rect 113920 269929 113978 269963
rect 113920 269895 113932 269929
rect 113966 269895 113978 269929
rect 113920 269861 113978 269895
rect 113920 269827 113932 269861
rect 113966 269827 113978 269861
rect 113920 269793 113978 269827
rect 113920 269759 113932 269793
rect 113966 269759 113978 269793
rect 113920 269725 113978 269759
rect 113920 269691 113932 269725
rect 113966 269691 113978 269725
rect 113920 269657 113978 269691
rect 113920 269623 113932 269657
rect 113966 269623 113978 269657
rect 113920 269589 113978 269623
rect 113920 269555 113932 269589
rect 113966 269555 113978 269589
rect 113920 269521 113978 269555
rect 113920 269487 113932 269521
rect 113966 269487 113978 269521
rect 113920 269453 113978 269487
rect 113920 269419 113932 269453
rect 113966 269419 113978 269453
rect 113920 269385 113978 269419
rect 113920 269351 113932 269385
rect 113966 269351 113978 269385
rect 113920 269317 113978 269351
rect 113920 269283 113932 269317
rect 113966 269283 113978 269317
rect 113920 269249 113978 269283
rect 113920 269215 113932 269249
rect 113966 269215 113978 269249
rect 113920 269181 113978 269215
rect 113920 269147 113932 269181
rect 113966 269147 113978 269181
rect 113920 269124 113978 269147
rect 114102 270201 114160 270224
rect 114102 270167 114114 270201
rect 114148 270167 114160 270201
rect 114102 270133 114160 270167
rect 114102 270099 114114 270133
rect 114148 270099 114160 270133
rect 114102 270065 114160 270099
rect 114102 270031 114114 270065
rect 114148 270031 114160 270065
rect 114102 269997 114160 270031
rect 114102 269963 114114 269997
rect 114148 269963 114160 269997
rect 114102 269929 114160 269963
rect 114102 269895 114114 269929
rect 114148 269895 114160 269929
rect 114102 269861 114160 269895
rect 114102 269827 114114 269861
rect 114148 269827 114160 269861
rect 114102 269793 114160 269827
rect 114102 269759 114114 269793
rect 114148 269759 114160 269793
rect 114102 269725 114160 269759
rect 114102 269691 114114 269725
rect 114148 269691 114160 269725
rect 114102 269657 114160 269691
rect 114102 269623 114114 269657
rect 114148 269623 114160 269657
rect 114102 269589 114160 269623
rect 114102 269555 114114 269589
rect 114148 269555 114160 269589
rect 114102 269521 114160 269555
rect 114102 269487 114114 269521
rect 114148 269487 114160 269521
rect 114102 269453 114160 269487
rect 114102 269419 114114 269453
rect 114148 269419 114160 269453
rect 114102 269385 114160 269419
rect 114102 269351 114114 269385
rect 114148 269351 114160 269385
rect 114102 269317 114160 269351
rect 114102 269283 114114 269317
rect 114148 269283 114160 269317
rect 114102 269249 114160 269283
rect 114102 269215 114114 269249
rect 114148 269215 114160 269249
rect 114102 269181 114160 269215
rect 114102 269147 114114 269181
rect 114148 269147 114160 269181
rect 114102 269124 114160 269147
rect 114320 270201 114378 270224
rect 114320 270167 114332 270201
rect 114366 270167 114378 270201
rect 114320 270133 114378 270167
rect 114320 270099 114332 270133
rect 114366 270099 114378 270133
rect 114320 270065 114378 270099
rect 114320 270031 114332 270065
rect 114366 270031 114378 270065
rect 114320 269997 114378 270031
rect 114320 269963 114332 269997
rect 114366 269963 114378 269997
rect 114320 269929 114378 269963
rect 114320 269895 114332 269929
rect 114366 269895 114378 269929
rect 114320 269861 114378 269895
rect 114320 269827 114332 269861
rect 114366 269827 114378 269861
rect 114320 269793 114378 269827
rect 114320 269759 114332 269793
rect 114366 269759 114378 269793
rect 114320 269725 114378 269759
rect 114320 269691 114332 269725
rect 114366 269691 114378 269725
rect 114320 269657 114378 269691
rect 114320 269623 114332 269657
rect 114366 269623 114378 269657
rect 114320 269589 114378 269623
rect 114320 269555 114332 269589
rect 114366 269555 114378 269589
rect 114320 269521 114378 269555
rect 114320 269487 114332 269521
rect 114366 269487 114378 269521
rect 114320 269453 114378 269487
rect 114320 269419 114332 269453
rect 114366 269419 114378 269453
rect 114320 269385 114378 269419
rect 114320 269351 114332 269385
rect 114366 269351 114378 269385
rect 114320 269317 114378 269351
rect 114320 269283 114332 269317
rect 114366 269283 114378 269317
rect 114320 269249 114378 269283
rect 114320 269215 114332 269249
rect 114366 269215 114378 269249
rect 114320 269181 114378 269215
rect 114320 269147 114332 269181
rect 114366 269147 114378 269181
rect 114320 269124 114378 269147
rect 114502 270201 114560 270224
rect 114502 270167 114514 270201
rect 114548 270167 114560 270201
rect 114502 270133 114560 270167
rect 114502 270099 114514 270133
rect 114548 270099 114560 270133
rect 114502 270065 114560 270099
rect 114502 270031 114514 270065
rect 114548 270031 114560 270065
rect 114502 269997 114560 270031
rect 114502 269963 114514 269997
rect 114548 269963 114560 269997
rect 114502 269929 114560 269963
rect 114502 269895 114514 269929
rect 114548 269895 114560 269929
rect 114502 269861 114560 269895
rect 114502 269827 114514 269861
rect 114548 269827 114560 269861
rect 114502 269793 114560 269827
rect 114502 269759 114514 269793
rect 114548 269759 114560 269793
rect 114502 269725 114560 269759
rect 114502 269691 114514 269725
rect 114548 269691 114560 269725
rect 114502 269657 114560 269691
rect 114502 269623 114514 269657
rect 114548 269623 114560 269657
rect 114502 269589 114560 269623
rect 114502 269555 114514 269589
rect 114548 269555 114560 269589
rect 114502 269521 114560 269555
rect 114502 269487 114514 269521
rect 114548 269487 114560 269521
rect 114502 269453 114560 269487
rect 114502 269419 114514 269453
rect 114548 269419 114560 269453
rect 114502 269385 114560 269419
rect 114502 269351 114514 269385
rect 114548 269351 114560 269385
rect 114502 269317 114560 269351
rect 114502 269283 114514 269317
rect 114548 269283 114560 269317
rect 114502 269249 114560 269283
rect 114502 269215 114514 269249
rect 114548 269215 114560 269249
rect 114502 269181 114560 269215
rect 114502 269147 114514 269181
rect 114548 269147 114560 269181
rect 114502 269124 114560 269147
rect 114720 270201 114778 270224
rect 114720 270167 114732 270201
rect 114766 270167 114778 270201
rect 114720 270133 114778 270167
rect 114720 270099 114732 270133
rect 114766 270099 114778 270133
rect 114720 270065 114778 270099
rect 114720 270031 114732 270065
rect 114766 270031 114778 270065
rect 114720 269997 114778 270031
rect 114720 269963 114732 269997
rect 114766 269963 114778 269997
rect 114720 269929 114778 269963
rect 114720 269895 114732 269929
rect 114766 269895 114778 269929
rect 114720 269861 114778 269895
rect 114720 269827 114732 269861
rect 114766 269827 114778 269861
rect 114720 269793 114778 269827
rect 114720 269759 114732 269793
rect 114766 269759 114778 269793
rect 114720 269725 114778 269759
rect 114720 269691 114732 269725
rect 114766 269691 114778 269725
rect 114720 269657 114778 269691
rect 114720 269623 114732 269657
rect 114766 269623 114778 269657
rect 114720 269589 114778 269623
rect 114720 269555 114732 269589
rect 114766 269555 114778 269589
rect 114720 269521 114778 269555
rect 114720 269487 114732 269521
rect 114766 269487 114778 269521
rect 114720 269453 114778 269487
rect 114720 269419 114732 269453
rect 114766 269419 114778 269453
rect 114720 269385 114778 269419
rect 114720 269351 114732 269385
rect 114766 269351 114778 269385
rect 114720 269317 114778 269351
rect 114720 269283 114732 269317
rect 114766 269283 114778 269317
rect 114720 269249 114778 269283
rect 114720 269215 114732 269249
rect 114766 269215 114778 269249
rect 114720 269181 114778 269215
rect 114720 269147 114732 269181
rect 114766 269147 114778 269181
rect 114720 269124 114778 269147
rect 114902 270201 114960 270224
rect 114902 270167 114914 270201
rect 114948 270167 114960 270201
rect 114902 270133 114960 270167
rect 114902 270099 114914 270133
rect 114948 270099 114960 270133
rect 114902 270065 114960 270099
rect 114902 270031 114914 270065
rect 114948 270031 114960 270065
rect 114902 269997 114960 270031
rect 114902 269963 114914 269997
rect 114948 269963 114960 269997
rect 114902 269929 114960 269963
rect 114902 269895 114914 269929
rect 114948 269895 114960 269929
rect 114902 269861 114960 269895
rect 114902 269827 114914 269861
rect 114948 269827 114960 269861
rect 114902 269793 114960 269827
rect 114902 269759 114914 269793
rect 114948 269759 114960 269793
rect 114902 269725 114960 269759
rect 114902 269691 114914 269725
rect 114948 269691 114960 269725
rect 114902 269657 114960 269691
rect 114902 269623 114914 269657
rect 114948 269623 114960 269657
rect 114902 269589 114960 269623
rect 114902 269555 114914 269589
rect 114948 269555 114960 269589
rect 114902 269521 114960 269555
rect 114902 269487 114914 269521
rect 114948 269487 114960 269521
rect 114902 269453 114960 269487
rect 114902 269419 114914 269453
rect 114948 269419 114960 269453
rect 114902 269385 114960 269419
rect 114902 269351 114914 269385
rect 114948 269351 114960 269385
rect 114902 269317 114960 269351
rect 114902 269283 114914 269317
rect 114948 269283 114960 269317
rect 114902 269249 114960 269283
rect 114902 269215 114914 269249
rect 114948 269215 114960 269249
rect 114902 269181 114960 269215
rect 114902 269147 114914 269181
rect 114948 269147 114960 269181
rect 114902 269124 114960 269147
rect 115120 270201 115178 270224
rect 115120 270167 115132 270201
rect 115166 270167 115178 270201
rect 115120 270133 115178 270167
rect 115120 270099 115132 270133
rect 115166 270099 115178 270133
rect 115120 270065 115178 270099
rect 115120 270031 115132 270065
rect 115166 270031 115178 270065
rect 115120 269997 115178 270031
rect 115120 269963 115132 269997
rect 115166 269963 115178 269997
rect 115120 269929 115178 269963
rect 115120 269895 115132 269929
rect 115166 269895 115178 269929
rect 115120 269861 115178 269895
rect 115120 269827 115132 269861
rect 115166 269827 115178 269861
rect 115120 269793 115178 269827
rect 115120 269759 115132 269793
rect 115166 269759 115178 269793
rect 115120 269725 115178 269759
rect 115120 269691 115132 269725
rect 115166 269691 115178 269725
rect 115120 269657 115178 269691
rect 115120 269623 115132 269657
rect 115166 269623 115178 269657
rect 115120 269589 115178 269623
rect 115120 269555 115132 269589
rect 115166 269555 115178 269589
rect 115120 269521 115178 269555
rect 115120 269487 115132 269521
rect 115166 269487 115178 269521
rect 115120 269453 115178 269487
rect 115120 269419 115132 269453
rect 115166 269419 115178 269453
rect 115120 269385 115178 269419
rect 115120 269351 115132 269385
rect 115166 269351 115178 269385
rect 115120 269317 115178 269351
rect 115120 269283 115132 269317
rect 115166 269283 115178 269317
rect 115120 269249 115178 269283
rect 115120 269215 115132 269249
rect 115166 269215 115178 269249
rect 115120 269181 115178 269215
rect 115120 269147 115132 269181
rect 115166 269147 115178 269181
rect 115120 269124 115178 269147
rect 115302 270201 115360 270224
rect 115302 270167 115314 270201
rect 115348 270167 115360 270201
rect 115302 270133 115360 270167
rect 115302 270099 115314 270133
rect 115348 270099 115360 270133
rect 115302 270065 115360 270099
rect 115302 270031 115314 270065
rect 115348 270031 115360 270065
rect 115302 269997 115360 270031
rect 115302 269963 115314 269997
rect 115348 269963 115360 269997
rect 115302 269929 115360 269963
rect 115302 269895 115314 269929
rect 115348 269895 115360 269929
rect 115302 269861 115360 269895
rect 115302 269827 115314 269861
rect 115348 269827 115360 269861
rect 115302 269793 115360 269827
rect 115302 269759 115314 269793
rect 115348 269759 115360 269793
rect 115302 269725 115360 269759
rect 115302 269691 115314 269725
rect 115348 269691 115360 269725
rect 115302 269657 115360 269691
rect 115302 269623 115314 269657
rect 115348 269623 115360 269657
rect 115302 269589 115360 269623
rect 115302 269555 115314 269589
rect 115348 269555 115360 269589
rect 115302 269521 115360 269555
rect 115302 269487 115314 269521
rect 115348 269487 115360 269521
rect 115302 269453 115360 269487
rect 115302 269419 115314 269453
rect 115348 269419 115360 269453
rect 115302 269385 115360 269419
rect 115302 269351 115314 269385
rect 115348 269351 115360 269385
rect 115302 269317 115360 269351
rect 115302 269283 115314 269317
rect 115348 269283 115360 269317
rect 115302 269249 115360 269283
rect 115302 269215 115314 269249
rect 115348 269215 115360 269249
rect 115302 269181 115360 269215
rect 115302 269147 115314 269181
rect 115348 269147 115360 269181
rect 115302 269124 115360 269147
rect 115520 270201 115578 270224
rect 115520 270167 115532 270201
rect 115566 270167 115578 270201
rect 115520 270133 115578 270167
rect 115520 270099 115532 270133
rect 115566 270099 115578 270133
rect 115520 270065 115578 270099
rect 115520 270031 115532 270065
rect 115566 270031 115578 270065
rect 115520 269997 115578 270031
rect 115520 269963 115532 269997
rect 115566 269963 115578 269997
rect 115520 269929 115578 269963
rect 115520 269895 115532 269929
rect 115566 269895 115578 269929
rect 115520 269861 115578 269895
rect 115520 269827 115532 269861
rect 115566 269827 115578 269861
rect 115520 269793 115578 269827
rect 115520 269759 115532 269793
rect 115566 269759 115578 269793
rect 115520 269725 115578 269759
rect 115520 269691 115532 269725
rect 115566 269691 115578 269725
rect 115520 269657 115578 269691
rect 115520 269623 115532 269657
rect 115566 269623 115578 269657
rect 115520 269589 115578 269623
rect 115520 269555 115532 269589
rect 115566 269555 115578 269589
rect 115520 269521 115578 269555
rect 115520 269487 115532 269521
rect 115566 269487 115578 269521
rect 115520 269453 115578 269487
rect 115520 269419 115532 269453
rect 115566 269419 115578 269453
rect 115520 269385 115578 269419
rect 115520 269351 115532 269385
rect 115566 269351 115578 269385
rect 115520 269317 115578 269351
rect 115520 269283 115532 269317
rect 115566 269283 115578 269317
rect 115520 269249 115578 269283
rect 115520 269215 115532 269249
rect 115566 269215 115578 269249
rect 115520 269181 115578 269215
rect 115520 269147 115532 269181
rect 115566 269147 115578 269181
rect 115520 269124 115578 269147
rect 115702 270201 115760 270224
rect 115702 270167 115714 270201
rect 115748 270167 115760 270201
rect 115702 270133 115760 270167
rect 115702 270099 115714 270133
rect 115748 270099 115760 270133
rect 115702 270065 115760 270099
rect 115702 270031 115714 270065
rect 115748 270031 115760 270065
rect 115702 269997 115760 270031
rect 115702 269963 115714 269997
rect 115748 269963 115760 269997
rect 115702 269929 115760 269963
rect 115702 269895 115714 269929
rect 115748 269895 115760 269929
rect 115702 269861 115760 269895
rect 115702 269827 115714 269861
rect 115748 269827 115760 269861
rect 115702 269793 115760 269827
rect 115702 269759 115714 269793
rect 115748 269759 115760 269793
rect 115702 269725 115760 269759
rect 115702 269691 115714 269725
rect 115748 269691 115760 269725
rect 115702 269657 115760 269691
rect 115702 269623 115714 269657
rect 115748 269623 115760 269657
rect 115702 269589 115760 269623
rect 115702 269555 115714 269589
rect 115748 269555 115760 269589
rect 115702 269521 115760 269555
rect 115702 269487 115714 269521
rect 115748 269487 115760 269521
rect 115702 269453 115760 269487
rect 115702 269419 115714 269453
rect 115748 269419 115760 269453
rect 115702 269385 115760 269419
rect 115702 269351 115714 269385
rect 115748 269351 115760 269385
rect 115702 269317 115760 269351
rect 115702 269283 115714 269317
rect 115748 269283 115760 269317
rect 115702 269249 115760 269283
rect 115702 269215 115714 269249
rect 115748 269215 115760 269249
rect 115702 269181 115760 269215
rect 115702 269147 115714 269181
rect 115748 269147 115760 269181
rect 115702 269124 115760 269147
rect 115920 270201 115978 270224
rect 115920 270167 115932 270201
rect 115966 270167 115978 270201
rect 115920 270133 115978 270167
rect 115920 270099 115932 270133
rect 115966 270099 115978 270133
rect 115920 270065 115978 270099
rect 115920 270031 115932 270065
rect 115966 270031 115978 270065
rect 115920 269997 115978 270031
rect 115920 269963 115932 269997
rect 115966 269963 115978 269997
rect 115920 269929 115978 269963
rect 115920 269895 115932 269929
rect 115966 269895 115978 269929
rect 115920 269861 115978 269895
rect 115920 269827 115932 269861
rect 115966 269827 115978 269861
rect 115920 269793 115978 269827
rect 115920 269759 115932 269793
rect 115966 269759 115978 269793
rect 115920 269725 115978 269759
rect 115920 269691 115932 269725
rect 115966 269691 115978 269725
rect 115920 269657 115978 269691
rect 115920 269623 115932 269657
rect 115966 269623 115978 269657
rect 115920 269589 115978 269623
rect 115920 269555 115932 269589
rect 115966 269555 115978 269589
rect 115920 269521 115978 269555
rect 115920 269487 115932 269521
rect 115966 269487 115978 269521
rect 115920 269453 115978 269487
rect 115920 269419 115932 269453
rect 115966 269419 115978 269453
rect 115920 269385 115978 269419
rect 115920 269351 115932 269385
rect 115966 269351 115978 269385
rect 115920 269317 115978 269351
rect 115920 269283 115932 269317
rect 115966 269283 115978 269317
rect 115920 269249 115978 269283
rect 115920 269215 115932 269249
rect 115966 269215 115978 269249
rect 115920 269181 115978 269215
rect 115920 269147 115932 269181
rect 115966 269147 115978 269181
rect 115920 269124 115978 269147
rect 116102 270201 116160 270224
rect 116102 270167 116114 270201
rect 116148 270167 116160 270201
rect 116102 270133 116160 270167
rect 116102 270099 116114 270133
rect 116148 270099 116160 270133
rect 116102 270065 116160 270099
rect 116102 270031 116114 270065
rect 116148 270031 116160 270065
rect 116102 269997 116160 270031
rect 116102 269963 116114 269997
rect 116148 269963 116160 269997
rect 116102 269929 116160 269963
rect 116102 269895 116114 269929
rect 116148 269895 116160 269929
rect 116102 269861 116160 269895
rect 116102 269827 116114 269861
rect 116148 269827 116160 269861
rect 116102 269793 116160 269827
rect 116102 269759 116114 269793
rect 116148 269759 116160 269793
rect 116102 269725 116160 269759
rect 116102 269691 116114 269725
rect 116148 269691 116160 269725
rect 116102 269657 116160 269691
rect 116102 269623 116114 269657
rect 116148 269623 116160 269657
rect 116102 269589 116160 269623
rect 116102 269555 116114 269589
rect 116148 269555 116160 269589
rect 116102 269521 116160 269555
rect 116102 269487 116114 269521
rect 116148 269487 116160 269521
rect 116102 269453 116160 269487
rect 116102 269419 116114 269453
rect 116148 269419 116160 269453
rect 116102 269385 116160 269419
rect 116102 269351 116114 269385
rect 116148 269351 116160 269385
rect 116102 269317 116160 269351
rect 116102 269283 116114 269317
rect 116148 269283 116160 269317
rect 116102 269249 116160 269283
rect 116102 269215 116114 269249
rect 116148 269215 116160 269249
rect 116102 269181 116160 269215
rect 116102 269147 116114 269181
rect 116148 269147 116160 269181
rect 116102 269124 116160 269147
rect 116320 270201 116378 270224
rect 116320 270167 116332 270201
rect 116366 270167 116378 270201
rect 116320 270133 116378 270167
rect 116320 270099 116332 270133
rect 116366 270099 116378 270133
rect 116320 270065 116378 270099
rect 116320 270031 116332 270065
rect 116366 270031 116378 270065
rect 116320 269997 116378 270031
rect 116320 269963 116332 269997
rect 116366 269963 116378 269997
rect 116320 269929 116378 269963
rect 116320 269895 116332 269929
rect 116366 269895 116378 269929
rect 116320 269861 116378 269895
rect 116320 269827 116332 269861
rect 116366 269827 116378 269861
rect 116320 269793 116378 269827
rect 116320 269759 116332 269793
rect 116366 269759 116378 269793
rect 116320 269725 116378 269759
rect 116320 269691 116332 269725
rect 116366 269691 116378 269725
rect 116320 269657 116378 269691
rect 116320 269623 116332 269657
rect 116366 269623 116378 269657
rect 116320 269589 116378 269623
rect 116320 269555 116332 269589
rect 116366 269555 116378 269589
rect 116320 269521 116378 269555
rect 116320 269487 116332 269521
rect 116366 269487 116378 269521
rect 116320 269453 116378 269487
rect 116320 269419 116332 269453
rect 116366 269419 116378 269453
rect 116320 269385 116378 269419
rect 116320 269351 116332 269385
rect 116366 269351 116378 269385
rect 116320 269317 116378 269351
rect 116320 269283 116332 269317
rect 116366 269283 116378 269317
rect 116320 269249 116378 269283
rect 116320 269215 116332 269249
rect 116366 269215 116378 269249
rect 116320 269181 116378 269215
rect 116320 269147 116332 269181
rect 116366 269147 116378 269181
rect 116320 269124 116378 269147
rect 116502 270201 116560 270224
rect 116502 270167 116514 270201
rect 116548 270167 116560 270201
rect 116502 270133 116560 270167
rect 116502 270099 116514 270133
rect 116548 270099 116560 270133
rect 116502 270065 116560 270099
rect 116502 270031 116514 270065
rect 116548 270031 116560 270065
rect 116502 269997 116560 270031
rect 116502 269963 116514 269997
rect 116548 269963 116560 269997
rect 116502 269929 116560 269963
rect 116502 269895 116514 269929
rect 116548 269895 116560 269929
rect 116502 269861 116560 269895
rect 116502 269827 116514 269861
rect 116548 269827 116560 269861
rect 116502 269793 116560 269827
rect 116502 269759 116514 269793
rect 116548 269759 116560 269793
rect 116502 269725 116560 269759
rect 116502 269691 116514 269725
rect 116548 269691 116560 269725
rect 116502 269657 116560 269691
rect 116502 269623 116514 269657
rect 116548 269623 116560 269657
rect 116502 269589 116560 269623
rect 116502 269555 116514 269589
rect 116548 269555 116560 269589
rect 116502 269521 116560 269555
rect 116502 269487 116514 269521
rect 116548 269487 116560 269521
rect 116502 269453 116560 269487
rect 116502 269419 116514 269453
rect 116548 269419 116560 269453
rect 116502 269385 116560 269419
rect 116502 269351 116514 269385
rect 116548 269351 116560 269385
rect 116502 269317 116560 269351
rect 116502 269283 116514 269317
rect 116548 269283 116560 269317
rect 116502 269249 116560 269283
rect 116502 269215 116514 269249
rect 116548 269215 116560 269249
rect 116502 269181 116560 269215
rect 116502 269147 116514 269181
rect 116548 269147 116560 269181
rect 116502 269124 116560 269147
rect 116720 270201 116778 270224
rect 116720 270167 116732 270201
rect 116766 270167 116778 270201
rect 116720 270133 116778 270167
rect 116720 270099 116732 270133
rect 116766 270099 116778 270133
rect 116720 270065 116778 270099
rect 116720 270031 116732 270065
rect 116766 270031 116778 270065
rect 116720 269997 116778 270031
rect 116720 269963 116732 269997
rect 116766 269963 116778 269997
rect 116720 269929 116778 269963
rect 116720 269895 116732 269929
rect 116766 269895 116778 269929
rect 116720 269861 116778 269895
rect 116720 269827 116732 269861
rect 116766 269827 116778 269861
rect 116720 269793 116778 269827
rect 116720 269759 116732 269793
rect 116766 269759 116778 269793
rect 116720 269725 116778 269759
rect 116720 269691 116732 269725
rect 116766 269691 116778 269725
rect 116720 269657 116778 269691
rect 116720 269623 116732 269657
rect 116766 269623 116778 269657
rect 116720 269589 116778 269623
rect 116720 269555 116732 269589
rect 116766 269555 116778 269589
rect 116720 269521 116778 269555
rect 116720 269487 116732 269521
rect 116766 269487 116778 269521
rect 116720 269453 116778 269487
rect 116720 269419 116732 269453
rect 116766 269419 116778 269453
rect 116720 269385 116778 269419
rect 116720 269351 116732 269385
rect 116766 269351 116778 269385
rect 116720 269317 116778 269351
rect 116720 269283 116732 269317
rect 116766 269283 116778 269317
rect 116720 269249 116778 269283
rect 116720 269215 116732 269249
rect 116766 269215 116778 269249
rect 116720 269181 116778 269215
rect 116720 269147 116732 269181
rect 116766 269147 116778 269181
rect 116720 269124 116778 269147
rect 116902 270201 116960 270224
rect 116902 270167 116914 270201
rect 116948 270167 116960 270201
rect 116902 270133 116960 270167
rect 116902 270099 116914 270133
rect 116948 270099 116960 270133
rect 116902 270065 116960 270099
rect 116902 270031 116914 270065
rect 116948 270031 116960 270065
rect 116902 269997 116960 270031
rect 116902 269963 116914 269997
rect 116948 269963 116960 269997
rect 116902 269929 116960 269963
rect 116902 269895 116914 269929
rect 116948 269895 116960 269929
rect 116902 269861 116960 269895
rect 116902 269827 116914 269861
rect 116948 269827 116960 269861
rect 116902 269793 116960 269827
rect 116902 269759 116914 269793
rect 116948 269759 116960 269793
rect 116902 269725 116960 269759
rect 116902 269691 116914 269725
rect 116948 269691 116960 269725
rect 116902 269657 116960 269691
rect 116902 269623 116914 269657
rect 116948 269623 116960 269657
rect 116902 269589 116960 269623
rect 116902 269555 116914 269589
rect 116948 269555 116960 269589
rect 116902 269521 116960 269555
rect 116902 269487 116914 269521
rect 116948 269487 116960 269521
rect 116902 269453 116960 269487
rect 116902 269419 116914 269453
rect 116948 269419 116960 269453
rect 116902 269385 116960 269419
rect 116902 269351 116914 269385
rect 116948 269351 116960 269385
rect 116902 269317 116960 269351
rect 116902 269283 116914 269317
rect 116948 269283 116960 269317
rect 116902 269249 116960 269283
rect 116902 269215 116914 269249
rect 116948 269215 116960 269249
rect 116902 269181 116960 269215
rect 116902 269147 116914 269181
rect 116948 269147 116960 269181
rect 116902 269124 116960 269147
rect 117120 270201 117178 270224
rect 117120 270167 117132 270201
rect 117166 270167 117178 270201
rect 117120 270133 117178 270167
rect 117120 270099 117132 270133
rect 117166 270099 117178 270133
rect 117120 270065 117178 270099
rect 117120 270031 117132 270065
rect 117166 270031 117178 270065
rect 117120 269997 117178 270031
rect 117120 269963 117132 269997
rect 117166 269963 117178 269997
rect 117120 269929 117178 269963
rect 117120 269895 117132 269929
rect 117166 269895 117178 269929
rect 117120 269861 117178 269895
rect 117120 269827 117132 269861
rect 117166 269827 117178 269861
rect 117120 269793 117178 269827
rect 117120 269759 117132 269793
rect 117166 269759 117178 269793
rect 117120 269725 117178 269759
rect 117120 269691 117132 269725
rect 117166 269691 117178 269725
rect 117120 269657 117178 269691
rect 117120 269623 117132 269657
rect 117166 269623 117178 269657
rect 117120 269589 117178 269623
rect 117120 269555 117132 269589
rect 117166 269555 117178 269589
rect 117120 269521 117178 269555
rect 117120 269487 117132 269521
rect 117166 269487 117178 269521
rect 117120 269453 117178 269487
rect 117120 269419 117132 269453
rect 117166 269419 117178 269453
rect 117120 269385 117178 269419
rect 117120 269351 117132 269385
rect 117166 269351 117178 269385
rect 117120 269317 117178 269351
rect 117120 269283 117132 269317
rect 117166 269283 117178 269317
rect 117120 269249 117178 269283
rect 117120 269215 117132 269249
rect 117166 269215 117178 269249
rect 117120 269181 117178 269215
rect 117120 269147 117132 269181
rect 117166 269147 117178 269181
rect 117120 269124 117178 269147
rect 117302 270201 117360 270224
rect 117302 270167 117314 270201
rect 117348 270167 117360 270201
rect 117302 270133 117360 270167
rect 117302 270099 117314 270133
rect 117348 270099 117360 270133
rect 117302 270065 117360 270099
rect 117302 270031 117314 270065
rect 117348 270031 117360 270065
rect 117302 269997 117360 270031
rect 117302 269963 117314 269997
rect 117348 269963 117360 269997
rect 117302 269929 117360 269963
rect 117302 269895 117314 269929
rect 117348 269895 117360 269929
rect 117302 269861 117360 269895
rect 117302 269827 117314 269861
rect 117348 269827 117360 269861
rect 117302 269793 117360 269827
rect 117302 269759 117314 269793
rect 117348 269759 117360 269793
rect 117302 269725 117360 269759
rect 117302 269691 117314 269725
rect 117348 269691 117360 269725
rect 117302 269657 117360 269691
rect 117302 269623 117314 269657
rect 117348 269623 117360 269657
rect 117302 269589 117360 269623
rect 117302 269555 117314 269589
rect 117348 269555 117360 269589
rect 117302 269521 117360 269555
rect 117302 269487 117314 269521
rect 117348 269487 117360 269521
rect 117302 269453 117360 269487
rect 117302 269419 117314 269453
rect 117348 269419 117360 269453
rect 117302 269385 117360 269419
rect 117302 269351 117314 269385
rect 117348 269351 117360 269385
rect 117302 269317 117360 269351
rect 117302 269283 117314 269317
rect 117348 269283 117360 269317
rect 117302 269249 117360 269283
rect 117302 269215 117314 269249
rect 117348 269215 117360 269249
rect 117302 269181 117360 269215
rect 117302 269147 117314 269181
rect 117348 269147 117360 269181
rect 117302 269124 117360 269147
rect 117520 270201 117578 270224
rect 117520 270167 117532 270201
rect 117566 270167 117578 270201
rect 117520 270133 117578 270167
rect 117520 270099 117532 270133
rect 117566 270099 117578 270133
rect 117520 270065 117578 270099
rect 117520 270031 117532 270065
rect 117566 270031 117578 270065
rect 117520 269997 117578 270031
rect 117520 269963 117532 269997
rect 117566 269963 117578 269997
rect 117520 269929 117578 269963
rect 117520 269895 117532 269929
rect 117566 269895 117578 269929
rect 117520 269861 117578 269895
rect 117520 269827 117532 269861
rect 117566 269827 117578 269861
rect 117520 269793 117578 269827
rect 117520 269759 117532 269793
rect 117566 269759 117578 269793
rect 117520 269725 117578 269759
rect 117520 269691 117532 269725
rect 117566 269691 117578 269725
rect 117520 269657 117578 269691
rect 117520 269623 117532 269657
rect 117566 269623 117578 269657
rect 117520 269589 117578 269623
rect 117520 269555 117532 269589
rect 117566 269555 117578 269589
rect 117520 269521 117578 269555
rect 117520 269487 117532 269521
rect 117566 269487 117578 269521
rect 117520 269453 117578 269487
rect 117520 269419 117532 269453
rect 117566 269419 117578 269453
rect 117520 269385 117578 269419
rect 117520 269351 117532 269385
rect 117566 269351 117578 269385
rect 117520 269317 117578 269351
rect 117520 269283 117532 269317
rect 117566 269283 117578 269317
rect 117520 269249 117578 269283
rect 117520 269215 117532 269249
rect 117566 269215 117578 269249
rect 117520 269181 117578 269215
rect 117520 269147 117532 269181
rect 117566 269147 117578 269181
rect 117520 269124 117578 269147
rect 117702 270201 117760 270224
rect 117702 270167 117714 270201
rect 117748 270167 117760 270201
rect 117702 270133 117760 270167
rect 117702 270099 117714 270133
rect 117748 270099 117760 270133
rect 117702 270065 117760 270099
rect 117702 270031 117714 270065
rect 117748 270031 117760 270065
rect 117702 269997 117760 270031
rect 117702 269963 117714 269997
rect 117748 269963 117760 269997
rect 117702 269929 117760 269963
rect 117702 269895 117714 269929
rect 117748 269895 117760 269929
rect 117702 269861 117760 269895
rect 117702 269827 117714 269861
rect 117748 269827 117760 269861
rect 117702 269793 117760 269827
rect 117702 269759 117714 269793
rect 117748 269759 117760 269793
rect 117702 269725 117760 269759
rect 117702 269691 117714 269725
rect 117748 269691 117760 269725
rect 117702 269657 117760 269691
rect 117702 269623 117714 269657
rect 117748 269623 117760 269657
rect 117702 269589 117760 269623
rect 117702 269555 117714 269589
rect 117748 269555 117760 269589
rect 117702 269521 117760 269555
rect 117702 269487 117714 269521
rect 117748 269487 117760 269521
rect 117702 269453 117760 269487
rect 117702 269419 117714 269453
rect 117748 269419 117760 269453
rect 117702 269385 117760 269419
rect 117702 269351 117714 269385
rect 117748 269351 117760 269385
rect 117702 269317 117760 269351
rect 117702 269283 117714 269317
rect 117748 269283 117760 269317
rect 117702 269249 117760 269283
rect 117702 269215 117714 269249
rect 117748 269215 117760 269249
rect 117702 269181 117760 269215
rect 117702 269147 117714 269181
rect 117748 269147 117760 269181
rect 117702 269124 117760 269147
rect 117920 270201 117978 270224
rect 117920 270167 117932 270201
rect 117966 270167 117978 270201
rect 117920 270133 117978 270167
rect 117920 270099 117932 270133
rect 117966 270099 117978 270133
rect 117920 270065 117978 270099
rect 117920 270031 117932 270065
rect 117966 270031 117978 270065
rect 117920 269997 117978 270031
rect 117920 269963 117932 269997
rect 117966 269963 117978 269997
rect 117920 269929 117978 269963
rect 117920 269895 117932 269929
rect 117966 269895 117978 269929
rect 117920 269861 117978 269895
rect 117920 269827 117932 269861
rect 117966 269827 117978 269861
rect 117920 269793 117978 269827
rect 117920 269759 117932 269793
rect 117966 269759 117978 269793
rect 117920 269725 117978 269759
rect 117920 269691 117932 269725
rect 117966 269691 117978 269725
rect 117920 269657 117978 269691
rect 117920 269623 117932 269657
rect 117966 269623 117978 269657
rect 117920 269589 117978 269623
rect 117920 269555 117932 269589
rect 117966 269555 117978 269589
rect 117920 269521 117978 269555
rect 117920 269487 117932 269521
rect 117966 269487 117978 269521
rect 117920 269453 117978 269487
rect 117920 269419 117932 269453
rect 117966 269419 117978 269453
rect 117920 269385 117978 269419
rect 117920 269351 117932 269385
rect 117966 269351 117978 269385
rect 117920 269317 117978 269351
rect 117920 269283 117932 269317
rect 117966 269283 117978 269317
rect 117920 269249 117978 269283
rect 117920 269215 117932 269249
rect 117966 269215 117978 269249
rect 117920 269181 117978 269215
rect 117920 269147 117932 269181
rect 117966 269147 117978 269181
rect 117920 269124 117978 269147
rect 118102 270201 118160 270224
rect 118102 270167 118114 270201
rect 118148 270167 118160 270201
rect 118102 270133 118160 270167
rect 118102 270099 118114 270133
rect 118148 270099 118160 270133
rect 118102 270065 118160 270099
rect 118102 270031 118114 270065
rect 118148 270031 118160 270065
rect 118102 269997 118160 270031
rect 118102 269963 118114 269997
rect 118148 269963 118160 269997
rect 118102 269929 118160 269963
rect 118102 269895 118114 269929
rect 118148 269895 118160 269929
rect 118102 269861 118160 269895
rect 118102 269827 118114 269861
rect 118148 269827 118160 269861
rect 118102 269793 118160 269827
rect 118102 269759 118114 269793
rect 118148 269759 118160 269793
rect 118102 269725 118160 269759
rect 118102 269691 118114 269725
rect 118148 269691 118160 269725
rect 118102 269657 118160 269691
rect 118102 269623 118114 269657
rect 118148 269623 118160 269657
rect 118102 269589 118160 269623
rect 118102 269555 118114 269589
rect 118148 269555 118160 269589
rect 118102 269521 118160 269555
rect 118102 269487 118114 269521
rect 118148 269487 118160 269521
rect 118102 269453 118160 269487
rect 118102 269419 118114 269453
rect 118148 269419 118160 269453
rect 118102 269385 118160 269419
rect 118102 269351 118114 269385
rect 118148 269351 118160 269385
rect 118102 269317 118160 269351
rect 118102 269283 118114 269317
rect 118148 269283 118160 269317
rect 118102 269249 118160 269283
rect 118102 269215 118114 269249
rect 118148 269215 118160 269249
rect 118102 269181 118160 269215
rect 118102 269147 118114 269181
rect 118148 269147 118160 269181
rect 118102 269124 118160 269147
rect 118320 270201 118378 270224
rect 118320 270167 118332 270201
rect 118366 270167 118378 270201
rect 118320 270133 118378 270167
rect 118320 270099 118332 270133
rect 118366 270099 118378 270133
rect 118320 270065 118378 270099
rect 118320 270031 118332 270065
rect 118366 270031 118378 270065
rect 118320 269997 118378 270031
rect 118320 269963 118332 269997
rect 118366 269963 118378 269997
rect 118320 269929 118378 269963
rect 118320 269895 118332 269929
rect 118366 269895 118378 269929
rect 118320 269861 118378 269895
rect 118320 269827 118332 269861
rect 118366 269827 118378 269861
rect 118320 269793 118378 269827
rect 118320 269759 118332 269793
rect 118366 269759 118378 269793
rect 118320 269725 118378 269759
rect 118320 269691 118332 269725
rect 118366 269691 118378 269725
rect 118320 269657 118378 269691
rect 118320 269623 118332 269657
rect 118366 269623 118378 269657
rect 118320 269589 118378 269623
rect 118320 269555 118332 269589
rect 118366 269555 118378 269589
rect 118320 269521 118378 269555
rect 118320 269487 118332 269521
rect 118366 269487 118378 269521
rect 118320 269453 118378 269487
rect 118320 269419 118332 269453
rect 118366 269419 118378 269453
rect 118320 269385 118378 269419
rect 118320 269351 118332 269385
rect 118366 269351 118378 269385
rect 118320 269317 118378 269351
rect 118320 269283 118332 269317
rect 118366 269283 118378 269317
rect 118320 269249 118378 269283
rect 118320 269215 118332 269249
rect 118366 269215 118378 269249
rect 118320 269181 118378 269215
rect 118320 269147 118332 269181
rect 118366 269147 118378 269181
rect 118320 269124 118378 269147
rect 118502 270201 118560 270224
rect 118502 270167 118514 270201
rect 118548 270167 118560 270201
rect 118502 270133 118560 270167
rect 118502 270099 118514 270133
rect 118548 270099 118560 270133
rect 118502 270065 118560 270099
rect 118502 270031 118514 270065
rect 118548 270031 118560 270065
rect 118502 269997 118560 270031
rect 118502 269963 118514 269997
rect 118548 269963 118560 269997
rect 118502 269929 118560 269963
rect 118502 269895 118514 269929
rect 118548 269895 118560 269929
rect 118502 269861 118560 269895
rect 118502 269827 118514 269861
rect 118548 269827 118560 269861
rect 118502 269793 118560 269827
rect 118502 269759 118514 269793
rect 118548 269759 118560 269793
rect 118502 269725 118560 269759
rect 118502 269691 118514 269725
rect 118548 269691 118560 269725
rect 118502 269657 118560 269691
rect 118502 269623 118514 269657
rect 118548 269623 118560 269657
rect 118502 269589 118560 269623
rect 118502 269555 118514 269589
rect 118548 269555 118560 269589
rect 118502 269521 118560 269555
rect 118502 269487 118514 269521
rect 118548 269487 118560 269521
rect 118502 269453 118560 269487
rect 118502 269419 118514 269453
rect 118548 269419 118560 269453
rect 118502 269385 118560 269419
rect 118502 269351 118514 269385
rect 118548 269351 118560 269385
rect 118502 269317 118560 269351
rect 118502 269283 118514 269317
rect 118548 269283 118560 269317
rect 118502 269249 118560 269283
rect 118502 269215 118514 269249
rect 118548 269215 118560 269249
rect 118502 269181 118560 269215
rect 118502 269147 118514 269181
rect 118548 269147 118560 269181
rect 118502 269124 118560 269147
rect 118720 270201 118778 270224
rect 118720 270167 118732 270201
rect 118766 270167 118778 270201
rect 118720 270133 118778 270167
rect 118720 270099 118732 270133
rect 118766 270099 118778 270133
rect 118720 270065 118778 270099
rect 118720 270031 118732 270065
rect 118766 270031 118778 270065
rect 118720 269997 118778 270031
rect 118720 269963 118732 269997
rect 118766 269963 118778 269997
rect 118720 269929 118778 269963
rect 118720 269895 118732 269929
rect 118766 269895 118778 269929
rect 118720 269861 118778 269895
rect 118720 269827 118732 269861
rect 118766 269827 118778 269861
rect 118720 269793 118778 269827
rect 118720 269759 118732 269793
rect 118766 269759 118778 269793
rect 118720 269725 118778 269759
rect 118720 269691 118732 269725
rect 118766 269691 118778 269725
rect 118720 269657 118778 269691
rect 118720 269623 118732 269657
rect 118766 269623 118778 269657
rect 118720 269589 118778 269623
rect 118720 269555 118732 269589
rect 118766 269555 118778 269589
rect 118720 269521 118778 269555
rect 118720 269487 118732 269521
rect 118766 269487 118778 269521
rect 118720 269453 118778 269487
rect 118720 269419 118732 269453
rect 118766 269419 118778 269453
rect 118720 269385 118778 269419
rect 118720 269351 118732 269385
rect 118766 269351 118778 269385
rect 118720 269317 118778 269351
rect 118720 269283 118732 269317
rect 118766 269283 118778 269317
rect 118720 269249 118778 269283
rect 118720 269215 118732 269249
rect 118766 269215 118778 269249
rect 118720 269181 118778 269215
rect 118720 269147 118732 269181
rect 118766 269147 118778 269181
rect 118720 269124 118778 269147
rect 122894 274847 122952 274862
rect 122894 274813 122906 274847
rect 122940 274813 122952 274847
rect 122894 274779 122952 274813
rect 122894 274745 122906 274779
rect 122940 274745 122952 274779
rect 122894 274711 122952 274745
rect 122894 274677 122906 274711
rect 122940 274677 122952 274711
rect 122894 274662 122952 274677
rect 123952 274847 124010 274862
rect 123952 274813 123964 274847
rect 123998 274813 124010 274847
rect 123952 274779 124010 274813
rect 123952 274745 123964 274779
rect 123998 274745 124010 274779
rect 123952 274711 124010 274745
rect 123952 274677 123964 274711
rect 123998 274677 124010 274711
rect 123952 274662 124010 274677
rect 122219 274249 122277 274278
rect 122219 274215 122231 274249
rect 122265 274215 122277 274249
rect 122219 274181 122277 274215
rect 122219 274147 122231 274181
rect 122265 274147 122277 274181
rect 122219 274113 122277 274147
rect 122219 274079 122231 274113
rect 122265 274079 122277 274113
rect 122219 274045 122277 274079
rect 122219 274011 122231 274045
rect 122265 274011 122277 274045
rect 122219 273977 122277 274011
rect 122219 273943 122231 273977
rect 122265 273943 122277 273977
rect 122219 273909 122277 273943
rect 122219 273875 122231 273909
rect 122265 273875 122277 273909
rect 122219 273841 122277 273875
rect 122219 273807 122231 273841
rect 122265 273807 122277 273841
rect 122219 273778 122277 273807
rect 122477 274249 122535 274278
rect 122477 274215 122489 274249
rect 122523 274215 122535 274249
rect 122477 274181 122535 274215
rect 122477 274147 122489 274181
rect 122523 274147 122535 274181
rect 122477 274113 122535 274147
rect 122477 274079 122489 274113
rect 122523 274079 122535 274113
rect 122477 274045 122535 274079
rect 122477 274011 122489 274045
rect 122523 274011 122535 274045
rect 122477 273977 122535 274011
rect 122477 273943 122489 273977
rect 122523 273943 122535 273977
rect 122477 273909 122535 273943
rect 122477 273875 122489 273909
rect 122523 273875 122535 273909
rect 122477 273841 122535 273875
rect 122477 273807 122489 273841
rect 122523 273807 122535 273841
rect 122477 273778 122535 273807
rect 122635 274249 122693 274278
rect 122635 274215 122647 274249
rect 122681 274215 122693 274249
rect 122635 274181 122693 274215
rect 122635 274147 122647 274181
rect 122681 274147 122693 274181
rect 122635 274113 122693 274147
rect 122635 274079 122647 274113
rect 122681 274079 122693 274113
rect 122635 274045 122693 274079
rect 122635 274011 122647 274045
rect 122681 274011 122693 274045
rect 122635 273977 122693 274011
rect 122635 273943 122647 273977
rect 122681 273943 122693 273977
rect 122635 273909 122693 273943
rect 122635 273875 122647 273909
rect 122681 273875 122693 273909
rect 122635 273841 122693 273875
rect 122635 273807 122647 273841
rect 122681 273807 122693 273841
rect 122635 273778 122693 273807
rect 122893 274249 122951 274278
rect 122893 274215 122905 274249
rect 122939 274215 122951 274249
rect 122893 274181 122951 274215
rect 122893 274147 122905 274181
rect 122939 274147 122951 274181
rect 122893 274113 122951 274147
rect 122893 274079 122905 274113
rect 122939 274079 122951 274113
rect 122893 274045 122951 274079
rect 122893 274011 122905 274045
rect 122939 274011 122951 274045
rect 122893 273977 122951 274011
rect 122893 273943 122905 273977
rect 122939 273943 122951 273977
rect 122893 273909 122951 273943
rect 122893 273875 122905 273909
rect 122939 273875 122951 273909
rect 122893 273841 122951 273875
rect 122893 273807 122905 273841
rect 122939 273807 122951 273841
rect 122893 273778 122951 273807
rect 123051 274249 123109 274278
rect 123051 274215 123063 274249
rect 123097 274215 123109 274249
rect 123051 274181 123109 274215
rect 123051 274147 123063 274181
rect 123097 274147 123109 274181
rect 123051 274113 123109 274147
rect 123051 274079 123063 274113
rect 123097 274079 123109 274113
rect 123051 274045 123109 274079
rect 123051 274011 123063 274045
rect 123097 274011 123109 274045
rect 123051 273977 123109 274011
rect 123051 273943 123063 273977
rect 123097 273943 123109 273977
rect 123051 273909 123109 273943
rect 123051 273875 123063 273909
rect 123097 273875 123109 273909
rect 123051 273841 123109 273875
rect 123051 273807 123063 273841
rect 123097 273807 123109 273841
rect 123051 273778 123109 273807
rect 123309 274249 123367 274278
rect 123309 274215 123321 274249
rect 123355 274215 123367 274249
rect 123309 274181 123367 274215
rect 123309 274147 123321 274181
rect 123355 274147 123367 274181
rect 123309 274113 123367 274147
rect 123309 274079 123321 274113
rect 123355 274079 123367 274113
rect 123309 274045 123367 274079
rect 123309 274011 123321 274045
rect 123355 274011 123367 274045
rect 123309 273977 123367 274011
rect 123309 273943 123321 273977
rect 123355 273943 123367 273977
rect 123309 273909 123367 273943
rect 123309 273875 123321 273909
rect 123355 273875 123367 273909
rect 123309 273841 123367 273875
rect 123309 273807 123321 273841
rect 123355 273807 123367 273841
rect 123309 273778 123367 273807
rect 123467 274249 123525 274278
rect 123467 274215 123479 274249
rect 123513 274215 123525 274249
rect 123467 274181 123525 274215
rect 123467 274147 123479 274181
rect 123513 274147 123525 274181
rect 123467 274113 123525 274147
rect 123467 274079 123479 274113
rect 123513 274079 123525 274113
rect 123467 274045 123525 274079
rect 123467 274011 123479 274045
rect 123513 274011 123525 274045
rect 123467 273977 123525 274011
rect 123467 273943 123479 273977
rect 123513 273943 123525 273977
rect 123467 273909 123525 273943
rect 123467 273875 123479 273909
rect 123513 273875 123525 273909
rect 123467 273841 123525 273875
rect 123467 273807 123479 273841
rect 123513 273807 123525 273841
rect 123467 273778 123525 273807
rect 123725 274249 123783 274278
rect 123725 274215 123737 274249
rect 123771 274215 123783 274249
rect 123725 274181 123783 274215
rect 123725 274147 123737 274181
rect 123771 274147 123783 274181
rect 123725 274113 123783 274147
rect 123725 274079 123737 274113
rect 123771 274079 123783 274113
rect 123725 274045 123783 274079
rect 123725 274011 123737 274045
rect 123771 274011 123783 274045
rect 123725 273977 123783 274011
rect 123725 273943 123737 273977
rect 123771 273943 123783 273977
rect 123725 273909 123783 273943
rect 123725 273875 123737 273909
rect 123771 273875 123783 273909
rect 123725 273841 123783 273875
rect 123725 273807 123737 273841
rect 123771 273807 123783 273841
rect 123725 273778 123783 273807
rect 123883 274249 123941 274278
rect 123883 274215 123895 274249
rect 123929 274215 123941 274249
rect 123883 274181 123941 274215
rect 123883 274147 123895 274181
rect 123929 274147 123941 274181
rect 123883 274113 123941 274147
rect 123883 274079 123895 274113
rect 123929 274079 123941 274113
rect 123883 274045 123941 274079
rect 123883 274011 123895 274045
rect 123929 274011 123941 274045
rect 123883 273977 123941 274011
rect 123883 273943 123895 273977
rect 123929 273943 123941 273977
rect 123883 273909 123941 273943
rect 123883 273875 123895 273909
rect 123929 273875 123941 273909
rect 123883 273841 123941 273875
rect 123883 273807 123895 273841
rect 123929 273807 123941 273841
rect 123883 273778 123941 273807
rect 124141 274249 124199 274278
rect 124141 274215 124153 274249
rect 124187 274215 124199 274249
rect 124141 274181 124199 274215
rect 124141 274147 124153 274181
rect 124187 274147 124199 274181
rect 124141 274113 124199 274147
rect 124141 274079 124153 274113
rect 124187 274079 124199 274113
rect 124141 274045 124199 274079
rect 124141 274011 124153 274045
rect 124187 274011 124199 274045
rect 124141 273977 124199 274011
rect 124141 273943 124153 273977
rect 124187 273943 124199 273977
rect 124141 273909 124199 273943
rect 124141 273875 124153 273909
rect 124187 273875 124199 273909
rect 124141 273841 124199 273875
rect 124141 273807 124153 273841
rect 124187 273807 124199 273841
rect 124141 273778 124199 273807
rect 124299 274249 124357 274278
rect 124299 274215 124311 274249
rect 124345 274215 124357 274249
rect 124299 274181 124357 274215
rect 124299 274147 124311 274181
rect 124345 274147 124357 274181
rect 124299 274113 124357 274147
rect 124299 274079 124311 274113
rect 124345 274079 124357 274113
rect 124299 274045 124357 274079
rect 124299 274011 124311 274045
rect 124345 274011 124357 274045
rect 124299 273977 124357 274011
rect 124299 273943 124311 273977
rect 124345 273943 124357 273977
rect 124299 273909 124357 273943
rect 124299 273875 124311 273909
rect 124345 273875 124357 273909
rect 124299 273841 124357 273875
rect 124299 273807 124311 273841
rect 124345 273807 124357 273841
rect 124299 273778 124357 273807
rect 124557 274249 124615 274278
rect 124557 274215 124569 274249
rect 124603 274215 124615 274249
rect 124557 274181 124615 274215
rect 124557 274147 124569 274181
rect 124603 274147 124615 274181
rect 124557 274113 124615 274147
rect 124557 274079 124569 274113
rect 124603 274079 124615 274113
rect 124557 274045 124615 274079
rect 124557 274011 124569 274045
rect 124603 274011 124615 274045
rect 124557 273977 124615 274011
rect 124557 273943 124569 273977
rect 124603 273943 124615 273977
rect 124557 273909 124615 273943
rect 124557 273875 124569 273909
rect 124603 273875 124615 273909
rect 124557 273841 124615 273875
rect 124557 273807 124569 273841
rect 124603 273807 124615 273841
rect 124557 273778 124615 273807
rect 124192 272566 124692 272578
rect 124192 272532 124221 272566
rect 124255 272532 124289 272566
rect 124323 272532 124357 272566
rect 124391 272532 124425 272566
rect 124459 272532 124493 272566
rect 124527 272532 124561 272566
rect 124595 272532 124629 272566
rect 124663 272532 124692 272566
rect 124192 272520 124692 272532
rect 124192 272308 124692 272320
rect 124192 272274 124221 272308
rect 124255 272274 124289 272308
rect 124323 272274 124357 272308
rect 124391 272274 124425 272308
rect 124459 272274 124493 272308
rect 124527 272274 124561 272308
rect 124595 272274 124629 272308
rect 124663 272274 124692 272308
rect 124192 272262 124692 272274
rect 124192 272150 124692 272162
rect 124192 272116 124221 272150
rect 124255 272116 124289 272150
rect 124323 272116 124357 272150
rect 124391 272116 124425 272150
rect 124459 272116 124493 272150
rect 124527 272116 124561 272150
rect 124595 272116 124629 272150
rect 124663 272116 124692 272150
rect 124192 272104 124692 272116
rect 124192 271892 124692 271904
rect 124192 271858 124221 271892
rect 124255 271858 124289 271892
rect 124323 271858 124357 271892
rect 124391 271858 124425 271892
rect 124459 271858 124493 271892
rect 124527 271858 124561 271892
rect 124595 271858 124629 271892
rect 124663 271858 124692 271892
rect 124192 271846 124692 271858
rect 124192 271734 124692 271746
rect 124192 271700 124221 271734
rect 124255 271700 124289 271734
rect 124323 271700 124357 271734
rect 124391 271700 124425 271734
rect 124459 271700 124493 271734
rect 124527 271700 124561 271734
rect 124595 271700 124629 271734
rect 124663 271700 124692 271734
rect 124192 271688 124692 271700
rect 124192 271476 124692 271488
rect 124192 271442 124221 271476
rect 124255 271442 124289 271476
rect 124323 271442 124357 271476
rect 124391 271442 124425 271476
rect 124459 271442 124493 271476
rect 124527 271442 124561 271476
rect 124595 271442 124629 271476
rect 124663 271442 124692 271476
rect 124192 271430 124692 271442
rect 124192 271318 124692 271330
rect 124192 271284 124221 271318
rect 124255 271284 124289 271318
rect 124323 271284 124357 271318
rect 124391 271284 124425 271318
rect 124459 271284 124493 271318
rect 124527 271284 124561 271318
rect 124595 271284 124629 271318
rect 124663 271284 124692 271318
rect 124192 271272 124692 271284
rect 124192 271060 124692 271072
rect 124192 271026 124221 271060
rect 124255 271026 124289 271060
rect 124323 271026 124357 271060
rect 124391 271026 124425 271060
rect 124459 271026 124493 271060
rect 124527 271026 124561 271060
rect 124595 271026 124629 271060
rect 124663 271026 124692 271060
rect 124192 271014 124692 271026
rect 124192 270902 124692 270914
rect 124192 270868 124221 270902
rect 124255 270868 124289 270902
rect 124323 270868 124357 270902
rect 124391 270868 124425 270902
rect 124459 270868 124493 270902
rect 124527 270868 124561 270902
rect 124595 270868 124629 270902
rect 124663 270868 124692 270902
rect 124192 270856 124692 270868
rect 124192 270644 124692 270656
rect 124192 270610 124221 270644
rect 124255 270610 124289 270644
rect 124323 270610 124357 270644
rect 124391 270610 124425 270644
rect 124459 270610 124493 270644
rect 124527 270610 124561 270644
rect 124595 270610 124629 270644
rect 124663 270610 124692 270644
rect 124192 270598 124692 270610
rect 124192 270486 124692 270498
rect 124192 270452 124221 270486
rect 124255 270452 124289 270486
rect 124323 270452 124357 270486
rect 124391 270452 124425 270486
rect 124459 270452 124493 270486
rect 124527 270452 124561 270486
rect 124595 270452 124629 270486
rect 124663 270452 124692 270486
rect 124192 270440 124692 270452
rect 124192 270228 124692 270240
rect 124192 270194 124221 270228
rect 124255 270194 124289 270228
rect 124323 270194 124357 270228
rect 124391 270194 124425 270228
rect 124459 270194 124493 270228
rect 124527 270194 124561 270228
rect 124595 270194 124629 270228
rect 124663 270194 124692 270228
rect 124192 270182 124692 270194
rect 124192 270070 124692 270082
rect 124192 270036 124221 270070
rect 124255 270036 124289 270070
rect 124323 270036 124357 270070
rect 124391 270036 124425 270070
rect 124459 270036 124493 270070
rect 124527 270036 124561 270070
rect 124595 270036 124629 270070
rect 124663 270036 124692 270070
rect 124192 270024 124692 270036
rect 124192 269812 124692 269824
rect 124192 269778 124221 269812
rect 124255 269778 124289 269812
rect 124323 269778 124357 269812
rect 124391 269778 124425 269812
rect 124459 269778 124493 269812
rect 124527 269778 124561 269812
rect 124595 269778 124629 269812
rect 124663 269778 124692 269812
rect 124192 269766 124692 269778
rect 124192 269654 124692 269666
rect 124192 269620 124221 269654
rect 124255 269620 124289 269654
rect 124323 269620 124357 269654
rect 124391 269620 124425 269654
rect 124459 269620 124493 269654
rect 124527 269620 124561 269654
rect 124595 269620 124629 269654
rect 124663 269620 124692 269654
rect 124192 269608 124692 269620
rect 124192 269396 124692 269408
rect 124192 269362 124221 269396
rect 124255 269362 124289 269396
rect 124323 269362 124357 269396
rect 124391 269362 124425 269396
rect 124459 269362 124493 269396
rect 124527 269362 124561 269396
rect 124595 269362 124629 269396
rect 124663 269362 124692 269396
rect 124192 269350 124692 269362
<< pdiff >>
rect 106368 279057 107582 279069
rect 106368 279023 106380 279057
rect 106414 279023 106448 279057
rect 106482 279023 106516 279057
rect 106550 279023 106584 279057
rect 106618 279023 106652 279057
rect 106686 279023 106720 279057
rect 106754 279023 106788 279057
rect 106822 279023 106856 279057
rect 106890 279023 106924 279057
rect 106958 279023 106992 279057
rect 107026 279023 107060 279057
rect 107094 279023 107128 279057
rect 107162 279023 107196 279057
rect 107230 279023 107264 279057
rect 107298 279023 107332 279057
rect 107366 279023 107400 279057
rect 107434 279023 107468 279057
rect 107502 279023 107536 279057
rect 107570 279023 107582 279057
rect 106368 279011 107582 279023
rect 106368 278745 107582 278757
rect 106368 278711 106380 278745
rect 106414 278711 106448 278745
rect 106482 278711 106516 278745
rect 106550 278711 106584 278745
rect 106618 278711 106652 278745
rect 106686 278711 106720 278745
rect 106754 278711 106788 278745
rect 106822 278711 106856 278745
rect 106890 278711 106924 278745
rect 106958 278711 106992 278745
rect 107026 278711 107060 278745
rect 107094 278711 107128 278745
rect 107162 278711 107196 278745
rect 107230 278711 107264 278745
rect 107298 278711 107332 278745
rect 107366 278711 107400 278745
rect 107434 278711 107468 278745
rect 107502 278711 107536 278745
rect 107570 278711 107582 278745
rect 106368 278699 107582 278711
rect 106368 278457 107582 278469
rect 106368 278423 106380 278457
rect 106414 278423 106448 278457
rect 106482 278423 106516 278457
rect 106550 278423 106584 278457
rect 106618 278423 106652 278457
rect 106686 278423 106720 278457
rect 106754 278423 106788 278457
rect 106822 278423 106856 278457
rect 106890 278423 106924 278457
rect 106958 278423 106992 278457
rect 107026 278423 107060 278457
rect 107094 278423 107128 278457
rect 107162 278423 107196 278457
rect 107230 278423 107264 278457
rect 107298 278423 107332 278457
rect 107366 278423 107400 278457
rect 107434 278423 107468 278457
rect 107502 278423 107536 278457
rect 107570 278423 107582 278457
rect 106368 278411 107582 278423
rect 106368 278145 107582 278157
rect 106368 278111 106380 278145
rect 106414 278111 106448 278145
rect 106482 278111 106516 278145
rect 106550 278111 106584 278145
rect 106618 278111 106652 278145
rect 106686 278111 106720 278145
rect 106754 278111 106788 278145
rect 106822 278111 106856 278145
rect 106890 278111 106924 278145
rect 106958 278111 106992 278145
rect 107026 278111 107060 278145
rect 107094 278111 107128 278145
rect 107162 278111 107196 278145
rect 107230 278111 107264 278145
rect 107298 278111 107332 278145
rect 107366 278111 107400 278145
rect 107434 278111 107468 278145
rect 107502 278111 107536 278145
rect 107570 278111 107582 278145
rect 106368 278099 107582 278111
rect 106491 277210 107525 277222
rect 106491 277176 106515 277210
rect 106549 277176 106583 277210
rect 106617 277176 106651 277210
rect 106685 277176 106719 277210
rect 106753 277176 106787 277210
rect 106821 277176 106855 277210
rect 106889 277176 106923 277210
rect 106957 277176 106991 277210
rect 107025 277176 107059 277210
rect 107093 277176 107127 277210
rect 107161 277176 107195 277210
rect 107229 277176 107263 277210
rect 107297 277176 107331 277210
rect 107365 277176 107399 277210
rect 107433 277176 107467 277210
rect 107501 277176 107525 277210
rect 106491 277164 107525 277176
rect 106491 277078 107525 277090
rect 106491 277044 106515 277078
rect 106549 277044 106583 277078
rect 106617 277044 106651 277078
rect 106685 277044 106719 277078
rect 106753 277044 106787 277078
rect 106821 277044 106855 277078
rect 106889 277044 106923 277078
rect 106957 277044 106991 277078
rect 107025 277044 107059 277078
rect 107093 277044 107127 277078
rect 107161 277044 107195 277078
rect 107229 277044 107263 277078
rect 107297 277044 107331 277078
rect 107365 277044 107399 277078
rect 107433 277044 107467 277078
rect 107501 277044 107525 277078
rect 106491 277032 107525 277044
rect 106951 275759 107129 275771
rect 106951 275725 106989 275759
rect 107023 275725 107057 275759
rect 107091 275725 107129 275759
rect 106951 275713 107129 275725
rect 107451 275759 107629 275771
rect 107451 275725 107489 275759
rect 107523 275725 107557 275759
rect 107591 275725 107629 275759
rect 107451 275713 107629 275725
rect 107951 275759 108129 275771
rect 107951 275725 107989 275759
rect 108023 275725 108057 275759
rect 108091 275725 108129 275759
rect 107951 275713 108129 275725
rect 108451 275759 108629 275771
rect 108451 275725 108489 275759
rect 108523 275725 108557 275759
rect 108591 275725 108629 275759
rect 108451 275713 108629 275725
rect 108951 275759 109129 275771
rect 108951 275725 108989 275759
rect 109023 275725 109057 275759
rect 109091 275725 109129 275759
rect 108951 275713 109129 275725
rect 109451 275759 109629 275771
rect 109451 275725 109489 275759
rect 109523 275725 109557 275759
rect 109591 275725 109629 275759
rect 109451 275713 109629 275725
rect 106951 274923 107129 274935
rect 106951 274889 106989 274923
rect 107023 274889 107057 274923
rect 107091 274889 107129 274923
rect 106951 274877 107129 274889
rect 107451 274923 107629 274935
rect 107451 274889 107489 274923
rect 107523 274889 107557 274923
rect 107591 274889 107629 274923
rect 107451 274877 107629 274889
rect 107951 274923 108129 274935
rect 107951 274889 107989 274923
rect 108023 274889 108057 274923
rect 108091 274889 108129 274923
rect 107951 274877 108129 274889
rect 108451 274923 108629 274935
rect 108451 274889 108489 274923
rect 108523 274889 108557 274923
rect 108591 274889 108629 274923
rect 108451 274877 108629 274889
rect 108951 274923 109129 274935
rect 108951 274889 108989 274923
rect 109023 274889 109057 274923
rect 109091 274889 109129 274923
rect 108951 274877 109129 274889
rect 109451 274923 109629 274935
rect 109451 274889 109489 274923
rect 109523 274889 109557 274923
rect 109591 274889 109629 274923
rect 109451 274877 109629 274889
rect 109240 272399 109440 272426
rect 109240 272365 109394 272399
rect 109428 272365 109440 272399
rect 109240 272331 109440 272365
rect 109240 272297 109394 272331
rect 109428 272297 109440 272331
rect 109240 272263 109440 272297
rect 109240 272229 109394 272263
rect 109428 272229 109440 272263
rect 109240 272195 109440 272229
rect 109240 272161 109394 272195
rect 109428 272161 109440 272195
rect 109240 272127 109440 272161
rect 109240 272093 109394 272127
rect 109428 272093 109440 272127
rect 109240 272059 109440 272093
rect 109240 272025 109394 272059
rect 109428 272025 109440 272059
rect 109240 271991 109440 272025
rect 109240 271957 109394 271991
rect 109428 271957 109440 271991
rect 109240 271923 109440 271957
rect 109240 271889 109394 271923
rect 109428 271889 109440 271923
rect 109240 271855 109440 271889
rect 109240 271821 109394 271855
rect 109428 271821 109440 271855
rect 109240 271787 109440 271821
rect 109240 271753 109394 271787
rect 109428 271753 109440 271787
rect 109240 271719 109440 271753
rect 109240 271685 109394 271719
rect 109428 271685 109440 271719
rect 109240 271651 109440 271685
rect 109240 271617 109394 271651
rect 109428 271617 109440 271651
rect 109240 271583 109440 271617
rect 109240 271549 109394 271583
rect 109428 271549 109440 271583
rect 109240 271515 109440 271549
rect 109240 271481 109394 271515
rect 109428 271481 109440 271515
rect 109240 271447 109440 271481
rect 109240 271413 109394 271447
rect 109428 271413 109440 271447
rect 109240 271379 109440 271413
rect 109240 271345 109394 271379
rect 109428 271345 109440 271379
rect 109240 271311 109440 271345
rect 109240 271277 109394 271311
rect 109428 271277 109440 271311
rect 109240 271243 109440 271277
rect 109240 271209 109394 271243
rect 109428 271209 109440 271243
rect 109240 271175 109440 271209
rect 109240 271141 109394 271175
rect 109428 271141 109440 271175
rect 109240 271107 109440 271141
rect 109240 271073 109394 271107
rect 109428 271073 109440 271107
rect 109240 271039 109440 271073
rect 109240 271005 109394 271039
rect 109428 271005 109440 271039
rect 109240 270971 109440 271005
rect 109240 270937 109394 270971
rect 109428 270937 109440 270971
rect 109240 270903 109440 270937
rect 109240 270869 109394 270903
rect 109428 270869 109440 270903
rect 109240 270835 109440 270869
rect 109240 270801 109394 270835
rect 109428 270801 109440 270835
rect 109240 270767 109440 270801
rect 109240 270733 109394 270767
rect 109428 270733 109440 270767
rect 109240 270706 109440 270733
rect 109510 272399 109710 272426
rect 109510 272365 109522 272399
rect 109556 272365 109710 272399
rect 109510 272331 109710 272365
rect 109510 272297 109522 272331
rect 109556 272297 109710 272331
rect 109510 272263 109710 272297
rect 109510 272229 109522 272263
rect 109556 272229 109710 272263
rect 109510 272195 109710 272229
rect 109510 272161 109522 272195
rect 109556 272161 109710 272195
rect 109510 272127 109710 272161
rect 109510 272093 109522 272127
rect 109556 272093 109710 272127
rect 109510 272059 109710 272093
rect 109510 272025 109522 272059
rect 109556 272025 109710 272059
rect 109510 271991 109710 272025
rect 109510 271957 109522 271991
rect 109556 271957 109710 271991
rect 109510 271923 109710 271957
rect 109510 271889 109522 271923
rect 109556 271889 109710 271923
rect 109510 271855 109710 271889
rect 109510 271821 109522 271855
rect 109556 271821 109710 271855
rect 109510 271787 109710 271821
rect 109510 271753 109522 271787
rect 109556 271753 109710 271787
rect 109510 271719 109710 271753
rect 109510 271685 109522 271719
rect 109556 271685 109710 271719
rect 109510 271651 109710 271685
rect 109510 271617 109522 271651
rect 109556 271617 109710 271651
rect 109510 271583 109710 271617
rect 109510 271549 109522 271583
rect 109556 271549 109710 271583
rect 109510 271515 109710 271549
rect 109510 271481 109522 271515
rect 109556 271481 109710 271515
rect 109510 271447 109710 271481
rect 109510 271413 109522 271447
rect 109556 271413 109710 271447
rect 109510 271379 109710 271413
rect 109510 271345 109522 271379
rect 109556 271345 109710 271379
rect 109510 271311 109710 271345
rect 109510 271277 109522 271311
rect 109556 271277 109710 271311
rect 109510 271243 109710 271277
rect 109510 271209 109522 271243
rect 109556 271209 109710 271243
rect 109510 271175 109710 271209
rect 109510 271141 109522 271175
rect 109556 271141 109710 271175
rect 109510 271107 109710 271141
rect 109510 271073 109522 271107
rect 109556 271073 109710 271107
rect 109510 271039 109710 271073
rect 109510 271005 109522 271039
rect 109556 271005 109710 271039
rect 109510 270971 109710 271005
rect 109510 270937 109522 270971
rect 109556 270937 109710 270971
rect 109510 270903 109710 270937
rect 109510 270869 109522 270903
rect 109556 270869 109710 270903
rect 109510 270835 109710 270869
rect 109510 270801 109522 270835
rect 109556 270801 109710 270835
rect 109510 270767 109710 270801
rect 109510 270733 109522 270767
rect 109556 270733 109710 270767
rect 109510 270706 109710 270733
rect 114657 280849 114857 280861
rect 114657 280815 114672 280849
rect 114706 280815 114740 280849
rect 114774 280815 114808 280849
rect 114842 280815 114857 280849
rect 114657 280803 114857 280815
rect 114657 280391 114857 280403
rect 114657 280357 114672 280391
rect 114706 280357 114740 280391
rect 114774 280357 114808 280391
rect 114842 280357 114857 280391
rect 114657 280345 114857 280357
rect 114657 280163 114857 280175
rect 114657 280129 114672 280163
rect 114706 280129 114740 280163
rect 114774 280129 114808 280163
rect 114842 280129 114857 280163
rect 114657 280117 114857 280129
rect 114657 279945 114857 279957
rect 114657 279911 114672 279945
rect 114706 279911 114740 279945
rect 114774 279911 114808 279945
rect 114842 279911 114857 279945
rect 114657 279899 114857 279911
rect 114657 279755 114857 279767
rect 114657 279721 114672 279755
rect 114706 279721 114740 279755
rect 114774 279721 114808 279755
rect 114842 279721 114857 279755
rect 114657 279709 114857 279721
rect 114657 279537 114857 279549
rect 114657 279503 114672 279537
rect 114706 279503 114740 279537
rect 114774 279503 114808 279537
rect 114842 279503 114857 279537
rect 114657 279491 114857 279503
rect 115348 280849 115548 280861
rect 115348 280815 115363 280849
rect 115397 280815 115431 280849
rect 115465 280815 115499 280849
rect 115533 280815 115548 280849
rect 115348 280803 115548 280815
rect 115348 280391 115548 280403
rect 115348 280357 115363 280391
rect 115397 280357 115431 280391
rect 115465 280357 115499 280391
rect 115533 280357 115548 280391
rect 115348 280345 115548 280357
rect 115348 280163 115548 280175
rect 115348 280129 115363 280163
rect 115397 280129 115431 280163
rect 115465 280129 115499 280163
rect 115533 280129 115548 280163
rect 115348 280117 115548 280129
rect 115348 279945 115548 279957
rect 115348 279911 115363 279945
rect 115397 279911 115431 279945
rect 115465 279911 115499 279945
rect 115533 279911 115548 279945
rect 115348 279899 115548 279911
rect 115348 279755 115548 279767
rect 115348 279721 115363 279755
rect 115397 279721 115431 279755
rect 115465 279721 115499 279755
rect 115533 279721 115548 279755
rect 115348 279709 115548 279721
rect 115348 279537 115548 279549
rect 115348 279503 115363 279537
rect 115397 279503 115431 279537
rect 115465 279503 115499 279537
rect 115533 279503 115548 279537
rect 115348 279491 115548 279503
rect 114657 279183 114857 279195
rect 114657 279149 114672 279183
rect 114706 279149 114740 279183
rect 114774 279149 114808 279183
rect 114842 279149 114857 279183
rect 114657 279137 114857 279149
rect 114657 278725 114857 278737
rect 114657 278691 114672 278725
rect 114706 278691 114740 278725
rect 114774 278691 114808 278725
rect 114842 278691 114857 278725
rect 114657 278679 114857 278691
rect 114657 278497 114857 278509
rect 114657 278463 114672 278497
rect 114706 278463 114740 278497
rect 114774 278463 114808 278497
rect 114842 278463 114857 278497
rect 114657 278451 114857 278463
rect 114657 278279 114857 278291
rect 114657 278245 114672 278279
rect 114706 278245 114740 278279
rect 114774 278245 114808 278279
rect 114842 278245 114857 278279
rect 114657 278233 114857 278245
rect 114657 278089 114857 278101
rect 114657 278055 114672 278089
rect 114706 278055 114740 278089
rect 114774 278055 114808 278089
rect 114842 278055 114857 278089
rect 114657 278043 114857 278055
rect 114657 277871 114857 277883
rect 114657 277837 114672 277871
rect 114706 277837 114740 277871
rect 114774 277837 114808 277871
rect 114842 277837 114857 277871
rect 114657 277825 114857 277837
rect 115348 279183 115548 279195
rect 115348 279149 115363 279183
rect 115397 279149 115431 279183
rect 115465 279149 115499 279183
rect 115533 279149 115548 279183
rect 115348 279137 115548 279149
rect 115348 278725 115548 278737
rect 115348 278691 115363 278725
rect 115397 278691 115431 278725
rect 115465 278691 115499 278725
rect 115533 278691 115548 278725
rect 115348 278679 115548 278691
rect 115348 278497 115548 278509
rect 115348 278463 115363 278497
rect 115397 278463 115431 278497
rect 115465 278463 115499 278497
rect 115533 278463 115548 278497
rect 115348 278451 115548 278463
rect 115348 278279 115548 278291
rect 115348 278245 115363 278279
rect 115397 278245 115431 278279
rect 115465 278245 115499 278279
rect 115533 278245 115548 278279
rect 115348 278233 115548 278245
rect 115348 278089 115548 278101
rect 115348 278055 115363 278089
rect 115397 278055 115431 278089
rect 115465 278055 115499 278089
rect 115533 278055 115548 278089
rect 115348 278043 115548 278055
rect 115348 277871 115548 277883
rect 115348 277837 115363 277871
rect 115397 277837 115431 277871
rect 115465 277837 115499 277871
rect 115533 277837 115548 277871
rect 115348 277825 115548 277837
rect 114657 277517 114857 277529
rect 114657 277483 114672 277517
rect 114706 277483 114740 277517
rect 114774 277483 114808 277517
rect 114842 277483 114857 277517
rect 114657 277471 114857 277483
rect 114657 277059 114857 277071
rect 114657 277025 114672 277059
rect 114706 277025 114740 277059
rect 114774 277025 114808 277059
rect 114842 277025 114857 277059
rect 114657 277013 114857 277025
rect 114657 276831 114857 276843
rect 114657 276797 114672 276831
rect 114706 276797 114740 276831
rect 114774 276797 114808 276831
rect 114842 276797 114857 276831
rect 114657 276785 114857 276797
rect 114657 276613 114857 276625
rect 114657 276579 114672 276613
rect 114706 276579 114740 276613
rect 114774 276579 114808 276613
rect 114842 276579 114857 276613
rect 114657 276567 114857 276579
rect 114657 276423 114857 276435
rect 114657 276389 114672 276423
rect 114706 276389 114740 276423
rect 114774 276389 114808 276423
rect 114842 276389 114857 276423
rect 114657 276377 114857 276389
rect 114657 276205 114857 276217
rect 114657 276171 114672 276205
rect 114706 276171 114740 276205
rect 114774 276171 114808 276205
rect 114842 276171 114857 276205
rect 114657 276159 114857 276171
rect 115348 277517 115548 277529
rect 115348 277483 115363 277517
rect 115397 277483 115431 277517
rect 115465 277483 115499 277517
rect 115533 277483 115548 277517
rect 115348 277471 115548 277483
rect 115348 277059 115548 277071
rect 115348 277025 115363 277059
rect 115397 277025 115431 277059
rect 115465 277025 115499 277059
rect 115533 277025 115548 277059
rect 115348 277013 115548 277025
rect 115348 276831 115548 276843
rect 115348 276797 115363 276831
rect 115397 276797 115431 276831
rect 115465 276797 115499 276831
rect 115533 276797 115548 276831
rect 115348 276785 115548 276797
rect 115348 276613 115548 276625
rect 115348 276579 115363 276613
rect 115397 276579 115431 276613
rect 115465 276579 115499 276613
rect 115533 276579 115548 276613
rect 115348 276567 115548 276579
rect 115348 276423 115548 276435
rect 115348 276389 115363 276423
rect 115397 276389 115431 276423
rect 115465 276389 115499 276423
rect 115533 276389 115548 276423
rect 115348 276377 115548 276389
rect 115348 276205 115548 276217
rect 115348 276171 115363 276205
rect 115397 276171 115431 276205
rect 115465 276171 115499 276205
rect 115533 276171 115548 276205
rect 115348 276159 115548 276171
rect 114657 275851 114857 275863
rect 114657 275817 114672 275851
rect 114706 275817 114740 275851
rect 114774 275817 114808 275851
rect 114842 275817 114857 275851
rect 114657 275805 114857 275817
rect 114657 275393 114857 275405
rect 114657 275359 114672 275393
rect 114706 275359 114740 275393
rect 114774 275359 114808 275393
rect 114842 275359 114857 275393
rect 114657 275347 114857 275359
rect 114657 275165 114857 275177
rect 114657 275131 114672 275165
rect 114706 275131 114740 275165
rect 114774 275131 114808 275165
rect 114842 275131 114857 275165
rect 114657 275119 114857 275131
rect 114657 274947 114857 274959
rect 114657 274913 114672 274947
rect 114706 274913 114740 274947
rect 114774 274913 114808 274947
rect 114842 274913 114857 274947
rect 114657 274901 114857 274913
rect 114657 274757 114857 274769
rect 114657 274723 114672 274757
rect 114706 274723 114740 274757
rect 114774 274723 114808 274757
rect 114842 274723 114857 274757
rect 114657 274711 114857 274723
rect 114657 274539 114857 274551
rect 114657 274505 114672 274539
rect 114706 274505 114740 274539
rect 114774 274505 114808 274539
rect 114842 274505 114857 274539
rect 114657 274493 114857 274505
rect 115348 275851 115548 275863
rect 115348 275817 115363 275851
rect 115397 275817 115431 275851
rect 115465 275817 115499 275851
rect 115533 275817 115548 275851
rect 115348 275805 115548 275817
rect 115348 275393 115548 275405
rect 115348 275359 115363 275393
rect 115397 275359 115431 275393
rect 115465 275359 115499 275393
rect 115533 275359 115548 275393
rect 115348 275347 115548 275359
rect 115348 275165 115548 275177
rect 115348 275131 115363 275165
rect 115397 275131 115431 275165
rect 115465 275131 115499 275165
rect 115533 275131 115548 275165
rect 115348 275119 115548 275131
rect 115348 274947 115548 274959
rect 115348 274913 115363 274947
rect 115397 274913 115431 274947
rect 115465 274913 115499 274947
rect 115533 274913 115548 274947
rect 115348 274901 115548 274913
rect 115348 274757 115548 274769
rect 115348 274723 115363 274757
rect 115397 274723 115431 274757
rect 115465 274723 115499 274757
rect 115533 274723 115548 274757
rect 115348 274711 115548 274723
rect 115348 274539 115548 274551
rect 115348 274505 115363 274539
rect 115397 274505 115431 274539
rect 115465 274505 115499 274539
rect 115533 274505 115548 274539
rect 115348 274493 115548 274505
rect 114657 274185 114857 274197
rect 114657 274151 114672 274185
rect 114706 274151 114740 274185
rect 114774 274151 114808 274185
rect 114842 274151 114857 274185
rect 114657 274139 114857 274151
rect 114657 273727 114857 273739
rect 114657 273693 114672 273727
rect 114706 273693 114740 273727
rect 114774 273693 114808 273727
rect 114842 273693 114857 273727
rect 114657 273681 114857 273693
rect 114657 273499 114857 273511
rect 114657 273465 114672 273499
rect 114706 273465 114740 273499
rect 114774 273465 114808 273499
rect 114842 273465 114857 273499
rect 114657 273453 114857 273465
rect 114657 273281 114857 273293
rect 114657 273247 114672 273281
rect 114706 273247 114740 273281
rect 114774 273247 114808 273281
rect 114842 273247 114857 273281
rect 114657 273235 114857 273247
rect 114657 273091 114857 273103
rect 114657 273057 114672 273091
rect 114706 273057 114740 273091
rect 114774 273057 114808 273091
rect 114842 273057 114857 273091
rect 114657 273045 114857 273057
rect 114657 272873 114857 272885
rect 114657 272839 114672 272873
rect 114706 272839 114740 272873
rect 114774 272839 114808 272873
rect 114842 272839 114857 272873
rect 114657 272827 114857 272839
rect 115348 274185 115548 274197
rect 115348 274151 115363 274185
rect 115397 274151 115431 274185
rect 115465 274151 115499 274185
rect 115533 274151 115548 274185
rect 115348 274139 115548 274151
rect 115348 273727 115548 273739
rect 115348 273693 115363 273727
rect 115397 273693 115431 273727
rect 115465 273693 115499 273727
rect 115533 273693 115548 273727
rect 115348 273681 115548 273693
rect 115348 273499 115548 273511
rect 115348 273465 115363 273499
rect 115397 273465 115431 273499
rect 115465 273465 115499 273499
rect 115533 273465 115548 273499
rect 115348 273453 115548 273465
rect 115348 273281 115548 273293
rect 115348 273247 115363 273281
rect 115397 273247 115431 273281
rect 115465 273247 115499 273281
rect 115533 273247 115548 273281
rect 115348 273235 115548 273247
rect 115348 273091 115548 273103
rect 115348 273057 115363 273091
rect 115397 273057 115431 273091
rect 115465 273057 115499 273091
rect 115533 273057 115548 273091
rect 115348 273045 115548 273057
rect 115348 272873 115548 272885
rect 115348 272839 115363 272873
rect 115397 272839 115431 272873
rect 115465 272839 115499 272873
rect 115533 272839 115548 272873
rect 115348 272827 115548 272839
rect 112520 271291 112578 271306
rect 112520 271257 112532 271291
rect 112566 271257 112578 271291
rect 112520 271223 112578 271257
rect 112520 271189 112532 271223
rect 112566 271189 112578 271223
rect 112520 271155 112578 271189
rect 112520 271121 112532 271155
rect 112566 271121 112578 271155
rect 112520 271106 112578 271121
rect 112738 271291 112796 271306
rect 112738 271257 112750 271291
rect 112784 271257 112796 271291
rect 112738 271223 112796 271257
rect 112738 271189 112750 271223
rect 112784 271189 112796 271223
rect 112738 271155 112796 271189
rect 112738 271121 112750 271155
rect 112784 271121 112796 271155
rect 112738 271106 112796 271121
rect 112920 271291 112978 271306
rect 112920 271257 112932 271291
rect 112966 271257 112978 271291
rect 112920 271223 112978 271257
rect 112920 271189 112932 271223
rect 112966 271189 112978 271223
rect 112920 271155 112978 271189
rect 112920 271121 112932 271155
rect 112966 271121 112978 271155
rect 112920 271106 112978 271121
rect 113138 271291 113196 271306
rect 113138 271257 113150 271291
rect 113184 271257 113196 271291
rect 113138 271223 113196 271257
rect 113138 271189 113150 271223
rect 113184 271189 113196 271223
rect 113138 271155 113196 271189
rect 113138 271121 113150 271155
rect 113184 271121 113196 271155
rect 113138 271106 113196 271121
rect 113320 271291 113378 271306
rect 113320 271257 113332 271291
rect 113366 271257 113378 271291
rect 113320 271223 113378 271257
rect 113320 271189 113332 271223
rect 113366 271189 113378 271223
rect 113320 271155 113378 271189
rect 113320 271121 113332 271155
rect 113366 271121 113378 271155
rect 113320 271106 113378 271121
rect 113538 271291 113596 271306
rect 113538 271257 113550 271291
rect 113584 271257 113596 271291
rect 113538 271223 113596 271257
rect 113538 271189 113550 271223
rect 113584 271189 113596 271223
rect 113538 271155 113596 271189
rect 113538 271121 113550 271155
rect 113584 271121 113596 271155
rect 113538 271106 113596 271121
rect 113720 271291 113778 271306
rect 113720 271257 113732 271291
rect 113766 271257 113778 271291
rect 113720 271223 113778 271257
rect 113720 271189 113732 271223
rect 113766 271189 113778 271223
rect 113720 271155 113778 271189
rect 113720 271121 113732 271155
rect 113766 271121 113778 271155
rect 113720 271106 113778 271121
rect 113938 271291 113996 271306
rect 113938 271257 113950 271291
rect 113984 271257 113996 271291
rect 113938 271223 113996 271257
rect 113938 271189 113950 271223
rect 113984 271189 113996 271223
rect 113938 271155 113996 271189
rect 113938 271121 113950 271155
rect 113984 271121 113996 271155
rect 113938 271106 113996 271121
rect 114579 271262 114637 271277
rect 114579 271228 114591 271262
rect 114625 271228 114637 271262
rect 114579 271194 114637 271228
rect 114579 271160 114591 271194
rect 114625 271160 114637 271194
rect 114579 271126 114637 271160
rect 114579 271092 114591 271126
rect 114625 271092 114637 271126
rect 114579 271077 114637 271092
rect 114797 271262 114855 271277
rect 114797 271228 114809 271262
rect 114843 271228 114855 271262
rect 114797 271194 114855 271228
rect 114797 271160 114809 271194
rect 114843 271160 114855 271194
rect 114797 271126 114855 271160
rect 114797 271092 114809 271126
rect 114843 271092 114855 271126
rect 114797 271077 114855 271092
rect 114979 271262 115037 271277
rect 114979 271228 114991 271262
rect 115025 271228 115037 271262
rect 114979 271194 115037 271228
rect 114979 271160 114991 271194
rect 115025 271160 115037 271194
rect 114979 271126 115037 271160
rect 114979 271092 114991 271126
rect 115025 271092 115037 271126
rect 114979 271077 115037 271092
rect 115197 271262 115255 271277
rect 115197 271228 115209 271262
rect 115243 271228 115255 271262
rect 115197 271194 115255 271228
rect 115197 271160 115209 271194
rect 115243 271160 115255 271194
rect 115197 271126 115255 271160
rect 115197 271092 115209 271126
rect 115243 271092 115255 271126
rect 115197 271077 115255 271092
rect 120371 280604 120429 280637
rect 120371 280570 120383 280604
rect 120417 280570 120429 280604
rect 120371 280537 120429 280570
rect 120829 280604 120887 280637
rect 120829 280570 120841 280604
rect 120875 280570 120887 280604
rect 120829 280537 120887 280570
rect 121071 280604 121129 280637
rect 121071 280570 121083 280604
rect 121117 280570 121129 280604
rect 121071 280537 121129 280570
rect 121529 280604 121587 280637
rect 121529 280570 121541 280604
rect 121575 280570 121587 280604
rect 121529 280537 121587 280570
rect 120371 280224 120429 280253
rect 120371 280190 120383 280224
rect 120417 280190 120429 280224
rect 120371 280156 120429 280190
rect 120371 280122 120383 280156
rect 120417 280122 120429 280156
rect 120371 280088 120429 280122
rect 120371 280054 120383 280088
rect 120417 280054 120429 280088
rect 120371 280020 120429 280054
rect 120371 279986 120383 280020
rect 120417 279986 120429 280020
rect 120371 279952 120429 279986
rect 120371 279918 120383 279952
rect 120417 279918 120429 279952
rect 120371 279884 120429 279918
rect 120371 279850 120383 279884
rect 120417 279850 120429 279884
rect 120371 279816 120429 279850
rect 120371 279782 120383 279816
rect 120417 279782 120429 279816
rect 120371 279753 120429 279782
rect 120829 280224 120887 280253
rect 120829 280190 120841 280224
rect 120875 280190 120887 280224
rect 120829 280156 120887 280190
rect 120829 280122 120841 280156
rect 120875 280122 120887 280156
rect 120829 280088 120887 280122
rect 120829 280054 120841 280088
rect 120875 280054 120887 280088
rect 120829 280020 120887 280054
rect 120829 279986 120841 280020
rect 120875 279986 120887 280020
rect 120829 279952 120887 279986
rect 120829 279918 120841 279952
rect 120875 279918 120887 279952
rect 120829 279884 120887 279918
rect 120829 279850 120841 279884
rect 120875 279850 120887 279884
rect 120829 279816 120887 279850
rect 120829 279782 120841 279816
rect 120875 279782 120887 279816
rect 120829 279753 120887 279782
rect 121071 280224 121129 280253
rect 121071 280190 121083 280224
rect 121117 280190 121129 280224
rect 121071 280156 121129 280190
rect 121071 280122 121083 280156
rect 121117 280122 121129 280156
rect 121071 280088 121129 280122
rect 121071 280054 121083 280088
rect 121117 280054 121129 280088
rect 121071 280020 121129 280054
rect 121071 279986 121083 280020
rect 121117 279986 121129 280020
rect 121071 279952 121129 279986
rect 121071 279918 121083 279952
rect 121117 279918 121129 279952
rect 121071 279884 121129 279918
rect 121071 279850 121083 279884
rect 121117 279850 121129 279884
rect 121071 279816 121129 279850
rect 121071 279782 121083 279816
rect 121117 279782 121129 279816
rect 121071 279753 121129 279782
rect 121529 280224 121587 280253
rect 121529 280190 121541 280224
rect 121575 280190 121587 280224
rect 121529 280156 121587 280190
rect 121529 280122 121541 280156
rect 121575 280122 121587 280156
rect 121529 280088 121587 280122
rect 121529 280054 121541 280088
rect 121575 280054 121587 280088
rect 121529 280020 121587 280054
rect 121529 279986 121541 280020
rect 121575 279986 121587 280020
rect 121529 279952 121587 279986
rect 121529 279918 121541 279952
rect 121575 279918 121587 279952
rect 121529 279884 121587 279918
rect 121529 279850 121541 279884
rect 121575 279850 121587 279884
rect 121529 279816 121587 279850
rect 121529 279782 121541 279816
rect 121575 279782 121587 279816
rect 121529 279753 121587 279782
rect 120371 279440 120429 279469
rect 120371 279406 120383 279440
rect 120417 279406 120429 279440
rect 120371 279372 120429 279406
rect 120371 279338 120383 279372
rect 120417 279338 120429 279372
rect 120371 279304 120429 279338
rect 120371 279270 120383 279304
rect 120417 279270 120429 279304
rect 120371 279236 120429 279270
rect 120371 279202 120383 279236
rect 120417 279202 120429 279236
rect 120371 279168 120429 279202
rect 120371 279134 120383 279168
rect 120417 279134 120429 279168
rect 120371 279100 120429 279134
rect 120371 279066 120383 279100
rect 120417 279066 120429 279100
rect 120371 279032 120429 279066
rect 120371 278998 120383 279032
rect 120417 278998 120429 279032
rect 120371 278969 120429 278998
rect 120829 279440 120887 279469
rect 120829 279406 120841 279440
rect 120875 279406 120887 279440
rect 120829 279372 120887 279406
rect 120829 279338 120841 279372
rect 120875 279338 120887 279372
rect 120829 279304 120887 279338
rect 120829 279270 120841 279304
rect 120875 279270 120887 279304
rect 120829 279236 120887 279270
rect 120829 279202 120841 279236
rect 120875 279202 120887 279236
rect 120829 279168 120887 279202
rect 120829 279134 120841 279168
rect 120875 279134 120887 279168
rect 120829 279100 120887 279134
rect 120829 279066 120841 279100
rect 120875 279066 120887 279100
rect 120829 279032 120887 279066
rect 120829 278998 120841 279032
rect 120875 278998 120887 279032
rect 120829 278969 120887 278998
rect 121071 279440 121129 279469
rect 121071 279406 121083 279440
rect 121117 279406 121129 279440
rect 121071 279372 121129 279406
rect 121071 279338 121083 279372
rect 121117 279338 121129 279372
rect 121071 279304 121129 279338
rect 121071 279270 121083 279304
rect 121117 279270 121129 279304
rect 121071 279236 121129 279270
rect 121071 279202 121083 279236
rect 121117 279202 121129 279236
rect 121071 279168 121129 279202
rect 121071 279134 121083 279168
rect 121117 279134 121129 279168
rect 121071 279100 121129 279134
rect 121071 279066 121083 279100
rect 121117 279066 121129 279100
rect 121071 279032 121129 279066
rect 121071 278998 121083 279032
rect 121117 278998 121129 279032
rect 121071 278969 121129 278998
rect 121529 279440 121587 279469
rect 121529 279406 121541 279440
rect 121575 279406 121587 279440
rect 121529 279372 121587 279406
rect 121529 279338 121541 279372
rect 121575 279338 121587 279372
rect 121529 279304 121587 279338
rect 121529 279270 121541 279304
rect 121575 279270 121587 279304
rect 121529 279236 121587 279270
rect 121529 279202 121541 279236
rect 121575 279202 121587 279236
rect 121529 279168 121587 279202
rect 121529 279134 121541 279168
rect 121575 279134 121587 279168
rect 121529 279100 121587 279134
rect 121529 279066 121541 279100
rect 121575 279066 121587 279100
rect 121529 279032 121587 279066
rect 121529 278998 121541 279032
rect 121575 278998 121587 279032
rect 121529 278969 121587 278998
rect 122298 280394 122356 280423
rect 122298 280360 122310 280394
rect 122344 280360 122356 280394
rect 122298 280326 122356 280360
rect 122298 280292 122310 280326
rect 122344 280292 122356 280326
rect 122298 280258 122356 280292
rect 122298 280224 122310 280258
rect 122344 280224 122356 280258
rect 122298 280190 122356 280224
rect 122298 280156 122310 280190
rect 122344 280156 122356 280190
rect 122298 280122 122356 280156
rect 122298 280088 122310 280122
rect 122344 280088 122356 280122
rect 122298 280054 122356 280088
rect 122298 280020 122310 280054
rect 122344 280020 122356 280054
rect 122298 279986 122356 280020
rect 122298 279952 122310 279986
rect 122344 279952 122356 279986
rect 122298 279923 122356 279952
rect 122756 280394 122814 280423
rect 122756 280360 122768 280394
rect 122802 280360 122814 280394
rect 122756 280326 122814 280360
rect 122756 280292 122768 280326
rect 122802 280292 122814 280326
rect 122756 280258 122814 280292
rect 122756 280224 122768 280258
rect 122802 280224 122814 280258
rect 122756 280190 122814 280224
rect 122756 280156 122768 280190
rect 122802 280156 122814 280190
rect 122756 280122 122814 280156
rect 122756 280088 122768 280122
rect 122802 280088 122814 280122
rect 122756 280054 122814 280088
rect 122756 280020 122768 280054
rect 122802 280020 122814 280054
rect 122756 279986 122814 280020
rect 122756 279952 122768 279986
rect 122802 279952 122814 279986
rect 122756 279923 122814 279952
rect 122998 280394 123056 280423
rect 122998 280360 123010 280394
rect 123044 280360 123056 280394
rect 122998 280326 123056 280360
rect 122998 280292 123010 280326
rect 123044 280292 123056 280326
rect 122998 280258 123056 280292
rect 122998 280224 123010 280258
rect 123044 280224 123056 280258
rect 122998 280190 123056 280224
rect 122998 280156 123010 280190
rect 123044 280156 123056 280190
rect 122998 280122 123056 280156
rect 122998 280088 123010 280122
rect 123044 280088 123056 280122
rect 122998 280054 123056 280088
rect 122998 280020 123010 280054
rect 123044 280020 123056 280054
rect 122998 279986 123056 280020
rect 122998 279952 123010 279986
rect 123044 279952 123056 279986
rect 122998 279923 123056 279952
rect 123456 280394 123514 280423
rect 123456 280360 123468 280394
rect 123502 280360 123514 280394
rect 123456 280326 123514 280360
rect 123456 280292 123468 280326
rect 123502 280292 123514 280326
rect 123456 280258 123514 280292
rect 123456 280224 123468 280258
rect 123502 280224 123514 280258
rect 123456 280190 123514 280224
rect 123456 280156 123468 280190
rect 123502 280156 123514 280190
rect 123456 280122 123514 280156
rect 123456 280088 123468 280122
rect 123502 280088 123514 280122
rect 123456 280054 123514 280088
rect 123456 280020 123468 280054
rect 123502 280020 123514 280054
rect 123456 279986 123514 280020
rect 123456 279952 123468 279986
rect 123502 279952 123514 279986
rect 123456 279923 123514 279952
rect 122298 279610 122356 279639
rect 122298 279576 122310 279610
rect 122344 279576 122356 279610
rect 122298 279542 122356 279576
rect 122298 279508 122310 279542
rect 122344 279508 122356 279542
rect 122298 279474 122356 279508
rect 122298 279440 122310 279474
rect 122344 279440 122356 279474
rect 122298 279406 122356 279440
rect 122298 279372 122310 279406
rect 122344 279372 122356 279406
rect 122298 279338 122356 279372
rect 122298 279304 122310 279338
rect 122344 279304 122356 279338
rect 122298 279270 122356 279304
rect 122298 279236 122310 279270
rect 122344 279236 122356 279270
rect 122298 279202 122356 279236
rect 122298 279168 122310 279202
rect 122344 279168 122356 279202
rect 122298 279139 122356 279168
rect 122756 279610 122814 279639
rect 122756 279576 122768 279610
rect 122802 279576 122814 279610
rect 122756 279542 122814 279576
rect 122756 279508 122768 279542
rect 122802 279508 122814 279542
rect 122756 279474 122814 279508
rect 122756 279440 122768 279474
rect 122802 279440 122814 279474
rect 122756 279406 122814 279440
rect 122756 279372 122768 279406
rect 122802 279372 122814 279406
rect 122756 279338 122814 279372
rect 122756 279304 122768 279338
rect 122802 279304 122814 279338
rect 122756 279270 122814 279304
rect 122756 279236 122768 279270
rect 122802 279236 122814 279270
rect 122756 279202 122814 279236
rect 122756 279168 122768 279202
rect 122802 279168 122814 279202
rect 122756 279139 122814 279168
rect 122998 279610 123056 279639
rect 122998 279576 123010 279610
rect 123044 279576 123056 279610
rect 122998 279542 123056 279576
rect 122998 279508 123010 279542
rect 123044 279508 123056 279542
rect 122998 279474 123056 279508
rect 122998 279440 123010 279474
rect 123044 279440 123056 279474
rect 122998 279406 123056 279440
rect 122998 279372 123010 279406
rect 123044 279372 123056 279406
rect 122998 279338 123056 279372
rect 122998 279304 123010 279338
rect 123044 279304 123056 279338
rect 122998 279270 123056 279304
rect 122998 279236 123010 279270
rect 123044 279236 123056 279270
rect 122998 279202 123056 279236
rect 122998 279168 123010 279202
rect 123044 279168 123056 279202
rect 122998 279139 123056 279168
rect 123456 279610 123514 279639
rect 123456 279576 123468 279610
rect 123502 279576 123514 279610
rect 123456 279542 123514 279576
rect 123456 279508 123468 279542
rect 123502 279508 123514 279542
rect 123456 279474 123514 279508
rect 123456 279440 123468 279474
rect 123502 279440 123514 279474
rect 123456 279406 123514 279440
rect 123456 279372 123468 279406
rect 123502 279372 123514 279406
rect 123456 279338 123514 279372
rect 123456 279304 123468 279338
rect 123502 279304 123514 279338
rect 123456 279270 123514 279304
rect 123456 279236 123468 279270
rect 123502 279236 123514 279270
rect 123456 279202 123514 279236
rect 123456 279168 123468 279202
rect 123502 279168 123514 279202
rect 123456 279139 123514 279168
rect 120371 278656 120429 278685
rect 120371 278622 120383 278656
rect 120417 278622 120429 278656
rect 120371 278588 120429 278622
rect 120371 278554 120383 278588
rect 120417 278554 120429 278588
rect 120371 278520 120429 278554
rect 120371 278486 120383 278520
rect 120417 278486 120429 278520
rect 120371 278452 120429 278486
rect 120371 278418 120383 278452
rect 120417 278418 120429 278452
rect 120371 278384 120429 278418
rect 120371 278350 120383 278384
rect 120417 278350 120429 278384
rect 120371 278316 120429 278350
rect 120371 278282 120383 278316
rect 120417 278282 120429 278316
rect 120371 278248 120429 278282
rect 120371 278214 120383 278248
rect 120417 278214 120429 278248
rect 120371 278185 120429 278214
rect 120829 278656 120887 278685
rect 120829 278622 120841 278656
rect 120875 278622 120887 278656
rect 120829 278588 120887 278622
rect 120829 278554 120841 278588
rect 120875 278554 120887 278588
rect 120829 278520 120887 278554
rect 120829 278486 120841 278520
rect 120875 278486 120887 278520
rect 120829 278452 120887 278486
rect 120829 278418 120841 278452
rect 120875 278418 120887 278452
rect 120829 278384 120887 278418
rect 120829 278350 120841 278384
rect 120875 278350 120887 278384
rect 120829 278316 120887 278350
rect 120829 278282 120841 278316
rect 120875 278282 120887 278316
rect 120829 278248 120887 278282
rect 120829 278214 120841 278248
rect 120875 278214 120887 278248
rect 120829 278185 120887 278214
rect 121071 278656 121129 278685
rect 121071 278622 121083 278656
rect 121117 278622 121129 278656
rect 121071 278588 121129 278622
rect 121071 278554 121083 278588
rect 121117 278554 121129 278588
rect 121071 278520 121129 278554
rect 121071 278486 121083 278520
rect 121117 278486 121129 278520
rect 121071 278452 121129 278486
rect 121071 278418 121083 278452
rect 121117 278418 121129 278452
rect 121071 278384 121129 278418
rect 121071 278350 121083 278384
rect 121117 278350 121129 278384
rect 121071 278316 121129 278350
rect 121071 278282 121083 278316
rect 121117 278282 121129 278316
rect 121071 278248 121129 278282
rect 121071 278214 121083 278248
rect 121117 278214 121129 278248
rect 121071 278185 121129 278214
rect 121529 278656 121587 278685
rect 121529 278622 121541 278656
rect 121575 278622 121587 278656
rect 121529 278588 121587 278622
rect 121529 278554 121541 278588
rect 121575 278554 121587 278588
rect 121529 278520 121587 278554
rect 121529 278486 121541 278520
rect 121575 278486 121587 278520
rect 121529 278452 121587 278486
rect 121529 278418 121541 278452
rect 121575 278418 121587 278452
rect 121529 278384 121587 278418
rect 121529 278350 121541 278384
rect 121575 278350 121587 278384
rect 121529 278316 121587 278350
rect 121529 278282 121541 278316
rect 121575 278282 121587 278316
rect 121529 278248 121587 278282
rect 121529 278214 121541 278248
rect 121575 278214 121587 278248
rect 121529 278185 121587 278214
rect 120371 277872 120429 277901
rect 120371 277838 120383 277872
rect 120417 277838 120429 277872
rect 120371 277804 120429 277838
rect 120371 277770 120383 277804
rect 120417 277770 120429 277804
rect 120371 277736 120429 277770
rect 120371 277702 120383 277736
rect 120417 277702 120429 277736
rect 120371 277668 120429 277702
rect 120371 277634 120383 277668
rect 120417 277634 120429 277668
rect 120371 277600 120429 277634
rect 120371 277566 120383 277600
rect 120417 277566 120429 277600
rect 120371 277532 120429 277566
rect 120371 277498 120383 277532
rect 120417 277498 120429 277532
rect 120371 277464 120429 277498
rect 120371 277430 120383 277464
rect 120417 277430 120429 277464
rect 120371 277401 120429 277430
rect 120829 277872 120887 277901
rect 120829 277838 120841 277872
rect 120875 277838 120887 277872
rect 120829 277804 120887 277838
rect 120829 277770 120841 277804
rect 120875 277770 120887 277804
rect 120829 277736 120887 277770
rect 120829 277702 120841 277736
rect 120875 277702 120887 277736
rect 120829 277668 120887 277702
rect 120829 277634 120841 277668
rect 120875 277634 120887 277668
rect 120829 277600 120887 277634
rect 120829 277566 120841 277600
rect 120875 277566 120887 277600
rect 120829 277532 120887 277566
rect 120829 277498 120841 277532
rect 120875 277498 120887 277532
rect 120829 277464 120887 277498
rect 120829 277430 120841 277464
rect 120875 277430 120887 277464
rect 120829 277401 120887 277430
rect 121071 277872 121129 277901
rect 121071 277838 121083 277872
rect 121117 277838 121129 277872
rect 121071 277804 121129 277838
rect 121071 277770 121083 277804
rect 121117 277770 121129 277804
rect 121071 277736 121129 277770
rect 121071 277702 121083 277736
rect 121117 277702 121129 277736
rect 121071 277668 121129 277702
rect 121071 277634 121083 277668
rect 121117 277634 121129 277668
rect 121071 277600 121129 277634
rect 121071 277566 121083 277600
rect 121117 277566 121129 277600
rect 121071 277532 121129 277566
rect 121071 277498 121083 277532
rect 121117 277498 121129 277532
rect 121071 277464 121129 277498
rect 121071 277430 121083 277464
rect 121117 277430 121129 277464
rect 121071 277401 121129 277430
rect 121529 277872 121587 277901
rect 121529 277838 121541 277872
rect 121575 277838 121587 277872
rect 121529 277804 121587 277838
rect 121529 277770 121541 277804
rect 121575 277770 121587 277804
rect 121529 277736 121587 277770
rect 121529 277702 121541 277736
rect 121575 277702 121587 277736
rect 121529 277668 121587 277702
rect 121529 277634 121541 277668
rect 121575 277634 121587 277668
rect 121529 277600 121587 277634
rect 121529 277566 121541 277600
rect 121575 277566 121587 277600
rect 121529 277532 121587 277566
rect 121529 277498 121541 277532
rect 121575 277498 121587 277532
rect 121529 277464 121587 277498
rect 121529 277430 121541 277464
rect 121575 277430 121587 277464
rect 121529 277401 121587 277430
rect 120371 277088 120429 277117
rect 120371 277054 120383 277088
rect 120417 277054 120429 277088
rect 120371 277020 120429 277054
rect 120371 276986 120383 277020
rect 120417 276986 120429 277020
rect 120371 276952 120429 276986
rect 120371 276918 120383 276952
rect 120417 276918 120429 276952
rect 120371 276884 120429 276918
rect 120371 276850 120383 276884
rect 120417 276850 120429 276884
rect 120371 276816 120429 276850
rect 120371 276782 120383 276816
rect 120417 276782 120429 276816
rect 120371 276748 120429 276782
rect 120371 276714 120383 276748
rect 120417 276714 120429 276748
rect 120371 276680 120429 276714
rect 120371 276646 120383 276680
rect 120417 276646 120429 276680
rect 120371 276617 120429 276646
rect 120829 277088 120887 277117
rect 120829 277054 120841 277088
rect 120875 277054 120887 277088
rect 120829 277020 120887 277054
rect 120829 276986 120841 277020
rect 120875 276986 120887 277020
rect 120829 276952 120887 276986
rect 120829 276918 120841 276952
rect 120875 276918 120887 276952
rect 120829 276884 120887 276918
rect 120829 276850 120841 276884
rect 120875 276850 120887 276884
rect 120829 276816 120887 276850
rect 120829 276782 120841 276816
rect 120875 276782 120887 276816
rect 120829 276748 120887 276782
rect 120829 276714 120841 276748
rect 120875 276714 120887 276748
rect 120829 276680 120887 276714
rect 120829 276646 120841 276680
rect 120875 276646 120887 276680
rect 120829 276617 120887 276646
rect 121071 277088 121129 277117
rect 121071 277054 121083 277088
rect 121117 277054 121129 277088
rect 121071 277020 121129 277054
rect 121071 276986 121083 277020
rect 121117 276986 121129 277020
rect 121071 276952 121129 276986
rect 121071 276918 121083 276952
rect 121117 276918 121129 276952
rect 121071 276884 121129 276918
rect 121071 276850 121083 276884
rect 121117 276850 121129 276884
rect 121071 276816 121129 276850
rect 121071 276782 121083 276816
rect 121117 276782 121129 276816
rect 121071 276748 121129 276782
rect 121071 276714 121083 276748
rect 121117 276714 121129 276748
rect 121071 276680 121129 276714
rect 121071 276646 121083 276680
rect 121117 276646 121129 276680
rect 121071 276617 121129 276646
rect 121529 277088 121587 277117
rect 121529 277054 121541 277088
rect 121575 277054 121587 277088
rect 121529 277020 121587 277054
rect 121529 276986 121541 277020
rect 121575 276986 121587 277020
rect 121529 276952 121587 276986
rect 121529 276918 121541 276952
rect 121575 276918 121587 276952
rect 121529 276884 121587 276918
rect 121529 276850 121541 276884
rect 121575 276850 121587 276884
rect 121529 276816 121587 276850
rect 121529 276782 121541 276816
rect 121575 276782 121587 276816
rect 121529 276748 121587 276782
rect 121529 276714 121541 276748
rect 121575 276714 121587 276748
rect 121529 276680 121587 276714
rect 121529 276646 121541 276680
rect 121575 276646 121587 276680
rect 121529 276617 121587 276646
rect 120371 276304 120429 276333
rect 120371 276270 120383 276304
rect 120417 276270 120429 276304
rect 120371 276236 120429 276270
rect 120371 276202 120383 276236
rect 120417 276202 120429 276236
rect 120371 276168 120429 276202
rect 120371 276134 120383 276168
rect 120417 276134 120429 276168
rect 120371 276100 120429 276134
rect 120371 276066 120383 276100
rect 120417 276066 120429 276100
rect 120371 276032 120429 276066
rect 120371 275998 120383 276032
rect 120417 275998 120429 276032
rect 120371 275964 120429 275998
rect 120371 275930 120383 275964
rect 120417 275930 120429 275964
rect 120371 275896 120429 275930
rect 120371 275862 120383 275896
rect 120417 275862 120429 275896
rect 120371 275833 120429 275862
rect 120829 276304 120887 276333
rect 120829 276270 120841 276304
rect 120875 276270 120887 276304
rect 120829 276236 120887 276270
rect 120829 276202 120841 276236
rect 120875 276202 120887 276236
rect 120829 276168 120887 276202
rect 120829 276134 120841 276168
rect 120875 276134 120887 276168
rect 120829 276100 120887 276134
rect 120829 276066 120841 276100
rect 120875 276066 120887 276100
rect 120829 276032 120887 276066
rect 120829 275998 120841 276032
rect 120875 275998 120887 276032
rect 120829 275964 120887 275998
rect 120829 275930 120841 275964
rect 120875 275930 120887 275964
rect 120829 275896 120887 275930
rect 120829 275862 120841 275896
rect 120875 275862 120887 275896
rect 120829 275833 120887 275862
rect 121071 276304 121129 276333
rect 121071 276270 121083 276304
rect 121117 276270 121129 276304
rect 121071 276236 121129 276270
rect 121071 276202 121083 276236
rect 121117 276202 121129 276236
rect 121071 276168 121129 276202
rect 121071 276134 121083 276168
rect 121117 276134 121129 276168
rect 121071 276100 121129 276134
rect 121071 276066 121083 276100
rect 121117 276066 121129 276100
rect 121071 276032 121129 276066
rect 121071 275998 121083 276032
rect 121117 275998 121129 276032
rect 121071 275964 121129 275998
rect 121071 275930 121083 275964
rect 121117 275930 121129 275964
rect 121071 275896 121129 275930
rect 121071 275862 121083 275896
rect 121117 275862 121129 275896
rect 121071 275833 121129 275862
rect 121529 276304 121587 276333
rect 121529 276270 121541 276304
rect 121575 276270 121587 276304
rect 121529 276236 121587 276270
rect 121529 276202 121541 276236
rect 121575 276202 121587 276236
rect 121529 276168 121587 276202
rect 121529 276134 121541 276168
rect 121575 276134 121587 276168
rect 121529 276100 121587 276134
rect 121529 276066 121541 276100
rect 121575 276066 121587 276100
rect 121529 276032 121587 276066
rect 121529 275998 121541 276032
rect 121575 275998 121587 276032
rect 121529 275964 121587 275998
rect 121529 275930 121541 275964
rect 121575 275930 121587 275964
rect 121529 275896 121587 275930
rect 121529 275862 121541 275896
rect 121575 275862 121587 275896
rect 121529 275833 121587 275862
rect 120371 275520 120429 275549
rect 120371 275486 120383 275520
rect 120417 275486 120429 275520
rect 120371 275452 120429 275486
rect 120371 275418 120383 275452
rect 120417 275418 120429 275452
rect 120371 275384 120429 275418
rect 120371 275350 120383 275384
rect 120417 275350 120429 275384
rect 120371 275316 120429 275350
rect 120371 275282 120383 275316
rect 120417 275282 120429 275316
rect 120371 275248 120429 275282
rect 120371 275214 120383 275248
rect 120417 275214 120429 275248
rect 120371 275180 120429 275214
rect 120371 275146 120383 275180
rect 120417 275146 120429 275180
rect 120371 275112 120429 275146
rect 120371 275078 120383 275112
rect 120417 275078 120429 275112
rect 120371 275049 120429 275078
rect 120829 275520 120887 275549
rect 120829 275486 120841 275520
rect 120875 275486 120887 275520
rect 120829 275452 120887 275486
rect 120829 275418 120841 275452
rect 120875 275418 120887 275452
rect 120829 275384 120887 275418
rect 120829 275350 120841 275384
rect 120875 275350 120887 275384
rect 120829 275316 120887 275350
rect 120829 275282 120841 275316
rect 120875 275282 120887 275316
rect 120829 275248 120887 275282
rect 120829 275214 120841 275248
rect 120875 275214 120887 275248
rect 120829 275180 120887 275214
rect 120829 275146 120841 275180
rect 120875 275146 120887 275180
rect 120829 275112 120887 275146
rect 120829 275078 120841 275112
rect 120875 275078 120887 275112
rect 120829 275049 120887 275078
rect 121071 275520 121129 275549
rect 121071 275486 121083 275520
rect 121117 275486 121129 275520
rect 121071 275452 121129 275486
rect 121071 275418 121083 275452
rect 121117 275418 121129 275452
rect 121071 275384 121129 275418
rect 121071 275350 121083 275384
rect 121117 275350 121129 275384
rect 121071 275316 121129 275350
rect 121071 275282 121083 275316
rect 121117 275282 121129 275316
rect 121071 275248 121129 275282
rect 121071 275214 121083 275248
rect 121117 275214 121129 275248
rect 121071 275180 121129 275214
rect 121071 275146 121083 275180
rect 121117 275146 121129 275180
rect 121071 275112 121129 275146
rect 121071 275078 121083 275112
rect 121117 275078 121129 275112
rect 121071 275049 121129 275078
rect 121529 275520 121587 275549
rect 121529 275486 121541 275520
rect 121575 275486 121587 275520
rect 121529 275452 121587 275486
rect 121529 275418 121541 275452
rect 121575 275418 121587 275452
rect 121529 275384 121587 275418
rect 121529 275350 121541 275384
rect 121575 275350 121587 275384
rect 121529 275316 121587 275350
rect 121529 275282 121541 275316
rect 121575 275282 121587 275316
rect 121529 275248 121587 275282
rect 121529 275214 121541 275248
rect 121575 275214 121587 275248
rect 121529 275180 121587 275214
rect 121529 275146 121541 275180
rect 121575 275146 121587 275180
rect 121529 275112 121587 275146
rect 121529 275078 121541 275112
rect 121575 275078 121587 275112
rect 121529 275049 121587 275078
rect 122356 278250 122414 278266
rect 122356 278216 122368 278250
rect 122402 278216 122414 278250
rect 122356 278182 122414 278216
rect 122356 278148 122368 278182
rect 122402 278148 122414 278182
rect 122356 278114 122414 278148
rect 122356 278080 122368 278114
rect 122402 278080 122414 278114
rect 122356 278046 122414 278080
rect 122356 278012 122368 278046
rect 122402 278012 122414 278046
rect 122356 277978 122414 278012
rect 122356 277944 122368 277978
rect 122402 277944 122414 277978
rect 122356 277910 122414 277944
rect 122356 277876 122368 277910
rect 122402 277876 122414 277910
rect 122356 277842 122414 277876
rect 122356 277808 122368 277842
rect 122402 277808 122414 277842
rect 122356 277792 122414 277808
rect 123290 278250 123348 278266
rect 123290 278216 123302 278250
rect 123336 278216 123348 278250
rect 123290 278182 123348 278216
rect 123290 278148 123302 278182
rect 123336 278148 123348 278182
rect 123290 278114 123348 278148
rect 123290 278080 123302 278114
rect 123336 278080 123348 278114
rect 123290 278046 123348 278080
rect 123290 278012 123302 278046
rect 123336 278012 123348 278046
rect 123290 277978 123348 278012
rect 123290 277944 123302 277978
rect 123336 277944 123348 277978
rect 123290 277910 123348 277944
rect 123290 277876 123302 277910
rect 123336 277876 123348 277910
rect 123290 277842 123348 277876
rect 123290 277808 123302 277842
rect 123336 277808 123348 277842
rect 123290 277792 123348 277808
rect 123598 278060 123656 278080
rect 123598 278026 123610 278060
rect 123644 278026 123656 278060
rect 123598 277992 123656 278026
rect 123598 277958 123610 277992
rect 123644 277958 123656 277992
rect 123598 277924 123656 277958
rect 123598 277890 123610 277924
rect 123644 277890 123656 277924
rect 123598 277856 123656 277890
rect 123598 277822 123610 277856
rect 123644 277822 123656 277856
rect 123598 277788 123656 277822
rect 123598 277754 123610 277788
rect 123644 277754 123656 277788
rect 123598 277720 123656 277754
rect 123598 277686 123610 277720
rect 123644 277686 123656 277720
rect 123598 277652 123656 277686
rect 123598 277618 123610 277652
rect 123644 277618 123656 277652
rect 123598 277584 123656 277618
rect 123598 277550 123610 277584
rect 123644 277550 123656 277584
rect 123598 277516 123656 277550
rect 122358 277467 122416 277500
rect 122358 277433 122370 277467
rect 122404 277433 122416 277467
rect 122358 277400 122416 277433
rect 123216 277467 123274 277500
rect 123216 277433 123228 277467
rect 123262 277433 123274 277467
rect 123216 277400 123274 277433
rect 123598 277482 123610 277516
rect 123644 277482 123656 277516
rect 123598 277448 123656 277482
rect 123598 277414 123610 277448
rect 123644 277414 123656 277448
rect 123598 277394 123656 277414
rect 124210 278060 124268 278080
rect 124210 278026 124222 278060
rect 124256 278026 124268 278060
rect 124210 277992 124268 278026
rect 124210 277958 124222 277992
rect 124256 277958 124268 277992
rect 124210 277924 124268 277958
rect 124210 277890 124222 277924
rect 124256 277890 124268 277924
rect 124210 277856 124268 277890
rect 124210 277822 124222 277856
rect 124256 277822 124268 277856
rect 124210 277788 124268 277822
rect 124210 277754 124222 277788
rect 124256 277754 124268 277788
rect 124210 277720 124268 277754
rect 124210 277686 124222 277720
rect 124256 277686 124268 277720
rect 124210 277652 124268 277686
rect 124210 277618 124222 277652
rect 124256 277618 124268 277652
rect 124210 277584 124268 277618
rect 124210 277550 124222 277584
rect 124256 277550 124268 277584
rect 124210 277516 124268 277550
rect 124210 277482 124222 277516
rect 124256 277482 124268 277516
rect 124210 277448 124268 277482
rect 124210 277414 124222 277448
rect 124256 277414 124268 277448
rect 124210 277394 124268 277414
rect 122380 276631 122438 276668
rect 122380 276597 122392 276631
rect 122426 276597 122438 276631
rect 122380 276563 122438 276597
rect 122380 276529 122392 276563
rect 122426 276529 122438 276563
rect 122380 276492 122438 276529
rect 123832 276631 123890 276668
rect 123832 276597 123844 276631
rect 123878 276597 123890 276631
rect 123832 276563 123890 276597
rect 123832 276529 123844 276563
rect 123878 276529 123890 276563
rect 123832 276492 123890 276529
rect 122466 275857 122866 275869
rect 122466 275823 122479 275857
rect 122513 275823 122547 275857
rect 122581 275823 122615 275857
rect 122649 275823 122683 275857
rect 122717 275823 122751 275857
rect 122785 275823 122819 275857
rect 122853 275823 122866 275857
rect 122466 275811 122866 275823
rect 123102 275857 123502 275869
rect 123102 275823 123115 275857
rect 123149 275823 123183 275857
rect 123217 275823 123251 275857
rect 123285 275823 123319 275857
rect 123353 275823 123387 275857
rect 123421 275823 123455 275857
rect 123489 275823 123502 275857
rect 123102 275811 123502 275823
rect 123738 275857 124138 275869
rect 123738 275823 123751 275857
rect 123785 275823 123819 275857
rect 123853 275823 123887 275857
rect 123921 275823 123955 275857
rect 123989 275823 124023 275857
rect 124057 275823 124091 275857
rect 124125 275823 124138 275857
rect 123738 275811 124138 275823
rect 124374 275857 124774 275869
rect 124374 275823 124387 275857
rect 124421 275823 124455 275857
rect 124489 275823 124523 275857
rect 124557 275823 124591 275857
rect 124625 275823 124659 275857
rect 124693 275823 124727 275857
rect 124761 275823 124774 275857
rect 124374 275811 124774 275823
rect 122466 275699 122866 275711
rect 122466 275665 122479 275699
rect 122513 275665 122547 275699
rect 122581 275665 122615 275699
rect 122649 275665 122683 275699
rect 122717 275665 122751 275699
rect 122785 275665 122819 275699
rect 122853 275665 122866 275699
rect 122466 275653 122866 275665
rect 123102 275699 123502 275711
rect 123102 275665 123115 275699
rect 123149 275665 123183 275699
rect 123217 275665 123251 275699
rect 123285 275665 123319 275699
rect 123353 275665 123387 275699
rect 123421 275665 123455 275699
rect 123489 275665 123502 275699
rect 123102 275653 123502 275665
rect 123738 275699 124138 275711
rect 123738 275665 123751 275699
rect 123785 275665 123819 275699
rect 123853 275665 123887 275699
rect 123921 275665 123955 275699
rect 123989 275665 124023 275699
rect 124057 275665 124091 275699
rect 124125 275665 124138 275699
rect 123738 275653 124138 275665
rect 124374 275699 124774 275711
rect 124374 275665 124387 275699
rect 124421 275665 124455 275699
rect 124489 275665 124523 275699
rect 124557 275665 124591 275699
rect 124625 275665 124659 275699
rect 124693 275665 124727 275699
rect 124761 275665 124774 275699
rect 124374 275653 124774 275665
rect 120371 274736 120429 274765
rect 120371 274702 120383 274736
rect 120417 274702 120429 274736
rect 120371 274668 120429 274702
rect 120371 274634 120383 274668
rect 120417 274634 120429 274668
rect 120371 274600 120429 274634
rect 120371 274566 120383 274600
rect 120417 274566 120429 274600
rect 120371 274532 120429 274566
rect 120371 274498 120383 274532
rect 120417 274498 120429 274532
rect 120371 274464 120429 274498
rect 120371 274430 120383 274464
rect 120417 274430 120429 274464
rect 120371 274396 120429 274430
rect 120371 274362 120383 274396
rect 120417 274362 120429 274396
rect 120371 274328 120429 274362
rect 120371 274294 120383 274328
rect 120417 274294 120429 274328
rect 120371 274265 120429 274294
rect 120829 274736 120887 274765
rect 120829 274702 120841 274736
rect 120875 274702 120887 274736
rect 120829 274668 120887 274702
rect 120829 274634 120841 274668
rect 120875 274634 120887 274668
rect 120829 274600 120887 274634
rect 120829 274566 120841 274600
rect 120875 274566 120887 274600
rect 120829 274532 120887 274566
rect 120829 274498 120841 274532
rect 120875 274498 120887 274532
rect 120829 274464 120887 274498
rect 120829 274430 120841 274464
rect 120875 274430 120887 274464
rect 120829 274396 120887 274430
rect 120829 274362 120841 274396
rect 120875 274362 120887 274396
rect 120829 274328 120887 274362
rect 120829 274294 120841 274328
rect 120875 274294 120887 274328
rect 120829 274265 120887 274294
rect 121071 274736 121129 274765
rect 121071 274702 121083 274736
rect 121117 274702 121129 274736
rect 121071 274668 121129 274702
rect 121071 274634 121083 274668
rect 121117 274634 121129 274668
rect 121071 274600 121129 274634
rect 121071 274566 121083 274600
rect 121117 274566 121129 274600
rect 121071 274532 121129 274566
rect 121071 274498 121083 274532
rect 121117 274498 121129 274532
rect 121071 274464 121129 274498
rect 121071 274430 121083 274464
rect 121117 274430 121129 274464
rect 121071 274396 121129 274430
rect 121071 274362 121083 274396
rect 121117 274362 121129 274396
rect 121071 274328 121129 274362
rect 121071 274294 121083 274328
rect 121117 274294 121129 274328
rect 121071 274265 121129 274294
rect 121529 274736 121587 274765
rect 121529 274702 121541 274736
rect 121575 274702 121587 274736
rect 121529 274668 121587 274702
rect 121529 274634 121541 274668
rect 121575 274634 121587 274668
rect 121529 274600 121587 274634
rect 121529 274566 121541 274600
rect 121575 274566 121587 274600
rect 121529 274532 121587 274566
rect 121529 274498 121541 274532
rect 121575 274498 121587 274532
rect 121529 274464 121587 274498
rect 121529 274430 121541 274464
rect 121575 274430 121587 274464
rect 121529 274396 121587 274430
rect 121529 274362 121541 274396
rect 121575 274362 121587 274396
rect 121529 274328 121587 274362
rect 121529 274294 121541 274328
rect 121575 274294 121587 274328
rect 121529 274265 121587 274294
rect 120371 273952 120429 273981
rect 120371 273918 120383 273952
rect 120417 273918 120429 273952
rect 120371 273884 120429 273918
rect 120371 273850 120383 273884
rect 120417 273850 120429 273884
rect 120371 273816 120429 273850
rect 120371 273782 120383 273816
rect 120417 273782 120429 273816
rect 120371 273748 120429 273782
rect 120371 273714 120383 273748
rect 120417 273714 120429 273748
rect 120371 273680 120429 273714
rect 120371 273646 120383 273680
rect 120417 273646 120429 273680
rect 120371 273612 120429 273646
rect 120371 273578 120383 273612
rect 120417 273578 120429 273612
rect 120371 273544 120429 273578
rect 120371 273510 120383 273544
rect 120417 273510 120429 273544
rect 120371 273481 120429 273510
rect 120829 273952 120887 273981
rect 120829 273918 120841 273952
rect 120875 273918 120887 273952
rect 120829 273884 120887 273918
rect 120829 273850 120841 273884
rect 120875 273850 120887 273884
rect 120829 273816 120887 273850
rect 120829 273782 120841 273816
rect 120875 273782 120887 273816
rect 120829 273748 120887 273782
rect 120829 273714 120841 273748
rect 120875 273714 120887 273748
rect 120829 273680 120887 273714
rect 120829 273646 120841 273680
rect 120875 273646 120887 273680
rect 120829 273612 120887 273646
rect 120829 273578 120841 273612
rect 120875 273578 120887 273612
rect 120829 273544 120887 273578
rect 120829 273510 120841 273544
rect 120875 273510 120887 273544
rect 120829 273481 120887 273510
rect 121071 273952 121129 273981
rect 121071 273918 121083 273952
rect 121117 273918 121129 273952
rect 121071 273884 121129 273918
rect 121071 273850 121083 273884
rect 121117 273850 121129 273884
rect 121071 273816 121129 273850
rect 121071 273782 121083 273816
rect 121117 273782 121129 273816
rect 121071 273748 121129 273782
rect 121071 273714 121083 273748
rect 121117 273714 121129 273748
rect 121071 273680 121129 273714
rect 121071 273646 121083 273680
rect 121117 273646 121129 273680
rect 121071 273612 121129 273646
rect 121071 273578 121083 273612
rect 121117 273578 121129 273612
rect 121071 273544 121129 273578
rect 121071 273510 121083 273544
rect 121117 273510 121129 273544
rect 121071 273481 121129 273510
rect 121529 273952 121587 273981
rect 121529 273918 121541 273952
rect 121575 273918 121587 273952
rect 121529 273884 121587 273918
rect 121529 273850 121541 273884
rect 121575 273850 121587 273884
rect 121529 273816 121587 273850
rect 121529 273782 121541 273816
rect 121575 273782 121587 273816
rect 121529 273748 121587 273782
rect 121529 273714 121541 273748
rect 121575 273714 121587 273748
rect 121529 273680 121587 273714
rect 121529 273646 121541 273680
rect 121575 273646 121587 273680
rect 121529 273612 121587 273646
rect 121529 273578 121541 273612
rect 121575 273578 121587 273612
rect 121529 273544 121587 273578
rect 121529 273510 121541 273544
rect 121575 273510 121587 273544
rect 121529 273481 121587 273510
rect 120371 273168 120429 273197
rect 120371 273134 120383 273168
rect 120417 273134 120429 273168
rect 120371 273100 120429 273134
rect 120371 273066 120383 273100
rect 120417 273066 120429 273100
rect 120371 273032 120429 273066
rect 120371 272998 120383 273032
rect 120417 272998 120429 273032
rect 120371 272964 120429 272998
rect 120371 272930 120383 272964
rect 120417 272930 120429 272964
rect 120371 272896 120429 272930
rect 120371 272862 120383 272896
rect 120417 272862 120429 272896
rect 120371 272828 120429 272862
rect 120371 272794 120383 272828
rect 120417 272794 120429 272828
rect 120371 272760 120429 272794
rect 120371 272726 120383 272760
rect 120417 272726 120429 272760
rect 120371 272697 120429 272726
rect 120829 273168 120887 273197
rect 120829 273134 120841 273168
rect 120875 273134 120887 273168
rect 120829 273100 120887 273134
rect 120829 273066 120841 273100
rect 120875 273066 120887 273100
rect 120829 273032 120887 273066
rect 120829 272998 120841 273032
rect 120875 272998 120887 273032
rect 120829 272964 120887 272998
rect 120829 272930 120841 272964
rect 120875 272930 120887 272964
rect 120829 272896 120887 272930
rect 120829 272862 120841 272896
rect 120875 272862 120887 272896
rect 120829 272828 120887 272862
rect 120829 272794 120841 272828
rect 120875 272794 120887 272828
rect 120829 272760 120887 272794
rect 120829 272726 120841 272760
rect 120875 272726 120887 272760
rect 120829 272697 120887 272726
rect 121071 273168 121129 273197
rect 121071 273134 121083 273168
rect 121117 273134 121129 273168
rect 121071 273100 121129 273134
rect 121071 273066 121083 273100
rect 121117 273066 121129 273100
rect 121071 273032 121129 273066
rect 121071 272998 121083 273032
rect 121117 272998 121129 273032
rect 121071 272964 121129 272998
rect 121071 272930 121083 272964
rect 121117 272930 121129 272964
rect 121071 272896 121129 272930
rect 121071 272862 121083 272896
rect 121117 272862 121129 272896
rect 121071 272828 121129 272862
rect 121071 272794 121083 272828
rect 121117 272794 121129 272828
rect 121071 272760 121129 272794
rect 121071 272726 121083 272760
rect 121117 272726 121129 272760
rect 121071 272697 121129 272726
rect 121529 273168 121587 273197
rect 121529 273134 121541 273168
rect 121575 273134 121587 273168
rect 121529 273100 121587 273134
rect 121529 273066 121541 273100
rect 121575 273066 121587 273100
rect 121529 273032 121587 273066
rect 121529 272998 121541 273032
rect 121575 272998 121587 273032
rect 121529 272964 121587 272998
rect 121529 272930 121541 272964
rect 121575 272930 121587 272964
rect 121529 272896 121587 272930
rect 121529 272862 121541 272896
rect 121575 272862 121587 272896
rect 121529 272828 121587 272862
rect 121529 272794 121541 272828
rect 121575 272794 121587 272828
rect 121529 272760 121587 272794
rect 121529 272726 121541 272760
rect 121575 272726 121587 272760
rect 121529 272697 121587 272726
rect 120371 272384 120429 272413
rect 120371 272350 120383 272384
rect 120417 272350 120429 272384
rect 120371 272316 120429 272350
rect 120371 272282 120383 272316
rect 120417 272282 120429 272316
rect 120371 272248 120429 272282
rect 120371 272214 120383 272248
rect 120417 272214 120429 272248
rect 120371 272180 120429 272214
rect 120371 272146 120383 272180
rect 120417 272146 120429 272180
rect 120371 272112 120429 272146
rect 120371 272078 120383 272112
rect 120417 272078 120429 272112
rect 120371 272044 120429 272078
rect 120371 272010 120383 272044
rect 120417 272010 120429 272044
rect 120371 271976 120429 272010
rect 120371 271942 120383 271976
rect 120417 271942 120429 271976
rect 120371 271913 120429 271942
rect 120829 272384 120887 272413
rect 120829 272350 120841 272384
rect 120875 272350 120887 272384
rect 120829 272316 120887 272350
rect 120829 272282 120841 272316
rect 120875 272282 120887 272316
rect 120829 272248 120887 272282
rect 120829 272214 120841 272248
rect 120875 272214 120887 272248
rect 120829 272180 120887 272214
rect 120829 272146 120841 272180
rect 120875 272146 120887 272180
rect 120829 272112 120887 272146
rect 120829 272078 120841 272112
rect 120875 272078 120887 272112
rect 120829 272044 120887 272078
rect 120829 272010 120841 272044
rect 120875 272010 120887 272044
rect 120829 271976 120887 272010
rect 120829 271942 120841 271976
rect 120875 271942 120887 271976
rect 120829 271913 120887 271942
rect 121071 272384 121129 272413
rect 121071 272350 121083 272384
rect 121117 272350 121129 272384
rect 121071 272316 121129 272350
rect 121071 272282 121083 272316
rect 121117 272282 121129 272316
rect 121071 272248 121129 272282
rect 121071 272214 121083 272248
rect 121117 272214 121129 272248
rect 121071 272180 121129 272214
rect 121071 272146 121083 272180
rect 121117 272146 121129 272180
rect 121071 272112 121129 272146
rect 121071 272078 121083 272112
rect 121117 272078 121129 272112
rect 121071 272044 121129 272078
rect 121071 272010 121083 272044
rect 121117 272010 121129 272044
rect 121071 271976 121129 272010
rect 121071 271942 121083 271976
rect 121117 271942 121129 271976
rect 121071 271913 121129 271942
rect 121529 272384 121587 272413
rect 121529 272350 121541 272384
rect 121575 272350 121587 272384
rect 121529 272316 121587 272350
rect 121529 272282 121541 272316
rect 121575 272282 121587 272316
rect 121529 272248 121587 272282
rect 121529 272214 121541 272248
rect 121575 272214 121587 272248
rect 121529 272180 121587 272214
rect 121529 272146 121541 272180
rect 121575 272146 121587 272180
rect 121529 272112 121587 272146
rect 121529 272078 121541 272112
rect 121575 272078 121587 272112
rect 121529 272044 121587 272078
rect 121529 272010 121541 272044
rect 121575 272010 121587 272044
rect 121529 271976 121587 272010
rect 121529 271942 121541 271976
rect 121575 271942 121587 271976
rect 121529 271913 121587 271942
rect 120371 271600 120429 271629
rect 120371 271566 120383 271600
rect 120417 271566 120429 271600
rect 120371 271532 120429 271566
rect 120371 271498 120383 271532
rect 120417 271498 120429 271532
rect 120371 271464 120429 271498
rect 120371 271430 120383 271464
rect 120417 271430 120429 271464
rect 120371 271396 120429 271430
rect 120371 271362 120383 271396
rect 120417 271362 120429 271396
rect 120371 271328 120429 271362
rect 120371 271294 120383 271328
rect 120417 271294 120429 271328
rect 120371 271260 120429 271294
rect 120371 271226 120383 271260
rect 120417 271226 120429 271260
rect 120371 271192 120429 271226
rect 120371 271158 120383 271192
rect 120417 271158 120429 271192
rect 120371 271129 120429 271158
rect 120829 271600 120887 271629
rect 120829 271566 120841 271600
rect 120875 271566 120887 271600
rect 120829 271532 120887 271566
rect 120829 271498 120841 271532
rect 120875 271498 120887 271532
rect 120829 271464 120887 271498
rect 120829 271430 120841 271464
rect 120875 271430 120887 271464
rect 120829 271396 120887 271430
rect 120829 271362 120841 271396
rect 120875 271362 120887 271396
rect 120829 271328 120887 271362
rect 120829 271294 120841 271328
rect 120875 271294 120887 271328
rect 120829 271260 120887 271294
rect 120829 271226 120841 271260
rect 120875 271226 120887 271260
rect 120829 271192 120887 271226
rect 120829 271158 120841 271192
rect 120875 271158 120887 271192
rect 120829 271129 120887 271158
rect 121071 271600 121129 271629
rect 121071 271566 121083 271600
rect 121117 271566 121129 271600
rect 121071 271532 121129 271566
rect 121071 271498 121083 271532
rect 121117 271498 121129 271532
rect 121071 271464 121129 271498
rect 121071 271430 121083 271464
rect 121117 271430 121129 271464
rect 121071 271396 121129 271430
rect 121071 271362 121083 271396
rect 121117 271362 121129 271396
rect 121071 271328 121129 271362
rect 121071 271294 121083 271328
rect 121117 271294 121129 271328
rect 121071 271260 121129 271294
rect 121071 271226 121083 271260
rect 121117 271226 121129 271260
rect 121071 271192 121129 271226
rect 121071 271158 121083 271192
rect 121117 271158 121129 271192
rect 121071 271129 121129 271158
rect 121529 271600 121587 271629
rect 121529 271566 121541 271600
rect 121575 271566 121587 271600
rect 121529 271532 121587 271566
rect 121529 271498 121541 271532
rect 121575 271498 121587 271532
rect 121529 271464 121587 271498
rect 121529 271430 121541 271464
rect 121575 271430 121587 271464
rect 121529 271396 121587 271430
rect 121529 271362 121541 271396
rect 121575 271362 121587 271396
rect 121529 271328 121587 271362
rect 121529 271294 121541 271328
rect 121575 271294 121587 271328
rect 121529 271260 121587 271294
rect 121529 271226 121541 271260
rect 121575 271226 121587 271260
rect 121529 271192 121587 271226
rect 121529 271158 121541 271192
rect 121575 271158 121587 271192
rect 121529 271129 121587 271158
rect 120371 270816 120429 270845
rect 120371 270782 120383 270816
rect 120417 270782 120429 270816
rect 120371 270748 120429 270782
rect 120371 270714 120383 270748
rect 120417 270714 120429 270748
rect 120371 270680 120429 270714
rect 120371 270646 120383 270680
rect 120417 270646 120429 270680
rect 120371 270612 120429 270646
rect 120371 270578 120383 270612
rect 120417 270578 120429 270612
rect 120371 270544 120429 270578
rect 120371 270510 120383 270544
rect 120417 270510 120429 270544
rect 120371 270476 120429 270510
rect 120371 270442 120383 270476
rect 120417 270442 120429 270476
rect 120371 270408 120429 270442
rect 120371 270374 120383 270408
rect 120417 270374 120429 270408
rect 120371 270345 120429 270374
rect 120829 270816 120887 270845
rect 120829 270782 120841 270816
rect 120875 270782 120887 270816
rect 120829 270748 120887 270782
rect 120829 270714 120841 270748
rect 120875 270714 120887 270748
rect 120829 270680 120887 270714
rect 120829 270646 120841 270680
rect 120875 270646 120887 270680
rect 120829 270612 120887 270646
rect 120829 270578 120841 270612
rect 120875 270578 120887 270612
rect 120829 270544 120887 270578
rect 120829 270510 120841 270544
rect 120875 270510 120887 270544
rect 120829 270476 120887 270510
rect 120829 270442 120841 270476
rect 120875 270442 120887 270476
rect 120829 270408 120887 270442
rect 120829 270374 120841 270408
rect 120875 270374 120887 270408
rect 120829 270345 120887 270374
rect 121071 270816 121129 270845
rect 121071 270782 121083 270816
rect 121117 270782 121129 270816
rect 121071 270748 121129 270782
rect 121071 270714 121083 270748
rect 121117 270714 121129 270748
rect 121071 270680 121129 270714
rect 121071 270646 121083 270680
rect 121117 270646 121129 270680
rect 121071 270612 121129 270646
rect 121071 270578 121083 270612
rect 121117 270578 121129 270612
rect 121071 270544 121129 270578
rect 121071 270510 121083 270544
rect 121117 270510 121129 270544
rect 121071 270476 121129 270510
rect 121071 270442 121083 270476
rect 121117 270442 121129 270476
rect 121071 270408 121129 270442
rect 121071 270374 121083 270408
rect 121117 270374 121129 270408
rect 121071 270345 121129 270374
rect 121529 270816 121587 270845
rect 121529 270782 121541 270816
rect 121575 270782 121587 270816
rect 121529 270748 121587 270782
rect 121529 270714 121541 270748
rect 121575 270714 121587 270748
rect 121529 270680 121587 270714
rect 121529 270646 121541 270680
rect 121575 270646 121587 270680
rect 121529 270612 121587 270646
rect 121529 270578 121541 270612
rect 121575 270578 121587 270612
rect 121529 270544 121587 270578
rect 121529 270510 121541 270544
rect 121575 270510 121587 270544
rect 121529 270476 121587 270510
rect 121529 270442 121541 270476
rect 121575 270442 121587 270476
rect 121529 270408 121587 270442
rect 121529 270374 121541 270408
rect 121575 270374 121587 270408
rect 121529 270345 121587 270374
rect 120371 270032 120429 270061
rect 120371 269998 120383 270032
rect 120417 269998 120429 270032
rect 120371 269964 120429 269998
rect 120371 269930 120383 269964
rect 120417 269930 120429 269964
rect 120371 269896 120429 269930
rect 120371 269862 120383 269896
rect 120417 269862 120429 269896
rect 120371 269828 120429 269862
rect 120371 269794 120383 269828
rect 120417 269794 120429 269828
rect 120371 269760 120429 269794
rect 120371 269726 120383 269760
rect 120417 269726 120429 269760
rect 120371 269692 120429 269726
rect 120371 269658 120383 269692
rect 120417 269658 120429 269692
rect 120371 269624 120429 269658
rect 120371 269590 120383 269624
rect 120417 269590 120429 269624
rect 120371 269561 120429 269590
rect 120829 270032 120887 270061
rect 120829 269998 120841 270032
rect 120875 269998 120887 270032
rect 120829 269964 120887 269998
rect 120829 269930 120841 269964
rect 120875 269930 120887 269964
rect 120829 269896 120887 269930
rect 120829 269862 120841 269896
rect 120875 269862 120887 269896
rect 120829 269828 120887 269862
rect 120829 269794 120841 269828
rect 120875 269794 120887 269828
rect 120829 269760 120887 269794
rect 120829 269726 120841 269760
rect 120875 269726 120887 269760
rect 120829 269692 120887 269726
rect 120829 269658 120841 269692
rect 120875 269658 120887 269692
rect 120829 269624 120887 269658
rect 120829 269590 120841 269624
rect 120875 269590 120887 269624
rect 120829 269561 120887 269590
rect 121071 270032 121129 270061
rect 121071 269998 121083 270032
rect 121117 269998 121129 270032
rect 121071 269964 121129 269998
rect 121071 269930 121083 269964
rect 121117 269930 121129 269964
rect 121071 269896 121129 269930
rect 121071 269862 121083 269896
rect 121117 269862 121129 269896
rect 121071 269828 121129 269862
rect 121071 269794 121083 269828
rect 121117 269794 121129 269828
rect 121071 269760 121129 269794
rect 121071 269726 121083 269760
rect 121117 269726 121129 269760
rect 121071 269692 121129 269726
rect 121071 269658 121083 269692
rect 121117 269658 121129 269692
rect 121071 269624 121129 269658
rect 121071 269590 121083 269624
rect 121117 269590 121129 269624
rect 121071 269561 121129 269590
rect 121529 270032 121587 270061
rect 121529 269998 121541 270032
rect 121575 269998 121587 270032
rect 121529 269964 121587 269998
rect 121529 269930 121541 269964
rect 121575 269930 121587 269964
rect 121529 269896 121587 269930
rect 121529 269862 121541 269896
rect 121575 269862 121587 269896
rect 121529 269828 121587 269862
rect 121529 269794 121541 269828
rect 121575 269794 121587 269828
rect 121529 269760 121587 269794
rect 121529 269726 121541 269760
rect 121575 269726 121587 269760
rect 121529 269692 121587 269726
rect 121529 269658 121541 269692
rect 121575 269658 121587 269692
rect 121529 269624 121587 269658
rect 121529 269590 121541 269624
rect 121575 269590 121587 269624
rect 121529 269561 121587 269590
rect 120371 269244 120429 269277
rect 120371 269210 120383 269244
rect 120417 269210 120429 269244
rect 120371 269177 120429 269210
rect 120829 269244 120887 269277
rect 120829 269210 120841 269244
rect 120875 269210 120887 269244
rect 120829 269177 120887 269210
rect 121071 269244 121129 269277
rect 121071 269210 121083 269244
rect 121117 269210 121129 269244
rect 121071 269177 121129 269210
rect 121529 269244 121587 269277
rect 121529 269210 121541 269244
rect 121575 269210 121587 269244
rect 121529 269177 121587 269210
rect 122067 272780 122125 272813
rect 122067 272746 122079 272780
rect 122113 272746 122125 272780
rect 122067 272713 122125 272746
rect 122525 272780 122583 272813
rect 122525 272746 122537 272780
rect 122571 272746 122583 272780
rect 122525 272713 122583 272746
rect 122767 272780 122825 272813
rect 122767 272746 122779 272780
rect 122813 272746 122825 272780
rect 122767 272713 122825 272746
rect 123225 272780 123283 272813
rect 123225 272746 123237 272780
rect 123271 272746 123283 272780
rect 123225 272713 123283 272746
rect 122067 272400 122125 272429
rect 122067 272366 122079 272400
rect 122113 272366 122125 272400
rect 122067 272332 122125 272366
rect 122067 272298 122079 272332
rect 122113 272298 122125 272332
rect 122067 272264 122125 272298
rect 122067 272230 122079 272264
rect 122113 272230 122125 272264
rect 122067 272196 122125 272230
rect 122067 272162 122079 272196
rect 122113 272162 122125 272196
rect 122067 272128 122125 272162
rect 122067 272094 122079 272128
rect 122113 272094 122125 272128
rect 122067 272060 122125 272094
rect 122067 272026 122079 272060
rect 122113 272026 122125 272060
rect 122067 271992 122125 272026
rect 122067 271958 122079 271992
rect 122113 271958 122125 271992
rect 122067 271929 122125 271958
rect 122525 272400 122583 272429
rect 122525 272366 122537 272400
rect 122571 272366 122583 272400
rect 122525 272332 122583 272366
rect 122525 272298 122537 272332
rect 122571 272298 122583 272332
rect 122525 272264 122583 272298
rect 122525 272230 122537 272264
rect 122571 272230 122583 272264
rect 122525 272196 122583 272230
rect 122525 272162 122537 272196
rect 122571 272162 122583 272196
rect 122525 272128 122583 272162
rect 122525 272094 122537 272128
rect 122571 272094 122583 272128
rect 122525 272060 122583 272094
rect 122525 272026 122537 272060
rect 122571 272026 122583 272060
rect 122525 271992 122583 272026
rect 122525 271958 122537 271992
rect 122571 271958 122583 271992
rect 122525 271929 122583 271958
rect 122767 272400 122825 272429
rect 122767 272366 122779 272400
rect 122813 272366 122825 272400
rect 122767 272332 122825 272366
rect 122767 272298 122779 272332
rect 122813 272298 122825 272332
rect 122767 272264 122825 272298
rect 122767 272230 122779 272264
rect 122813 272230 122825 272264
rect 122767 272196 122825 272230
rect 122767 272162 122779 272196
rect 122813 272162 122825 272196
rect 122767 272128 122825 272162
rect 122767 272094 122779 272128
rect 122813 272094 122825 272128
rect 122767 272060 122825 272094
rect 122767 272026 122779 272060
rect 122813 272026 122825 272060
rect 122767 271992 122825 272026
rect 122767 271958 122779 271992
rect 122813 271958 122825 271992
rect 122767 271929 122825 271958
rect 123225 272400 123283 272429
rect 123225 272366 123237 272400
rect 123271 272366 123283 272400
rect 123225 272332 123283 272366
rect 123225 272298 123237 272332
rect 123271 272298 123283 272332
rect 123225 272264 123283 272298
rect 123225 272230 123237 272264
rect 123271 272230 123283 272264
rect 123225 272196 123283 272230
rect 123225 272162 123237 272196
rect 123271 272162 123283 272196
rect 123225 272128 123283 272162
rect 123225 272094 123237 272128
rect 123271 272094 123283 272128
rect 123225 272060 123283 272094
rect 123225 272026 123237 272060
rect 123271 272026 123283 272060
rect 123225 271992 123283 272026
rect 123225 271958 123237 271992
rect 123271 271958 123283 271992
rect 123225 271929 123283 271958
rect 122067 271616 122125 271645
rect 122067 271582 122079 271616
rect 122113 271582 122125 271616
rect 122067 271548 122125 271582
rect 122067 271514 122079 271548
rect 122113 271514 122125 271548
rect 122067 271480 122125 271514
rect 122067 271446 122079 271480
rect 122113 271446 122125 271480
rect 122067 271412 122125 271446
rect 122067 271378 122079 271412
rect 122113 271378 122125 271412
rect 122067 271344 122125 271378
rect 122067 271310 122079 271344
rect 122113 271310 122125 271344
rect 122067 271276 122125 271310
rect 122067 271242 122079 271276
rect 122113 271242 122125 271276
rect 122067 271208 122125 271242
rect 122067 271174 122079 271208
rect 122113 271174 122125 271208
rect 122067 271145 122125 271174
rect 122525 271616 122583 271645
rect 122525 271582 122537 271616
rect 122571 271582 122583 271616
rect 122525 271548 122583 271582
rect 122525 271514 122537 271548
rect 122571 271514 122583 271548
rect 122525 271480 122583 271514
rect 122525 271446 122537 271480
rect 122571 271446 122583 271480
rect 122525 271412 122583 271446
rect 122525 271378 122537 271412
rect 122571 271378 122583 271412
rect 122525 271344 122583 271378
rect 122525 271310 122537 271344
rect 122571 271310 122583 271344
rect 122525 271276 122583 271310
rect 122525 271242 122537 271276
rect 122571 271242 122583 271276
rect 122525 271208 122583 271242
rect 122525 271174 122537 271208
rect 122571 271174 122583 271208
rect 122525 271145 122583 271174
rect 122767 271616 122825 271645
rect 122767 271582 122779 271616
rect 122813 271582 122825 271616
rect 122767 271548 122825 271582
rect 122767 271514 122779 271548
rect 122813 271514 122825 271548
rect 122767 271480 122825 271514
rect 122767 271446 122779 271480
rect 122813 271446 122825 271480
rect 122767 271412 122825 271446
rect 122767 271378 122779 271412
rect 122813 271378 122825 271412
rect 122767 271344 122825 271378
rect 122767 271310 122779 271344
rect 122813 271310 122825 271344
rect 122767 271276 122825 271310
rect 122767 271242 122779 271276
rect 122813 271242 122825 271276
rect 122767 271208 122825 271242
rect 122767 271174 122779 271208
rect 122813 271174 122825 271208
rect 122767 271145 122825 271174
rect 123225 271616 123283 271645
rect 123225 271582 123237 271616
rect 123271 271582 123283 271616
rect 123225 271548 123283 271582
rect 123225 271514 123237 271548
rect 123271 271514 123283 271548
rect 123225 271480 123283 271514
rect 123225 271446 123237 271480
rect 123271 271446 123283 271480
rect 123225 271412 123283 271446
rect 123225 271378 123237 271412
rect 123271 271378 123283 271412
rect 123225 271344 123283 271378
rect 123225 271310 123237 271344
rect 123271 271310 123283 271344
rect 123225 271276 123283 271310
rect 123225 271242 123237 271276
rect 123271 271242 123283 271276
rect 123225 271208 123283 271242
rect 123225 271174 123237 271208
rect 123271 271174 123283 271208
rect 123225 271145 123283 271174
rect 122067 270832 122125 270861
rect 122067 270798 122079 270832
rect 122113 270798 122125 270832
rect 122067 270764 122125 270798
rect 122067 270730 122079 270764
rect 122113 270730 122125 270764
rect 122067 270696 122125 270730
rect 122067 270662 122079 270696
rect 122113 270662 122125 270696
rect 122067 270628 122125 270662
rect 122067 270594 122079 270628
rect 122113 270594 122125 270628
rect 122067 270560 122125 270594
rect 122067 270526 122079 270560
rect 122113 270526 122125 270560
rect 122067 270492 122125 270526
rect 122067 270458 122079 270492
rect 122113 270458 122125 270492
rect 122067 270424 122125 270458
rect 122067 270390 122079 270424
rect 122113 270390 122125 270424
rect 122067 270361 122125 270390
rect 122525 270832 122583 270861
rect 122525 270798 122537 270832
rect 122571 270798 122583 270832
rect 122525 270764 122583 270798
rect 122525 270730 122537 270764
rect 122571 270730 122583 270764
rect 122525 270696 122583 270730
rect 122525 270662 122537 270696
rect 122571 270662 122583 270696
rect 122525 270628 122583 270662
rect 122525 270594 122537 270628
rect 122571 270594 122583 270628
rect 122525 270560 122583 270594
rect 122525 270526 122537 270560
rect 122571 270526 122583 270560
rect 122525 270492 122583 270526
rect 122525 270458 122537 270492
rect 122571 270458 122583 270492
rect 122525 270424 122583 270458
rect 122525 270390 122537 270424
rect 122571 270390 122583 270424
rect 122525 270361 122583 270390
rect 122767 270832 122825 270861
rect 122767 270798 122779 270832
rect 122813 270798 122825 270832
rect 122767 270764 122825 270798
rect 122767 270730 122779 270764
rect 122813 270730 122825 270764
rect 122767 270696 122825 270730
rect 122767 270662 122779 270696
rect 122813 270662 122825 270696
rect 122767 270628 122825 270662
rect 122767 270594 122779 270628
rect 122813 270594 122825 270628
rect 122767 270560 122825 270594
rect 122767 270526 122779 270560
rect 122813 270526 122825 270560
rect 122767 270492 122825 270526
rect 122767 270458 122779 270492
rect 122813 270458 122825 270492
rect 122767 270424 122825 270458
rect 122767 270390 122779 270424
rect 122813 270390 122825 270424
rect 122767 270361 122825 270390
rect 123225 270832 123283 270861
rect 123225 270798 123237 270832
rect 123271 270798 123283 270832
rect 123225 270764 123283 270798
rect 123225 270730 123237 270764
rect 123271 270730 123283 270764
rect 123225 270696 123283 270730
rect 123225 270662 123237 270696
rect 123271 270662 123283 270696
rect 123225 270628 123283 270662
rect 123225 270594 123237 270628
rect 123271 270594 123283 270628
rect 123225 270560 123283 270594
rect 123225 270526 123237 270560
rect 123271 270526 123283 270560
rect 123225 270492 123283 270526
rect 123225 270458 123237 270492
rect 123271 270458 123283 270492
rect 123225 270424 123283 270458
rect 123225 270390 123237 270424
rect 123271 270390 123283 270424
rect 123225 270361 123283 270390
rect 122067 270048 122125 270077
rect 122067 270014 122079 270048
rect 122113 270014 122125 270048
rect 122067 269980 122125 270014
rect 122067 269946 122079 269980
rect 122113 269946 122125 269980
rect 122067 269912 122125 269946
rect 122067 269878 122079 269912
rect 122113 269878 122125 269912
rect 122067 269844 122125 269878
rect 122067 269810 122079 269844
rect 122113 269810 122125 269844
rect 122067 269776 122125 269810
rect 122067 269742 122079 269776
rect 122113 269742 122125 269776
rect 122067 269708 122125 269742
rect 122067 269674 122079 269708
rect 122113 269674 122125 269708
rect 122067 269640 122125 269674
rect 122067 269606 122079 269640
rect 122113 269606 122125 269640
rect 122067 269577 122125 269606
rect 122525 270048 122583 270077
rect 122525 270014 122537 270048
rect 122571 270014 122583 270048
rect 122525 269980 122583 270014
rect 122525 269946 122537 269980
rect 122571 269946 122583 269980
rect 122525 269912 122583 269946
rect 122525 269878 122537 269912
rect 122571 269878 122583 269912
rect 122525 269844 122583 269878
rect 122525 269810 122537 269844
rect 122571 269810 122583 269844
rect 122525 269776 122583 269810
rect 122525 269742 122537 269776
rect 122571 269742 122583 269776
rect 122525 269708 122583 269742
rect 122525 269674 122537 269708
rect 122571 269674 122583 269708
rect 122525 269640 122583 269674
rect 122525 269606 122537 269640
rect 122571 269606 122583 269640
rect 122525 269577 122583 269606
rect 122767 270048 122825 270077
rect 122767 270014 122779 270048
rect 122813 270014 122825 270048
rect 122767 269980 122825 270014
rect 122767 269946 122779 269980
rect 122813 269946 122825 269980
rect 122767 269912 122825 269946
rect 122767 269878 122779 269912
rect 122813 269878 122825 269912
rect 122767 269844 122825 269878
rect 122767 269810 122779 269844
rect 122813 269810 122825 269844
rect 122767 269776 122825 269810
rect 122767 269742 122779 269776
rect 122813 269742 122825 269776
rect 122767 269708 122825 269742
rect 122767 269674 122779 269708
rect 122813 269674 122825 269708
rect 122767 269640 122825 269674
rect 122767 269606 122779 269640
rect 122813 269606 122825 269640
rect 122767 269577 122825 269606
rect 123225 270048 123283 270077
rect 123225 270014 123237 270048
rect 123271 270014 123283 270048
rect 123225 269980 123283 270014
rect 123225 269946 123237 269980
rect 123271 269946 123283 269980
rect 123225 269912 123283 269946
rect 123225 269878 123237 269912
rect 123271 269878 123283 269912
rect 123225 269844 123283 269878
rect 123225 269810 123237 269844
rect 123271 269810 123283 269844
rect 123225 269776 123283 269810
rect 123225 269742 123237 269776
rect 123271 269742 123283 269776
rect 123225 269708 123283 269742
rect 123225 269674 123237 269708
rect 123271 269674 123283 269708
rect 123225 269640 123283 269674
rect 123225 269606 123237 269640
rect 123271 269606 123283 269640
rect 123225 269577 123283 269606
rect 122067 269260 122125 269293
rect 122067 269226 122079 269260
rect 122113 269226 122125 269260
rect 122067 269193 122125 269226
rect 122525 269260 122583 269293
rect 122525 269226 122537 269260
rect 122571 269226 122583 269260
rect 122525 269193 122583 269226
rect 122767 269260 122825 269293
rect 122767 269226 122779 269260
rect 122813 269226 122825 269260
rect 122767 269193 122825 269226
rect 123225 269260 123283 269293
rect 123225 269226 123237 269260
rect 123271 269226 123283 269260
rect 123225 269193 123283 269226
<< ndiffc >>
rect 106311 280762 106345 280796
rect 106311 280694 106345 280728
rect 106311 280626 106345 280660
rect 106311 280558 106345 280592
rect 106311 280490 106345 280524
rect 106311 280422 106345 280456
rect 106311 280354 106345 280388
rect 106311 280286 106345 280320
rect 106311 280218 106345 280252
rect 106311 280150 106345 280184
rect 106311 280082 106345 280116
rect 106311 280014 106345 280048
rect 106311 279946 106345 279980
rect 106311 279878 106345 279912
rect 106311 279810 106345 279844
rect 106501 280762 106535 280796
rect 106501 280694 106535 280728
rect 106501 280626 106535 280660
rect 106501 280558 106535 280592
rect 106501 280490 106535 280524
rect 106501 280422 106535 280456
rect 106501 280354 106535 280388
rect 106501 280286 106535 280320
rect 106501 280218 106535 280252
rect 106501 280150 106535 280184
rect 106501 280082 106535 280116
rect 106501 280014 106535 280048
rect 106501 279946 106535 279980
rect 106501 279878 106535 279912
rect 106501 279810 106535 279844
rect 106711 280762 106745 280796
rect 106711 280694 106745 280728
rect 106711 280626 106745 280660
rect 106711 280558 106745 280592
rect 106711 280490 106745 280524
rect 106711 280422 106745 280456
rect 106711 280354 106745 280388
rect 106711 280286 106745 280320
rect 106711 280218 106745 280252
rect 106711 280150 106745 280184
rect 106711 280082 106745 280116
rect 106711 280014 106745 280048
rect 106711 279946 106745 279980
rect 106711 279878 106745 279912
rect 106711 279810 106745 279844
rect 106901 280762 106935 280796
rect 106901 280694 106935 280728
rect 106901 280626 106935 280660
rect 106901 280558 106935 280592
rect 106901 280490 106935 280524
rect 106901 280422 106935 280456
rect 106901 280354 106935 280388
rect 106901 280286 106935 280320
rect 106901 280218 106935 280252
rect 106901 280150 106935 280184
rect 106901 280082 106935 280116
rect 106901 280014 106935 280048
rect 106901 279946 106935 279980
rect 106901 279878 106935 279912
rect 106901 279810 106935 279844
rect 107111 280762 107145 280796
rect 107111 280694 107145 280728
rect 107111 280626 107145 280660
rect 107111 280558 107145 280592
rect 107111 280490 107145 280524
rect 107111 280422 107145 280456
rect 107111 280354 107145 280388
rect 107111 280286 107145 280320
rect 107111 280218 107145 280252
rect 107111 280150 107145 280184
rect 107111 280082 107145 280116
rect 107111 280014 107145 280048
rect 107111 279946 107145 279980
rect 107111 279878 107145 279912
rect 107111 279810 107145 279844
rect 107301 280762 107335 280796
rect 107301 280694 107335 280728
rect 107301 280626 107335 280660
rect 107301 280558 107335 280592
rect 107301 280490 107335 280524
rect 107301 280422 107335 280456
rect 107301 280354 107335 280388
rect 107301 280286 107335 280320
rect 107301 280218 107335 280252
rect 107301 280150 107335 280184
rect 107301 280082 107335 280116
rect 107301 280014 107335 280048
rect 107301 279946 107335 279980
rect 107301 279878 107335 279912
rect 107301 279810 107335 279844
rect 107511 280762 107545 280796
rect 107511 280694 107545 280728
rect 107511 280626 107545 280660
rect 107511 280558 107545 280592
rect 107511 280490 107545 280524
rect 107511 280422 107545 280456
rect 107511 280354 107545 280388
rect 107511 280286 107545 280320
rect 107511 280218 107545 280252
rect 107511 280150 107545 280184
rect 107511 280082 107545 280116
rect 107511 280014 107545 280048
rect 107511 279946 107545 279980
rect 107511 279878 107545 279912
rect 107511 279810 107545 279844
rect 107701 280762 107735 280796
rect 107701 280694 107735 280728
rect 107701 280626 107735 280660
rect 107701 280558 107735 280592
rect 107701 280490 107735 280524
rect 107701 280422 107735 280456
rect 107701 280354 107735 280388
rect 107701 280286 107735 280320
rect 107701 280218 107735 280252
rect 107701 280150 107735 280184
rect 107701 280082 107735 280116
rect 107701 280014 107735 280048
rect 107701 279946 107735 279980
rect 107701 279878 107735 279912
rect 107701 279810 107735 279844
rect 107911 280762 107945 280796
rect 107911 280694 107945 280728
rect 107911 280626 107945 280660
rect 107911 280558 107945 280592
rect 107911 280490 107945 280524
rect 107911 280422 107945 280456
rect 107911 280354 107945 280388
rect 107911 280286 107945 280320
rect 107911 280218 107945 280252
rect 107911 280150 107945 280184
rect 107911 280082 107945 280116
rect 107911 280014 107945 280048
rect 107911 279946 107945 279980
rect 107911 279878 107945 279912
rect 107911 279810 107945 279844
rect 108101 280762 108135 280796
rect 108101 280694 108135 280728
rect 108101 280626 108135 280660
rect 108101 280558 108135 280592
rect 108101 280490 108135 280524
rect 108101 280422 108135 280456
rect 108101 280354 108135 280388
rect 108101 280286 108135 280320
rect 108101 280218 108135 280252
rect 108101 280150 108135 280184
rect 108101 280082 108135 280116
rect 108101 280014 108135 280048
rect 108101 279946 108135 279980
rect 108101 279878 108135 279912
rect 108101 279810 108135 279844
rect 108311 280762 108345 280796
rect 108311 280694 108345 280728
rect 108311 280626 108345 280660
rect 108311 280558 108345 280592
rect 108311 280490 108345 280524
rect 108311 280422 108345 280456
rect 108311 280354 108345 280388
rect 108311 280286 108345 280320
rect 108311 280218 108345 280252
rect 108311 280150 108345 280184
rect 108311 280082 108345 280116
rect 108311 280014 108345 280048
rect 108311 279946 108345 279980
rect 108311 279878 108345 279912
rect 108311 279810 108345 279844
rect 108501 280762 108535 280796
rect 108501 280694 108535 280728
rect 108501 280626 108535 280660
rect 108501 280558 108535 280592
rect 108501 280490 108535 280524
rect 108501 280422 108535 280456
rect 108501 280354 108535 280388
rect 108501 280286 108535 280320
rect 108501 280218 108535 280252
rect 108501 280150 108535 280184
rect 108501 280082 108535 280116
rect 108501 280014 108535 280048
rect 108501 279946 108535 279980
rect 108501 279878 108535 279912
rect 108501 279810 108535 279844
rect 108711 280762 108745 280796
rect 108711 280694 108745 280728
rect 108711 280626 108745 280660
rect 108711 280558 108745 280592
rect 108711 280490 108745 280524
rect 108711 280422 108745 280456
rect 108711 280354 108745 280388
rect 108711 280286 108745 280320
rect 108711 280218 108745 280252
rect 108711 280150 108745 280184
rect 108711 280082 108745 280116
rect 108711 280014 108745 280048
rect 108711 279946 108745 279980
rect 108711 279878 108745 279912
rect 108711 279810 108745 279844
rect 108901 280762 108935 280796
rect 108901 280694 108935 280728
rect 108901 280626 108935 280660
rect 108901 280558 108935 280592
rect 108901 280490 108935 280524
rect 108901 280422 108935 280456
rect 108901 280354 108935 280388
rect 108901 280286 108935 280320
rect 108901 280218 108935 280252
rect 108901 280150 108935 280184
rect 108901 280082 108935 280116
rect 108901 280014 108935 280048
rect 108901 279946 108935 279980
rect 108901 279878 108935 279912
rect 108901 279810 108935 279844
rect 109111 280762 109145 280796
rect 109111 280694 109145 280728
rect 109111 280626 109145 280660
rect 109111 280558 109145 280592
rect 109111 280490 109145 280524
rect 109111 280422 109145 280456
rect 109111 280354 109145 280388
rect 109111 280286 109145 280320
rect 109111 280218 109145 280252
rect 109111 280150 109145 280184
rect 109111 280082 109145 280116
rect 109111 280014 109145 280048
rect 109111 279946 109145 279980
rect 109111 279878 109145 279912
rect 109111 279810 109145 279844
rect 109301 280762 109335 280796
rect 109301 280694 109335 280728
rect 109301 280626 109335 280660
rect 109301 280558 109335 280592
rect 109301 280490 109335 280524
rect 109301 280422 109335 280456
rect 109301 280354 109335 280388
rect 109301 280286 109335 280320
rect 109301 280218 109335 280252
rect 109301 280150 109335 280184
rect 109301 280082 109335 280116
rect 109301 280014 109335 280048
rect 109301 279946 109335 279980
rect 109301 279878 109335 279912
rect 109301 279810 109335 279844
rect 109511 280762 109545 280796
rect 109511 280694 109545 280728
rect 109511 280626 109545 280660
rect 109511 280558 109545 280592
rect 109511 280490 109545 280524
rect 109511 280422 109545 280456
rect 109511 280354 109545 280388
rect 109511 280286 109545 280320
rect 109511 280218 109545 280252
rect 109511 280150 109545 280184
rect 109511 280082 109545 280116
rect 109511 280014 109545 280048
rect 109511 279946 109545 279980
rect 109511 279878 109545 279912
rect 109511 279810 109545 279844
rect 109701 280762 109735 280796
rect 109701 280694 109735 280728
rect 109701 280626 109735 280660
rect 109701 280558 109735 280592
rect 109701 280490 109735 280524
rect 109701 280422 109735 280456
rect 109701 280354 109735 280388
rect 109701 280286 109735 280320
rect 109701 280218 109735 280252
rect 109701 280150 109735 280184
rect 109701 280082 109735 280116
rect 109701 280014 109735 280048
rect 109701 279946 109735 279980
rect 109701 279878 109735 279912
rect 109701 279810 109735 279844
rect 109911 280762 109945 280796
rect 109911 280694 109945 280728
rect 109911 280626 109945 280660
rect 109911 280558 109945 280592
rect 109911 280490 109945 280524
rect 109911 280422 109945 280456
rect 109911 280354 109945 280388
rect 109911 280286 109945 280320
rect 109911 280218 109945 280252
rect 109911 280150 109945 280184
rect 109911 280082 109945 280116
rect 109911 280014 109945 280048
rect 109911 279946 109945 279980
rect 109911 279878 109945 279912
rect 109911 279810 109945 279844
rect 110101 280762 110135 280796
rect 110101 280694 110135 280728
rect 110101 280626 110135 280660
rect 110101 280558 110135 280592
rect 110101 280490 110135 280524
rect 110101 280422 110135 280456
rect 110101 280354 110135 280388
rect 110101 280286 110135 280320
rect 110101 280218 110135 280252
rect 110101 280150 110135 280184
rect 110101 280082 110135 280116
rect 110101 280014 110135 280048
rect 110101 279946 110135 279980
rect 110101 279878 110135 279912
rect 110101 279810 110135 279844
rect 109731 278951 109765 278985
rect 109731 278883 109765 278917
rect 109731 278815 109765 278849
rect 109731 278747 109765 278781
rect 109731 278679 109765 278713
rect 109731 278611 109765 278645
rect 109731 278543 109765 278577
rect 109731 278475 109765 278509
rect 109731 278407 109765 278441
rect 109731 278339 109765 278373
rect 109731 278271 109765 278305
rect 109731 278203 109765 278237
rect 109731 278135 109765 278169
rect 109731 278067 109765 278101
rect 109731 277999 109765 278033
rect 110075 278951 110109 278985
rect 110075 278883 110109 278917
rect 110075 278815 110109 278849
rect 110075 278747 110109 278781
rect 110075 278679 110109 278713
rect 110075 278611 110109 278645
rect 110075 278543 110109 278577
rect 110075 278475 110109 278509
rect 110075 278407 110109 278441
rect 110075 278339 110109 278373
rect 110075 278271 110109 278305
rect 110075 278203 110109 278237
rect 110075 278135 110109 278169
rect 110075 278067 110109 278101
rect 110075 277999 110109 278033
rect 109731 277695 109765 277729
rect 109731 277627 109765 277661
rect 109731 277559 109765 277593
rect 109731 277491 109765 277525
rect 109731 277423 109765 277457
rect 109731 277355 109765 277389
rect 109731 277287 109765 277321
rect 109731 277219 109765 277253
rect 109731 277151 109765 277185
rect 109731 277083 109765 277117
rect 109731 277015 109765 277049
rect 109731 276947 109765 276981
rect 109731 276879 109765 276913
rect 109731 276811 109765 276845
rect 109731 276743 109765 276777
rect 110075 277695 110109 277729
rect 110075 277627 110109 277661
rect 110075 277559 110109 277593
rect 110075 277491 110109 277525
rect 110075 277423 110109 277457
rect 110075 277355 110109 277389
rect 110075 277287 110109 277321
rect 110075 277219 110109 277253
rect 110075 277151 110109 277185
rect 110075 277083 110109 277117
rect 110075 277015 110109 277049
rect 110075 276947 110109 276981
rect 110075 276879 110109 276913
rect 110075 276811 110109 276845
rect 110075 276743 110109 276777
rect 107413 272026 107447 272060
rect 106935 271906 106969 271940
rect 106935 271838 106969 271872
rect 107203 271906 107237 271940
rect 107203 271838 107237 271872
rect 107413 271958 107447 271992
rect 107413 271890 107447 271924
rect 107413 271822 107447 271856
rect 107413 271754 107447 271788
rect 108091 272026 108125 272060
rect 108091 271958 108125 271992
rect 108091 271890 108125 271924
rect 108091 271822 108125 271856
rect 108091 271754 108125 271788
rect 107212 271501 107246 271535
rect 107280 271501 107314 271535
rect 107348 271501 107382 271535
rect 107416 271501 107450 271535
rect 107484 271501 107518 271535
rect 107552 271501 107586 271535
rect 107620 271501 107654 271535
rect 107688 271501 107722 271535
rect 107756 271501 107790 271535
rect 107824 271501 107858 271535
rect 107892 271501 107926 271535
rect 107960 271501 107994 271535
rect 108028 271501 108062 271535
rect 108096 271501 108130 271535
rect 108164 271501 108198 271535
rect 108232 271501 108266 271535
rect 108300 271501 108334 271535
rect 107212 271265 107246 271299
rect 107280 271265 107314 271299
rect 107348 271265 107382 271299
rect 107416 271265 107450 271299
rect 107484 271265 107518 271299
rect 107552 271265 107586 271299
rect 107620 271265 107654 271299
rect 107688 271265 107722 271299
rect 107756 271265 107790 271299
rect 107824 271265 107858 271299
rect 107892 271265 107926 271299
rect 107960 271265 107994 271299
rect 108028 271265 108062 271299
rect 108096 271265 108130 271299
rect 108164 271265 108198 271299
rect 108232 271265 108266 271299
rect 108300 271265 108334 271299
rect 107212 271131 107246 271165
rect 107280 271131 107314 271165
rect 107348 271131 107382 271165
rect 107416 271131 107450 271165
rect 107484 271131 107518 271165
rect 107552 271131 107586 271165
rect 107620 271131 107654 271165
rect 107688 271131 107722 271165
rect 107756 271131 107790 271165
rect 107824 271131 107858 271165
rect 107892 271131 107926 271165
rect 107960 271131 107994 271165
rect 108028 271131 108062 271165
rect 108096 271131 108130 271165
rect 108164 271131 108198 271165
rect 108232 271131 108266 271165
rect 108300 271131 108334 271165
rect 107212 270895 107246 270929
rect 107280 270895 107314 270929
rect 107348 270895 107382 270929
rect 107416 270895 107450 270929
rect 107484 270895 107518 270929
rect 107552 270895 107586 270929
rect 107620 270895 107654 270929
rect 107688 270895 107722 270929
rect 107756 270895 107790 270929
rect 107824 270895 107858 270929
rect 107892 270895 107926 270929
rect 107960 270895 107994 270929
rect 108028 270895 108062 270929
rect 108096 270895 108130 270929
rect 108164 270895 108198 270929
rect 108232 270895 108266 270929
rect 108300 270895 108334 270929
rect 111547 280832 111581 280866
rect 111615 280832 111649 280866
rect 111683 280832 111717 280866
rect 111751 280832 111785 280866
rect 111819 280832 111853 280866
rect 111887 280832 111921 280866
rect 111955 280832 111989 280866
rect 112023 280832 112057 280866
rect 112091 280832 112125 280866
rect 112159 280832 112193 280866
rect 112227 280832 112261 280866
rect 112295 280832 112329 280866
rect 112363 280832 112397 280866
rect 112431 280832 112465 280866
rect 112499 280832 112533 280866
rect 112567 280832 112601 280866
rect 112993 280840 113027 280874
rect 113061 280840 113095 280874
rect 113129 280840 113163 280874
rect 113197 280840 113231 280874
rect 113265 280840 113299 280874
rect 113333 280840 113367 280874
rect 113401 280840 113435 280874
rect 113469 280840 113503 280874
rect 113537 280840 113571 280874
rect 113605 280840 113639 280874
rect 113673 280840 113707 280874
rect 113741 280840 113775 280874
rect 113809 280840 113843 280874
rect 113877 280840 113911 280874
rect 113945 280840 113979 280874
rect 114013 280840 114047 280874
rect 111547 280614 111581 280648
rect 111615 280614 111649 280648
rect 111683 280614 111717 280648
rect 111751 280614 111785 280648
rect 111819 280614 111853 280648
rect 111887 280614 111921 280648
rect 111955 280614 111989 280648
rect 112023 280614 112057 280648
rect 112091 280614 112125 280648
rect 112159 280614 112193 280648
rect 112227 280614 112261 280648
rect 112295 280614 112329 280648
rect 112363 280614 112397 280648
rect 112431 280614 112465 280648
rect 112499 280614 112533 280648
rect 112567 280614 112601 280648
rect 112993 280582 113027 280616
rect 113061 280582 113095 280616
rect 113129 280582 113163 280616
rect 113197 280582 113231 280616
rect 113265 280582 113299 280616
rect 113333 280582 113367 280616
rect 113401 280582 113435 280616
rect 113469 280582 113503 280616
rect 113537 280582 113571 280616
rect 113605 280582 113639 280616
rect 113673 280582 113707 280616
rect 113741 280582 113775 280616
rect 113809 280582 113843 280616
rect 113877 280582 113911 280616
rect 113945 280582 113979 280616
rect 114013 280582 114047 280616
rect 111547 280472 111581 280506
rect 111615 280472 111649 280506
rect 111683 280472 111717 280506
rect 111751 280472 111785 280506
rect 111819 280472 111853 280506
rect 111887 280472 111921 280506
rect 111955 280472 111989 280506
rect 112023 280472 112057 280506
rect 112091 280472 112125 280506
rect 112159 280472 112193 280506
rect 112227 280472 112261 280506
rect 112295 280472 112329 280506
rect 112363 280472 112397 280506
rect 112431 280472 112465 280506
rect 112499 280472 112533 280506
rect 112567 280472 112601 280506
rect 112993 280416 113027 280450
rect 113061 280416 113095 280450
rect 113129 280416 113163 280450
rect 113197 280416 113231 280450
rect 113265 280416 113299 280450
rect 113333 280416 113367 280450
rect 113401 280416 113435 280450
rect 113469 280416 113503 280450
rect 113537 280416 113571 280450
rect 113605 280416 113639 280450
rect 113673 280416 113707 280450
rect 113741 280416 113775 280450
rect 113809 280416 113843 280450
rect 113877 280416 113911 280450
rect 113945 280416 113979 280450
rect 114013 280416 114047 280450
rect 111547 280254 111581 280288
rect 111615 280254 111649 280288
rect 111683 280254 111717 280288
rect 111751 280254 111785 280288
rect 111819 280254 111853 280288
rect 111887 280254 111921 280288
rect 111955 280254 111989 280288
rect 112023 280254 112057 280288
rect 112091 280254 112125 280288
rect 112159 280254 112193 280288
rect 112227 280254 112261 280288
rect 112295 280254 112329 280288
rect 112363 280254 112397 280288
rect 112431 280254 112465 280288
rect 112499 280254 112533 280288
rect 112567 280254 112601 280288
rect 112993 280158 113027 280192
rect 113061 280158 113095 280192
rect 113129 280158 113163 280192
rect 113197 280158 113231 280192
rect 113265 280158 113299 280192
rect 113333 280158 113367 280192
rect 113401 280158 113435 280192
rect 113469 280158 113503 280192
rect 113537 280158 113571 280192
rect 113605 280158 113639 280192
rect 113673 280158 113707 280192
rect 113741 280158 113775 280192
rect 113809 280158 113843 280192
rect 113877 280158 113911 280192
rect 113945 280158 113979 280192
rect 114013 280158 114047 280192
rect 111547 280112 111581 280146
rect 111615 280112 111649 280146
rect 111683 280112 111717 280146
rect 111751 280112 111785 280146
rect 111819 280112 111853 280146
rect 111887 280112 111921 280146
rect 111955 280112 111989 280146
rect 112023 280112 112057 280146
rect 112091 280112 112125 280146
rect 112159 280112 112193 280146
rect 112227 280112 112261 280146
rect 112295 280112 112329 280146
rect 112363 280112 112397 280146
rect 112431 280112 112465 280146
rect 112499 280112 112533 280146
rect 112567 280112 112601 280146
rect 113023 280014 113057 280048
rect 113091 280014 113125 280048
rect 113159 280014 113193 280048
rect 113227 280014 113261 280048
rect 113295 280014 113329 280048
rect 113363 280014 113397 280048
rect 113431 280014 113465 280048
rect 113499 280014 113533 280048
rect 113567 280014 113601 280048
rect 113635 280014 113669 280048
rect 113703 280014 113737 280048
rect 113771 280014 113805 280048
rect 113839 280014 113873 280048
rect 113907 280014 113941 280048
rect 113975 280014 114009 280048
rect 114043 280014 114077 280048
rect 111547 279894 111581 279928
rect 111615 279894 111649 279928
rect 111683 279894 111717 279928
rect 111751 279894 111785 279928
rect 111819 279894 111853 279928
rect 111887 279894 111921 279928
rect 111955 279894 111989 279928
rect 112023 279894 112057 279928
rect 112091 279894 112125 279928
rect 112159 279894 112193 279928
rect 112227 279894 112261 279928
rect 112295 279894 112329 279928
rect 112363 279894 112397 279928
rect 112431 279894 112465 279928
rect 112499 279894 112533 279928
rect 112567 279894 112601 279928
rect 113023 279876 113057 279910
rect 113091 279876 113125 279910
rect 113159 279876 113193 279910
rect 113227 279876 113261 279910
rect 113295 279876 113329 279910
rect 113363 279876 113397 279910
rect 113431 279876 113465 279910
rect 113499 279876 113533 279910
rect 113567 279876 113601 279910
rect 113635 279876 113669 279910
rect 113703 279876 113737 279910
rect 113771 279876 113805 279910
rect 113839 279876 113873 279910
rect 113907 279876 113941 279910
rect 113975 279876 114009 279910
rect 114043 279876 114077 279910
rect 111547 279752 111581 279786
rect 111615 279752 111649 279786
rect 111683 279752 111717 279786
rect 111751 279752 111785 279786
rect 111819 279752 111853 279786
rect 111887 279752 111921 279786
rect 111955 279752 111989 279786
rect 112023 279752 112057 279786
rect 112091 279752 112125 279786
rect 112159 279752 112193 279786
rect 112227 279752 112261 279786
rect 112295 279752 112329 279786
rect 112363 279752 112397 279786
rect 112431 279752 112465 279786
rect 112499 279752 112533 279786
rect 112567 279752 112601 279786
rect 113023 279716 113057 279750
rect 113091 279716 113125 279750
rect 113159 279716 113193 279750
rect 113227 279716 113261 279750
rect 113295 279716 113329 279750
rect 113363 279716 113397 279750
rect 113431 279716 113465 279750
rect 113499 279716 113533 279750
rect 113567 279716 113601 279750
rect 113635 279716 113669 279750
rect 113703 279716 113737 279750
rect 113771 279716 113805 279750
rect 113839 279716 113873 279750
rect 113907 279716 113941 279750
rect 113975 279716 114009 279750
rect 114043 279716 114077 279750
rect 111547 279534 111581 279568
rect 111615 279534 111649 279568
rect 111683 279534 111717 279568
rect 111751 279534 111785 279568
rect 111819 279534 111853 279568
rect 111887 279534 111921 279568
rect 111955 279534 111989 279568
rect 112023 279534 112057 279568
rect 112091 279534 112125 279568
rect 112159 279534 112193 279568
rect 112227 279534 112261 279568
rect 112295 279534 112329 279568
rect 112363 279534 112397 279568
rect 112431 279534 112465 279568
rect 112499 279534 112533 279568
rect 112567 279534 112601 279568
rect 113023 279578 113057 279612
rect 113091 279578 113125 279612
rect 113159 279578 113193 279612
rect 113227 279578 113261 279612
rect 113295 279578 113329 279612
rect 113363 279578 113397 279612
rect 113431 279578 113465 279612
rect 113499 279578 113533 279612
rect 113567 279578 113601 279612
rect 113635 279578 113669 279612
rect 113703 279578 113737 279612
rect 113771 279578 113805 279612
rect 113839 279578 113873 279612
rect 113907 279578 113941 279612
rect 113975 279578 114009 279612
rect 114043 279578 114077 279612
rect 116158 280840 116192 280874
rect 116226 280840 116260 280874
rect 116294 280840 116328 280874
rect 116362 280840 116396 280874
rect 116430 280840 116464 280874
rect 116498 280840 116532 280874
rect 116566 280840 116600 280874
rect 116634 280840 116668 280874
rect 116702 280840 116736 280874
rect 116770 280840 116804 280874
rect 116838 280840 116872 280874
rect 116906 280840 116940 280874
rect 116974 280840 117008 280874
rect 117042 280840 117076 280874
rect 117110 280840 117144 280874
rect 117178 280840 117212 280874
rect 117604 280832 117638 280866
rect 117672 280832 117706 280866
rect 117740 280832 117774 280866
rect 117808 280832 117842 280866
rect 117876 280832 117910 280866
rect 117944 280832 117978 280866
rect 118012 280832 118046 280866
rect 118080 280832 118114 280866
rect 118148 280832 118182 280866
rect 118216 280832 118250 280866
rect 118284 280832 118318 280866
rect 118352 280832 118386 280866
rect 118420 280832 118454 280866
rect 118488 280832 118522 280866
rect 118556 280832 118590 280866
rect 118624 280832 118658 280866
rect 116158 280582 116192 280616
rect 116226 280582 116260 280616
rect 116294 280582 116328 280616
rect 116362 280582 116396 280616
rect 116430 280582 116464 280616
rect 116498 280582 116532 280616
rect 116566 280582 116600 280616
rect 116634 280582 116668 280616
rect 116702 280582 116736 280616
rect 116770 280582 116804 280616
rect 116838 280582 116872 280616
rect 116906 280582 116940 280616
rect 116974 280582 117008 280616
rect 117042 280582 117076 280616
rect 117110 280582 117144 280616
rect 117178 280582 117212 280616
rect 117604 280614 117638 280648
rect 117672 280614 117706 280648
rect 117740 280614 117774 280648
rect 117808 280614 117842 280648
rect 117876 280614 117910 280648
rect 117944 280614 117978 280648
rect 118012 280614 118046 280648
rect 118080 280614 118114 280648
rect 118148 280614 118182 280648
rect 118216 280614 118250 280648
rect 118284 280614 118318 280648
rect 118352 280614 118386 280648
rect 118420 280614 118454 280648
rect 118488 280614 118522 280648
rect 118556 280614 118590 280648
rect 118624 280614 118658 280648
rect 117604 280472 117638 280506
rect 117672 280472 117706 280506
rect 117740 280472 117774 280506
rect 117808 280472 117842 280506
rect 117876 280472 117910 280506
rect 117944 280472 117978 280506
rect 118012 280472 118046 280506
rect 118080 280472 118114 280506
rect 118148 280472 118182 280506
rect 118216 280472 118250 280506
rect 118284 280472 118318 280506
rect 118352 280472 118386 280506
rect 118420 280472 118454 280506
rect 118488 280472 118522 280506
rect 118556 280472 118590 280506
rect 118624 280472 118658 280506
rect 116158 280416 116192 280450
rect 116226 280416 116260 280450
rect 116294 280416 116328 280450
rect 116362 280416 116396 280450
rect 116430 280416 116464 280450
rect 116498 280416 116532 280450
rect 116566 280416 116600 280450
rect 116634 280416 116668 280450
rect 116702 280416 116736 280450
rect 116770 280416 116804 280450
rect 116838 280416 116872 280450
rect 116906 280416 116940 280450
rect 116974 280416 117008 280450
rect 117042 280416 117076 280450
rect 117110 280416 117144 280450
rect 117178 280416 117212 280450
rect 117604 280254 117638 280288
rect 117672 280254 117706 280288
rect 117740 280254 117774 280288
rect 117808 280254 117842 280288
rect 117876 280254 117910 280288
rect 117944 280254 117978 280288
rect 118012 280254 118046 280288
rect 118080 280254 118114 280288
rect 118148 280254 118182 280288
rect 118216 280254 118250 280288
rect 118284 280254 118318 280288
rect 118352 280254 118386 280288
rect 118420 280254 118454 280288
rect 118488 280254 118522 280288
rect 118556 280254 118590 280288
rect 118624 280254 118658 280288
rect 116158 280158 116192 280192
rect 116226 280158 116260 280192
rect 116294 280158 116328 280192
rect 116362 280158 116396 280192
rect 116430 280158 116464 280192
rect 116498 280158 116532 280192
rect 116566 280158 116600 280192
rect 116634 280158 116668 280192
rect 116702 280158 116736 280192
rect 116770 280158 116804 280192
rect 116838 280158 116872 280192
rect 116906 280158 116940 280192
rect 116974 280158 117008 280192
rect 117042 280158 117076 280192
rect 117110 280158 117144 280192
rect 117178 280158 117212 280192
rect 117604 280112 117638 280146
rect 117672 280112 117706 280146
rect 117740 280112 117774 280146
rect 117808 280112 117842 280146
rect 117876 280112 117910 280146
rect 117944 280112 117978 280146
rect 118012 280112 118046 280146
rect 118080 280112 118114 280146
rect 118148 280112 118182 280146
rect 118216 280112 118250 280146
rect 118284 280112 118318 280146
rect 118352 280112 118386 280146
rect 118420 280112 118454 280146
rect 118488 280112 118522 280146
rect 118556 280112 118590 280146
rect 118624 280112 118658 280146
rect 116128 280014 116162 280048
rect 116196 280014 116230 280048
rect 116264 280014 116298 280048
rect 116332 280014 116366 280048
rect 116400 280014 116434 280048
rect 116468 280014 116502 280048
rect 116536 280014 116570 280048
rect 116604 280014 116638 280048
rect 116672 280014 116706 280048
rect 116740 280014 116774 280048
rect 116808 280014 116842 280048
rect 116876 280014 116910 280048
rect 116944 280014 116978 280048
rect 117012 280014 117046 280048
rect 117080 280014 117114 280048
rect 117148 280014 117182 280048
rect 116128 279876 116162 279910
rect 116196 279876 116230 279910
rect 116264 279876 116298 279910
rect 116332 279876 116366 279910
rect 116400 279876 116434 279910
rect 116468 279876 116502 279910
rect 116536 279876 116570 279910
rect 116604 279876 116638 279910
rect 116672 279876 116706 279910
rect 116740 279876 116774 279910
rect 116808 279876 116842 279910
rect 116876 279876 116910 279910
rect 116944 279876 116978 279910
rect 117012 279876 117046 279910
rect 117080 279876 117114 279910
rect 117148 279876 117182 279910
rect 117604 279894 117638 279928
rect 117672 279894 117706 279928
rect 117740 279894 117774 279928
rect 117808 279894 117842 279928
rect 117876 279894 117910 279928
rect 117944 279894 117978 279928
rect 118012 279894 118046 279928
rect 118080 279894 118114 279928
rect 118148 279894 118182 279928
rect 118216 279894 118250 279928
rect 118284 279894 118318 279928
rect 118352 279894 118386 279928
rect 118420 279894 118454 279928
rect 118488 279894 118522 279928
rect 118556 279894 118590 279928
rect 118624 279894 118658 279928
rect 116128 279716 116162 279750
rect 116196 279716 116230 279750
rect 116264 279716 116298 279750
rect 116332 279716 116366 279750
rect 116400 279716 116434 279750
rect 116468 279716 116502 279750
rect 116536 279716 116570 279750
rect 116604 279716 116638 279750
rect 116672 279716 116706 279750
rect 116740 279716 116774 279750
rect 116808 279716 116842 279750
rect 116876 279716 116910 279750
rect 116944 279716 116978 279750
rect 117012 279716 117046 279750
rect 117080 279716 117114 279750
rect 117148 279716 117182 279750
rect 117604 279752 117638 279786
rect 117672 279752 117706 279786
rect 117740 279752 117774 279786
rect 117808 279752 117842 279786
rect 117876 279752 117910 279786
rect 117944 279752 117978 279786
rect 118012 279752 118046 279786
rect 118080 279752 118114 279786
rect 118148 279752 118182 279786
rect 118216 279752 118250 279786
rect 118284 279752 118318 279786
rect 118352 279752 118386 279786
rect 118420 279752 118454 279786
rect 118488 279752 118522 279786
rect 118556 279752 118590 279786
rect 118624 279752 118658 279786
rect 116128 279578 116162 279612
rect 116196 279578 116230 279612
rect 116264 279578 116298 279612
rect 116332 279578 116366 279612
rect 116400 279578 116434 279612
rect 116468 279578 116502 279612
rect 116536 279578 116570 279612
rect 116604 279578 116638 279612
rect 116672 279578 116706 279612
rect 116740 279578 116774 279612
rect 116808 279578 116842 279612
rect 116876 279578 116910 279612
rect 116944 279578 116978 279612
rect 117012 279578 117046 279612
rect 117080 279578 117114 279612
rect 117148 279578 117182 279612
rect 117604 279534 117638 279568
rect 117672 279534 117706 279568
rect 117740 279534 117774 279568
rect 117808 279534 117842 279568
rect 117876 279534 117910 279568
rect 117944 279534 117978 279568
rect 118012 279534 118046 279568
rect 118080 279534 118114 279568
rect 118148 279534 118182 279568
rect 118216 279534 118250 279568
rect 118284 279534 118318 279568
rect 118352 279534 118386 279568
rect 118420 279534 118454 279568
rect 118488 279534 118522 279568
rect 118556 279534 118590 279568
rect 118624 279534 118658 279568
rect 111547 279166 111581 279200
rect 111615 279166 111649 279200
rect 111683 279166 111717 279200
rect 111751 279166 111785 279200
rect 111819 279166 111853 279200
rect 111887 279166 111921 279200
rect 111955 279166 111989 279200
rect 112023 279166 112057 279200
rect 112091 279166 112125 279200
rect 112159 279166 112193 279200
rect 112227 279166 112261 279200
rect 112295 279166 112329 279200
rect 112363 279166 112397 279200
rect 112431 279166 112465 279200
rect 112499 279166 112533 279200
rect 112567 279166 112601 279200
rect 112993 279174 113027 279208
rect 113061 279174 113095 279208
rect 113129 279174 113163 279208
rect 113197 279174 113231 279208
rect 113265 279174 113299 279208
rect 113333 279174 113367 279208
rect 113401 279174 113435 279208
rect 113469 279174 113503 279208
rect 113537 279174 113571 279208
rect 113605 279174 113639 279208
rect 113673 279174 113707 279208
rect 113741 279174 113775 279208
rect 113809 279174 113843 279208
rect 113877 279174 113911 279208
rect 113945 279174 113979 279208
rect 114013 279174 114047 279208
rect 111547 278948 111581 278982
rect 111615 278948 111649 278982
rect 111683 278948 111717 278982
rect 111751 278948 111785 278982
rect 111819 278948 111853 278982
rect 111887 278948 111921 278982
rect 111955 278948 111989 278982
rect 112023 278948 112057 278982
rect 112091 278948 112125 278982
rect 112159 278948 112193 278982
rect 112227 278948 112261 278982
rect 112295 278948 112329 278982
rect 112363 278948 112397 278982
rect 112431 278948 112465 278982
rect 112499 278948 112533 278982
rect 112567 278948 112601 278982
rect 112993 278916 113027 278950
rect 113061 278916 113095 278950
rect 113129 278916 113163 278950
rect 113197 278916 113231 278950
rect 113265 278916 113299 278950
rect 113333 278916 113367 278950
rect 113401 278916 113435 278950
rect 113469 278916 113503 278950
rect 113537 278916 113571 278950
rect 113605 278916 113639 278950
rect 113673 278916 113707 278950
rect 113741 278916 113775 278950
rect 113809 278916 113843 278950
rect 113877 278916 113911 278950
rect 113945 278916 113979 278950
rect 114013 278916 114047 278950
rect 111547 278806 111581 278840
rect 111615 278806 111649 278840
rect 111683 278806 111717 278840
rect 111751 278806 111785 278840
rect 111819 278806 111853 278840
rect 111887 278806 111921 278840
rect 111955 278806 111989 278840
rect 112023 278806 112057 278840
rect 112091 278806 112125 278840
rect 112159 278806 112193 278840
rect 112227 278806 112261 278840
rect 112295 278806 112329 278840
rect 112363 278806 112397 278840
rect 112431 278806 112465 278840
rect 112499 278806 112533 278840
rect 112567 278806 112601 278840
rect 112993 278750 113027 278784
rect 113061 278750 113095 278784
rect 113129 278750 113163 278784
rect 113197 278750 113231 278784
rect 113265 278750 113299 278784
rect 113333 278750 113367 278784
rect 113401 278750 113435 278784
rect 113469 278750 113503 278784
rect 113537 278750 113571 278784
rect 113605 278750 113639 278784
rect 113673 278750 113707 278784
rect 113741 278750 113775 278784
rect 113809 278750 113843 278784
rect 113877 278750 113911 278784
rect 113945 278750 113979 278784
rect 114013 278750 114047 278784
rect 111547 278588 111581 278622
rect 111615 278588 111649 278622
rect 111683 278588 111717 278622
rect 111751 278588 111785 278622
rect 111819 278588 111853 278622
rect 111887 278588 111921 278622
rect 111955 278588 111989 278622
rect 112023 278588 112057 278622
rect 112091 278588 112125 278622
rect 112159 278588 112193 278622
rect 112227 278588 112261 278622
rect 112295 278588 112329 278622
rect 112363 278588 112397 278622
rect 112431 278588 112465 278622
rect 112499 278588 112533 278622
rect 112567 278588 112601 278622
rect 112993 278492 113027 278526
rect 113061 278492 113095 278526
rect 113129 278492 113163 278526
rect 113197 278492 113231 278526
rect 113265 278492 113299 278526
rect 113333 278492 113367 278526
rect 113401 278492 113435 278526
rect 113469 278492 113503 278526
rect 113537 278492 113571 278526
rect 113605 278492 113639 278526
rect 113673 278492 113707 278526
rect 113741 278492 113775 278526
rect 113809 278492 113843 278526
rect 113877 278492 113911 278526
rect 113945 278492 113979 278526
rect 114013 278492 114047 278526
rect 111547 278446 111581 278480
rect 111615 278446 111649 278480
rect 111683 278446 111717 278480
rect 111751 278446 111785 278480
rect 111819 278446 111853 278480
rect 111887 278446 111921 278480
rect 111955 278446 111989 278480
rect 112023 278446 112057 278480
rect 112091 278446 112125 278480
rect 112159 278446 112193 278480
rect 112227 278446 112261 278480
rect 112295 278446 112329 278480
rect 112363 278446 112397 278480
rect 112431 278446 112465 278480
rect 112499 278446 112533 278480
rect 112567 278446 112601 278480
rect 113023 278348 113057 278382
rect 113091 278348 113125 278382
rect 113159 278348 113193 278382
rect 113227 278348 113261 278382
rect 113295 278348 113329 278382
rect 113363 278348 113397 278382
rect 113431 278348 113465 278382
rect 113499 278348 113533 278382
rect 113567 278348 113601 278382
rect 113635 278348 113669 278382
rect 113703 278348 113737 278382
rect 113771 278348 113805 278382
rect 113839 278348 113873 278382
rect 113907 278348 113941 278382
rect 113975 278348 114009 278382
rect 114043 278348 114077 278382
rect 111547 278228 111581 278262
rect 111615 278228 111649 278262
rect 111683 278228 111717 278262
rect 111751 278228 111785 278262
rect 111819 278228 111853 278262
rect 111887 278228 111921 278262
rect 111955 278228 111989 278262
rect 112023 278228 112057 278262
rect 112091 278228 112125 278262
rect 112159 278228 112193 278262
rect 112227 278228 112261 278262
rect 112295 278228 112329 278262
rect 112363 278228 112397 278262
rect 112431 278228 112465 278262
rect 112499 278228 112533 278262
rect 112567 278228 112601 278262
rect 113023 278210 113057 278244
rect 113091 278210 113125 278244
rect 113159 278210 113193 278244
rect 113227 278210 113261 278244
rect 113295 278210 113329 278244
rect 113363 278210 113397 278244
rect 113431 278210 113465 278244
rect 113499 278210 113533 278244
rect 113567 278210 113601 278244
rect 113635 278210 113669 278244
rect 113703 278210 113737 278244
rect 113771 278210 113805 278244
rect 113839 278210 113873 278244
rect 113907 278210 113941 278244
rect 113975 278210 114009 278244
rect 114043 278210 114077 278244
rect 111547 278086 111581 278120
rect 111615 278086 111649 278120
rect 111683 278086 111717 278120
rect 111751 278086 111785 278120
rect 111819 278086 111853 278120
rect 111887 278086 111921 278120
rect 111955 278086 111989 278120
rect 112023 278086 112057 278120
rect 112091 278086 112125 278120
rect 112159 278086 112193 278120
rect 112227 278086 112261 278120
rect 112295 278086 112329 278120
rect 112363 278086 112397 278120
rect 112431 278086 112465 278120
rect 112499 278086 112533 278120
rect 112567 278086 112601 278120
rect 113023 278050 113057 278084
rect 113091 278050 113125 278084
rect 113159 278050 113193 278084
rect 113227 278050 113261 278084
rect 113295 278050 113329 278084
rect 113363 278050 113397 278084
rect 113431 278050 113465 278084
rect 113499 278050 113533 278084
rect 113567 278050 113601 278084
rect 113635 278050 113669 278084
rect 113703 278050 113737 278084
rect 113771 278050 113805 278084
rect 113839 278050 113873 278084
rect 113907 278050 113941 278084
rect 113975 278050 114009 278084
rect 114043 278050 114077 278084
rect 111547 277868 111581 277902
rect 111615 277868 111649 277902
rect 111683 277868 111717 277902
rect 111751 277868 111785 277902
rect 111819 277868 111853 277902
rect 111887 277868 111921 277902
rect 111955 277868 111989 277902
rect 112023 277868 112057 277902
rect 112091 277868 112125 277902
rect 112159 277868 112193 277902
rect 112227 277868 112261 277902
rect 112295 277868 112329 277902
rect 112363 277868 112397 277902
rect 112431 277868 112465 277902
rect 112499 277868 112533 277902
rect 112567 277868 112601 277902
rect 113023 277912 113057 277946
rect 113091 277912 113125 277946
rect 113159 277912 113193 277946
rect 113227 277912 113261 277946
rect 113295 277912 113329 277946
rect 113363 277912 113397 277946
rect 113431 277912 113465 277946
rect 113499 277912 113533 277946
rect 113567 277912 113601 277946
rect 113635 277912 113669 277946
rect 113703 277912 113737 277946
rect 113771 277912 113805 277946
rect 113839 277912 113873 277946
rect 113907 277912 113941 277946
rect 113975 277912 114009 277946
rect 114043 277912 114077 277946
rect 116158 279174 116192 279208
rect 116226 279174 116260 279208
rect 116294 279174 116328 279208
rect 116362 279174 116396 279208
rect 116430 279174 116464 279208
rect 116498 279174 116532 279208
rect 116566 279174 116600 279208
rect 116634 279174 116668 279208
rect 116702 279174 116736 279208
rect 116770 279174 116804 279208
rect 116838 279174 116872 279208
rect 116906 279174 116940 279208
rect 116974 279174 117008 279208
rect 117042 279174 117076 279208
rect 117110 279174 117144 279208
rect 117178 279174 117212 279208
rect 117604 279166 117638 279200
rect 117672 279166 117706 279200
rect 117740 279166 117774 279200
rect 117808 279166 117842 279200
rect 117876 279166 117910 279200
rect 117944 279166 117978 279200
rect 118012 279166 118046 279200
rect 118080 279166 118114 279200
rect 118148 279166 118182 279200
rect 118216 279166 118250 279200
rect 118284 279166 118318 279200
rect 118352 279166 118386 279200
rect 118420 279166 118454 279200
rect 118488 279166 118522 279200
rect 118556 279166 118590 279200
rect 118624 279166 118658 279200
rect 116158 278916 116192 278950
rect 116226 278916 116260 278950
rect 116294 278916 116328 278950
rect 116362 278916 116396 278950
rect 116430 278916 116464 278950
rect 116498 278916 116532 278950
rect 116566 278916 116600 278950
rect 116634 278916 116668 278950
rect 116702 278916 116736 278950
rect 116770 278916 116804 278950
rect 116838 278916 116872 278950
rect 116906 278916 116940 278950
rect 116974 278916 117008 278950
rect 117042 278916 117076 278950
rect 117110 278916 117144 278950
rect 117178 278916 117212 278950
rect 117604 278948 117638 278982
rect 117672 278948 117706 278982
rect 117740 278948 117774 278982
rect 117808 278948 117842 278982
rect 117876 278948 117910 278982
rect 117944 278948 117978 278982
rect 118012 278948 118046 278982
rect 118080 278948 118114 278982
rect 118148 278948 118182 278982
rect 118216 278948 118250 278982
rect 118284 278948 118318 278982
rect 118352 278948 118386 278982
rect 118420 278948 118454 278982
rect 118488 278948 118522 278982
rect 118556 278948 118590 278982
rect 118624 278948 118658 278982
rect 117604 278806 117638 278840
rect 117672 278806 117706 278840
rect 117740 278806 117774 278840
rect 117808 278806 117842 278840
rect 117876 278806 117910 278840
rect 117944 278806 117978 278840
rect 118012 278806 118046 278840
rect 118080 278806 118114 278840
rect 118148 278806 118182 278840
rect 118216 278806 118250 278840
rect 118284 278806 118318 278840
rect 118352 278806 118386 278840
rect 118420 278806 118454 278840
rect 118488 278806 118522 278840
rect 118556 278806 118590 278840
rect 118624 278806 118658 278840
rect 116158 278750 116192 278784
rect 116226 278750 116260 278784
rect 116294 278750 116328 278784
rect 116362 278750 116396 278784
rect 116430 278750 116464 278784
rect 116498 278750 116532 278784
rect 116566 278750 116600 278784
rect 116634 278750 116668 278784
rect 116702 278750 116736 278784
rect 116770 278750 116804 278784
rect 116838 278750 116872 278784
rect 116906 278750 116940 278784
rect 116974 278750 117008 278784
rect 117042 278750 117076 278784
rect 117110 278750 117144 278784
rect 117178 278750 117212 278784
rect 117604 278588 117638 278622
rect 117672 278588 117706 278622
rect 117740 278588 117774 278622
rect 117808 278588 117842 278622
rect 117876 278588 117910 278622
rect 117944 278588 117978 278622
rect 118012 278588 118046 278622
rect 118080 278588 118114 278622
rect 118148 278588 118182 278622
rect 118216 278588 118250 278622
rect 118284 278588 118318 278622
rect 118352 278588 118386 278622
rect 118420 278588 118454 278622
rect 118488 278588 118522 278622
rect 118556 278588 118590 278622
rect 118624 278588 118658 278622
rect 116158 278492 116192 278526
rect 116226 278492 116260 278526
rect 116294 278492 116328 278526
rect 116362 278492 116396 278526
rect 116430 278492 116464 278526
rect 116498 278492 116532 278526
rect 116566 278492 116600 278526
rect 116634 278492 116668 278526
rect 116702 278492 116736 278526
rect 116770 278492 116804 278526
rect 116838 278492 116872 278526
rect 116906 278492 116940 278526
rect 116974 278492 117008 278526
rect 117042 278492 117076 278526
rect 117110 278492 117144 278526
rect 117178 278492 117212 278526
rect 117604 278446 117638 278480
rect 117672 278446 117706 278480
rect 117740 278446 117774 278480
rect 117808 278446 117842 278480
rect 117876 278446 117910 278480
rect 117944 278446 117978 278480
rect 118012 278446 118046 278480
rect 118080 278446 118114 278480
rect 118148 278446 118182 278480
rect 118216 278446 118250 278480
rect 118284 278446 118318 278480
rect 118352 278446 118386 278480
rect 118420 278446 118454 278480
rect 118488 278446 118522 278480
rect 118556 278446 118590 278480
rect 118624 278446 118658 278480
rect 116128 278348 116162 278382
rect 116196 278348 116230 278382
rect 116264 278348 116298 278382
rect 116332 278348 116366 278382
rect 116400 278348 116434 278382
rect 116468 278348 116502 278382
rect 116536 278348 116570 278382
rect 116604 278348 116638 278382
rect 116672 278348 116706 278382
rect 116740 278348 116774 278382
rect 116808 278348 116842 278382
rect 116876 278348 116910 278382
rect 116944 278348 116978 278382
rect 117012 278348 117046 278382
rect 117080 278348 117114 278382
rect 117148 278348 117182 278382
rect 116128 278210 116162 278244
rect 116196 278210 116230 278244
rect 116264 278210 116298 278244
rect 116332 278210 116366 278244
rect 116400 278210 116434 278244
rect 116468 278210 116502 278244
rect 116536 278210 116570 278244
rect 116604 278210 116638 278244
rect 116672 278210 116706 278244
rect 116740 278210 116774 278244
rect 116808 278210 116842 278244
rect 116876 278210 116910 278244
rect 116944 278210 116978 278244
rect 117012 278210 117046 278244
rect 117080 278210 117114 278244
rect 117148 278210 117182 278244
rect 117604 278228 117638 278262
rect 117672 278228 117706 278262
rect 117740 278228 117774 278262
rect 117808 278228 117842 278262
rect 117876 278228 117910 278262
rect 117944 278228 117978 278262
rect 118012 278228 118046 278262
rect 118080 278228 118114 278262
rect 118148 278228 118182 278262
rect 118216 278228 118250 278262
rect 118284 278228 118318 278262
rect 118352 278228 118386 278262
rect 118420 278228 118454 278262
rect 118488 278228 118522 278262
rect 118556 278228 118590 278262
rect 118624 278228 118658 278262
rect 116128 278050 116162 278084
rect 116196 278050 116230 278084
rect 116264 278050 116298 278084
rect 116332 278050 116366 278084
rect 116400 278050 116434 278084
rect 116468 278050 116502 278084
rect 116536 278050 116570 278084
rect 116604 278050 116638 278084
rect 116672 278050 116706 278084
rect 116740 278050 116774 278084
rect 116808 278050 116842 278084
rect 116876 278050 116910 278084
rect 116944 278050 116978 278084
rect 117012 278050 117046 278084
rect 117080 278050 117114 278084
rect 117148 278050 117182 278084
rect 117604 278086 117638 278120
rect 117672 278086 117706 278120
rect 117740 278086 117774 278120
rect 117808 278086 117842 278120
rect 117876 278086 117910 278120
rect 117944 278086 117978 278120
rect 118012 278086 118046 278120
rect 118080 278086 118114 278120
rect 118148 278086 118182 278120
rect 118216 278086 118250 278120
rect 118284 278086 118318 278120
rect 118352 278086 118386 278120
rect 118420 278086 118454 278120
rect 118488 278086 118522 278120
rect 118556 278086 118590 278120
rect 118624 278086 118658 278120
rect 116128 277912 116162 277946
rect 116196 277912 116230 277946
rect 116264 277912 116298 277946
rect 116332 277912 116366 277946
rect 116400 277912 116434 277946
rect 116468 277912 116502 277946
rect 116536 277912 116570 277946
rect 116604 277912 116638 277946
rect 116672 277912 116706 277946
rect 116740 277912 116774 277946
rect 116808 277912 116842 277946
rect 116876 277912 116910 277946
rect 116944 277912 116978 277946
rect 117012 277912 117046 277946
rect 117080 277912 117114 277946
rect 117148 277912 117182 277946
rect 117604 277868 117638 277902
rect 117672 277868 117706 277902
rect 117740 277868 117774 277902
rect 117808 277868 117842 277902
rect 117876 277868 117910 277902
rect 117944 277868 117978 277902
rect 118012 277868 118046 277902
rect 118080 277868 118114 277902
rect 118148 277868 118182 277902
rect 118216 277868 118250 277902
rect 118284 277868 118318 277902
rect 118352 277868 118386 277902
rect 118420 277868 118454 277902
rect 118488 277868 118522 277902
rect 118556 277868 118590 277902
rect 118624 277868 118658 277902
rect 111547 277500 111581 277534
rect 111615 277500 111649 277534
rect 111683 277500 111717 277534
rect 111751 277500 111785 277534
rect 111819 277500 111853 277534
rect 111887 277500 111921 277534
rect 111955 277500 111989 277534
rect 112023 277500 112057 277534
rect 112091 277500 112125 277534
rect 112159 277500 112193 277534
rect 112227 277500 112261 277534
rect 112295 277500 112329 277534
rect 112363 277500 112397 277534
rect 112431 277500 112465 277534
rect 112499 277500 112533 277534
rect 112567 277500 112601 277534
rect 112993 277508 113027 277542
rect 113061 277508 113095 277542
rect 113129 277508 113163 277542
rect 113197 277508 113231 277542
rect 113265 277508 113299 277542
rect 113333 277508 113367 277542
rect 113401 277508 113435 277542
rect 113469 277508 113503 277542
rect 113537 277508 113571 277542
rect 113605 277508 113639 277542
rect 113673 277508 113707 277542
rect 113741 277508 113775 277542
rect 113809 277508 113843 277542
rect 113877 277508 113911 277542
rect 113945 277508 113979 277542
rect 114013 277508 114047 277542
rect 111547 277282 111581 277316
rect 111615 277282 111649 277316
rect 111683 277282 111717 277316
rect 111751 277282 111785 277316
rect 111819 277282 111853 277316
rect 111887 277282 111921 277316
rect 111955 277282 111989 277316
rect 112023 277282 112057 277316
rect 112091 277282 112125 277316
rect 112159 277282 112193 277316
rect 112227 277282 112261 277316
rect 112295 277282 112329 277316
rect 112363 277282 112397 277316
rect 112431 277282 112465 277316
rect 112499 277282 112533 277316
rect 112567 277282 112601 277316
rect 112993 277250 113027 277284
rect 113061 277250 113095 277284
rect 113129 277250 113163 277284
rect 113197 277250 113231 277284
rect 113265 277250 113299 277284
rect 113333 277250 113367 277284
rect 113401 277250 113435 277284
rect 113469 277250 113503 277284
rect 113537 277250 113571 277284
rect 113605 277250 113639 277284
rect 113673 277250 113707 277284
rect 113741 277250 113775 277284
rect 113809 277250 113843 277284
rect 113877 277250 113911 277284
rect 113945 277250 113979 277284
rect 114013 277250 114047 277284
rect 111547 277140 111581 277174
rect 111615 277140 111649 277174
rect 111683 277140 111717 277174
rect 111751 277140 111785 277174
rect 111819 277140 111853 277174
rect 111887 277140 111921 277174
rect 111955 277140 111989 277174
rect 112023 277140 112057 277174
rect 112091 277140 112125 277174
rect 112159 277140 112193 277174
rect 112227 277140 112261 277174
rect 112295 277140 112329 277174
rect 112363 277140 112397 277174
rect 112431 277140 112465 277174
rect 112499 277140 112533 277174
rect 112567 277140 112601 277174
rect 112993 277084 113027 277118
rect 113061 277084 113095 277118
rect 113129 277084 113163 277118
rect 113197 277084 113231 277118
rect 113265 277084 113299 277118
rect 113333 277084 113367 277118
rect 113401 277084 113435 277118
rect 113469 277084 113503 277118
rect 113537 277084 113571 277118
rect 113605 277084 113639 277118
rect 113673 277084 113707 277118
rect 113741 277084 113775 277118
rect 113809 277084 113843 277118
rect 113877 277084 113911 277118
rect 113945 277084 113979 277118
rect 114013 277084 114047 277118
rect 111547 276922 111581 276956
rect 111615 276922 111649 276956
rect 111683 276922 111717 276956
rect 111751 276922 111785 276956
rect 111819 276922 111853 276956
rect 111887 276922 111921 276956
rect 111955 276922 111989 276956
rect 112023 276922 112057 276956
rect 112091 276922 112125 276956
rect 112159 276922 112193 276956
rect 112227 276922 112261 276956
rect 112295 276922 112329 276956
rect 112363 276922 112397 276956
rect 112431 276922 112465 276956
rect 112499 276922 112533 276956
rect 112567 276922 112601 276956
rect 112993 276826 113027 276860
rect 113061 276826 113095 276860
rect 113129 276826 113163 276860
rect 113197 276826 113231 276860
rect 113265 276826 113299 276860
rect 113333 276826 113367 276860
rect 113401 276826 113435 276860
rect 113469 276826 113503 276860
rect 113537 276826 113571 276860
rect 113605 276826 113639 276860
rect 113673 276826 113707 276860
rect 113741 276826 113775 276860
rect 113809 276826 113843 276860
rect 113877 276826 113911 276860
rect 113945 276826 113979 276860
rect 114013 276826 114047 276860
rect 111547 276780 111581 276814
rect 111615 276780 111649 276814
rect 111683 276780 111717 276814
rect 111751 276780 111785 276814
rect 111819 276780 111853 276814
rect 111887 276780 111921 276814
rect 111955 276780 111989 276814
rect 112023 276780 112057 276814
rect 112091 276780 112125 276814
rect 112159 276780 112193 276814
rect 112227 276780 112261 276814
rect 112295 276780 112329 276814
rect 112363 276780 112397 276814
rect 112431 276780 112465 276814
rect 112499 276780 112533 276814
rect 112567 276780 112601 276814
rect 113023 276682 113057 276716
rect 113091 276682 113125 276716
rect 113159 276682 113193 276716
rect 113227 276682 113261 276716
rect 113295 276682 113329 276716
rect 113363 276682 113397 276716
rect 113431 276682 113465 276716
rect 113499 276682 113533 276716
rect 113567 276682 113601 276716
rect 113635 276682 113669 276716
rect 113703 276682 113737 276716
rect 113771 276682 113805 276716
rect 113839 276682 113873 276716
rect 113907 276682 113941 276716
rect 113975 276682 114009 276716
rect 114043 276682 114077 276716
rect 111547 276562 111581 276596
rect 111615 276562 111649 276596
rect 111683 276562 111717 276596
rect 111751 276562 111785 276596
rect 111819 276562 111853 276596
rect 111887 276562 111921 276596
rect 111955 276562 111989 276596
rect 112023 276562 112057 276596
rect 112091 276562 112125 276596
rect 112159 276562 112193 276596
rect 112227 276562 112261 276596
rect 112295 276562 112329 276596
rect 112363 276562 112397 276596
rect 112431 276562 112465 276596
rect 112499 276562 112533 276596
rect 112567 276562 112601 276596
rect 113023 276544 113057 276578
rect 113091 276544 113125 276578
rect 113159 276544 113193 276578
rect 113227 276544 113261 276578
rect 113295 276544 113329 276578
rect 113363 276544 113397 276578
rect 113431 276544 113465 276578
rect 113499 276544 113533 276578
rect 113567 276544 113601 276578
rect 113635 276544 113669 276578
rect 113703 276544 113737 276578
rect 113771 276544 113805 276578
rect 113839 276544 113873 276578
rect 113907 276544 113941 276578
rect 113975 276544 114009 276578
rect 114043 276544 114077 276578
rect 111547 276420 111581 276454
rect 111615 276420 111649 276454
rect 111683 276420 111717 276454
rect 111751 276420 111785 276454
rect 111819 276420 111853 276454
rect 111887 276420 111921 276454
rect 111955 276420 111989 276454
rect 112023 276420 112057 276454
rect 112091 276420 112125 276454
rect 112159 276420 112193 276454
rect 112227 276420 112261 276454
rect 112295 276420 112329 276454
rect 112363 276420 112397 276454
rect 112431 276420 112465 276454
rect 112499 276420 112533 276454
rect 112567 276420 112601 276454
rect 113023 276384 113057 276418
rect 113091 276384 113125 276418
rect 113159 276384 113193 276418
rect 113227 276384 113261 276418
rect 113295 276384 113329 276418
rect 113363 276384 113397 276418
rect 113431 276384 113465 276418
rect 113499 276384 113533 276418
rect 113567 276384 113601 276418
rect 113635 276384 113669 276418
rect 113703 276384 113737 276418
rect 113771 276384 113805 276418
rect 113839 276384 113873 276418
rect 113907 276384 113941 276418
rect 113975 276384 114009 276418
rect 114043 276384 114077 276418
rect 111547 276202 111581 276236
rect 111615 276202 111649 276236
rect 111683 276202 111717 276236
rect 111751 276202 111785 276236
rect 111819 276202 111853 276236
rect 111887 276202 111921 276236
rect 111955 276202 111989 276236
rect 112023 276202 112057 276236
rect 112091 276202 112125 276236
rect 112159 276202 112193 276236
rect 112227 276202 112261 276236
rect 112295 276202 112329 276236
rect 112363 276202 112397 276236
rect 112431 276202 112465 276236
rect 112499 276202 112533 276236
rect 112567 276202 112601 276236
rect 113023 276246 113057 276280
rect 113091 276246 113125 276280
rect 113159 276246 113193 276280
rect 113227 276246 113261 276280
rect 113295 276246 113329 276280
rect 113363 276246 113397 276280
rect 113431 276246 113465 276280
rect 113499 276246 113533 276280
rect 113567 276246 113601 276280
rect 113635 276246 113669 276280
rect 113703 276246 113737 276280
rect 113771 276246 113805 276280
rect 113839 276246 113873 276280
rect 113907 276246 113941 276280
rect 113975 276246 114009 276280
rect 114043 276246 114077 276280
rect 116158 277508 116192 277542
rect 116226 277508 116260 277542
rect 116294 277508 116328 277542
rect 116362 277508 116396 277542
rect 116430 277508 116464 277542
rect 116498 277508 116532 277542
rect 116566 277508 116600 277542
rect 116634 277508 116668 277542
rect 116702 277508 116736 277542
rect 116770 277508 116804 277542
rect 116838 277508 116872 277542
rect 116906 277508 116940 277542
rect 116974 277508 117008 277542
rect 117042 277508 117076 277542
rect 117110 277508 117144 277542
rect 117178 277508 117212 277542
rect 117604 277500 117638 277534
rect 117672 277500 117706 277534
rect 117740 277500 117774 277534
rect 117808 277500 117842 277534
rect 117876 277500 117910 277534
rect 117944 277500 117978 277534
rect 118012 277500 118046 277534
rect 118080 277500 118114 277534
rect 118148 277500 118182 277534
rect 118216 277500 118250 277534
rect 118284 277500 118318 277534
rect 118352 277500 118386 277534
rect 118420 277500 118454 277534
rect 118488 277500 118522 277534
rect 118556 277500 118590 277534
rect 118624 277500 118658 277534
rect 116158 277250 116192 277284
rect 116226 277250 116260 277284
rect 116294 277250 116328 277284
rect 116362 277250 116396 277284
rect 116430 277250 116464 277284
rect 116498 277250 116532 277284
rect 116566 277250 116600 277284
rect 116634 277250 116668 277284
rect 116702 277250 116736 277284
rect 116770 277250 116804 277284
rect 116838 277250 116872 277284
rect 116906 277250 116940 277284
rect 116974 277250 117008 277284
rect 117042 277250 117076 277284
rect 117110 277250 117144 277284
rect 117178 277250 117212 277284
rect 117604 277282 117638 277316
rect 117672 277282 117706 277316
rect 117740 277282 117774 277316
rect 117808 277282 117842 277316
rect 117876 277282 117910 277316
rect 117944 277282 117978 277316
rect 118012 277282 118046 277316
rect 118080 277282 118114 277316
rect 118148 277282 118182 277316
rect 118216 277282 118250 277316
rect 118284 277282 118318 277316
rect 118352 277282 118386 277316
rect 118420 277282 118454 277316
rect 118488 277282 118522 277316
rect 118556 277282 118590 277316
rect 118624 277282 118658 277316
rect 117604 277140 117638 277174
rect 117672 277140 117706 277174
rect 117740 277140 117774 277174
rect 117808 277140 117842 277174
rect 117876 277140 117910 277174
rect 117944 277140 117978 277174
rect 118012 277140 118046 277174
rect 118080 277140 118114 277174
rect 118148 277140 118182 277174
rect 118216 277140 118250 277174
rect 118284 277140 118318 277174
rect 118352 277140 118386 277174
rect 118420 277140 118454 277174
rect 118488 277140 118522 277174
rect 118556 277140 118590 277174
rect 118624 277140 118658 277174
rect 116158 277084 116192 277118
rect 116226 277084 116260 277118
rect 116294 277084 116328 277118
rect 116362 277084 116396 277118
rect 116430 277084 116464 277118
rect 116498 277084 116532 277118
rect 116566 277084 116600 277118
rect 116634 277084 116668 277118
rect 116702 277084 116736 277118
rect 116770 277084 116804 277118
rect 116838 277084 116872 277118
rect 116906 277084 116940 277118
rect 116974 277084 117008 277118
rect 117042 277084 117076 277118
rect 117110 277084 117144 277118
rect 117178 277084 117212 277118
rect 117604 276922 117638 276956
rect 117672 276922 117706 276956
rect 117740 276922 117774 276956
rect 117808 276922 117842 276956
rect 117876 276922 117910 276956
rect 117944 276922 117978 276956
rect 118012 276922 118046 276956
rect 118080 276922 118114 276956
rect 118148 276922 118182 276956
rect 118216 276922 118250 276956
rect 118284 276922 118318 276956
rect 118352 276922 118386 276956
rect 118420 276922 118454 276956
rect 118488 276922 118522 276956
rect 118556 276922 118590 276956
rect 118624 276922 118658 276956
rect 116158 276826 116192 276860
rect 116226 276826 116260 276860
rect 116294 276826 116328 276860
rect 116362 276826 116396 276860
rect 116430 276826 116464 276860
rect 116498 276826 116532 276860
rect 116566 276826 116600 276860
rect 116634 276826 116668 276860
rect 116702 276826 116736 276860
rect 116770 276826 116804 276860
rect 116838 276826 116872 276860
rect 116906 276826 116940 276860
rect 116974 276826 117008 276860
rect 117042 276826 117076 276860
rect 117110 276826 117144 276860
rect 117178 276826 117212 276860
rect 117604 276780 117638 276814
rect 117672 276780 117706 276814
rect 117740 276780 117774 276814
rect 117808 276780 117842 276814
rect 117876 276780 117910 276814
rect 117944 276780 117978 276814
rect 118012 276780 118046 276814
rect 118080 276780 118114 276814
rect 118148 276780 118182 276814
rect 118216 276780 118250 276814
rect 118284 276780 118318 276814
rect 118352 276780 118386 276814
rect 118420 276780 118454 276814
rect 118488 276780 118522 276814
rect 118556 276780 118590 276814
rect 118624 276780 118658 276814
rect 116128 276682 116162 276716
rect 116196 276682 116230 276716
rect 116264 276682 116298 276716
rect 116332 276682 116366 276716
rect 116400 276682 116434 276716
rect 116468 276682 116502 276716
rect 116536 276682 116570 276716
rect 116604 276682 116638 276716
rect 116672 276682 116706 276716
rect 116740 276682 116774 276716
rect 116808 276682 116842 276716
rect 116876 276682 116910 276716
rect 116944 276682 116978 276716
rect 117012 276682 117046 276716
rect 117080 276682 117114 276716
rect 117148 276682 117182 276716
rect 116128 276544 116162 276578
rect 116196 276544 116230 276578
rect 116264 276544 116298 276578
rect 116332 276544 116366 276578
rect 116400 276544 116434 276578
rect 116468 276544 116502 276578
rect 116536 276544 116570 276578
rect 116604 276544 116638 276578
rect 116672 276544 116706 276578
rect 116740 276544 116774 276578
rect 116808 276544 116842 276578
rect 116876 276544 116910 276578
rect 116944 276544 116978 276578
rect 117012 276544 117046 276578
rect 117080 276544 117114 276578
rect 117148 276544 117182 276578
rect 117604 276562 117638 276596
rect 117672 276562 117706 276596
rect 117740 276562 117774 276596
rect 117808 276562 117842 276596
rect 117876 276562 117910 276596
rect 117944 276562 117978 276596
rect 118012 276562 118046 276596
rect 118080 276562 118114 276596
rect 118148 276562 118182 276596
rect 118216 276562 118250 276596
rect 118284 276562 118318 276596
rect 118352 276562 118386 276596
rect 118420 276562 118454 276596
rect 118488 276562 118522 276596
rect 118556 276562 118590 276596
rect 118624 276562 118658 276596
rect 116128 276384 116162 276418
rect 116196 276384 116230 276418
rect 116264 276384 116298 276418
rect 116332 276384 116366 276418
rect 116400 276384 116434 276418
rect 116468 276384 116502 276418
rect 116536 276384 116570 276418
rect 116604 276384 116638 276418
rect 116672 276384 116706 276418
rect 116740 276384 116774 276418
rect 116808 276384 116842 276418
rect 116876 276384 116910 276418
rect 116944 276384 116978 276418
rect 117012 276384 117046 276418
rect 117080 276384 117114 276418
rect 117148 276384 117182 276418
rect 117604 276420 117638 276454
rect 117672 276420 117706 276454
rect 117740 276420 117774 276454
rect 117808 276420 117842 276454
rect 117876 276420 117910 276454
rect 117944 276420 117978 276454
rect 118012 276420 118046 276454
rect 118080 276420 118114 276454
rect 118148 276420 118182 276454
rect 118216 276420 118250 276454
rect 118284 276420 118318 276454
rect 118352 276420 118386 276454
rect 118420 276420 118454 276454
rect 118488 276420 118522 276454
rect 118556 276420 118590 276454
rect 118624 276420 118658 276454
rect 116128 276246 116162 276280
rect 116196 276246 116230 276280
rect 116264 276246 116298 276280
rect 116332 276246 116366 276280
rect 116400 276246 116434 276280
rect 116468 276246 116502 276280
rect 116536 276246 116570 276280
rect 116604 276246 116638 276280
rect 116672 276246 116706 276280
rect 116740 276246 116774 276280
rect 116808 276246 116842 276280
rect 116876 276246 116910 276280
rect 116944 276246 116978 276280
rect 117012 276246 117046 276280
rect 117080 276246 117114 276280
rect 117148 276246 117182 276280
rect 117604 276202 117638 276236
rect 117672 276202 117706 276236
rect 117740 276202 117774 276236
rect 117808 276202 117842 276236
rect 117876 276202 117910 276236
rect 117944 276202 117978 276236
rect 118012 276202 118046 276236
rect 118080 276202 118114 276236
rect 118148 276202 118182 276236
rect 118216 276202 118250 276236
rect 118284 276202 118318 276236
rect 118352 276202 118386 276236
rect 118420 276202 118454 276236
rect 118488 276202 118522 276236
rect 118556 276202 118590 276236
rect 118624 276202 118658 276236
rect 111547 275834 111581 275868
rect 111615 275834 111649 275868
rect 111683 275834 111717 275868
rect 111751 275834 111785 275868
rect 111819 275834 111853 275868
rect 111887 275834 111921 275868
rect 111955 275834 111989 275868
rect 112023 275834 112057 275868
rect 112091 275834 112125 275868
rect 112159 275834 112193 275868
rect 112227 275834 112261 275868
rect 112295 275834 112329 275868
rect 112363 275834 112397 275868
rect 112431 275834 112465 275868
rect 112499 275834 112533 275868
rect 112567 275834 112601 275868
rect 112993 275842 113027 275876
rect 113061 275842 113095 275876
rect 113129 275842 113163 275876
rect 113197 275842 113231 275876
rect 113265 275842 113299 275876
rect 113333 275842 113367 275876
rect 113401 275842 113435 275876
rect 113469 275842 113503 275876
rect 113537 275842 113571 275876
rect 113605 275842 113639 275876
rect 113673 275842 113707 275876
rect 113741 275842 113775 275876
rect 113809 275842 113843 275876
rect 113877 275842 113911 275876
rect 113945 275842 113979 275876
rect 114013 275842 114047 275876
rect 111547 275616 111581 275650
rect 111615 275616 111649 275650
rect 111683 275616 111717 275650
rect 111751 275616 111785 275650
rect 111819 275616 111853 275650
rect 111887 275616 111921 275650
rect 111955 275616 111989 275650
rect 112023 275616 112057 275650
rect 112091 275616 112125 275650
rect 112159 275616 112193 275650
rect 112227 275616 112261 275650
rect 112295 275616 112329 275650
rect 112363 275616 112397 275650
rect 112431 275616 112465 275650
rect 112499 275616 112533 275650
rect 112567 275616 112601 275650
rect 112993 275584 113027 275618
rect 113061 275584 113095 275618
rect 113129 275584 113163 275618
rect 113197 275584 113231 275618
rect 113265 275584 113299 275618
rect 113333 275584 113367 275618
rect 113401 275584 113435 275618
rect 113469 275584 113503 275618
rect 113537 275584 113571 275618
rect 113605 275584 113639 275618
rect 113673 275584 113707 275618
rect 113741 275584 113775 275618
rect 113809 275584 113843 275618
rect 113877 275584 113911 275618
rect 113945 275584 113979 275618
rect 114013 275584 114047 275618
rect 111547 275474 111581 275508
rect 111615 275474 111649 275508
rect 111683 275474 111717 275508
rect 111751 275474 111785 275508
rect 111819 275474 111853 275508
rect 111887 275474 111921 275508
rect 111955 275474 111989 275508
rect 112023 275474 112057 275508
rect 112091 275474 112125 275508
rect 112159 275474 112193 275508
rect 112227 275474 112261 275508
rect 112295 275474 112329 275508
rect 112363 275474 112397 275508
rect 112431 275474 112465 275508
rect 112499 275474 112533 275508
rect 112567 275474 112601 275508
rect 112993 275418 113027 275452
rect 113061 275418 113095 275452
rect 113129 275418 113163 275452
rect 113197 275418 113231 275452
rect 113265 275418 113299 275452
rect 113333 275418 113367 275452
rect 113401 275418 113435 275452
rect 113469 275418 113503 275452
rect 113537 275418 113571 275452
rect 113605 275418 113639 275452
rect 113673 275418 113707 275452
rect 113741 275418 113775 275452
rect 113809 275418 113843 275452
rect 113877 275418 113911 275452
rect 113945 275418 113979 275452
rect 114013 275418 114047 275452
rect 111547 275256 111581 275290
rect 111615 275256 111649 275290
rect 111683 275256 111717 275290
rect 111751 275256 111785 275290
rect 111819 275256 111853 275290
rect 111887 275256 111921 275290
rect 111955 275256 111989 275290
rect 112023 275256 112057 275290
rect 112091 275256 112125 275290
rect 112159 275256 112193 275290
rect 112227 275256 112261 275290
rect 112295 275256 112329 275290
rect 112363 275256 112397 275290
rect 112431 275256 112465 275290
rect 112499 275256 112533 275290
rect 112567 275256 112601 275290
rect 112993 275160 113027 275194
rect 113061 275160 113095 275194
rect 113129 275160 113163 275194
rect 113197 275160 113231 275194
rect 113265 275160 113299 275194
rect 113333 275160 113367 275194
rect 113401 275160 113435 275194
rect 113469 275160 113503 275194
rect 113537 275160 113571 275194
rect 113605 275160 113639 275194
rect 113673 275160 113707 275194
rect 113741 275160 113775 275194
rect 113809 275160 113843 275194
rect 113877 275160 113911 275194
rect 113945 275160 113979 275194
rect 114013 275160 114047 275194
rect 111547 275114 111581 275148
rect 111615 275114 111649 275148
rect 111683 275114 111717 275148
rect 111751 275114 111785 275148
rect 111819 275114 111853 275148
rect 111887 275114 111921 275148
rect 111955 275114 111989 275148
rect 112023 275114 112057 275148
rect 112091 275114 112125 275148
rect 112159 275114 112193 275148
rect 112227 275114 112261 275148
rect 112295 275114 112329 275148
rect 112363 275114 112397 275148
rect 112431 275114 112465 275148
rect 112499 275114 112533 275148
rect 112567 275114 112601 275148
rect 113023 275016 113057 275050
rect 113091 275016 113125 275050
rect 113159 275016 113193 275050
rect 113227 275016 113261 275050
rect 113295 275016 113329 275050
rect 113363 275016 113397 275050
rect 113431 275016 113465 275050
rect 113499 275016 113533 275050
rect 113567 275016 113601 275050
rect 113635 275016 113669 275050
rect 113703 275016 113737 275050
rect 113771 275016 113805 275050
rect 113839 275016 113873 275050
rect 113907 275016 113941 275050
rect 113975 275016 114009 275050
rect 114043 275016 114077 275050
rect 111547 274896 111581 274930
rect 111615 274896 111649 274930
rect 111683 274896 111717 274930
rect 111751 274896 111785 274930
rect 111819 274896 111853 274930
rect 111887 274896 111921 274930
rect 111955 274896 111989 274930
rect 112023 274896 112057 274930
rect 112091 274896 112125 274930
rect 112159 274896 112193 274930
rect 112227 274896 112261 274930
rect 112295 274896 112329 274930
rect 112363 274896 112397 274930
rect 112431 274896 112465 274930
rect 112499 274896 112533 274930
rect 112567 274896 112601 274930
rect 113023 274878 113057 274912
rect 113091 274878 113125 274912
rect 113159 274878 113193 274912
rect 113227 274878 113261 274912
rect 113295 274878 113329 274912
rect 113363 274878 113397 274912
rect 113431 274878 113465 274912
rect 113499 274878 113533 274912
rect 113567 274878 113601 274912
rect 113635 274878 113669 274912
rect 113703 274878 113737 274912
rect 113771 274878 113805 274912
rect 113839 274878 113873 274912
rect 113907 274878 113941 274912
rect 113975 274878 114009 274912
rect 114043 274878 114077 274912
rect 111547 274754 111581 274788
rect 111615 274754 111649 274788
rect 111683 274754 111717 274788
rect 111751 274754 111785 274788
rect 111819 274754 111853 274788
rect 111887 274754 111921 274788
rect 111955 274754 111989 274788
rect 112023 274754 112057 274788
rect 112091 274754 112125 274788
rect 112159 274754 112193 274788
rect 112227 274754 112261 274788
rect 112295 274754 112329 274788
rect 112363 274754 112397 274788
rect 112431 274754 112465 274788
rect 112499 274754 112533 274788
rect 112567 274754 112601 274788
rect 113023 274718 113057 274752
rect 113091 274718 113125 274752
rect 113159 274718 113193 274752
rect 113227 274718 113261 274752
rect 113295 274718 113329 274752
rect 113363 274718 113397 274752
rect 113431 274718 113465 274752
rect 113499 274718 113533 274752
rect 113567 274718 113601 274752
rect 113635 274718 113669 274752
rect 113703 274718 113737 274752
rect 113771 274718 113805 274752
rect 113839 274718 113873 274752
rect 113907 274718 113941 274752
rect 113975 274718 114009 274752
rect 114043 274718 114077 274752
rect 111547 274536 111581 274570
rect 111615 274536 111649 274570
rect 111683 274536 111717 274570
rect 111751 274536 111785 274570
rect 111819 274536 111853 274570
rect 111887 274536 111921 274570
rect 111955 274536 111989 274570
rect 112023 274536 112057 274570
rect 112091 274536 112125 274570
rect 112159 274536 112193 274570
rect 112227 274536 112261 274570
rect 112295 274536 112329 274570
rect 112363 274536 112397 274570
rect 112431 274536 112465 274570
rect 112499 274536 112533 274570
rect 112567 274536 112601 274570
rect 113023 274580 113057 274614
rect 113091 274580 113125 274614
rect 113159 274580 113193 274614
rect 113227 274580 113261 274614
rect 113295 274580 113329 274614
rect 113363 274580 113397 274614
rect 113431 274580 113465 274614
rect 113499 274580 113533 274614
rect 113567 274580 113601 274614
rect 113635 274580 113669 274614
rect 113703 274580 113737 274614
rect 113771 274580 113805 274614
rect 113839 274580 113873 274614
rect 113907 274580 113941 274614
rect 113975 274580 114009 274614
rect 114043 274580 114077 274614
rect 116158 275842 116192 275876
rect 116226 275842 116260 275876
rect 116294 275842 116328 275876
rect 116362 275842 116396 275876
rect 116430 275842 116464 275876
rect 116498 275842 116532 275876
rect 116566 275842 116600 275876
rect 116634 275842 116668 275876
rect 116702 275842 116736 275876
rect 116770 275842 116804 275876
rect 116838 275842 116872 275876
rect 116906 275842 116940 275876
rect 116974 275842 117008 275876
rect 117042 275842 117076 275876
rect 117110 275842 117144 275876
rect 117178 275842 117212 275876
rect 117604 275834 117638 275868
rect 117672 275834 117706 275868
rect 117740 275834 117774 275868
rect 117808 275834 117842 275868
rect 117876 275834 117910 275868
rect 117944 275834 117978 275868
rect 118012 275834 118046 275868
rect 118080 275834 118114 275868
rect 118148 275834 118182 275868
rect 118216 275834 118250 275868
rect 118284 275834 118318 275868
rect 118352 275834 118386 275868
rect 118420 275834 118454 275868
rect 118488 275834 118522 275868
rect 118556 275834 118590 275868
rect 118624 275834 118658 275868
rect 116158 275584 116192 275618
rect 116226 275584 116260 275618
rect 116294 275584 116328 275618
rect 116362 275584 116396 275618
rect 116430 275584 116464 275618
rect 116498 275584 116532 275618
rect 116566 275584 116600 275618
rect 116634 275584 116668 275618
rect 116702 275584 116736 275618
rect 116770 275584 116804 275618
rect 116838 275584 116872 275618
rect 116906 275584 116940 275618
rect 116974 275584 117008 275618
rect 117042 275584 117076 275618
rect 117110 275584 117144 275618
rect 117178 275584 117212 275618
rect 117604 275616 117638 275650
rect 117672 275616 117706 275650
rect 117740 275616 117774 275650
rect 117808 275616 117842 275650
rect 117876 275616 117910 275650
rect 117944 275616 117978 275650
rect 118012 275616 118046 275650
rect 118080 275616 118114 275650
rect 118148 275616 118182 275650
rect 118216 275616 118250 275650
rect 118284 275616 118318 275650
rect 118352 275616 118386 275650
rect 118420 275616 118454 275650
rect 118488 275616 118522 275650
rect 118556 275616 118590 275650
rect 118624 275616 118658 275650
rect 117604 275474 117638 275508
rect 117672 275474 117706 275508
rect 117740 275474 117774 275508
rect 117808 275474 117842 275508
rect 117876 275474 117910 275508
rect 117944 275474 117978 275508
rect 118012 275474 118046 275508
rect 118080 275474 118114 275508
rect 118148 275474 118182 275508
rect 118216 275474 118250 275508
rect 118284 275474 118318 275508
rect 118352 275474 118386 275508
rect 118420 275474 118454 275508
rect 118488 275474 118522 275508
rect 118556 275474 118590 275508
rect 118624 275474 118658 275508
rect 116158 275418 116192 275452
rect 116226 275418 116260 275452
rect 116294 275418 116328 275452
rect 116362 275418 116396 275452
rect 116430 275418 116464 275452
rect 116498 275418 116532 275452
rect 116566 275418 116600 275452
rect 116634 275418 116668 275452
rect 116702 275418 116736 275452
rect 116770 275418 116804 275452
rect 116838 275418 116872 275452
rect 116906 275418 116940 275452
rect 116974 275418 117008 275452
rect 117042 275418 117076 275452
rect 117110 275418 117144 275452
rect 117178 275418 117212 275452
rect 117604 275256 117638 275290
rect 117672 275256 117706 275290
rect 117740 275256 117774 275290
rect 117808 275256 117842 275290
rect 117876 275256 117910 275290
rect 117944 275256 117978 275290
rect 118012 275256 118046 275290
rect 118080 275256 118114 275290
rect 118148 275256 118182 275290
rect 118216 275256 118250 275290
rect 118284 275256 118318 275290
rect 118352 275256 118386 275290
rect 118420 275256 118454 275290
rect 118488 275256 118522 275290
rect 118556 275256 118590 275290
rect 118624 275256 118658 275290
rect 116158 275160 116192 275194
rect 116226 275160 116260 275194
rect 116294 275160 116328 275194
rect 116362 275160 116396 275194
rect 116430 275160 116464 275194
rect 116498 275160 116532 275194
rect 116566 275160 116600 275194
rect 116634 275160 116668 275194
rect 116702 275160 116736 275194
rect 116770 275160 116804 275194
rect 116838 275160 116872 275194
rect 116906 275160 116940 275194
rect 116974 275160 117008 275194
rect 117042 275160 117076 275194
rect 117110 275160 117144 275194
rect 117178 275160 117212 275194
rect 117604 275114 117638 275148
rect 117672 275114 117706 275148
rect 117740 275114 117774 275148
rect 117808 275114 117842 275148
rect 117876 275114 117910 275148
rect 117944 275114 117978 275148
rect 118012 275114 118046 275148
rect 118080 275114 118114 275148
rect 118148 275114 118182 275148
rect 118216 275114 118250 275148
rect 118284 275114 118318 275148
rect 118352 275114 118386 275148
rect 118420 275114 118454 275148
rect 118488 275114 118522 275148
rect 118556 275114 118590 275148
rect 118624 275114 118658 275148
rect 116128 275016 116162 275050
rect 116196 275016 116230 275050
rect 116264 275016 116298 275050
rect 116332 275016 116366 275050
rect 116400 275016 116434 275050
rect 116468 275016 116502 275050
rect 116536 275016 116570 275050
rect 116604 275016 116638 275050
rect 116672 275016 116706 275050
rect 116740 275016 116774 275050
rect 116808 275016 116842 275050
rect 116876 275016 116910 275050
rect 116944 275016 116978 275050
rect 117012 275016 117046 275050
rect 117080 275016 117114 275050
rect 117148 275016 117182 275050
rect 116128 274878 116162 274912
rect 116196 274878 116230 274912
rect 116264 274878 116298 274912
rect 116332 274878 116366 274912
rect 116400 274878 116434 274912
rect 116468 274878 116502 274912
rect 116536 274878 116570 274912
rect 116604 274878 116638 274912
rect 116672 274878 116706 274912
rect 116740 274878 116774 274912
rect 116808 274878 116842 274912
rect 116876 274878 116910 274912
rect 116944 274878 116978 274912
rect 117012 274878 117046 274912
rect 117080 274878 117114 274912
rect 117148 274878 117182 274912
rect 117604 274896 117638 274930
rect 117672 274896 117706 274930
rect 117740 274896 117774 274930
rect 117808 274896 117842 274930
rect 117876 274896 117910 274930
rect 117944 274896 117978 274930
rect 118012 274896 118046 274930
rect 118080 274896 118114 274930
rect 118148 274896 118182 274930
rect 118216 274896 118250 274930
rect 118284 274896 118318 274930
rect 118352 274896 118386 274930
rect 118420 274896 118454 274930
rect 118488 274896 118522 274930
rect 118556 274896 118590 274930
rect 118624 274896 118658 274930
rect 116128 274718 116162 274752
rect 116196 274718 116230 274752
rect 116264 274718 116298 274752
rect 116332 274718 116366 274752
rect 116400 274718 116434 274752
rect 116468 274718 116502 274752
rect 116536 274718 116570 274752
rect 116604 274718 116638 274752
rect 116672 274718 116706 274752
rect 116740 274718 116774 274752
rect 116808 274718 116842 274752
rect 116876 274718 116910 274752
rect 116944 274718 116978 274752
rect 117012 274718 117046 274752
rect 117080 274718 117114 274752
rect 117148 274718 117182 274752
rect 117604 274754 117638 274788
rect 117672 274754 117706 274788
rect 117740 274754 117774 274788
rect 117808 274754 117842 274788
rect 117876 274754 117910 274788
rect 117944 274754 117978 274788
rect 118012 274754 118046 274788
rect 118080 274754 118114 274788
rect 118148 274754 118182 274788
rect 118216 274754 118250 274788
rect 118284 274754 118318 274788
rect 118352 274754 118386 274788
rect 118420 274754 118454 274788
rect 118488 274754 118522 274788
rect 118556 274754 118590 274788
rect 118624 274754 118658 274788
rect 116128 274580 116162 274614
rect 116196 274580 116230 274614
rect 116264 274580 116298 274614
rect 116332 274580 116366 274614
rect 116400 274580 116434 274614
rect 116468 274580 116502 274614
rect 116536 274580 116570 274614
rect 116604 274580 116638 274614
rect 116672 274580 116706 274614
rect 116740 274580 116774 274614
rect 116808 274580 116842 274614
rect 116876 274580 116910 274614
rect 116944 274580 116978 274614
rect 117012 274580 117046 274614
rect 117080 274580 117114 274614
rect 117148 274580 117182 274614
rect 117604 274536 117638 274570
rect 117672 274536 117706 274570
rect 117740 274536 117774 274570
rect 117808 274536 117842 274570
rect 117876 274536 117910 274570
rect 117944 274536 117978 274570
rect 118012 274536 118046 274570
rect 118080 274536 118114 274570
rect 118148 274536 118182 274570
rect 118216 274536 118250 274570
rect 118284 274536 118318 274570
rect 118352 274536 118386 274570
rect 118420 274536 118454 274570
rect 118488 274536 118522 274570
rect 118556 274536 118590 274570
rect 118624 274536 118658 274570
rect 111547 274168 111581 274202
rect 111615 274168 111649 274202
rect 111683 274168 111717 274202
rect 111751 274168 111785 274202
rect 111819 274168 111853 274202
rect 111887 274168 111921 274202
rect 111955 274168 111989 274202
rect 112023 274168 112057 274202
rect 112091 274168 112125 274202
rect 112159 274168 112193 274202
rect 112227 274168 112261 274202
rect 112295 274168 112329 274202
rect 112363 274168 112397 274202
rect 112431 274168 112465 274202
rect 112499 274168 112533 274202
rect 112567 274168 112601 274202
rect 112993 274176 113027 274210
rect 113061 274176 113095 274210
rect 113129 274176 113163 274210
rect 113197 274176 113231 274210
rect 113265 274176 113299 274210
rect 113333 274176 113367 274210
rect 113401 274176 113435 274210
rect 113469 274176 113503 274210
rect 113537 274176 113571 274210
rect 113605 274176 113639 274210
rect 113673 274176 113707 274210
rect 113741 274176 113775 274210
rect 113809 274176 113843 274210
rect 113877 274176 113911 274210
rect 113945 274176 113979 274210
rect 114013 274176 114047 274210
rect 111547 273950 111581 273984
rect 111615 273950 111649 273984
rect 111683 273950 111717 273984
rect 111751 273950 111785 273984
rect 111819 273950 111853 273984
rect 111887 273950 111921 273984
rect 111955 273950 111989 273984
rect 112023 273950 112057 273984
rect 112091 273950 112125 273984
rect 112159 273950 112193 273984
rect 112227 273950 112261 273984
rect 112295 273950 112329 273984
rect 112363 273950 112397 273984
rect 112431 273950 112465 273984
rect 112499 273950 112533 273984
rect 112567 273950 112601 273984
rect 112993 273918 113027 273952
rect 113061 273918 113095 273952
rect 113129 273918 113163 273952
rect 113197 273918 113231 273952
rect 113265 273918 113299 273952
rect 113333 273918 113367 273952
rect 113401 273918 113435 273952
rect 113469 273918 113503 273952
rect 113537 273918 113571 273952
rect 113605 273918 113639 273952
rect 113673 273918 113707 273952
rect 113741 273918 113775 273952
rect 113809 273918 113843 273952
rect 113877 273918 113911 273952
rect 113945 273918 113979 273952
rect 114013 273918 114047 273952
rect 111547 273808 111581 273842
rect 111615 273808 111649 273842
rect 111683 273808 111717 273842
rect 111751 273808 111785 273842
rect 111819 273808 111853 273842
rect 111887 273808 111921 273842
rect 111955 273808 111989 273842
rect 112023 273808 112057 273842
rect 112091 273808 112125 273842
rect 112159 273808 112193 273842
rect 112227 273808 112261 273842
rect 112295 273808 112329 273842
rect 112363 273808 112397 273842
rect 112431 273808 112465 273842
rect 112499 273808 112533 273842
rect 112567 273808 112601 273842
rect 112993 273752 113027 273786
rect 113061 273752 113095 273786
rect 113129 273752 113163 273786
rect 113197 273752 113231 273786
rect 113265 273752 113299 273786
rect 113333 273752 113367 273786
rect 113401 273752 113435 273786
rect 113469 273752 113503 273786
rect 113537 273752 113571 273786
rect 113605 273752 113639 273786
rect 113673 273752 113707 273786
rect 113741 273752 113775 273786
rect 113809 273752 113843 273786
rect 113877 273752 113911 273786
rect 113945 273752 113979 273786
rect 114013 273752 114047 273786
rect 111547 273590 111581 273624
rect 111615 273590 111649 273624
rect 111683 273590 111717 273624
rect 111751 273590 111785 273624
rect 111819 273590 111853 273624
rect 111887 273590 111921 273624
rect 111955 273590 111989 273624
rect 112023 273590 112057 273624
rect 112091 273590 112125 273624
rect 112159 273590 112193 273624
rect 112227 273590 112261 273624
rect 112295 273590 112329 273624
rect 112363 273590 112397 273624
rect 112431 273590 112465 273624
rect 112499 273590 112533 273624
rect 112567 273590 112601 273624
rect 112993 273494 113027 273528
rect 113061 273494 113095 273528
rect 113129 273494 113163 273528
rect 113197 273494 113231 273528
rect 113265 273494 113299 273528
rect 113333 273494 113367 273528
rect 113401 273494 113435 273528
rect 113469 273494 113503 273528
rect 113537 273494 113571 273528
rect 113605 273494 113639 273528
rect 113673 273494 113707 273528
rect 113741 273494 113775 273528
rect 113809 273494 113843 273528
rect 113877 273494 113911 273528
rect 113945 273494 113979 273528
rect 114013 273494 114047 273528
rect 111547 273448 111581 273482
rect 111615 273448 111649 273482
rect 111683 273448 111717 273482
rect 111751 273448 111785 273482
rect 111819 273448 111853 273482
rect 111887 273448 111921 273482
rect 111955 273448 111989 273482
rect 112023 273448 112057 273482
rect 112091 273448 112125 273482
rect 112159 273448 112193 273482
rect 112227 273448 112261 273482
rect 112295 273448 112329 273482
rect 112363 273448 112397 273482
rect 112431 273448 112465 273482
rect 112499 273448 112533 273482
rect 112567 273448 112601 273482
rect 113023 273350 113057 273384
rect 113091 273350 113125 273384
rect 113159 273350 113193 273384
rect 113227 273350 113261 273384
rect 113295 273350 113329 273384
rect 113363 273350 113397 273384
rect 113431 273350 113465 273384
rect 113499 273350 113533 273384
rect 113567 273350 113601 273384
rect 113635 273350 113669 273384
rect 113703 273350 113737 273384
rect 113771 273350 113805 273384
rect 113839 273350 113873 273384
rect 113907 273350 113941 273384
rect 113975 273350 114009 273384
rect 114043 273350 114077 273384
rect 111547 273230 111581 273264
rect 111615 273230 111649 273264
rect 111683 273230 111717 273264
rect 111751 273230 111785 273264
rect 111819 273230 111853 273264
rect 111887 273230 111921 273264
rect 111955 273230 111989 273264
rect 112023 273230 112057 273264
rect 112091 273230 112125 273264
rect 112159 273230 112193 273264
rect 112227 273230 112261 273264
rect 112295 273230 112329 273264
rect 112363 273230 112397 273264
rect 112431 273230 112465 273264
rect 112499 273230 112533 273264
rect 112567 273230 112601 273264
rect 113023 273212 113057 273246
rect 113091 273212 113125 273246
rect 113159 273212 113193 273246
rect 113227 273212 113261 273246
rect 113295 273212 113329 273246
rect 113363 273212 113397 273246
rect 113431 273212 113465 273246
rect 113499 273212 113533 273246
rect 113567 273212 113601 273246
rect 113635 273212 113669 273246
rect 113703 273212 113737 273246
rect 113771 273212 113805 273246
rect 113839 273212 113873 273246
rect 113907 273212 113941 273246
rect 113975 273212 114009 273246
rect 114043 273212 114077 273246
rect 111547 273088 111581 273122
rect 111615 273088 111649 273122
rect 111683 273088 111717 273122
rect 111751 273088 111785 273122
rect 111819 273088 111853 273122
rect 111887 273088 111921 273122
rect 111955 273088 111989 273122
rect 112023 273088 112057 273122
rect 112091 273088 112125 273122
rect 112159 273088 112193 273122
rect 112227 273088 112261 273122
rect 112295 273088 112329 273122
rect 112363 273088 112397 273122
rect 112431 273088 112465 273122
rect 112499 273088 112533 273122
rect 112567 273088 112601 273122
rect 113023 273052 113057 273086
rect 113091 273052 113125 273086
rect 113159 273052 113193 273086
rect 113227 273052 113261 273086
rect 113295 273052 113329 273086
rect 113363 273052 113397 273086
rect 113431 273052 113465 273086
rect 113499 273052 113533 273086
rect 113567 273052 113601 273086
rect 113635 273052 113669 273086
rect 113703 273052 113737 273086
rect 113771 273052 113805 273086
rect 113839 273052 113873 273086
rect 113907 273052 113941 273086
rect 113975 273052 114009 273086
rect 114043 273052 114077 273086
rect 111547 272870 111581 272904
rect 111615 272870 111649 272904
rect 111683 272870 111717 272904
rect 111751 272870 111785 272904
rect 111819 272870 111853 272904
rect 111887 272870 111921 272904
rect 111955 272870 111989 272904
rect 112023 272870 112057 272904
rect 112091 272870 112125 272904
rect 112159 272870 112193 272904
rect 112227 272870 112261 272904
rect 112295 272870 112329 272904
rect 112363 272870 112397 272904
rect 112431 272870 112465 272904
rect 112499 272870 112533 272904
rect 112567 272870 112601 272904
rect 113023 272914 113057 272948
rect 113091 272914 113125 272948
rect 113159 272914 113193 272948
rect 113227 272914 113261 272948
rect 113295 272914 113329 272948
rect 113363 272914 113397 272948
rect 113431 272914 113465 272948
rect 113499 272914 113533 272948
rect 113567 272914 113601 272948
rect 113635 272914 113669 272948
rect 113703 272914 113737 272948
rect 113771 272914 113805 272948
rect 113839 272914 113873 272948
rect 113907 272914 113941 272948
rect 113975 272914 114009 272948
rect 114043 272914 114077 272948
rect 116158 274176 116192 274210
rect 116226 274176 116260 274210
rect 116294 274176 116328 274210
rect 116362 274176 116396 274210
rect 116430 274176 116464 274210
rect 116498 274176 116532 274210
rect 116566 274176 116600 274210
rect 116634 274176 116668 274210
rect 116702 274176 116736 274210
rect 116770 274176 116804 274210
rect 116838 274176 116872 274210
rect 116906 274176 116940 274210
rect 116974 274176 117008 274210
rect 117042 274176 117076 274210
rect 117110 274176 117144 274210
rect 117178 274176 117212 274210
rect 117604 274168 117638 274202
rect 117672 274168 117706 274202
rect 117740 274168 117774 274202
rect 117808 274168 117842 274202
rect 117876 274168 117910 274202
rect 117944 274168 117978 274202
rect 118012 274168 118046 274202
rect 118080 274168 118114 274202
rect 118148 274168 118182 274202
rect 118216 274168 118250 274202
rect 118284 274168 118318 274202
rect 118352 274168 118386 274202
rect 118420 274168 118454 274202
rect 118488 274168 118522 274202
rect 118556 274168 118590 274202
rect 118624 274168 118658 274202
rect 116158 273918 116192 273952
rect 116226 273918 116260 273952
rect 116294 273918 116328 273952
rect 116362 273918 116396 273952
rect 116430 273918 116464 273952
rect 116498 273918 116532 273952
rect 116566 273918 116600 273952
rect 116634 273918 116668 273952
rect 116702 273918 116736 273952
rect 116770 273918 116804 273952
rect 116838 273918 116872 273952
rect 116906 273918 116940 273952
rect 116974 273918 117008 273952
rect 117042 273918 117076 273952
rect 117110 273918 117144 273952
rect 117178 273918 117212 273952
rect 117604 273950 117638 273984
rect 117672 273950 117706 273984
rect 117740 273950 117774 273984
rect 117808 273950 117842 273984
rect 117876 273950 117910 273984
rect 117944 273950 117978 273984
rect 118012 273950 118046 273984
rect 118080 273950 118114 273984
rect 118148 273950 118182 273984
rect 118216 273950 118250 273984
rect 118284 273950 118318 273984
rect 118352 273950 118386 273984
rect 118420 273950 118454 273984
rect 118488 273950 118522 273984
rect 118556 273950 118590 273984
rect 118624 273950 118658 273984
rect 117604 273808 117638 273842
rect 117672 273808 117706 273842
rect 117740 273808 117774 273842
rect 117808 273808 117842 273842
rect 117876 273808 117910 273842
rect 117944 273808 117978 273842
rect 118012 273808 118046 273842
rect 118080 273808 118114 273842
rect 118148 273808 118182 273842
rect 118216 273808 118250 273842
rect 118284 273808 118318 273842
rect 118352 273808 118386 273842
rect 118420 273808 118454 273842
rect 118488 273808 118522 273842
rect 118556 273808 118590 273842
rect 118624 273808 118658 273842
rect 116158 273752 116192 273786
rect 116226 273752 116260 273786
rect 116294 273752 116328 273786
rect 116362 273752 116396 273786
rect 116430 273752 116464 273786
rect 116498 273752 116532 273786
rect 116566 273752 116600 273786
rect 116634 273752 116668 273786
rect 116702 273752 116736 273786
rect 116770 273752 116804 273786
rect 116838 273752 116872 273786
rect 116906 273752 116940 273786
rect 116974 273752 117008 273786
rect 117042 273752 117076 273786
rect 117110 273752 117144 273786
rect 117178 273752 117212 273786
rect 117604 273590 117638 273624
rect 117672 273590 117706 273624
rect 117740 273590 117774 273624
rect 117808 273590 117842 273624
rect 117876 273590 117910 273624
rect 117944 273590 117978 273624
rect 118012 273590 118046 273624
rect 118080 273590 118114 273624
rect 118148 273590 118182 273624
rect 118216 273590 118250 273624
rect 118284 273590 118318 273624
rect 118352 273590 118386 273624
rect 118420 273590 118454 273624
rect 118488 273590 118522 273624
rect 118556 273590 118590 273624
rect 118624 273590 118658 273624
rect 116158 273494 116192 273528
rect 116226 273494 116260 273528
rect 116294 273494 116328 273528
rect 116362 273494 116396 273528
rect 116430 273494 116464 273528
rect 116498 273494 116532 273528
rect 116566 273494 116600 273528
rect 116634 273494 116668 273528
rect 116702 273494 116736 273528
rect 116770 273494 116804 273528
rect 116838 273494 116872 273528
rect 116906 273494 116940 273528
rect 116974 273494 117008 273528
rect 117042 273494 117076 273528
rect 117110 273494 117144 273528
rect 117178 273494 117212 273528
rect 117604 273448 117638 273482
rect 117672 273448 117706 273482
rect 117740 273448 117774 273482
rect 117808 273448 117842 273482
rect 117876 273448 117910 273482
rect 117944 273448 117978 273482
rect 118012 273448 118046 273482
rect 118080 273448 118114 273482
rect 118148 273448 118182 273482
rect 118216 273448 118250 273482
rect 118284 273448 118318 273482
rect 118352 273448 118386 273482
rect 118420 273448 118454 273482
rect 118488 273448 118522 273482
rect 118556 273448 118590 273482
rect 118624 273448 118658 273482
rect 116128 273350 116162 273384
rect 116196 273350 116230 273384
rect 116264 273350 116298 273384
rect 116332 273350 116366 273384
rect 116400 273350 116434 273384
rect 116468 273350 116502 273384
rect 116536 273350 116570 273384
rect 116604 273350 116638 273384
rect 116672 273350 116706 273384
rect 116740 273350 116774 273384
rect 116808 273350 116842 273384
rect 116876 273350 116910 273384
rect 116944 273350 116978 273384
rect 117012 273350 117046 273384
rect 117080 273350 117114 273384
rect 117148 273350 117182 273384
rect 116128 273212 116162 273246
rect 116196 273212 116230 273246
rect 116264 273212 116298 273246
rect 116332 273212 116366 273246
rect 116400 273212 116434 273246
rect 116468 273212 116502 273246
rect 116536 273212 116570 273246
rect 116604 273212 116638 273246
rect 116672 273212 116706 273246
rect 116740 273212 116774 273246
rect 116808 273212 116842 273246
rect 116876 273212 116910 273246
rect 116944 273212 116978 273246
rect 117012 273212 117046 273246
rect 117080 273212 117114 273246
rect 117148 273212 117182 273246
rect 117604 273230 117638 273264
rect 117672 273230 117706 273264
rect 117740 273230 117774 273264
rect 117808 273230 117842 273264
rect 117876 273230 117910 273264
rect 117944 273230 117978 273264
rect 118012 273230 118046 273264
rect 118080 273230 118114 273264
rect 118148 273230 118182 273264
rect 118216 273230 118250 273264
rect 118284 273230 118318 273264
rect 118352 273230 118386 273264
rect 118420 273230 118454 273264
rect 118488 273230 118522 273264
rect 118556 273230 118590 273264
rect 118624 273230 118658 273264
rect 116128 273052 116162 273086
rect 116196 273052 116230 273086
rect 116264 273052 116298 273086
rect 116332 273052 116366 273086
rect 116400 273052 116434 273086
rect 116468 273052 116502 273086
rect 116536 273052 116570 273086
rect 116604 273052 116638 273086
rect 116672 273052 116706 273086
rect 116740 273052 116774 273086
rect 116808 273052 116842 273086
rect 116876 273052 116910 273086
rect 116944 273052 116978 273086
rect 117012 273052 117046 273086
rect 117080 273052 117114 273086
rect 117148 273052 117182 273086
rect 117604 273088 117638 273122
rect 117672 273088 117706 273122
rect 117740 273088 117774 273122
rect 117808 273088 117842 273122
rect 117876 273088 117910 273122
rect 117944 273088 117978 273122
rect 118012 273088 118046 273122
rect 118080 273088 118114 273122
rect 118148 273088 118182 273122
rect 118216 273088 118250 273122
rect 118284 273088 118318 273122
rect 118352 273088 118386 273122
rect 118420 273088 118454 273122
rect 118488 273088 118522 273122
rect 118556 273088 118590 273122
rect 118624 273088 118658 273122
rect 116128 272914 116162 272948
rect 116196 272914 116230 272948
rect 116264 272914 116298 272948
rect 116332 272914 116366 272948
rect 116400 272914 116434 272948
rect 116468 272914 116502 272948
rect 116536 272914 116570 272948
rect 116604 272914 116638 272948
rect 116672 272914 116706 272948
rect 116740 272914 116774 272948
rect 116808 272914 116842 272948
rect 116876 272914 116910 272948
rect 116944 272914 116978 272948
rect 117012 272914 117046 272948
rect 117080 272914 117114 272948
rect 117148 272914 117182 272948
rect 117604 272870 117638 272904
rect 117672 272870 117706 272904
rect 117740 272870 117774 272904
rect 117808 272870 117842 272904
rect 117876 272870 117910 272904
rect 117944 272870 117978 272904
rect 118012 272870 118046 272904
rect 118080 272870 118114 272904
rect 118148 272870 118182 272904
rect 118216 272870 118250 272904
rect 118284 272870 118318 272904
rect 118352 272870 118386 272904
rect 118420 272870 118454 272904
rect 118488 272870 118522 272904
rect 118556 272870 118590 272904
rect 118624 272870 118658 272904
rect 115835 271867 115869 271901
rect 115835 271799 115869 271833
rect 115835 271731 115869 271765
rect 115835 271663 115869 271697
rect 115835 271595 115869 271629
rect 115835 271527 115869 271561
rect 115835 271459 115869 271493
rect 115835 271391 115869 271425
rect 115835 271323 115869 271357
rect 115835 271255 115869 271289
rect 115835 271187 115869 271221
rect 115835 271119 115869 271153
rect 115835 271051 115869 271085
rect 115835 270983 115869 271017
rect 115835 270915 115869 270949
rect 115835 270847 115869 270881
rect 116053 271867 116087 271901
rect 116053 271799 116087 271833
rect 116053 271731 116087 271765
rect 116053 271663 116087 271697
rect 116053 271595 116087 271629
rect 116053 271527 116087 271561
rect 116053 271459 116087 271493
rect 116053 271391 116087 271425
rect 116053 271323 116087 271357
rect 116053 271255 116087 271289
rect 116053 271187 116087 271221
rect 116053 271119 116087 271153
rect 116053 271051 116087 271085
rect 116053 270983 116087 271017
rect 116053 270915 116087 270949
rect 116053 270847 116087 270881
rect 116235 271867 116269 271901
rect 116235 271799 116269 271833
rect 116235 271731 116269 271765
rect 116235 271663 116269 271697
rect 116235 271595 116269 271629
rect 116235 271527 116269 271561
rect 116235 271459 116269 271493
rect 116235 271391 116269 271425
rect 116235 271323 116269 271357
rect 116235 271255 116269 271289
rect 116235 271187 116269 271221
rect 116235 271119 116269 271153
rect 116235 271051 116269 271085
rect 116235 270983 116269 271017
rect 116235 270915 116269 270949
rect 116235 270847 116269 270881
rect 116453 271867 116487 271901
rect 116453 271799 116487 271833
rect 116453 271731 116487 271765
rect 116453 271663 116487 271697
rect 116453 271595 116487 271629
rect 116453 271527 116487 271561
rect 116453 271459 116487 271493
rect 116453 271391 116487 271425
rect 116453 271323 116487 271357
rect 116453 271255 116487 271289
rect 116453 271187 116487 271221
rect 116453 271119 116487 271153
rect 116453 271051 116487 271085
rect 116453 270983 116487 271017
rect 116453 270915 116487 270949
rect 116453 270847 116487 270881
rect 116635 271867 116669 271901
rect 116635 271799 116669 271833
rect 116635 271731 116669 271765
rect 116635 271663 116669 271697
rect 116635 271595 116669 271629
rect 116635 271527 116669 271561
rect 116635 271459 116669 271493
rect 116635 271391 116669 271425
rect 116635 271323 116669 271357
rect 116635 271255 116669 271289
rect 116635 271187 116669 271221
rect 116635 271119 116669 271153
rect 116635 271051 116669 271085
rect 116635 270983 116669 271017
rect 116635 270915 116669 270949
rect 116635 270847 116669 270881
rect 116853 271867 116887 271901
rect 116853 271799 116887 271833
rect 116853 271731 116887 271765
rect 116853 271663 116887 271697
rect 116853 271595 116887 271629
rect 116853 271527 116887 271561
rect 116853 271459 116887 271493
rect 116853 271391 116887 271425
rect 116853 271323 116887 271357
rect 116853 271255 116887 271289
rect 116853 271187 116887 271221
rect 116853 271119 116887 271153
rect 116853 271051 116887 271085
rect 116853 270983 116887 271017
rect 116853 270915 116887 270949
rect 116853 270847 116887 270881
rect 117035 271867 117069 271901
rect 117035 271799 117069 271833
rect 117035 271731 117069 271765
rect 117035 271663 117069 271697
rect 117035 271595 117069 271629
rect 117035 271527 117069 271561
rect 117035 271459 117069 271493
rect 117035 271391 117069 271425
rect 117035 271323 117069 271357
rect 117035 271255 117069 271289
rect 117035 271187 117069 271221
rect 117035 271119 117069 271153
rect 117035 271051 117069 271085
rect 117035 270983 117069 271017
rect 117035 270915 117069 270949
rect 117035 270847 117069 270881
rect 117253 271867 117287 271901
rect 117253 271799 117287 271833
rect 117253 271731 117287 271765
rect 117253 271663 117287 271697
rect 117253 271595 117287 271629
rect 117253 271527 117287 271561
rect 117253 271459 117287 271493
rect 117253 271391 117287 271425
rect 117253 271323 117287 271357
rect 117253 271255 117287 271289
rect 117253 271187 117287 271221
rect 117253 271119 117287 271153
rect 117253 271051 117287 271085
rect 117253 270983 117287 271017
rect 117253 270915 117287 270949
rect 117253 270847 117287 270881
rect 117435 271867 117469 271901
rect 117435 271799 117469 271833
rect 117435 271731 117469 271765
rect 117435 271663 117469 271697
rect 117435 271595 117469 271629
rect 117435 271527 117469 271561
rect 117435 271459 117469 271493
rect 117435 271391 117469 271425
rect 117435 271323 117469 271357
rect 117435 271255 117469 271289
rect 117435 271187 117469 271221
rect 117435 271119 117469 271153
rect 117435 271051 117469 271085
rect 117435 270983 117469 271017
rect 117435 270915 117469 270949
rect 117435 270847 117469 270881
rect 117653 271867 117687 271901
rect 117653 271799 117687 271833
rect 117653 271731 117687 271765
rect 117653 271663 117687 271697
rect 117653 271595 117687 271629
rect 117653 271527 117687 271561
rect 117653 271459 117687 271493
rect 117653 271391 117687 271425
rect 117653 271323 117687 271357
rect 117653 271255 117687 271289
rect 117653 271187 117687 271221
rect 117653 271119 117687 271153
rect 117653 271051 117687 271085
rect 117653 270983 117687 271017
rect 117653 270915 117687 270949
rect 117653 270847 117687 270881
rect 117835 271867 117869 271901
rect 117835 271799 117869 271833
rect 117835 271731 117869 271765
rect 117835 271663 117869 271697
rect 117835 271595 117869 271629
rect 117835 271527 117869 271561
rect 117835 271459 117869 271493
rect 117835 271391 117869 271425
rect 117835 271323 117869 271357
rect 117835 271255 117869 271289
rect 117835 271187 117869 271221
rect 117835 271119 117869 271153
rect 117835 271051 117869 271085
rect 117835 270983 117869 271017
rect 117835 270915 117869 270949
rect 117835 270847 117869 270881
rect 118053 271867 118087 271901
rect 118053 271799 118087 271833
rect 118053 271731 118087 271765
rect 118053 271663 118087 271697
rect 118053 271595 118087 271629
rect 118053 271527 118087 271561
rect 118053 271459 118087 271493
rect 118053 271391 118087 271425
rect 118053 271323 118087 271357
rect 118053 271255 118087 271289
rect 118053 271187 118087 271221
rect 118053 271119 118087 271153
rect 118053 271051 118087 271085
rect 118053 270983 118087 271017
rect 118053 270915 118087 270949
rect 118053 270847 118087 270881
rect 118235 271867 118269 271901
rect 118235 271799 118269 271833
rect 118235 271731 118269 271765
rect 118235 271663 118269 271697
rect 118235 271595 118269 271629
rect 118235 271527 118269 271561
rect 118235 271459 118269 271493
rect 118235 271391 118269 271425
rect 118235 271323 118269 271357
rect 118235 271255 118269 271289
rect 118235 271187 118269 271221
rect 118235 271119 118269 271153
rect 118235 271051 118269 271085
rect 118235 270983 118269 271017
rect 118235 270915 118269 270949
rect 118235 270847 118269 270881
rect 118453 271867 118487 271901
rect 118453 271799 118487 271833
rect 118453 271731 118487 271765
rect 118453 271663 118487 271697
rect 118453 271595 118487 271629
rect 118453 271527 118487 271561
rect 118453 271459 118487 271493
rect 118453 271391 118487 271425
rect 118453 271323 118487 271357
rect 118453 271255 118487 271289
rect 118453 271187 118487 271221
rect 118453 271119 118487 271153
rect 118453 271051 118487 271085
rect 118453 270983 118487 271017
rect 118453 270915 118487 270949
rect 118453 270847 118487 270881
rect 118635 271867 118669 271901
rect 118635 271799 118669 271833
rect 118635 271731 118669 271765
rect 118635 271663 118669 271697
rect 118635 271595 118669 271629
rect 118635 271527 118669 271561
rect 118635 271459 118669 271493
rect 118635 271391 118669 271425
rect 118635 271323 118669 271357
rect 118635 271255 118669 271289
rect 118635 271187 118669 271221
rect 118635 271119 118669 271153
rect 118635 271051 118669 271085
rect 118635 270983 118669 271017
rect 118635 270915 118669 270949
rect 118635 270847 118669 270881
rect 118853 271867 118887 271901
rect 118853 271799 118887 271833
rect 118853 271731 118887 271765
rect 118853 271663 118887 271697
rect 118853 271595 118887 271629
rect 118853 271527 118887 271561
rect 118853 271459 118887 271493
rect 118853 271391 118887 271425
rect 118853 271323 118887 271357
rect 118853 271255 118887 271289
rect 118853 271187 118887 271221
rect 118853 271119 118887 271153
rect 118853 271051 118887 271085
rect 118853 270983 118887 271017
rect 118853 270915 118887 270949
rect 118853 270847 118887 270881
rect 112514 270167 112548 270201
rect 112514 270099 112548 270133
rect 112514 270031 112548 270065
rect 112514 269963 112548 269997
rect 112514 269895 112548 269929
rect 112514 269827 112548 269861
rect 112514 269759 112548 269793
rect 112514 269691 112548 269725
rect 112514 269623 112548 269657
rect 112514 269555 112548 269589
rect 112514 269487 112548 269521
rect 112514 269419 112548 269453
rect 112514 269351 112548 269385
rect 112514 269283 112548 269317
rect 112514 269215 112548 269249
rect 112514 269147 112548 269181
rect 112732 270167 112766 270201
rect 112732 270099 112766 270133
rect 112732 270031 112766 270065
rect 112732 269963 112766 269997
rect 112732 269895 112766 269929
rect 112732 269827 112766 269861
rect 112732 269759 112766 269793
rect 112732 269691 112766 269725
rect 112732 269623 112766 269657
rect 112732 269555 112766 269589
rect 112732 269487 112766 269521
rect 112732 269419 112766 269453
rect 112732 269351 112766 269385
rect 112732 269283 112766 269317
rect 112732 269215 112766 269249
rect 112732 269147 112766 269181
rect 112914 270167 112948 270201
rect 112914 270099 112948 270133
rect 112914 270031 112948 270065
rect 112914 269963 112948 269997
rect 112914 269895 112948 269929
rect 112914 269827 112948 269861
rect 112914 269759 112948 269793
rect 112914 269691 112948 269725
rect 112914 269623 112948 269657
rect 112914 269555 112948 269589
rect 112914 269487 112948 269521
rect 112914 269419 112948 269453
rect 112914 269351 112948 269385
rect 112914 269283 112948 269317
rect 112914 269215 112948 269249
rect 112914 269147 112948 269181
rect 113132 270167 113166 270201
rect 113132 270099 113166 270133
rect 113132 270031 113166 270065
rect 113132 269963 113166 269997
rect 113132 269895 113166 269929
rect 113132 269827 113166 269861
rect 113132 269759 113166 269793
rect 113132 269691 113166 269725
rect 113132 269623 113166 269657
rect 113132 269555 113166 269589
rect 113132 269487 113166 269521
rect 113132 269419 113166 269453
rect 113132 269351 113166 269385
rect 113132 269283 113166 269317
rect 113132 269215 113166 269249
rect 113132 269147 113166 269181
rect 113314 270167 113348 270201
rect 113314 270099 113348 270133
rect 113314 270031 113348 270065
rect 113314 269963 113348 269997
rect 113314 269895 113348 269929
rect 113314 269827 113348 269861
rect 113314 269759 113348 269793
rect 113314 269691 113348 269725
rect 113314 269623 113348 269657
rect 113314 269555 113348 269589
rect 113314 269487 113348 269521
rect 113314 269419 113348 269453
rect 113314 269351 113348 269385
rect 113314 269283 113348 269317
rect 113314 269215 113348 269249
rect 113314 269147 113348 269181
rect 113532 270167 113566 270201
rect 113532 270099 113566 270133
rect 113532 270031 113566 270065
rect 113532 269963 113566 269997
rect 113532 269895 113566 269929
rect 113532 269827 113566 269861
rect 113532 269759 113566 269793
rect 113532 269691 113566 269725
rect 113532 269623 113566 269657
rect 113532 269555 113566 269589
rect 113532 269487 113566 269521
rect 113532 269419 113566 269453
rect 113532 269351 113566 269385
rect 113532 269283 113566 269317
rect 113532 269215 113566 269249
rect 113532 269147 113566 269181
rect 113714 270167 113748 270201
rect 113714 270099 113748 270133
rect 113714 270031 113748 270065
rect 113714 269963 113748 269997
rect 113714 269895 113748 269929
rect 113714 269827 113748 269861
rect 113714 269759 113748 269793
rect 113714 269691 113748 269725
rect 113714 269623 113748 269657
rect 113714 269555 113748 269589
rect 113714 269487 113748 269521
rect 113714 269419 113748 269453
rect 113714 269351 113748 269385
rect 113714 269283 113748 269317
rect 113714 269215 113748 269249
rect 113714 269147 113748 269181
rect 113932 270167 113966 270201
rect 113932 270099 113966 270133
rect 113932 270031 113966 270065
rect 113932 269963 113966 269997
rect 113932 269895 113966 269929
rect 113932 269827 113966 269861
rect 113932 269759 113966 269793
rect 113932 269691 113966 269725
rect 113932 269623 113966 269657
rect 113932 269555 113966 269589
rect 113932 269487 113966 269521
rect 113932 269419 113966 269453
rect 113932 269351 113966 269385
rect 113932 269283 113966 269317
rect 113932 269215 113966 269249
rect 113932 269147 113966 269181
rect 114114 270167 114148 270201
rect 114114 270099 114148 270133
rect 114114 270031 114148 270065
rect 114114 269963 114148 269997
rect 114114 269895 114148 269929
rect 114114 269827 114148 269861
rect 114114 269759 114148 269793
rect 114114 269691 114148 269725
rect 114114 269623 114148 269657
rect 114114 269555 114148 269589
rect 114114 269487 114148 269521
rect 114114 269419 114148 269453
rect 114114 269351 114148 269385
rect 114114 269283 114148 269317
rect 114114 269215 114148 269249
rect 114114 269147 114148 269181
rect 114332 270167 114366 270201
rect 114332 270099 114366 270133
rect 114332 270031 114366 270065
rect 114332 269963 114366 269997
rect 114332 269895 114366 269929
rect 114332 269827 114366 269861
rect 114332 269759 114366 269793
rect 114332 269691 114366 269725
rect 114332 269623 114366 269657
rect 114332 269555 114366 269589
rect 114332 269487 114366 269521
rect 114332 269419 114366 269453
rect 114332 269351 114366 269385
rect 114332 269283 114366 269317
rect 114332 269215 114366 269249
rect 114332 269147 114366 269181
rect 114514 270167 114548 270201
rect 114514 270099 114548 270133
rect 114514 270031 114548 270065
rect 114514 269963 114548 269997
rect 114514 269895 114548 269929
rect 114514 269827 114548 269861
rect 114514 269759 114548 269793
rect 114514 269691 114548 269725
rect 114514 269623 114548 269657
rect 114514 269555 114548 269589
rect 114514 269487 114548 269521
rect 114514 269419 114548 269453
rect 114514 269351 114548 269385
rect 114514 269283 114548 269317
rect 114514 269215 114548 269249
rect 114514 269147 114548 269181
rect 114732 270167 114766 270201
rect 114732 270099 114766 270133
rect 114732 270031 114766 270065
rect 114732 269963 114766 269997
rect 114732 269895 114766 269929
rect 114732 269827 114766 269861
rect 114732 269759 114766 269793
rect 114732 269691 114766 269725
rect 114732 269623 114766 269657
rect 114732 269555 114766 269589
rect 114732 269487 114766 269521
rect 114732 269419 114766 269453
rect 114732 269351 114766 269385
rect 114732 269283 114766 269317
rect 114732 269215 114766 269249
rect 114732 269147 114766 269181
rect 114914 270167 114948 270201
rect 114914 270099 114948 270133
rect 114914 270031 114948 270065
rect 114914 269963 114948 269997
rect 114914 269895 114948 269929
rect 114914 269827 114948 269861
rect 114914 269759 114948 269793
rect 114914 269691 114948 269725
rect 114914 269623 114948 269657
rect 114914 269555 114948 269589
rect 114914 269487 114948 269521
rect 114914 269419 114948 269453
rect 114914 269351 114948 269385
rect 114914 269283 114948 269317
rect 114914 269215 114948 269249
rect 114914 269147 114948 269181
rect 115132 270167 115166 270201
rect 115132 270099 115166 270133
rect 115132 270031 115166 270065
rect 115132 269963 115166 269997
rect 115132 269895 115166 269929
rect 115132 269827 115166 269861
rect 115132 269759 115166 269793
rect 115132 269691 115166 269725
rect 115132 269623 115166 269657
rect 115132 269555 115166 269589
rect 115132 269487 115166 269521
rect 115132 269419 115166 269453
rect 115132 269351 115166 269385
rect 115132 269283 115166 269317
rect 115132 269215 115166 269249
rect 115132 269147 115166 269181
rect 115314 270167 115348 270201
rect 115314 270099 115348 270133
rect 115314 270031 115348 270065
rect 115314 269963 115348 269997
rect 115314 269895 115348 269929
rect 115314 269827 115348 269861
rect 115314 269759 115348 269793
rect 115314 269691 115348 269725
rect 115314 269623 115348 269657
rect 115314 269555 115348 269589
rect 115314 269487 115348 269521
rect 115314 269419 115348 269453
rect 115314 269351 115348 269385
rect 115314 269283 115348 269317
rect 115314 269215 115348 269249
rect 115314 269147 115348 269181
rect 115532 270167 115566 270201
rect 115532 270099 115566 270133
rect 115532 270031 115566 270065
rect 115532 269963 115566 269997
rect 115532 269895 115566 269929
rect 115532 269827 115566 269861
rect 115532 269759 115566 269793
rect 115532 269691 115566 269725
rect 115532 269623 115566 269657
rect 115532 269555 115566 269589
rect 115532 269487 115566 269521
rect 115532 269419 115566 269453
rect 115532 269351 115566 269385
rect 115532 269283 115566 269317
rect 115532 269215 115566 269249
rect 115532 269147 115566 269181
rect 115714 270167 115748 270201
rect 115714 270099 115748 270133
rect 115714 270031 115748 270065
rect 115714 269963 115748 269997
rect 115714 269895 115748 269929
rect 115714 269827 115748 269861
rect 115714 269759 115748 269793
rect 115714 269691 115748 269725
rect 115714 269623 115748 269657
rect 115714 269555 115748 269589
rect 115714 269487 115748 269521
rect 115714 269419 115748 269453
rect 115714 269351 115748 269385
rect 115714 269283 115748 269317
rect 115714 269215 115748 269249
rect 115714 269147 115748 269181
rect 115932 270167 115966 270201
rect 115932 270099 115966 270133
rect 115932 270031 115966 270065
rect 115932 269963 115966 269997
rect 115932 269895 115966 269929
rect 115932 269827 115966 269861
rect 115932 269759 115966 269793
rect 115932 269691 115966 269725
rect 115932 269623 115966 269657
rect 115932 269555 115966 269589
rect 115932 269487 115966 269521
rect 115932 269419 115966 269453
rect 115932 269351 115966 269385
rect 115932 269283 115966 269317
rect 115932 269215 115966 269249
rect 115932 269147 115966 269181
rect 116114 270167 116148 270201
rect 116114 270099 116148 270133
rect 116114 270031 116148 270065
rect 116114 269963 116148 269997
rect 116114 269895 116148 269929
rect 116114 269827 116148 269861
rect 116114 269759 116148 269793
rect 116114 269691 116148 269725
rect 116114 269623 116148 269657
rect 116114 269555 116148 269589
rect 116114 269487 116148 269521
rect 116114 269419 116148 269453
rect 116114 269351 116148 269385
rect 116114 269283 116148 269317
rect 116114 269215 116148 269249
rect 116114 269147 116148 269181
rect 116332 270167 116366 270201
rect 116332 270099 116366 270133
rect 116332 270031 116366 270065
rect 116332 269963 116366 269997
rect 116332 269895 116366 269929
rect 116332 269827 116366 269861
rect 116332 269759 116366 269793
rect 116332 269691 116366 269725
rect 116332 269623 116366 269657
rect 116332 269555 116366 269589
rect 116332 269487 116366 269521
rect 116332 269419 116366 269453
rect 116332 269351 116366 269385
rect 116332 269283 116366 269317
rect 116332 269215 116366 269249
rect 116332 269147 116366 269181
rect 116514 270167 116548 270201
rect 116514 270099 116548 270133
rect 116514 270031 116548 270065
rect 116514 269963 116548 269997
rect 116514 269895 116548 269929
rect 116514 269827 116548 269861
rect 116514 269759 116548 269793
rect 116514 269691 116548 269725
rect 116514 269623 116548 269657
rect 116514 269555 116548 269589
rect 116514 269487 116548 269521
rect 116514 269419 116548 269453
rect 116514 269351 116548 269385
rect 116514 269283 116548 269317
rect 116514 269215 116548 269249
rect 116514 269147 116548 269181
rect 116732 270167 116766 270201
rect 116732 270099 116766 270133
rect 116732 270031 116766 270065
rect 116732 269963 116766 269997
rect 116732 269895 116766 269929
rect 116732 269827 116766 269861
rect 116732 269759 116766 269793
rect 116732 269691 116766 269725
rect 116732 269623 116766 269657
rect 116732 269555 116766 269589
rect 116732 269487 116766 269521
rect 116732 269419 116766 269453
rect 116732 269351 116766 269385
rect 116732 269283 116766 269317
rect 116732 269215 116766 269249
rect 116732 269147 116766 269181
rect 116914 270167 116948 270201
rect 116914 270099 116948 270133
rect 116914 270031 116948 270065
rect 116914 269963 116948 269997
rect 116914 269895 116948 269929
rect 116914 269827 116948 269861
rect 116914 269759 116948 269793
rect 116914 269691 116948 269725
rect 116914 269623 116948 269657
rect 116914 269555 116948 269589
rect 116914 269487 116948 269521
rect 116914 269419 116948 269453
rect 116914 269351 116948 269385
rect 116914 269283 116948 269317
rect 116914 269215 116948 269249
rect 116914 269147 116948 269181
rect 117132 270167 117166 270201
rect 117132 270099 117166 270133
rect 117132 270031 117166 270065
rect 117132 269963 117166 269997
rect 117132 269895 117166 269929
rect 117132 269827 117166 269861
rect 117132 269759 117166 269793
rect 117132 269691 117166 269725
rect 117132 269623 117166 269657
rect 117132 269555 117166 269589
rect 117132 269487 117166 269521
rect 117132 269419 117166 269453
rect 117132 269351 117166 269385
rect 117132 269283 117166 269317
rect 117132 269215 117166 269249
rect 117132 269147 117166 269181
rect 117314 270167 117348 270201
rect 117314 270099 117348 270133
rect 117314 270031 117348 270065
rect 117314 269963 117348 269997
rect 117314 269895 117348 269929
rect 117314 269827 117348 269861
rect 117314 269759 117348 269793
rect 117314 269691 117348 269725
rect 117314 269623 117348 269657
rect 117314 269555 117348 269589
rect 117314 269487 117348 269521
rect 117314 269419 117348 269453
rect 117314 269351 117348 269385
rect 117314 269283 117348 269317
rect 117314 269215 117348 269249
rect 117314 269147 117348 269181
rect 117532 270167 117566 270201
rect 117532 270099 117566 270133
rect 117532 270031 117566 270065
rect 117532 269963 117566 269997
rect 117532 269895 117566 269929
rect 117532 269827 117566 269861
rect 117532 269759 117566 269793
rect 117532 269691 117566 269725
rect 117532 269623 117566 269657
rect 117532 269555 117566 269589
rect 117532 269487 117566 269521
rect 117532 269419 117566 269453
rect 117532 269351 117566 269385
rect 117532 269283 117566 269317
rect 117532 269215 117566 269249
rect 117532 269147 117566 269181
rect 117714 270167 117748 270201
rect 117714 270099 117748 270133
rect 117714 270031 117748 270065
rect 117714 269963 117748 269997
rect 117714 269895 117748 269929
rect 117714 269827 117748 269861
rect 117714 269759 117748 269793
rect 117714 269691 117748 269725
rect 117714 269623 117748 269657
rect 117714 269555 117748 269589
rect 117714 269487 117748 269521
rect 117714 269419 117748 269453
rect 117714 269351 117748 269385
rect 117714 269283 117748 269317
rect 117714 269215 117748 269249
rect 117714 269147 117748 269181
rect 117932 270167 117966 270201
rect 117932 270099 117966 270133
rect 117932 270031 117966 270065
rect 117932 269963 117966 269997
rect 117932 269895 117966 269929
rect 117932 269827 117966 269861
rect 117932 269759 117966 269793
rect 117932 269691 117966 269725
rect 117932 269623 117966 269657
rect 117932 269555 117966 269589
rect 117932 269487 117966 269521
rect 117932 269419 117966 269453
rect 117932 269351 117966 269385
rect 117932 269283 117966 269317
rect 117932 269215 117966 269249
rect 117932 269147 117966 269181
rect 118114 270167 118148 270201
rect 118114 270099 118148 270133
rect 118114 270031 118148 270065
rect 118114 269963 118148 269997
rect 118114 269895 118148 269929
rect 118114 269827 118148 269861
rect 118114 269759 118148 269793
rect 118114 269691 118148 269725
rect 118114 269623 118148 269657
rect 118114 269555 118148 269589
rect 118114 269487 118148 269521
rect 118114 269419 118148 269453
rect 118114 269351 118148 269385
rect 118114 269283 118148 269317
rect 118114 269215 118148 269249
rect 118114 269147 118148 269181
rect 118332 270167 118366 270201
rect 118332 270099 118366 270133
rect 118332 270031 118366 270065
rect 118332 269963 118366 269997
rect 118332 269895 118366 269929
rect 118332 269827 118366 269861
rect 118332 269759 118366 269793
rect 118332 269691 118366 269725
rect 118332 269623 118366 269657
rect 118332 269555 118366 269589
rect 118332 269487 118366 269521
rect 118332 269419 118366 269453
rect 118332 269351 118366 269385
rect 118332 269283 118366 269317
rect 118332 269215 118366 269249
rect 118332 269147 118366 269181
rect 118514 270167 118548 270201
rect 118514 270099 118548 270133
rect 118514 270031 118548 270065
rect 118514 269963 118548 269997
rect 118514 269895 118548 269929
rect 118514 269827 118548 269861
rect 118514 269759 118548 269793
rect 118514 269691 118548 269725
rect 118514 269623 118548 269657
rect 118514 269555 118548 269589
rect 118514 269487 118548 269521
rect 118514 269419 118548 269453
rect 118514 269351 118548 269385
rect 118514 269283 118548 269317
rect 118514 269215 118548 269249
rect 118514 269147 118548 269181
rect 118732 270167 118766 270201
rect 118732 270099 118766 270133
rect 118732 270031 118766 270065
rect 118732 269963 118766 269997
rect 118732 269895 118766 269929
rect 118732 269827 118766 269861
rect 118732 269759 118766 269793
rect 118732 269691 118766 269725
rect 118732 269623 118766 269657
rect 118732 269555 118766 269589
rect 118732 269487 118766 269521
rect 118732 269419 118766 269453
rect 118732 269351 118766 269385
rect 118732 269283 118766 269317
rect 118732 269215 118766 269249
rect 118732 269147 118766 269181
rect 122906 274813 122940 274847
rect 122906 274745 122940 274779
rect 122906 274677 122940 274711
rect 123964 274813 123998 274847
rect 123964 274745 123998 274779
rect 123964 274677 123998 274711
rect 122231 274215 122265 274249
rect 122231 274147 122265 274181
rect 122231 274079 122265 274113
rect 122231 274011 122265 274045
rect 122231 273943 122265 273977
rect 122231 273875 122265 273909
rect 122231 273807 122265 273841
rect 122489 274215 122523 274249
rect 122489 274147 122523 274181
rect 122489 274079 122523 274113
rect 122489 274011 122523 274045
rect 122489 273943 122523 273977
rect 122489 273875 122523 273909
rect 122489 273807 122523 273841
rect 122647 274215 122681 274249
rect 122647 274147 122681 274181
rect 122647 274079 122681 274113
rect 122647 274011 122681 274045
rect 122647 273943 122681 273977
rect 122647 273875 122681 273909
rect 122647 273807 122681 273841
rect 122905 274215 122939 274249
rect 122905 274147 122939 274181
rect 122905 274079 122939 274113
rect 122905 274011 122939 274045
rect 122905 273943 122939 273977
rect 122905 273875 122939 273909
rect 122905 273807 122939 273841
rect 123063 274215 123097 274249
rect 123063 274147 123097 274181
rect 123063 274079 123097 274113
rect 123063 274011 123097 274045
rect 123063 273943 123097 273977
rect 123063 273875 123097 273909
rect 123063 273807 123097 273841
rect 123321 274215 123355 274249
rect 123321 274147 123355 274181
rect 123321 274079 123355 274113
rect 123321 274011 123355 274045
rect 123321 273943 123355 273977
rect 123321 273875 123355 273909
rect 123321 273807 123355 273841
rect 123479 274215 123513 274249
rect 123479 274147 123513 274181
rect 123479 274079 123513 274113
rect 123479 274011 123513 274045
rect 123479 273943 123513 273977
rect 123479 273875 123513 273909
rect 123479 273807 123513 273841
rect 123737 274215 123771 274249
rect 123737 274147 123771 274181
rect 123737 274079 123771 274113
rect 123737 274011 123771 274045
rect 123737 273943 123771 273977
rect 123737 273875 123771 273909
rect 123737 273807 123771 273841
rect 123895 274215 123929 274249
rect 123895 274147 123929 274181
rect 123895 274079 123929 274113
rect 123895 274011 123929 274045
rect 123895 273943 123929 273977
rect 123895 273875 123929 273909
rect 123895 273807 123929 273841
rect 124153 274215 124187 274249
rect 124153 274147 124187 274181
rect 124153 274079 124187 274113
rect 124153 274011 124187 274045
rect 124153 273943 124187 273977
rect 124153 273875 124187 273909
rect 124153 273807 124187 273841
rect 124311 274215 124345 274249
rect 124311 274147 124345 274181
rect 124311 274079 124345 274113
rect 124311 274011 124345 274045
rect 124311 273943 124345 273977
rect 124311 273875 124345 273909
rect 124311 273807 124345 273841
rect 124569 274215 124603 274249
rect 124569 274147 124603 274181
rect 124569 274079 124603 274113
rect 124569 274011 124603 274045
rect 124569 273943 124603 273977
rect 124569 273875 124603 273909
rect 124569 273807 124603 273841
rect 124221 272532 124255 272566
rect 124289 272532 124323 272566
rect 124357 272532 124391 272566
rect 124425 272532 124459 272566
rect 124493 272532 124527 272566
rect 124561 272532 124595 272566
rect 124629 272532 124663 272566
rect 124221 272274 124255 272308
rect 124289 272274 124323 272308
rect 124357 272274 124391 272308
rect 124425 272274 124459 272308
rect 124493 272274 124527 272308
rect 124561 272274 124595 272308
rect 124629 272274 124663 272308
rect 124221 272116 124255 272150
rect 124289 272116 124323 272150
rect 124357 272116 124391 272150
rect 124425 272116 124459 272150
rect 124493 272116 124527 272150
rect 124561 272116 124595 272150
rect 124629 272116 124663 272150
rect 124221 271858 124255 271892
rect 124289 271858 124323 271892
rect 124357 271858 124391 271892
rect 124425 271858 124459 271892
rect 124493 271858 124527 271892
rect 124561 271858 124595 271892
rect 124629 271858 124663 271892
rect 124221 271700 124255 271734
rect 124289 271700 124323 271734
rect 124357 271700 124391 271734
rect 124425 271700 124459 271734
rect 124493 271700 124527 271734
rect 124561 271700 124595 271734
rect 124629 271700 124663 271734
rect 124221 271442 124255 271476
rect 124289 271442 124323 271476
rect 124357 271442 124391 271476
rect 124425 271442 124459 271476
rect 124493 271442 124527 271476
rect 124561 271442 124595 271476
rect 124629 271442 124663 271476
rect 124221 271284 124255 271318
rect 124289 271284 124323 271318
rect 124357 271284 124391 271318
rect 124425 271284 124459 271318
rect 124493 271284 124527 271318
rect 124561 271284 124595 271318
rect 124629 271284 124663 271318
rect 124221 271026 124255 271060
rect 124289 271026 124323 271060
rect 124357 271026 124391 271060
rect 124425 271026 124459 271060
rect 124493 271026 124527 271060
rect 124561 271026 124595 271060
rect 124629 271026 124663 271060
rect 124221 270868 124255 270902
rect 124289 270868 124323 270902
rect 124357 270868 124391 270902
rect 124425 270868 124459 270902
rect 124493 270868 124527 270902
rect 124561 270868 124595 270902
rect 124629 270868 124663 270902
rect 124221 270610 124255 270644
rect 124289 270610 124323 270644
rect 124357 270610 124391 270644
rect 124425 270610 124459 270644
rect 124493 270610 124527 270644
rect 124561 270610 124595 270644
rect 124629 270610 124663 270644
rect 124221 270452 124255 270486
rect 124289 270452 124323 270486
rect 124357 270452 124391 270486
rect 124425 270452 124459 270486
rect 124493 270452 124527 270486
rect 124561 270452 124595 270486
rect 124629 270452 124663 270486
rect 124221 270194 124255 270228
rect 124289 270194 124323 270228
rect 124357 270194 124391 270228
rect 124425 270194 124459 270228
rect 124493 270194 124527 270228
rect 124561 270194 124595 270228
rect 124629 270194 124663 270228
rect 124221 270036 124255 270070
rect 124289 270036 124323 270070
rect 124357 270036 124391 270070
rect 124425 270036 124459 270070
rect 124493 270036 124527 270070
rect 124561 270036 124595 270070
rect 124629 270036 124663 270070
rect 124221 269778 124255 269812
rect 124289 269778 124323 269812
rect 124357 269778 124391 269812
rect 124425 269778 124459 269812
rect 124493 269778 124527 269812
rect 124561 269778 124595 269812
rect 124629 269778 124663 269812
rect 124221 269620 124255 269654
rect 124289 269620 124323 269654
rect 124357 269620 124391 269654
rect 124425 269620 124459 269654
rect 124493 269620 124527 269654
rect 124561 269620 124595 269654
rect 124629 269620 124663 269654
rect 124221 269362 124255 269396
rect 124289 269362 124323 269396
rect 124357 269362 124391 269396
rect 124425 269362 124459 269396
rect 124493 269362 124527 269396
rect 124561 269362 124595 269396
rect 124629 269362 124663 269396
<< pdiffc >>
rect 106380 279023 106414 279057
rect 106448 279023 106482 279057
rect 106516 279023 106550 279057
rect 106584 279023 106618 279057
rect 106652 279023 106686 279057
rect 106720 279023 106754 279057
rect 106788 279023 106822 279057
rect 106856 279023 106890 279057
rect 106924 279023 106958 279057
rect 106992 279023 107026 279057
rect 107060 279023 107094 279057
rect 107128 279023 107162 279057
rect 107196 279023 107230 279057
rect 107264 279023 107298 279057
rect 107332 279023 107366 279057
rect 107400 279023 107434 279057
rect 107468 279023 107502 279057
rect 107536 279023 107570 279057
rect 106380 278711 106414 278745
rect 106448 278711 106482 278745
rect 106516 278711 106550 278745
rect 106584 278711 106618 278745
rect 106652 278711 106686 278745
rect 106720 278711 106754 278745
rect 106788 278711 106822 278745
rect 106856 278711 106890 278745
rect 106924 278711 106958 278745
rect 106992 278711 107026 278745
rect 107060 278711 107094 278745
rect 107128 278711 107162 278745
rect 107196 278711 107230 278745
rect 107264 278711 107298 278745
rect 107332 278711 107366 278745
rect 107400 278711 107434 278745
rect 107468 278711 107502 278745
rect 107536 278711 107570 278745
rect 106380 278423 106414 278457
rect 106448 278423 106482 278457
rect 106516 278423 106550 278457
rect 106584 278423 106618 278457
rect 106652 278423 106686 278457
rect 106720 278423 106754 278457
rect 106788 278423 106822 278457
rect 106856 278423 106890 278457
rect 106924 278423 106958 278457
rect 106992 278423 107026 278457
rect 107060 278423 107094 278457
rect 107128 278423 107162 278457
rect 107196 278423 107230 278457
rect 107264 278423 107298 278457
rect 107332 278423 107366 278457
rect 107400 278423 107434 278457
rect 107468 278423 107502 278457
rect 107536 278423 107570 278457
rect 106380 278111 106414 278145
rect 106448 278111 106482 278145
rect 106516 278111 106550 278145
rect 106584 278111 106618 278145
rect 106652 278111 106686 278145
rect 106720 278111 106754 278145
rect 106788 278111 106822 278145
rect 106856 278111 106890 278145
rect 106924 278111 106958 278145
rect 106992 278111 107026 278145
rect 107060 278111 107094 278145
rect 107128 278111 107162 278145
rect 107196 278111 107230 278145
rect 107264 278111 107298 278145
rect 107332 278111 107366 278145
rect 107400 278111 107434 278145
rect 107468 278111 107502 278145
rect 107536 278111 107570 278145
rect 106515 277176 106549 277210
rect 106583 277176 106617 277210
rect 106651 277176 106685 277210
rect 106719 277176 106753 277210
rect 106787 277176 106821 277210
rect 106855 277176 106889 277210
rect 106923 277176 106957 277210
rect 106991 277176 107025 277210
rect 107059 277176 107093 277210
rect 107127 277176 107161 277210
rect 107195 277176 107229 277210
rect 107263 277176 107297 277210
rect 107331 277176 107365 277210
rect 107399 277176 107433 277210
rect 107467 277176 107501 277210
rect 106515 277044 106549 277078
rect 106583 277044 106617 277078
rect 106651 277044 106685 277078
rect 106719 277044 106753 277078
rect 106787 277044 106821 277078
rect 106855 277044 106889 277078
rect 106923 277044 106957 277078
rect 106991 277044 107025 277078
rect 107059 277044 107093 277078
rect 107127 277044 107161 277078
rect 107195 277044 107229 277078
rect 107263 277044 107297 277078
rect 107331 277044 107365 277078
rect 107399 277044 107433 277078
rect 107467 277044 107501 277078
rect 106989 275725 107023 275759
rect 107057 275725 107091 275759
rect 107489 275725 107523 275759
rect 107557 275725 107591 275759
rect 107989 275725 108023 275759
rect 108057 275725 108091 275759
rect 108489 275725 108523 275759
rect 108557 275725 108591 275759
rect 108989 275725 109023 275759
rect 109057 275725 109091 275759
rect 109489 275725 109523 275759
rect 109557 275725 109591 275759
rect 106989 274889 107023 274923
rect 107057 274889 107091 274923
rect 107489 274889 107523 274923
rect 107557 274889 107591 274923
rect 107989 274889 108023 274923
rect 108057 274889 108091 274923
rect 108489 274889 108523 274923
rect 108557 274889 108591 274923
rect 108989 274889 109023 274923
rect 109057 274889 109091 274923
rect 109489 274889 109523 274923
rect 109557 274889 109591 274923
rect 109394 272365 109428 272399
rect 109394 272297 109428 272331
rect 109394 272229 109428 272263
rect 109394 272161 109428 272195
rect 109394 272093 109428 272127
rect 109394 272025 109428 272059
rect 109394 271957 109428 271991
rect 109394 271889 109428 271923
rect 109394 271821 109428 271855
rect 109394 271753 109428 271787
rect 109394 271685 109428 271719
rect 109394 271617 109428 271651
rect 109394 271549 109428 271583
rect 109394 271481 109428 271515
rect 109394 271413 109428 271447
rect 109394 271345 109428 271379
rect 109394 271277 109428 271311
rect 109394 271209 109428 271243
rect 109394 271141 109428 271175
rect 109394 271073 109428 271107
rect 109394 271005 109428 271039
rect 109394 270937 109428 270971
rect 109394 270869 109428 270903
rect 109394 270801 109428 270835
rect 109394 270733 109428 270767
rect 109522 272365 109556 272399
rect 109522 272297 109556 272331
rect 109522 272229 109556 272263
rect 109522 272161 109556 272195
rect 109522 272093 109556 272127
rect 109522 272025 109556 272059
rect 109522 271957 109556 271991
rect 109522 271889 109556 271923
rect 109522 271821 109556 271855
rect 109522 271753 109556 271787
rect 109522 271685 109556 271719
rect 109522 271617 109556 271651
rect 109522 271549 109556 271583
rect 109522 271481 109556 271515
rect 109522 271413 109556 271447
rect 109522 271345 109556 271379
rect 109522 271277 109556 271311
rect 109522 271209 109556 271243
rect 109522 271141 109556 271175
rect 109522 271073 109556 271107
rect 109522 271005 109556 271039
rect 109522 270937 109556 270971
rect 109522 270869 109556 270903
rect 109522 270801 109556 270835
rect 109522 270733 109556 270767
rect 114672 280815 114706 280849
rect 114740 280815 114774 280849
rect 114808 280815 114842 280849
rect 114672 280357 114706 280391
rect 114740 280357 114774 280391
rect 114808 280357 114842 280391
rect 114672 280129 114706 280163
rect 114740 280129 114774 280163
rect 114808 280129 114842 280163
rect 114672 279911 114706 279945
rect 114740 279911 114774 279945
rect 114808 279911 114842 279945
rect 114672 279721 114706 279755
rect 114740 279721 114774 279755
rect 114808 279721 114842 279755
rect 114672 279503 114706 279537
rect 114740 279503 114774 279537
rect 114808 279503 114842 279537
rect 115363 280815 115397 280849
rect 115431 280815 115465 280849
rect 115499 280815 115533 280849
rect 115363 280357 115397 280391
rect 115431 280357 115465 280391
rect 115499 280357 115533 280391
rect 115363 280129 115397 280163
rect 115431 280129 115465 280163
rect 115499 280129 115533 280163
rect 115363 279911 115397 279945
rect 115431 279911 115465 279945
rect 115499 279911 115533 279945
rect 115363 279721 115397 279755
rect 115431 279721 115465 279755
rect 115499 279721 115533 279755
rect 115363 279503 115397 279537
rect 115431 279503 115465 279537
rect 115499 279503 115533 279537
rect 114672 279149 114706 279183
rect 114740 279149 114774 279183
rect 114808 279149 114842 279183
rect 114672 278691 114706 278725
rect 114740 278691 114774 278725
rect 114808 278691 114842 278725
rect 114672 278463 114706 278497
rect 114740 278463 114774 278497
rect 114808 278463 114842 278497
rect 114672 278245 114706 278279
rect 114740 278245 114774 278279
rect 114808 278245 114842 278279
rect 114672 278055 114706 278089
rect 114740 278055 114774 278089
rect 114808 278055 114842 278089
rect 114672 277837 114706 277871
rect 114740 277837 114774 277871
rect 114808 277837 114842 277871
rect 115363 279149 115397 279183
rect 115431 279149 115465 279183
rect 115499 279149 115533 279183
rect 115363 278691 115397 278725
rect 115431 278691 115465 278725
rect 115499 278691 115533 278725
rect 115363 278463 115397 278497
rect 115431 278463 115465 278497
rect 115499 278463 115533 278497
rect 115363 278245 115397 278279
rect 115431 278245 115465 278279
rect 115499 278245 115533 278279
rect 115363 278055 115397 278089
rect 115431 278055 115465 278089
rect 115499 278055 115533 278089
rect 115363 277837 115397 277871
rect 115431 277837 115465 277871
rect 115499 277837 115533 277871
rect 114672 277483 114706 277517
rect 114740 277483 114774 277517
rect 114808 277483 114842 277517
rect 114672 277025 114706 277059
rect 114740 277025 114774 277059
rect 114808 277025 114842 277059
rect 114672 276797 114706 276831
rect 114740 276797 114774 276831
rect 114808 276797 114842 276831
rect 114672 276579 114706 276613
rect 114740 276579 114774 276613
rect 114808 276579 114842 276613
rect 114672 276389 114706 276423
rect 114740 276389 114774 276423
rect 114808 276389 114842 276423
rect 114672 276171 114706 276205
rect 114740 276171 114774 276205
rect 114808 276171 114842 276205
rect 115363 277483 115397 277517
rect 115431 277483 115465 277517
rect 115499 277483 115533 277517
rect 115363 277025 115397 277059
rect 115431 277025 115465 277059
rect 115499 277025 115533 277059
rect 115363 276797 115397 276831
rect 115431 276797 115465 276831
rect 115499 276797 115533 276831
rect 115363 276579 115397 276613
rect 115431 276579 115465 276613
rect 115499 276579 115533 276613
rect 115363 276389 115397 276423
rect 115431 276389 115465 276423
rect 115499 276389 115533 276423
rect 115363 276171 115397 276205
rect 115431 276171 115465 276205
rect 115499 276171 115533 276205
rect 114672 275817 114706 275851
rect 114740 275817 114774 275851
rect 114808 275817 114842 275851
rect 114672 275359 114706 275393
rect 114740 275359 114774 275393
rect 114808 275359 114842 275393
rect 114672 275131 114706 275165
rect 114740 275131 114774 275165
rect 114808 275131 114842 275165
rect 114672 274913 114706 274947
rect 114740 274913 114774 274947
rect 114808 274913 114842 274947
rect 114672 274723 114706 274757
rect 114740 274723 114774 274757
rect 114808 274723 114842 274757
rect 114672 274505 114706 274539
rect 114740 274505 114774 274539
rect 114808 274505 114842 274539
rect 115363 275817 115397 275851
rect 115431 275817 115465 275851
rect 115499 275817 115533 275851
rect 115363 275359 115397 275393
rect 115431 275359 115465 275393
rect 115499 275359 115533 275393
rect 115363 275131 115397 275165
rect 115431 275131 115465 275165
rect 115499 275131 115533 275165
rect 115363 274913 115397 274947
rect 115431 274913 115465 274947
rect 115499 274913 115533 274947
rect 115363 274723 115397 274757
rect 115431 274723 115465 274757
rect 115499 274723 115533 274757
rect 115363 274505 115397 274539
rect 115431 274505 115465 274539
rect 115499 274505 115533 274539
rect 114672 274151 114706 274185
rect 114740 274151 114774 274185
rect 114808 274151 114842 274185
rect 114672 273693 114706 273727
rect 114740 273693 114774 273727
rect 114808 273693 114842 273727
rect 114672 273465 114706 273499
rect 114740 273465 114774 273499
rect 114808 273465 114842 273499
rect 114672 273247 114706 273281
rect 114740 273247 114774 273281
rect 114808 273247 114842 273281
rect 114672 273057 114706 273091
rect 114740 273057 114774 273091
rect 114808 273057 114842 273091
rect 114672 272839 114706 272873
rect 114740 272839 114774 272873
rect 114808 272839 114842 272873
rect 115363 274151 115397 274185
rect 115431 274151 115465 274185
rect 115499 274151 115533 274185
rect 115363 273693 115397 273727
rect 115431 273693 115465 273727
rect 115499 273693 115533 273727
rect 115363 273465 115397 273499
rect 115431 273465 115465 273499
rect 115499 273465 115533 273499
rect 115363 273247 115397 273281
rect 115431 273247 115465 273281
rect 115499 273247 115533 273281
rect 115363 273057 115397 273091
rect 115431 273057 115465 273091
rect 115499 273057 115533 273091
rect 115363 272839 115397 272873
rect 115431 272839 115465 272873
rect 115499 272839 115533 272873
rect 112532 271257 112566 271291
rect 112532 271189 112566 271223
rect 112532 271121 112566 271155
rect 112750 271257 112784 271291
rect 112750 271189 112784 271223
rect 112750 271121 112784 271155
rect 112932 271257 112966 271291
rect 112932 271189 112966 271223
rect 112932 271121 112966 271155
rect 113150 271257 113184 271291
rect 113150 271189 113184 271223
rect 113150 271121 113184 271155
rect 113332 271257 113366 271291
rect 113332 271189 113366 271223
rect 113332 271121 113366 271155
rect 113550 271257 113584 271291
rect 113550 271189 113584 271223
rect 113550 271121 113584 271155
rect 113732 271257 113766 271291
rect 113732 271189 113766 271223
rect 113732 271121 113766 271155
rect 113950 271257 113984 271291
rect 113950 271189 113984 271223
rect 113950 271121 113984 271155
rect 114591 271228 114625 271262
rect 114591 271160 114625 271194
rect 114591 271092 114625 271126
rect 114809 271228 114843 271262
rect 114809 271160 114843 271194
rect 114809 271092 114843 271126
rect 114991 271228 115025 271262
rect 114991 271160 115025 271194
rect 114991 271092 115025 271126
rect 115209 271228 115243 271262
rect 115209 271160 115243 271194
rect 115209 271092 115243 271126
rect 120383 280570 120417 280604
rect 120841 280570 120875 280604
rect 121083 280570 121117 280604
rect 121541 280570 121575 280604
rect 120383 280190 120417 280224
rect 120383 280122 120417 280156
rect 120383 280054 120417 280088
rect 120383 279986 120417 280020
rect 120383 279918 120417 279952
rect 120383 279850 120417 279884
rect 120383 279782 120417 279816
rect 120841 280190 120875 280224
rect 120841 280122 120875 280156
rect 120841 280054 120875 280088
rect 120841 279986 120875 280020
rect 120841 279918 120875 279952
rect 120841 279850 120875 279884
rect 120841 279782 120875 279816
rect 121083 280190 121117 280224
rect 121083 280122 121117 280156
rect 121083 280054 121117 280088
rect 121083 279986 121117 280020
rect 121083 279918 121117 279952
rect 121083 279850 121117 279884
rect 121083 279782 121117 279816
rect 121541 280190 121575 280224
rect 121541 280122 121575 280156
rect 121541 280054 121575 280088
rect 121541 279986 121575 280020
rect 121541 279918 121575 279952
rect 121541 279850 121575 279884
rect 121541 279782 121575 279816
rect 120383 279406 120417 279440
rect 120383 279338 120417 279372
rect 120383 279270 120417 279304
rect 120383 279202 120417 279236
rect 120383 279134 120417 279168
rect 120383 279066 120417 279100
rect 120383 278998 120417 279032
rect 120841 279406 120875 279440
rect 120841 279338 120875 279372
rect 120841 279270 120875 279304
rect 120841 279202 120875 279236
rect 120841 279134 120875 279168
rect 120841 279066 120875 279100
rect 120841 278998 120875 279032
rect 121083 279406 121117 279440
rect 121083 279338 121117 279372
rect 121083 279270 121117 279304
rect 121083 279202 121117 279236
rect 121083 279134 121117 279168
rect 121083 279066 121117 279100
rect 121083 278998 121117 279032
rect 121541 279406 121575 279440
rect 121541 279338 121575 279372
rect 121541 279270 121575 279304
rect 121541 279202 121575 279236
rect 121541 279134 121575 279168
rect 121541 279066 121575 279100
rect 121541 278998 121575 279032
rect 122310 280360 122344 280394
rect 122310 280292 122344 280326
rect 122310 280224 122344 280258
rect 122310 280156 122344 280190
rect 122310 280088 122344 280122
rect 122310 280020 122344 280054
rect 122310 279952 122344 279986
rect 122768 280360 122802 280394
rect 122768 280292 122802 280326
rect 122768 280224 122802 280258
rect 122768 280156 122802 280190
rect 122768 280088 122802 280122
rect 122768 280020 122802 280054
rect 122768 279952 122802 279986
rect 123010 280360 123044 280394
rect 123010 280292 123044 280326
rect 123010 280224 123044 280258
rect 123010 280156 123044 280190
rect 123010 280088 123044 280122
rect 123010 280020 123044 280054
rect 123010 279952 123044 279986
rect 123468 280360 123502 280394
rect 123468 280292 123502 280326
rect 123468 280224 123502 280258
rect 123468 280156 123502 280190
rect 123468 280088 123502 280122
rect 123468 280020 123502 280054
rect 123468 279952 123502 279986
rect 122310 279576 122344 279610
rect 122310 279508 122344 279542
rect 122310 279440 122344 279474
rect 122310 279372 122344 279406
rect 122310 279304 122344 279338
rect 122310 279236 122344 279270
rect 122310 279168 122344 279202
rect 122768 279576 122802 279610
rect 122768 279508 122802 279542
rect 122768 279440 122802 279474
rect 122768 279372 122802 279406
rect 122768 279304 122802 279338
rect 122768 279236 122802 279270
rect 122768 279168 122802 279202
rect 123010 279576 123044 279610
rect 123010 279508 123044 279542
rect 123010 279440 123044 279474
rect 123010 279372 123044 279406
rect 123010 279304 123044 279338
rect 123010 279236 123044 279270
rect 123010 279168 123044 279202
rect 123468 279576 123502 279610
rect 123468 279508 123502 279542
rect 123468 279440 123502 279474
rect 123468 279372 123502 279406
rect 123468 279304 123502 279338
rect 123468 279236 123502 279270
rect 123468 279168 123502 279202
rect 120383 278622 120417 278656
rect 120383 278554 120417 278588
rect 120383 278486 120417 278520
rect 120383 278418 120417 278452
rect 120383 278350 120417 278384
rect 120383 278282 120417 278316
rect 120383 278214 120417 278248
rect 120841 278622 120875 278656
rect 120841 278554 120875 278588
rect 120841 278486 120875 278520
rect 120841 278418 120875 278452
rect 120841 278350 120875 278384
rect 120841 278282 120875 278316
rect 120841 278214 120875 278248
rect 121083 278622 121117 278656
rect 121083 278554 121117 278588
rect 121083 278486 121117 278520
rect 121083 278418 121117 278452
rect 121083 278350 121117 278384
rect 121083 278282 121117 278316
rect 121083 278214 121117 278248
rect 121541 278622 121575 278656
rect 121541 278554 121575 278588
rect 121541 278486 121575 278520
rect 121541 278418 121575 278452
rect 121541 278350 121575 278384
rect 121541 278282 121575 278316
rect 121541 278214 121575 278248
rect 120383 277838 120417 277872
rect 120383 277770 120417 277804
rect 120383 277702 120417 277736
rect 120383 277634 120417 277668
rect 120383 277566 120417 277600
rect 120383 277498 120417 277532
rect 120383 277430 120417 277464
rect 120841 277838 120875 277872
rect 120841 277770 120875 277804
rect 120841 277702 120875 277736
rect 120841 277634 120875 277668
rect 120841 277566 120875 277600
rect 120841 277498 120875 277532
rect 120841 277430 120875 277464
rect 121083 277838 121117 277872
rect 121083 277770 121117 277804
rect 121083 277702 121117 277736
rect 121083 277634 121117 277668
rect 121083 277566 121117 277600
rect 121083 277498 121117 277532
rect 121083 277430 121117 277464
rect 121541 277838 121575 277872
rect 121541 277770 121575 277804
rect 121541 277702 121575 277736
rect 121541 277634 121575 277668
rect 121541 277566 121575 277600
rect 121541 277498 121575 277532
rect 121541 277430 121575 277464
rect 120383 277054 120417 277088
rect 120383 276986 120417 277020
rect 120383 276918 120417 276952
rect 120383 276850 120417 276884
rect 120383 276782 120417 276816
rect 120383 276714 120417 276748
rect 120383 276646 120417 276680
rect 120841 277054 120875 277088
rect 120841 276986 120875 277020
rect 120841 276918 120875 276952
rect 120841 276850 120875 276884
rect 120841 276782 120875 276816
rect 120841 276714 120875 276748
rect 120841 276646 120875 276680
rect 121083 277054 121117 277088
rect 121083 276986 121117 277020
rect 121083 276918 121117 276952
rect 121083 276850 121117 276884
rect 121083 276782 121117 276816
rect 121083 276714 121117 276748
rect 121083 276646 121117 276680
rect 121541 277054 121575 277088
rect 121541 276986 121575 277020
rect 121541 276918 121575 276952
rect 121541 276850 121575 276884
rect 121541 276782 121575 276816
rect 121541 276714 121575 276748
rect 121541 276646 121575 276680
rect 120383 276270 120417 276304
rect 120383 276202 120417 276236
rect 120383 276134 120417 276168
rect 120383 276066 120417 276100
rect 120383 275998 120417 276032
rect 120383 275930 120417 275964
rect 120383 275862 120417 275896
rect 120841 276270 120875 276304
rect 120841 276202 120875 276236
rect 120841 276134 120875 276168
rect 120841 276066 120875 276100
rect 120841 275998 120875 276032
rect 120841 275930 120875 275964
rect 120841 275862 120875 275896
rect 121083 276270 121117 276304
rect 121083 276202 121117 276236
rect 121083 276134 121117 276168
rect 121083 276066 121117 276100
rect 121083 275998 121117 276032
rect 121083 275930 121117 275964
rect 121083 275862 121117 275896
rect 121541 276270 121575 276304
rect 121541 276202 121575 276236
rect 121541 276134 121575 276168
rect 121541 276066 121575 276100
rect 121541 275998 121575 276032
rect 121541 275930 121575 275964
rect 121541 275862 121575 275896
rect 120383 275486 120417 275520
rect 120383 275418 120417 275452
rect 120383 275350 120417 275384
rect 120383 275282 120417 275316
rect 120383 275214 120417 275248
rect 120383 275146 120417 275180
rect 120383 275078 120417 275112
rect 120841 275486 120875 275520
rect 120841 275418 120875 275452
rect 120841 275350 120875 275384
rect 120841 275282 120875 275316
rect 120841 275214 120875 275248
rect 120841 275146 120875 275180
rect 120841 275078 120875 275112
rect 121083 275486 121117 275520
rect 121083 275418 121117 275452
rect 121083 275350 121117 275384
rect 121083 275282 121117 275316
rect 121083 275214 121117 275248
rect 121083 275146 121117 275180
rect 121083 275078 121117 275112
rect 121541 275486 121575 275520
rect 121541 275418 121575 275452
rect 121541 275350 121575 275384
rect 121541 275282 121575 275316
rect 121541 275214 121575 275248
rect 121541 275146 121575 275180
rect 121541 275078 121575 275112
rect 122368 278216 122402 278250
rect 122368 278148 122402 278182
rect 122368 278080 122402 278114
rect 122368 278012 122402 278046
rect 122368 277944 122402 277978
rect 122368 277876 122402 277910
rect 122368 277808 122402 277842
rect 123302 278216 123336 278250
rect 123302 278148 123336 278182
rect 123302 278080 123336 278114
rect 123302 278012 123336 278046
rect 123302 277944 123336 277978
rect 123302 277876 123336 277910
rect 123302 277808 123336 277842
rect 123610 278026 123644 278060
rect 123610 277958 123644 277992
rect 123610 277890 123644 277924
rect 123610 277822 123644 277856
rect 123610 277754 123644 277788
rect 123610 277686 123644 277720
rect 123610 277618 123644 277652
rect 123610 277550 123644 277584
rect 122370 277433 122404 277467
rect 123228 277433 123262 277467
rect 123610 277482 123644 277516
rect 123610 277414 123644 277448
rect 124222 278026 124256 278060
rect 124222 277958 124256 277992
rect 124222 277890 124256 277924
rect 124222 277822 124256 277856
rect 124222 277754 124256 277788
rect 124222 277686 124256 277720
rect 124222 277618 124256 277652
rect 124222 277550 124256 277584
rect 124222 277482 124256 277516
rect 124222 277414 124256 277448
rect 122392 276597 122426 276631
rect 122392 276529 122426 276563
rect 123844 276597 123878 276631
rect 123844 276529 123878 276563
rect 122479 275823 122513 275857
rect 122547 275823 122581 275857
rect 122615 275823 122649 275857
rect 122683 275823 122717 275857
rect 122751 275823 122785 275857
rect 122819 275823 122853 275857
rect 123115 275823 123149 275857
rect 123183 275823 123217 275857
rect 123251 275823 123285 275857
rect 123319 275823 123353 275857
rect 123387 275823 123421 275857
rect 123455 275823 123489 275857
rect 123751 275823 123785 275857
rect 123819 275823 123853 275857
rect 123887 275823 123921 275857
rect 123955 275823 123989 275857
rect 124023 275823 124057 275857
rect 124091 275823 124125 275857
rect 124387 275823 124421 275857
rect 124455 275823 124489 275857
rect 124523 275823 124557 275857
rect 124591 275823 124625 275857
rect 124659 275823 124693 275857
rect 124727 275823 124761 275857
rect 122479 275665 122513 275699
rect 122547 275665 122581 275699
rect 122615 275665 122649 275699
rect 122683 275665 122717 275699
rect 122751 275665 122785 275699
rect 122819 275665 122853 275699
rect 123115 275665 123149 275699
rect 123183 275665 123217 275699
rect 123251 275665 123285 275699
rect 123319 275665 123353 275699
rect 123387 275665 123421 275699
rect 123455 275665 123489 275699
rect 123751 275665 123785 275699
rect 123819 275665 123853 275699
rect 123887 275665 123921 275699
rect 123955 275665 123989 275699
rect 124023 275665 124057 275699
rect 124091 275665 124125 275699
rect 124387 275665 124421 275699
rect 124455 275665 124489 275699
rect 124523 275665 124557 275699
rect 124591 275665 124625 275699
rect 124659 275665 124693 275699
rect 124727 275665 124761 275699
rect 120383 274702 120417 274736
rect 120383 274634 120417 274668
rect 120383 274566 120417 274600
rect 120383 274498 120417 274532
rect 120383 274430 120417 274464
rect 120383 274362 120417 274396
rect 120383 274294 120417 274328
rect 120841 274702 120875 274736
rect 120841 274634 120875 274668
rect 120841 274566 120875 274600
rect 120841 274498 120875 274532
rect 120841 274430 120875 274464
rect 120841 274362 120875 274396
rect 120841 274294 120875 274328
rect 121083 274702 121117 274736
rect 121083 274634 121117 274668
rect 121083 274566 121117 274600
rect 121083 274498 121117 274532
rect 121083 274430 121117 274464
rect 121083 274362 121117 274396
rect 121083 274294 121117 274328
rect 121541 274702 121575 274736
rect 121541 274634 121575 274668
rect 121541 274566 121575 274600
rect 121541 274498 121575 274532
rect 121541 274430 121575 274464
rect 121541 274362 121575 274396
rect 121541 274294 121575 274328
rect 120383 273918 120417 273952
rect 120383 273850 120417 273884
rect 120383 273782 120417 273816
rect 120383 273714 120417 273748
rect 120383 273646 120417 273680
rect 120383 273578 120417 273612
rect 120383 273510 120417 273544
rect 120841 273918 120875 273952
rect 120841 273850 120875 273884
rect 120841 273782 120875 273816
rect 120841 273714 120875 273748
rect 120841 273646 120875 273680
rect 120841 273578 120875 273612
rect 120841 273510 120875 273544
rect 121083 273918 121117 273952
rect 121083 273850 121117 273884
rect 121083 273782 121117 273816
rect 121083 273714 121117 273748
rect 121083 273646 121117 273680
rect 121083 273578 121117 273612
rect 121083 273510 121117 273544
rect 121541 273918 121575 273952
rect 121541 273850 121575 273884
rect 121541 273782 121575 273816
rect 121541 273714 121575 273748
rect 121541 273646 121575 273680
rect 121541 273578 121575 273612
rect 121541 273510 121575 273544
rect 120383 273134 120417 273168
rect 120383 273066 120417 273100
rect 120383 272998 120417 273032
rect 120383 272930 120417 272964
rect 120383 272862 120417 272896
rect 120383 272794 120417 272828
rect 120383 272726 120417 272760
rect 120841 273134 120875 273168
rect 120841 273066 120875 273100
rect 120841 272998 120875 273032
rect 120841 272930 120875 272964
rect 120841 272862 120875 272896
rect 120841 272794 120875 272828
rect 120841 272726 120875 272760
rect 121083 273134 121117 273168
rect 121083 273066 121117 273100
rect 121083 272998 121117 273032
rect 121083 272930 121117 272964
rect 121083 272862 121117 272896
rect 121083 272794 121117 272828
rect 121083 272726 121117 272760
rect 121541 273134 121575 273168
rect 121541 273066 121575 273100
rect 121541 272998 121575 273032
rect 121541 272930 121575 272964
rect 121541 272862 121575 272896
rect 121541 272794 121575 272828
rect 121541 272726 121575 272760
rect 120383 272350 120417 272384
rect 120383 272282 120417 272316
rect 120383 272214 120417 272248
rect 120383 272146 120417 272180
rect 120383 272078 120417 272112
rect 120383 272010 120417 272044
rect 120383 271942 120417 271976
rect 120841 272350 120875 272384
rect 120841 272282 120875 272316
rect 120841 272214 120875 272248
rect 120841 272146 120875 272180
rect 120841 272078 120875 272112
rect 120841 272010 120875 272044
rect 120841 271942 120875 271976
rect 121083 272350 121117 272384
rect 121083 272282 121117 272316
rect 121083 272214 121117 272248
rect 121083 272146 121117 272180
rect 121083 272078 121117 272112
rect 121083 272010 121117 272044
rect 121083 271942 121117 271976
rect 121541 272350 121575 272384
rect 121541 272282 121575 272316
rect 121541 272214 121575 272248
rect 121541 272146 121575 272180
rect 121541 272078 121575 272112
rect 121541 272010 121575 272044
rect 121541 271942 121575 271976
rect 120383 271566 120417 271600
rect 120383 271498 120417 271532
rect 120383 271430 120417 271464
rect 120383 271362 120417 271396
rect 120383 271294 120417 271328
rect 120383 271226 120417 271260
rect 120383 271158 120417 271192
rect 120841 271566 120875 271600
rect 120841 271498 120875 271532
rect 120841 271430 120875 271464
rect 120841 271362 120875 271396
rect 120841 271294 120875 271328
rect 120841 271226 120875 271260
rect 120841 271158 120875 271192
rect 121083 271566 121117 271600
rect 121083 271498 121117 271532
rect 121083 271430 121117 271464
rect 121083 271362 121117 271396
rect 121083 271294 121117 271328
rect 121083 271226 121117 271260
rect 121083 271158 121117 271192
rect 121541 271566 121575 271600
rect 121541 271498 121575 271532
rect 121541 271430 121575 271464
rect 121541 271362 121575 271396
rect 121541 271294 121575 271328
rect 121541 271226 121575 271260
rect 121541 271158 121575 271192
rect 120383 270782 120417 270816
rect 120383 270714 120417 270748
rect 120383 270646 120417 270680
rect 120383 270578 120417 270612
rect 120383 270510 120417 270544
rect 120383 270442 120417 270476
rect 120383 270374 120417 270408
rect 120841 270782 120875 270816
rect 120841 270714 120875 270748
rect 120841 270646 120875 270680
rect 120841 270578 120875 270612
rect 120841 270510 120875 270544
rect 120841 270442 120875 270476
rect 120841 270374 120875 270408
rect 121083 270782 121117 270816
rect 121083 270714 121117 270748
rect 121083 270646 121117 270680
rect 121083 270578 121117 270612
rect 121083 270510 121117 270544
rect 121083 270442 121117 270476
rect 121083 270374 121117 270408
rect 121541 270782 121575 270816
rect 121541 270714 121575 270748
rect 121541 270646 121575 270680
rect 121541 270578 121575 270612
rect 121541 270510 121575 270544
rect 121541 270442 121575 270476
rect 121541 270374 121575 270408
rect 120383 269998 120417 270032
rect 120383 269930 120417 269964
rect 120383 269862 120417 269896
rect 120383 269794 120417 269828
rect 120383 269726 120417 269760
rect 120383 269658 120417 269692
rect 120383 269590 120417 269624
rect 120841 269998 120875 270032
rect 120841 269930 120875 269964
rect 120841 269862 120875 269896
rect 120841 269794 120875 269828
rect 120841 269726 120875 269760
rect 120841 269658 120875 269692
rect 120841 269590 120875 269624
rect 121083 269998 121117 270032
rect 121083 269930 121117 269964
rect 121083 269862 121117 269896
rect 121083 269794 121117 269828
rect 121083 269726 121117 269760
rect 121083 269658 121117 269692
rect 121083 269590 121117 269624
rect 121541 269998 121575 270032
rect 121541 269930 121575 269964
rect 121541 269862 121575 269896
rect 121541 269794 121575 269828
rect 121541 269726 121575 269760
rect 121541 269658 121575 269692
rect 121541 269590 121575 269624
rect 120383 269210 120417 269244
rect 120841 269210 120875 269244
rect 121083 269210 121117 269244
rect 121541 269210 121575 269244
rect 122079 272746 122113 272780
rect 122537 272746 122571 272780
rect 122779 272746 122813 272780
rect 123237 272746 123271 272780
rect 122079 272366 122113 272400
rect 122079 272298 122113 272332
rect 122079 272230 122113 272264
rect 122079 272162 122113 272196
rect 122079 272094 122113 272128
rect 122079 272026 122113 272060
rect 122079 271958 122113 271992
rect 122537 272366 122571 272400
rect 122537 272298 122571 272332
rect 122537 272230 122571 272264
rect 122537 272162 122571 272196
rect 122537 272094 122571 272128
rect 122537 272026 122571 272060
rect 122537 271958 122571 271992
rect 122779 272366 122813 272400
rect 122779 272298 122813 272332
rect 122779 272230 122813 272264
rect 122779 272162 122813 272196
rect 122779 272094 122813 272128
rect 122779 272026 122813 272060
rect 122779 271958 122813 271992
rect 123237 272366 123271 272400
rect 123237 272298 123271 272332
rect 123237 272230 123271 272264
rect 123237 272162 123271 272196
rect 123237 272094 123271 272128
rect 123237 272026 123271 272060
rect 123237 271958 123271 271992
rect 122079 271582 122113 271616
rect 122079 271514 122113 271548
rect 122079 271446 122113 271480
rect 122079 271378 122113 271412
rect 122079 271310 122113 271344
rect 122079 271242 122113 271276
rect 122079 271174 122113 271208
rect 122537 271582 122571 271616
rect 122537 271514 122571 271548
rect 122537 271446 122571 271480
rect 122537 271378 122571 271412
rect 122537 271310 122571 271344
rect 122537 271242 122571 271276
rect 122537 271174 122571 271208
rect 122779 271582 122813 271616
rect 122779 271514 122813 271548
rect 122779 271446 122813 271480
rect 122779 271378 122813 271412
rect 122779 271310 122813 271344
rect 122779 271242 122813 271276
rect 122779 271174 122813 271208
rect 123237 271582 123271 271616
rect 123237 271514 123271 271548
rect 123237 271446 123271 271480
rect 123237 271378 123271 271412
rect 123237 271310 123271 271344
rect 123237 271242 123271 271276
rect 123237 271174 123271 271208
rect 122079 270798 122113 270832
rect 122079 270730 122113 270764
rect 122079 270662 122113 270696
rect 122079 270594 122113 270628
rect 122079 270526 122113 270560
rect 122079 270458 122113 270492
rect 122079 270390 122113 270424
rect 122537 270798 122571 270832
rect 122537 270730 122571 270764
rect 122537 270662 122571 270696
rect 122537 270594 122571 270628
rect 122537 270526 122571 270560
rect 122537 270458 122571 270492
rect 122537 270390 122571 270424
rect 122779 270798 122813 270832
rect 122779 270730 122813 270764
rect 122779 270662 122813 270696
rect 122779 270594 122813 270628
rect 122779 270526 122813 270560
rect 122779 270458 122813 270492
rect 122779 270390 122813 270424
rect 123237 270798 123271 270832
rect 123237 270730 123271 270764
rect 123237 270662 123271 270696
rect 123237 270594 123271 270628
rect 123237 270526 123271 270560
rect 123237 270458 123271 270492
rect 123237 270390 123271 270424
rect 122079 270014 122113 270048
rect 122079 269946 122113 269980
rect 122079 269878 122113 269912
rect 122079 269810 122113 269844
rect 122079 269742 122113 269776
rect 122079 269674 122113 269708
rect 122079 269606 122113 269640
rect 122537 270014 122571 270048
rect 122537 269946 122571 269980
rect 122537 269878 122571 269912
rect 122537 269810 122571 269844
rect 122537 269742 122571 269776
rect 122537 269674 122571 269708
rect 122537 269606 122571 269640
rect 122779 270014 122813 270048
rect 122779 269946 122813 269980
rect 122779 269878 122813 269912
rect 122779 269810 122813 269844
rect 122779 269742 122813 269776
rect 122779 269674 122813 269708
rect 122779 269606 122813 269640
rect 123237 270014 123271 270048
rect 123237 269946 123271 269980
rect 123237 269878 123271 269912
rect 123237 269810 123271 269844
rect 123237 269742 123271 269776
rect 123237 269674 123271 269708
rect 123237 269606 123271 269640
rect 122079 269226 122113 269260
rect 122537 269226 122571 269260
rect 122779 269226 122813 269260
rect 123237 269226 123271 269260
<< psubdiff >>
rect 111046 281156 119159 281179
rect 111046 281122 111264 281156
rect 111298 281122 111332 281156
rect 111366 281122 111400 281156
rect 111434 281122 111468 281156
rect 111502 281122 111536 281156
rect 111570 281122 111604 281156
rect 111638 281122 111672 281156
rect 111706 281122 111740 281156
rect 111774 281122 111808 281156
rect 111842 281122 111876 281156
rect 111910 281122 111944 281156
rect 111978 281122 112012 281156
rect 112046 281122 112080 281156
rect 112114 281122 112148 281156
rect 112182 281122 112216 281156
rect 112250 281122 112284 281156
rect 112318 281122 112352 281156
rect 112386 281122 112420 281156
rect 112454 281122 112488 281156
rect 112522 281122 112556 281156
rect 112590 281122 112624 281156
rect 112658 281122 112692 281156
rect 112726 281122 112760 281156
rect 112794 281122 112828 281156
rect 112862 281122 112896 281156
rect 112930 281122 112964 281156
rect 112998 281122 113032 281156
rect 113066 281122 113100 281156
rect 113134 281122 113168 281156
rect 113202 281122 113236 281156
rect 113270 281122 113304 281156
rect 113338 281122 113372 281156
rect 113406 281122 113440 281156
rect 113474 281122 113508 281156
rect 113542 281122 113576 281156
rect 113610 281122 113644 281156
rect 113678 281122 113712 281156
rect 113746 281122 113780 281156
rect 113814 281122 113848 281156
rect 113882 281122 113916 281156
rect 113950 281122 113984 281156
rect 114018 281122 114052 281156
rect 114086 281122 114120 281156
rect 114154 281122 114188 281156
rect 114222 281122 114256 281156
rect 114290 281122 114324 281156
rect 114358 281122 114392 281156
rect 114426 281122 114460 281156
rect 114494 281122 114528 281156
rect 114562 281122 114596 281156
rect 114630 281122 114664 281156
rect 114698 281122 114732 281156
rect 114766 281122 114800 281156
rect 114834 281122 114868 281156
rect 114902 281122 114936 281156
rect 114970 281122 115004 281156
rect 115038 281122 115072 281156
rect 115106 281122 115140 281156
rect 115174 281122 115208 281156
rect 115242 281122 115276 281156
rect 115310 281122 115344 281156
rect 115378 281122 115412 281156
rect 115446 281122 115480 281156
rect 115514 281122 115548 281156
rect 115582 281122 115616 281156
rect 115650 281122 115684 281156
rect 115718 281122 115752 281156
rect 115786 281122 115820 281156
rect 115854 281122 115888 281156
rect 115922 281122 115956 281156
rect 115990 281122 116024 281156
rect 116058 281122 116092 281156
rect 116126 281122 116160 281156
rect 116194 281122 116228 281156
rect 116262 281122 116296 281156
rect 116330 281122 116364 281156
rect 116398 281122 116432 281156
rect 116466 281122 116500 281156
rect 116534 281122 116568 281156
rect 116602 281122 116636 281156
rect 116670 281122 116704 281156
rect 116738 281122 116772 281156
rect 116806 281122 116840 281156
rect 116874 281122 116908 281156
rect 116942 281122 116976 281156
rect 117010 281122 117044 281156
rect 117078 281122 117112 281156
rect 117146 281122 117180 281156
rect 117214 281122 117248 281156
rect 117282 281122 117316 281156
rect 117350 281122 117384 281156
rect 117418 281122 117452 281156
rect 117486 281122 117520 281156
rect 117554 281122 117588 281156
rect 117622 281122 117656 281156
rect 117690 281122 117724 281156
rect 117758 281122 117792 281156
rect 117826 281122 117860 281156
rect 117894 281122 117928 281156
rect 117962 281122 117996 281156
rect 118030 281122 118064 281156
rect 118098 281122 118132 281156
rect 118166 281122 118200 281156
rect 118234 281122 118268 281156
rect 118302 281122 118336 281156
rect 118370 281122 118404 281156
rect 118438 281122 118472 281156
rect 118506 281122 118540 281156
rect 118574 281122 118608 281156
rect 118642 281122 118676 281156
rect 118710 281122 118744 281156
rect 118778 281122 118812 281156
rect 118846 281122 119159 281156
rect 111046 281102 119159 281122
rect 105974 281045 106147 281065
rect 105974 281020 110313 281045
rect 105974 281017 106176 281020
rect 105974 280983 106000 281017
rect 106034 280986 106176 281017
rect 106210 280986 106244 281020
rect 106278 280986 106312 281020
rect 106346 280986 106380 281020
rect 106414 280986 106448 281020
rect 106482 280986 106516 281020
rect 106550 280986 106584 281020
rect 106618 280986 106652 281020
rect 106686 280986 106720 281020
rect 106754 280986 106788 281020
rect 106822 280986 106856 281020
rect 106890 280986 106924 281020
rect 106958 280986 106992 281020
rect 107026 280986 107060 281020
rect 107094 280986 107128 281020
rect 107162 280986 107196 281020
rect 107230 280986 107264 281020
rect 107298 280986 107332 281020
rect 107366 280986 107400 281020
rect 107434 280986 107468 281020
rect 107502 280986 107536 281020
rect 107570 280986 107604 281020
rect 107638 280986 107672 281020
rect 107706 280986 107740 281020
rect 107774 280986 107808 281020
rect 107842 280986 107876 281020
rect 107910 280986 107944 281020
rect 107978 280986 108012 281020
rect 108046 280986 108080 281020
rect 108114 280986 108148 281020
rect 108182 280986 108216 281020
rect 108250 280986 108284 281020
rect 108318 280986 108352 281020
rect 108386 280986 108420 281020
rect 108454 280986 108488 281020
rect 108522 280986 108556 281020
rect 108590 280986 108624 281020
rect 108658 280986 108692 281020
rect 108726 280986 108760 281020
rect 108794 280986 108828 281020
rect 108862 280986 108896 281020
rect 108930 280986 108964 281020
rect 108998 280986 109032 281020
rect 109066 280986 109100 281020
rect 109134 280986 109168 281020
rect 109202 280986 109236 281020
rect 109270 280986 109304 281020
rect 109338 280986 109372 281020
rect 109406 280986 109440 281020
rect 109474 280986 109508 281020
rect 109542 280986 109576 281020
rect 109610 280986 109644 281020
rect 109678 280986 109712 281020
rect 109746 280986 109780 281020
rect 109814 280986 109848 281020
rect 109882 280986 109916 281020
rect 109950 280986 109984 281020
rect 110018 280986 110052 281020
rect 110086 280986 110120 281020
rect 110154 280986 110188 281020
rect 110222 280986 110313 281020
rect 106034 280983 110313 280986
rect 105974 280961 110313 280983
rect 105974 280949 106207 280961
rect 105974 280915 106000 280949
rect 106034 280915 106207 280949
rect 105974 280881 106207 280915
rect 105974 280847 106000 280881
rect 106034 280859 106207 280881
rect 106034 280847 106149 280859
rect 105974 280825 106149 280847
rect 106183 280825 106207 280859
rect 105974 280813 106207 280825
rect 110231 280841 110313 280961
rect 105974 280779 106000 280813
rect 106034 280791 106207 280813
rect 106034 280779 106149 280791
rect 105974 280757 106149 280779
rect 106183 280757 106207 280791
rect 105974 280745 106207 280757
rect 105974 280711 106000 280745
rect 106034 280723 106207 280745
rect 106034 280711 106149 280723
rect 105974 280689 106149 280711
rect 106183 280689 106207 280723
rect 105974 280677 106207 280689
rect 105974 280643 106000 280677
rect 106034 280655 106207 280677
rect 106034 280643 106149 280655
rect 105974 280621 106149 280643
rect 106183 280621 106207 280655
rect 105974 280609 106207 280621
rect 105974 280575 106000 280609
rect 106034 280587 106207 280609
rect 106034 280575 106149 280587
rect 105974 280553 106149 280575
rect 106183 280553 106207 280587
rect 105974 280541 106207 280553
rect 105974 280507 106000 280541
rect 106034 280519 106207 280541
rect 106034 280507 106149 280519
rect 105974 280485 106149 280507
rect 106183 280485 106207 280519
rect 105974 280473 106207 280485
rect 105974 280439 106000 280473
rect 106034 280451 106207 280473
rect 106034 280439 106149 280451
rect 105974 280417 106149 280439
rect 106183 280417 106207 280451
rect 105974 280405 106207 280417
rect 105974 280371 106000 280405
rect 106034 280383 106207 280405
rect 106034 280371 106149 280383
rect 105974 280349 106149 280371
rect 106183 280349 106207 280383
rect 105974 280337 106207 280349
rect 105974 280303 106000 280337
rect 106034 280315 106207 280337
rect 106034 280303 106149 280315
rect 105974 280281 106149 280303
rect 106183 280281 106207 280315
rect 105974 280269 106207 280281
rect 105974 280235 106000 280269
rect 106034 280247 106207 280269
rect 106034 280235 106149 280247
rect 105974 280213 106149 280235
rect 106183 280213 106207 280247
rect 105974 280201 106207 280213
rect 105974 280167 106000 280201
rect 106034 280179 106207 280201
rect 106034 280167 106149 280179
rect 105974 280145 106149 280167
rect 106183 280145 106207 280179
rect 105974 280133 106207 280145
rect 105974 280099 106000 280133
rect 106034 280111 106207 280133
rect 106034 280099 106149 280111
rect 105974 280077 106149 280099
rect 106183 280077 106207 280111
rect 105974 280065 106207 280077
rect 105974 280031 106000 280065
rect 106034 280043 106207 280065
rect 106034 280031 106149 280043
rect 105974 280009 106149 280031
rect 106183 280009 106207 280043
rect 105974 279997 106207 280009
rect 105974 279963 106000 279997
rect 106034 279975 106207 279997
rect 106034 279963 106149 279975
rect 105974 279941 106149 279963
rect 106183 279941 106207 279975
rect 105974 279929 106207 279941
rect 105974 279895 106000 279929
rect 106034 279907 106207 279929
rect 106034 279895 106149 279907
rect 105974 279873 106149 279895
rect 106183 279873 106207 279907
rect 105974 279861 106207 279873
rect 105974 279827 106000 279861
rect 106034 279839 106207 279861
rect 106034 279827 106149 279839
rect 105974 279805 106149 279827
rect 106183 279805 106207 279839
rect 105974 279793 106207 279805
rect 110231 280807 110255 280841
rect 110289 280807 110313 280841
rect 110231 280773 110313 280807
rect 110231 280739 110255 280773
rect 110289 280739 110313 280773
rect 110231 280705 110313 280739
rect 110231 280671 110255 280705
rect 110289 280671 110313 280705
rect 110231 280637 110313 280671
rect 110231 280603 110255 280637
rect 110289 280603 110313 280637
rect 110231 280569 110313 280603
rect 110231 280535 110255 280569
rect 110289 280535 110313 280569
rect 110231 280501 110313 280535
rect 110231 280467 110255 280501
rect 110289 280467 110313 280501
rect 110231 280433 110313 280467
rect 110231 280399 110255 280433
rect 110289 280399 110313 280433
rect 110231 280365 110313 280399
rect 110231 280331 110255 280365
rect 110289 280331 110313 280365
rect 110231 280297 110313 280331
rect 110231 280263 110255 280297
rect 110289 280263 110313 280297
rect 110231 280229 110313 280263
rect 110231 280195 110255 280229
rect 110289 280195 110313 280229
rect 110231 280161 110313 280195
rect 110231 280127 110255 280161
rect 110289 280127 110313 280161
rect 110231 280093 110313 280127
rect 110231 280059 110255 280093
rect 110289 280059 110313 280093
rect 110231 280025 110313 280059
rect 110231 279991 110255 280025
rect 110289 279991 110313 280025
rect 110231 279957 110313 279991
rect 110231 279923 110255 279957
rect 110289 279923 110313 279957
rect 110231 279889 110313 279923
rect 110231 279855 110255 279889
rect 110289 279855 110313 279889
rect 110231 279821 110313 279855
rect 105974 279759 106000 279793
rect 106034 279771 106207 279793
rect 106034 279759 106149 279771
rect 105974 279737 106149 279759
rect 106183 279737 106207 279771
rect 105974 279725 106207 279737
rect 105974 279691 106000 279725
rect 106034 279691 106207 279725
rect 110231 279787 110255 279821
rect 110289 279787 110313 279821
rect 110231 279753 110313 279787
rect 110231 279719 110255 279753
rect 110289 279719 110313 279753
rect 105974 279657 106207 279691
rect 105974 279623 106000 279657
rect 106034 279625 106207 279657
rect 110231 279625 110313 279719
rect 106034 279623 110313 279625
rect 105974 279600 110313 279623
rect 105974 279589 106176 279600
rect 105974 279555 106000 279589
rect 106034 279566 106176 279589
rect 106210 279566 106244 279600
rect 106278 279566 106312 279600
rect 106346 279566 106380 279600
rect 106414 279566 106448 279600
rect 106482 279566 106516 279600
rect 106550 279566 106584 279600
rect 106618 279566 106652 279600
rect 106686 279566 106720 279600
rect 106754 279566 106788 279600
rect 106822 279566 106856 279600
rect 106890 279566 106924 279600
rect 106958 279566 106992 279600
rect 107026 279566 107060 279600
rect 107094 279566 107128 279600
rect 107162 279566 107196 279600
rect 107230 279566 107264 279600
rect 107298 279566 107332 279600
rect 107366 279566 107400 279600
rect 107434 279566 107468 279600
rect 107502 279566 107536 279600
rect 107570 279566 107604 279600
rect 107638 279566 107672 279600
rect 107706 279566 107740 279600
rect 107774 279566 107808 279600
rect 107842 279566 107876 279600
rect 107910 279566 107944 279600
rect 107978 279566 108012 279600
rect 108046 279566 108080 279600
rect 108114 279566 108148 279600
rect 108182 279566 108216 279600
rect 108250 279566 108284 279600
rect 108318 279566 108352 279600
rect 108386 279566 108420 279600
rect 108454 279566 108488 279600
rect 108522 279566 108556 279600
rect 108590 279566 108624 279600
rect 108658 279566 108692 279600
rect 108726 279566 108760 279600
rect 108794 279566 108828 279600
rect 108862 279566 108896 279600
rect 108930 279566 108964 279600
rect 108998 279566 109032 279600
rect 109066 279566 109100 279600
rect 109134 279566 109168 279600
rect 109202 279566 109236 279600
rect 109270 279566 109304 279600
rect 109338 279566 109372 279600
rect 109406 279566 109440 279600
rect 109474 279566 109508 279600
rect 109542 279566 109576 279600
rect 109610 279566 109644 279600
rect 109678 279566 109712 279600
rect 109746 279566 109780 279600
rect 109814 279566 109848 279600
rect 109882 279566 109916 279600
rect 109950 279566 109984 279600
rect 110018 279566 110052 279600
rect 110086 279566 110120 279600
rect 110154 279566 110188 279600
rect 110222 279566 110313 279600
rect 106034 279555 110313 279566
rect 105974 279541 110313 279555
rect 105974 279521 106060 279541
rect 105974 279487 106000 279521
rect 106034 279487 106060 279521
rect 105974 279453 106060 279487
rect 105974 279419 106000 279453
rect 106034 279419 106060 279453
rect 105974 279385 106060 279419
rect 105974 279351 106000 279385
rect 106034 279351 106060 279385
rect 105974 279317 106060 279351
rect 105974 279283 106000 279317
rect 106034 279283 106060 279317
rect 105974 279249 106060 279283
rect 105974 279215 106000 279249
rect 106034 279215 106060 279249
rect 105974 279181 106060 279215
rect 105974 279147 106000 279181
rect 106034 279147 106060 279181
rect 105974 279113 106060 279147
rect 105974 279079 106000 279113
rect 106034 279079 106060 279113
rect 105974 279045 106060 279079
rect 105974 279011 106000 279045
rect 106034 279011 106060 279045
rect 105974 278977 106060 279011
rect 105974 278943 106000 278977
rect 106034 278943 106060 278977
rect 105974 278909 106060 278943
rect 105974 278875 106000 278909
rect 106034 278875 106060 278909
rect 105974 278841 106060 278875
rect 105974 278807 106000 278841
rect 106034 278807 106060 278841
rect 105974 278773 106060 278807
rect 105974 278739 106000 278773
rect 106034 278739 106060 278773
rect 105974 278705 106060 278739
rect 105974 278671 106000 278705
rect 106034 278671 106060 278705
rect 105974 278637 106060 278671
rect 105974 278603 106000 278637
rect 106034 278603 106060 278637
rect 105974 278569 106060 278603
rect 105974 278535 106000 278569
rect 106034 278535 106060 278569
rect 105974 278501 106060 278535
rect 105974 278467 106000 278501
rect 106034 278467 106060 278501
rect 105974 278433 106060 278467
rect 105974 278399 106000 278433
rect 106034 278399 106060 278433
rect 105974 278365 106060 278399
rect 105974 278331 106000 278365
rect 106034 278331 106060 278365
rect 105974 278297 106060 278331
rect 105974 278263 106000 278297
rect 106034 278263 106060 278297
rect 105974 278229 106060 278263
rect 105974 278195 106000 278229
rect 106034 278195 106060 278229
rect 105974 278161 106060 278195
rect 105974 278127 106000 278161
rect 106034 278127 106060 278161
rect 105974 278093 106060 278127
rect 105974 278059 106000 278093
rect 106034 278059 106060 278093
rect 105974 278025 106060 278059
rect 105974 277991 106000 278025
rect 106034 277991 106060 278025
rect 105974 277957 106060 277991
rect 105974 277923 106000 277957
rect 106034 277923 106060 277957
rect 110053 279185 110187 279541
rect 109617 279151 109733 279185
rect 109767 279151 109801 279185
rect 109835 279151 109869 279185
rect 109903 279151 109937 279185
rect 109971 279151 110005 279185
rect 110039 279151 110073 279185
rect 110107 279151 110223 279185
rect 109617 279071 109651 279151
rect 109617 279003 109651 279037
rect 110189 279071 110223 279151
rect 109617 278935 109651 278969
rect 109617 278867 109651 278901
rect 109617 278799 109651 278833
rect 109617 278731 109651 278765
rect 109617 278663 109651 278697
rect 109617 278595 109651 278629
rect 109617 278527 109651 278561
rect 109617 278459 109651 278493
rect 109617 278391 109651 278425
rect 109617 278323 109651 278357
rect 109617 278255 109651 278289
rect 109617 278187 109651 278221
rect 109617 278119 109651 278153
rect 109617 278051 109651 278085
rect 109617 277983 109651 278017
rect 105974 277889 106060 277923
rect 105974 277855 106000 277889
rect 106034 277855 106060 277889
rect 105974 277821 106060 277855
rect 105974 277787 106000 277821
rect 106034 277787 106060 277821
rect 105974 277753 106060 277787
rect 105974 277719 106000 277753
rect 106034 277719 106060 277753
rect 105974 277685 106060 277719
rect 105974 277651 106000 277685
rect 106034 277651 106060 277685
rect 105974 277617 106060 277651
rect 105974 277583 106000 277617
rect 106034 277583 106060 277617
rect 105974 277549 106060 277583
rect 105974 277515 106000 277549
rect 106034 277515 106060 277549
rect 105974 277481 106060 277515
rect 105974 277447 106000 277481
rect 106034 277447 106060 277481
rect 105974 277413 106060 277447
rect 105974 277379 106000 277413
rect 106034 277379 106060 277413
rect 105974 277345 106060 277379
rect 105974 277311 106000 277345
rect 106034 277311 106060 277345
rect 110189 279003 110223 279037
rect 110189 278935 110223 278969
rect 110189 278867 110223 278901
rect 110189 278799 110223 278833
rect 110189 278731 110223 278765
rect 110189 278663 110223 278697
rect 110189 278595 110223 278629
rect 110189 278527 110223 278561
rect 110189 278459 110223 278493
rect 110189 278391 110223 278425
rect 110189 278323 110223 278357
rect 110189 278255 110223 278289
rect 110189 278187 110223 278221
rect 110189 278119 110223 278153
rect 110189 278051 110223 278085
rect 110189 277983 110223 278017
rect 109617 277915 109651 277949
rect 110189 277915 110223 277949
rect 109617 277847 109651 277881
rect 110189 277847 110223 277881
rect 109617 277779 109651 277813
rect 110189 277779 110223 277813
rect 109617 277711 109651 277745
rect 109617 277643 109651 277677
rect 109617 277575 109651 277609
rect 109617 277507 109651 277541
rect 109617 277439 109651 277473
rect 109617 277371 109651 277405
rect 105974 277277 106060 277311
rect 105974 277243 106000 277277
rect 106034 277243 106060 277277
rect 105974 277209 106060 277243
rect 105974 277175 106000 277209
rect 106034 277175 106060 277209
rect 105974 277141 106060 277175
rect 105974 277107 106000 277141
rect 106034 277107 106060 277141
rect 105974 277073 106060 277107
rect 105974 277039 106000 277073
rect 106034 277039 106060 277073
rect 105974 277005 106060 277039
rect 105974 276971 106000 277005
rect 106034 276971 106060 277005
rect 105974 276937 106060 276971
rect 105974 276903 106000 276937
rect 106034 276903 106060 276937
rect 109617 277303 109651 277337
rect 109617 277235 109651 277269
rect 109617 277167 109651 277201
rect 109617 277099 109651 277133
rect 109617 277031 109651 277065
rect 109617 276963 109651 276997
rect 105974 276869 106060 276903
rect 105974 276835 106000 276869
rect 106034 276835 106060 276869
rect 105974 276801 106060 276835
rect 105974 276767 106000 276801
rect 106034 276767 106060 276801
rect 105974 276733 106060 276767
rect 105974 276699 106000 276733
rect 106034 276699 106060 276733
rect 105974 276665 106060 276699
rect 105974 276631 106000 276665
rect 106034 276631 106060 276665
rect 105974 276597 106060 276631
rect 105974 276563 106000 276597
rect 106034 276563 106060 276597
rect 105974 276529 106060 276563
rect 109617 276895 109651 276929
rect 109617 276827 109651 276861
rect 109617 276759 109651 276793
rect 109617 276691 109651 276725
rect 110189 277711 110223 277745
rect 110189 277643 110223 277677
rect 110189 277575 110223 277609
rect 110189 277507 110223 277541
rect 110189 277439 110223 277473
rect 110189 277371 110223 277405
rect 110189 277303 110223 277337
rect 110189 277235 110223 277269
rect 110189 277167 110223 277201
rect 110189 277099 110223 277133
rect 110189 277031 110223 277065
rect 110189 276963 110223 276997
rect 110189 276895 110223 276929
rect 110189 276827 110223 276861
rect 110189 276759 110223 276793
rect 109617 276577 109651 276657
rect 110189 276691 110223 276725
rect 110189 276577 110223 276657
rect 109617 276543 109733 276577
rect 109767 276543 109801 276577
rect 109835 276543 109869 276577
rect 109903 276543 109937 276577
rect 109971 276543 110005 276577
rect 110039 276543 110073 276577
rect 110107 276548 110223 276577
rect 110107 276543 110224 276548
rect 105974 276495 106000 276529
rect 106034 276495 106060 276529
rect 105974 276461 106060 276495
rect 105974 276427 106000 276461
rect 106034 276427 106060 276461
rect 105974 276393 106060 276427
rect 105974 276359 106000 276393
rect 106034 276359 106060 276393
rect 105974 276325 106060 276359
rect 105974 276291 106000 276325
rect 106034 276291 106060 276325
rect 105974 276257 106060 276291
rect 105974 276223 106000 276257
rect 106034 276223 106060 276257
rect 105974 276189 106060 276223
rect 105974 276155 106000 276189
rect 106034 276155 106060 276189
rect 105974 276121 106060 276155
rect 105974 276087 106000 276121
rect 106034 276087 106060 276121
rect 105974 276053 106060 276087
rect 105974 276019 106000 276053
rect 106034 276019 106060 276053
rect 105974 275985 106060 276019
rect 105974 275951 106000 275985
rect 106034 275951 106060 275985
rect 105974 275917 106060 275951
rect 110145 276025 110224 276543
rect 110145 275991 110167 276025
rect 110201 275991 110224 276025
rect 110145 275957 110224 275991
rect 105974 275883 106000 275917
rect 106034 275883 106060 275917
rect 105974 275849 106060 275883
rect 105974 275815 106000 275849
rect 106034 275815 106060 275849
rect 105974 275781 106060 275815
rect 105974 275747 106000 275781
rect 106034 275747 106060 275781
rect 105974 275713 106060 275747
rect 105974 275679 106000 275713
rect 106034 275679 106060 275713
rect 105974 275645 106060 275679
rect 105974 275611 106000 275645
rect 106034 275611 106060 275645
rect 105974 275577 106060 275611
rect 105974 275543 106000 275577
rect 106034 275543 106060 275577
rect 105974 275509 106060 275543
rect 105974 275475 106000 275509
rect 106034 275475 106060 275509
rect 105974 275441 106060 275475
rect 105974 275407 106000 275441
rect 106034 275407 106060 275441
rect 105974 275373 106060 275407
rect 105974 275339 106000 275373
rect 106034 275339 106060 275373
rect 105974 275305 106060 275339
rect 105974 275271 106000 275305
rect 106034 275271 106060 275305
rect 105974 275237 106060 275271
rect 105974 275203 106000 275237
rect 106034 275203 106060 275237
rect 105974 275169 106060 275203
rect 105974 275135 106000 275169
rect 106034 275135 106060 275169
rect 105974 275101 106060 275135
rect 105974 275067 106000 275101
rect 106034 275067 106060 275101
rect 105974 275033 106060 275067
rect 105974 274999 106000 275033
rect 106034 274999 106060 275033
rect 105974 274965 106060 274999
rect 105974 274931 106000 274965
rect 106034 274931 106060 274965
rect 105974 274897 106060 274931
rect 105974 274863 106000 274897
rect 106034 274863 106060 274897
rect 105974 274829 106060 274863
rect 105974 274795 106000 274829
rect 106034 274795 106060 274829
rect 105974 274761 106060 274795
rect 105974 274727 106000 274761
rect 106034 274727 106060 274761
rect 105974 274693 106060 274727
rect 110145 275923 110167 275957
rect 110201 275923 110224 275957
rect 110145 275889 110224 275923
rect 110145 275855 110167 275889
rect 110201 275855 110224 275889
rect 110145 275821 110224 275855
rect 110145 275787 110167 275821
rect 110201 275787 110224 275821
rect 110145 275753 110224 275787
rect 110145 275719 110167 275753
rect 110201 275719 110224 275753
rect 110145 275685 110224 275719
rect 110145 275651 110167 275685
rect 110201 275651 110224 275685
rect 110145 275617 110224 275651
rect 110145 275583 110167 275617
rect 110201 275583 110224 275617
rect 110145 275549 110224 275583
rect 110145 275515 110167 275549
rect 110201 275515 110224 275549
rect 110145 275481 110224 275515
rect 110145 275447 110167 275481
rect 110201 275447 110224 275481
rect 110145 275413 110224 275447
rect 110145 275379 110167 275413
rect 110201 275379 110224 275413
rect 110145 275345 110224 275379
rect 110145 275311 110167 275345
rect 110201 275311 110224 275345
rect 110145 275277 110224 275311
rect 110145 275243 110167 275277
rect 110201 275243 110224 275277
rect 110145 275209 110224 275243
rect 110145 275175 110167 275209
rect 110201 275175 110224 275209
rect 110145 275141 110224 275175
rect 110145 275107 110167 275141
rect 110201 275107 110224 275141
rect 110145 275073 110224 275107
rect 110145 275039 110167 275073
rect 110201 275039 110224 275073
rect 110145 275005 110224 275039
rect 110145 274971 110167 275005
rect 110201 274971 110224 275005
rect 110145 274937 110224 274971
rect 110145 274903 110167 274937
rect 110201 274903 110224 274937
rect 110145 274869 110224 274903
rect 110145 274835 110167 274869
rect 110201 274835 110224 274869
rect 110145 274801 110224 274835
rect 110145 274767 110167 274801
rect 110201 274767 110224 274801
rect 110145 274733 110224 274767
rect 105974 274659 106000 274693
rect 106034 274659 106060 274693
rect 105974 274619 106060 274659
rect 110145 274699 110167 274733
rect 110201 274699 110224 274733
rect 110145 274619 110224 274699
rect 105974 274590 110224 274619
rect 105974 274556 106117 274590
rect 106151 274556 106185 274590
rect 106219 274556 106253 274590
rect 106287 274556 106321 274590
rect 106355 274556 106389 274590
rect 106423 274556 106457 274590
rect 106491 274556 106525 274590
rect 106559 274556 106593 274590
rect 106627 274556 106661 274590
rect 106695 274556 106729 274590
rect 106763 274556 106797 274590
rect 106831 274556 106865 274590
rect 106899 274556 106933 274590
rect 106967 274556 107001 274590
rect 107035 274556 107069 274590
rect 107103 274556 107137 274590
rect 107171 274556 107205 274590
rect 107239 274556 107273 274590
rect 107307 274556 107341 274590
rect 107375 274556 107409 274590
rect 107443 274556 107477 274590
rect 107511 274556 107545 274590
rect 107579 274556 107613 274590
rect 107647 274556 107681 274590
rect 107715 274556 107749 274590
rect 107783 274556 107817 274590
rect 107851 274556 107885 274590
rect 107919 274556 107953 274590
rect 107987 274556 108021 274590
rect 108055 274556 108089 274590
rect 108123 274556 108157 274590
rect 108191 274556 108225 274590
rect 108259 274556 108293 274590
rect 108327 274556 108361 274590
rect 108395 274556 108429 274590
rect 108463 274556 108497 274590
rect 108531 274556 108565 274590
rect 108599 274556 108633 274590
rect 108667 274556 108701 274590
rect 108735 274556 108769 274590
rect 108803 274556 108837 274590
rect 108871 274556 108905 274590
rect 108939 274556 108973 274590
rect 109007 274556 109041 274590
rect 109075 274556 109109 274590
rect 109143 274556 109177 274590
rect 109211 274556 109245 274590
rect 109279 274556 109313 274590
rect 109347 274556 109381 274590
rect 109415 274556 109449 274590
rect 109483 274556 109517 274590
rect 109551 274556 109585 274590
rect 109619 274556 109653 274590
rect 109687 274556 109721 274590
rect 109755 274556 109789 274590
rect 109823 274556 109857 274590
rect 109891 274556 109925 274590
rect 109959 274556 109993 274590
rect 110027 274556 110061 274590
rect 110095 274556 110129 274590
rect 110163 274556 110224 274590
rect 105974 274527 110224 274556
rect 106281 272923 110259 272951
rect 106281 272898 106595 272923
rect 106281 270212 106285 272898
rect 106455 272821 106595 272898
rect 109961 272898 110259 272923
rect 109961 272821 110085 272898
rect 106455 272786 110085 272821
rect 106455 270334 106459 272786
rect 106715 272350 108803 272367
rect 106715 272321 106848 272350
rect 106715 272287 106735 272321
rect 106769 272316 106848 272321
rect 106882 272316 106977 272350
rect 107011 272316 107045 272350
rect 107079 272316 107113 272350
rect 107147 272316 107181 272350
rect 107215 272316 107249 272350
rect 107283 272316 107317 272350
rect 107351 272316 107385 272350
rect 107419 272316 107453 272350
rect 107487 272316 107521 272350
rect 107555 272316 107589 272350
rect 107623 272316 107657 272350
rect 107691 272316 107725 272350
rect 107759 272316 107793 272350
rect 107827 272316 107861 272350
rect 107895 272316 107929 272350
rect 107963 272316 107997 272350
rect 108031 272316 108065 272350
rect 108099 272316 108133 272350
rect 108167 272316 108201 272350
rect 108235 272316 108269 272350
rect 108303 272316 108337 272350
rect 108371 272316 108405 272350
rect 108439 272316 108473 272350
rect 108507 272316 108541 272350
rect 108575 272316 108609 272350
rect 108643 272321 108803 272350
rect 108643 272316 108749 272321
rect 106769 272299 108749 272316
rect 106769 272287 106789 272299
rect 106715 272253 106789 272287
rect 106715 272219 106735 272253
rect 106769 272219 106789 272253
rect 106715 272185 106789 272219
rect 106715 272151 106735 272185
rect 106769 272151 106789 272185
rect 108729 272287 108749 272299
rect 108783 272287 108803 272321
rect 108729 272253 108803 272287
rect 108729 272219 108749 272253
rect 108783 272219 108803 272253
rect 108729 272185 108803 272219
rect 106715 272117 106789 272151
rect 106715 272083 106735 272117
rect 106769 272083 106789 272117
rect 106715 272049 106789 272083
rect 108729 272151 108749 272185
rect 108783 272151 108803 272185
rect 108729 272117 108803 272151
rect 108729 272083 108749 272117
rect 108783 272083 108803 272117
rect 106715 272015 106735 272049
rect 106769 272015 106789 272049
rect 106715 271981 106789 272015
rect 106715 271947 106735 271981
rect 106769 271947 106789 271981
rect 106715 271913 106789 271947
rect 106715 271879 106735 271913
rect 106769 271879 106789 271913
rect 106715 271845 106789 271879
rect 106715 271811 106735 271845
rect 106769 271811 106789 271845
rect 106715 271777 106789 271811
rect 106715 271743 106735 271777
rect 106769 271743 106789 271777
rect 106715 271709 106789 271743
rect 108729 272049 108803 272083
rect 108729 272015 108749 272049
rect 108783 272015 108803 272049
rect 108729 271981 108803 272015
rect 108729 271947 108749 271981
rect 108783 271947 108803 271981
rect 108729 271913 108803 271947
rect 108729 271879 108749 271913
rect 108783 271879 108803 271913
rect 108729 271845 108803 271879
rect 108729 271811 108749 271845
rect 108783 271811 108803 271845
rect 108729 271777 108803 271811
rect 108729 271743 108749 271777
rect 108783 271743 108803 271777
rect 106715 271675 106735 271709
rect 106769 271675 106789 271709
rect 106715 271641 106789 271675
rect 108729 271709 108803 271743
rect 108729 271675 108749 271709
rect 108783 271675 108803 271709
rect 106715 271607 106735 271641
rect 106769 271607 106789 271641
rect 106715 271573 106789 271607
rect 106715 271539 106735 271573
rect 106769 271539 106789 271573
rect 108729 271641 108803 271675
rect 108729 271607 108749 271641
rect 108783 271607 108803 271641
rect 108729 271573 108803 271607
rect 106715 271505 106789 271539
rect 106715 271471 106735 271505
rect 106769 271471 106789 271505
rect 108729 271539 108749 271573
rect 108783 271539 108803 271573
rect 108729 271505 108803 271539
rect 106715 271437 106789 271471
rect 106715 271403 106735 271437
rect 106769 271403 106789 271437
rect 106715 271369 106789 271403
rect 106715 271335 106735 271369
rect 106769 271335 106789 271369
rect 106715 271301 106789 271335
rect 108729 271471 108749 271505
rect 108783 271471 108803 271505
rect 108729 271437 108803 271471
rect 108729 271403 108749 271437
rect 108783 271403 108803 271437
rect 108729 271369 108803 271403
rect 108729 271335 108749 271369
rect 108783 271335 108803 271369
rect 106715 271267 106735 271301
rect 106769 271267 106789 271301
rect 106715 271233 106789 271267
rect 108729 271301 108803 271335
rect 108729 271267 108749 271301
rect 108783 271267 108803 271301
rect 106715 271199 106735 271233
rect 106769 271199 106789 271233
rect 106715 271165 106789 271199
rect 108729 271233 108803 271267
rect 108729 271199 108749 271233
rect 108783 271199 108803 271233
rect 106715 271131 106735 271165
rect 106769 271131 106789 271165
rect 106715 271097 106789 271131
rect 108729 271165 108803 271199
rect 108729 271131 108749 271165
rect 108783 271131 108803 271165
rect 106715 271063 106735 271097
rect 106769 271063 106789 271097
rect 106715 271029 106789 271063
rect 106715 270995 106735 271029
rect 106769 270995 106789 271029
rect 106715 270961 106789 270995
rect 106715 270927 106735 270961
rect 106769 270927 106789 270961
rect 108729 271097 108803 271131
rect 108729 271063 108749 271097
rect 108783 271063 108803 271097
rect 108729 271029 108803 271063
rect 108729 270995 108749 271029
rect 108783 270995 108803 271029
rect 108729 270961 108803 270995
rect 106715 270893 106789 270927
rect 106715 270859 106735 270893
rect 106769 270859 106789 270893
rect 108729 270927 108749 270961
rect 108783 270927 108803 270961
rect 108729 270893 108803 270927
rect 106715 270825 106789 270859
rect 106715 270791 106735 270825
rect 106769 270801 106789 270825
rect 108729 270859 108749 270893
rect 108783 270859 108803 270893
rect 108729 270825 108803 270859
rect 108729 270801 108749 270825
rect 106769 270791 108749 270801
rect 108783 270791 108803 270825
rect 106715 270784 108803 270791
rect 106715 270750 106875 270784
rect 106909 270750 106943 270784
rect 106977 270750 107011 270784
rect 107045 270750 107079 270784
rect 107113 270750 107147 270784
rect 107181 270750 107215 270784
rect 107249 270750 107283 270784
rect 107317 270750 107351 270784
rect 107385 270750 107419 270784
rect 107453 270750 107487 270784
rect 107521 270750 107555 270784
rect 107589 270750 107623 270784
rect 107657 270750 107691 270784
rect 107725 270750 107759 270784
rect 107793 270750 107827 270784
rect 107861 270750 107895 270784
rect 107929 270750 107963 270784
rect 107997 270750 108031 270784
rect 108065 270750 108099 270784
rect 108133 270750 108167 270784
rect 108201 270750 108235 270784
rect 108269 270750 108303 270784
rect 108337 270750 108371 270784
rect 108405 270750 108439 270784
rect 108473 270750 108507 270784
rect 108541 270750 108575 270784
rect 108609 270750 108643 270784
rect 108677 270750 108803 270784
rect 106715 270733 108803 270750
rect 110081 270334 110085 272786
rect 106455 270306 110085 270334
rect 106455 270212 106585 270306
rect 106281 270204 106585 270212
rect 109951 270212 110085 270306
rect 110255 270212 110259 272898
rect 111046 272704 111072 281102
rect 111174 281099 119031 281102
rect 111174 279425 111200 281099
rect 114235 280876 114353 280908
rect 114235 280774 114243 280876
rect 114345 280774 114353 280876
rect 114235 280742 114353 280774
rect 111174 279397 114266 279425
rect 111174 279363 111340 279397
rect 111374 279363 111408 279397
rect 111442 279363 111476 279397
rect 111510 279363 111544 279397
rect 111578 279363 111612 279397
rect 111646 279363 111680 279397
rect 111714 279363 111748 279397
rect 111782 279363 111816 279397
rect 111850 279363 111884 279397
rect 111918 279363 111952 279397
rect 111986 279363 112020 279397
rect 112054 279363 112088 279397
rect 112122 279363 112156 279397
rect 112190 279363 112224 279397
rect 112258 279363 112292 279397
rect 112326 279363 112360 279397
rect 112394 279363 112428 279397
rect 112462 279363 112496 279397
rect 112530 279363 112564 279397
rect 112598 279363 112632 279397
rect 112666 279363 112700 279397
rect 112734 279363 112768 279397
rect 112802 279363 112836 279397
rect 112870 279363 112904 279397
rect 112938 279363 112972 279397
rect 113006 279363 113040 279397
rect 113074 279363 113108 279397
rect 113142 279363 113176 279397
rect 113210 279363 113244 279397
rect 113278 279363 113312 279397
rect 113346 279363 113380 279397
rect 113414 279363 113448 279397
rect 113482 279363 113516 279397
rect 113550 279363 113584 279397
rect 113618 279363 113652 279397
rect 113686 279363 113720 279397
rect 113754 279363 113788 279397
rect 113822 279363 113856 279397
rect 113890 279363 113924 279397
rect 113958 279363 113992 279397
rect 114026 279363 114060 279397
rect 114094 279363 114128 279397
rect 114162 279363 114196 279397
rect 114230 279363 114266 279397
rect 115852 280876 115970 280908
rect 115852 280774 115860 280876
rect 115962 280774 115970 280876
rect 115852 280742 115970 280774
rect 119005 279425 119031 281099
rect 115939 279397 119031 279425
rect 111174 279335 114266 279363
rect 115939 279363 115975 279397
rect 116009 279363 116043 279397
rect 116077 279363 116111 279397
rect 116145 279363 116179 279397
rect 116213 279363 116247 279397
rect 116281 279363 116315 279397
rect 116349 279363 116383 279397
rect 116417 279363 116451 279397
rect 116485 279363 116519 279397
rect 116553 279363 116587 279397
rect 116621 279363 116655 279397
rect 116689 279363 116723 279397
rect 116757 279363 116791 279397
rect 116825 279363 116859 279397
rect 116893 279363 116927 279397
rect 116961 279363 116995 279397
rect 117029 279363 117063 279397
rect 117097 279363 117131 279397
rect 117165 279363 117199 279397
rect 117233 279363 117267 279397
rect 117301 279363 117335 279397
rect 117369 279363 117403 279397
rect 117437 279363 117471 279397
rect 117505 279363 117539 279397
rect 117573 279363 117607 279397
rect 117641 279363 117675 279397
rect 117709 279363 117743 279397
rect 117777 279363 117811 279397
rect 117845 279363 117879 279397
rect 117913 279363 117947 279397
rect 117981 279363 118015 279397
rect 118049 279363 118083 279397
rect 118117 279363 118151 279397
rect 118185 279363 118219 279397
rect 118253 279363 118287 279397
rect 118321 279363 118355 279397
rect 118389 279363 118423 279397
rect 118457 279363 118491 279397
rect 118525 279363 118559 279397
rect 118593 279363 118627 279397
rect 118661 279363 118695 279397
rect 118729 279363 118763 279397
rect 118797 279363 118831 279397
rect 118865 279363 119031 279397
rect 115939 279335 119031 279363
rect 111174 277759 111200 279335
rect 114235 279210 114353 279242
rect 114235 279108 114243 279210
rect 114345 279108 114353 279210
rect 114235 279076 114353 279108
rect 111174 277731 114266 277759
rect 111174 277697 111340 277731
rect 111374 277697 111408 277731
rect 111442 277697 111476 277731
rect 111510 277697 111544 277731
rect 111578 277697 111612 277731
rect 111646 277697 111680 277731
rect 111714 277697 111748 277731
rect 111782 277697 111816 277731
rect 111850 277697 111884 277731
rect 111918 277697 111952 277731
rect 111986 277697 112020 277731
rect 112054 277697 112088 277731
rect 112122 277697 112156 277731
rect 112190 277697 112224 277731
rect 112258 277697 112292 277731
rect 112326 277697 112360 277731
rect 112394 277697 112428 277731
rect 112462 277697 112496 277731
rect 112530 277697 112564 277731
rect 112598 277697 112632 277731
rect 112666 277697 112700 277731
rect 112734 277697 112768 277731
rect 112802 277697 112836 277731
rect 112870 277697 112904 277731
rect 112938 277697 112972 277731
rect 113006 277697 113040 277731
rect 113074 277697 113108 277731
rect 113142 277697 113176 277731
rect 113210 277697 113244 277731
rect 113278 277697 113312 277731
rect 113346 277697 113380 277731
rect 113414 277697 113448 277731
rect 113482 277697 113516 277731
rect 113550 277697 113584 277731
rect 113618 277697 113652 277731
rect 113686 277697 113720 277731
rect 113754 277697 113788 277731
rect 113822 277697 113856 277731
rect 113890 277697 113924 277731
rect 113958 277697 113992 277731
rect 114026 277697 114060 277731
rect 114094 277697 114128 277731
rect 114162 277697 114196 277731
rect 114230 277697 114266 277731
rect 115852 279210 115970 279242
rect 115852 279108 115860 279210
rect 115962 279108 115970 279210
rect 115852 279076 115970 279108
rect 119005 277759 119031 279335
rect 115939 277731 119031 277759
rect 111174 277669 114266 277697
rect 115939 277697 115975 277731
rect 116009 277697 116043 277731
rect 116077 277697 116111 277731
rect 116145 277697 116179 277731
rect 116213 277697 116247 277731
rect 116281 277697 116315 277731
rect 116349 277697 116383 277731
rect 116417 277697 116451 277731
rect 116485 277697 116519 277731
rect 116553 277697 116587 277731
rect 116621 277697 116655 277731
rect 116689 277697 116723 277731
rect 116757 277697 116791 277731
rect 116825 277697 116859 277731
rect 116893 277697 116927 277731
rect 116961 277697 116995 277731
rect 117029 277697 117063 277731
rect 117097 277697 117131 277731
rect 117165 277697 117199 277731
rect 117233 277697 117267 277731
rect 117301 277697 117335 277731
rect 117369 277697 117403 277731
rect 117437 277697 117471 277731
rect 117505 277697 117539 277731
rect 117573 277697 117607 277731
rect 117641 277697 117675 277731
rect 117709 277697 117743 277731
rect 117777 277697 117811 277731
rect 117845 277697 117879 277731
rect 117913 277697 117947 277731
rect 117981 277697 118015 277731
rect 118049 277697 118083 277731
rect 118117 277697 118151 277731
rect 118185 277697 118219 277731
rect 118253 277697 118287 277731
rect 118321 277697 118355 277731
rect 118389 277697 118423 277731
rect 118457 277697 118491 277731
rect 118525 277697 118559 277731
rect 118593 277697 118627 277731
rect 118661 277697 118695 277731
rect 118729 277697 118763 277731
rect 118797 277697 118831 277731
rect 118865 277697 119031 277731
rect 115939 277669 119031 277697
rect 111174 276093 111200 277669
rect 114235 277544 114353 277576
rect 114235 277442 114243 277544
rect 114345 277442 114353 277544
rect 114235 277410 114353 277442
rect 111174 276065 114266 276093
rect 111174 276031 111340 276065
rect 111374 276031 111408 276065
rect 111442 276031 111476 276065
rect 111510 276031 111544 276065
rect 111578 276031 111612 276065
rect 111646 276031 111680 276065
rect 111714 276031 111748 276065
rect 111782 276031 111816 276065
rect 111850 276031 111884 276065
rect 111918 276031 111952 276065
rect 111986 276031 112020 276065
rect 112054 276031 112088 276065
rect 112122 276031 112156 276065
rect 112190 276031 112224 276065
rect 112258 276031 112292 276065
rect 112326 276031 112360 276065
rect 112394 276031 112428 276065
rect 112462 276031 112496 276065
rect 112530 276031 112564 276065
rect 112598 276031 112632 276065
rect 112666 276031 112700 276065
rect 112734 276031 112768 276065
rect 112802 276031 112836 276065
rect 112870 276031 112904 276065
rect 112938 276031 112972 276065
rect 113006 276031 113040 276065
rect 113074 276031 113108 276065
rect 113142 276031 113176 276065
rect 113210 276031 113244 276065
rect 113278 276031 113312 276065
rect 113346 276031 113380 276065
rect 113414 276031 113448 276065
rect 113482 276031 113516 276065
rect 113550 276031 113584 276065
rect 113618 276031 113652 276065
rect 113686 276031 113720 276065
rect 113754 276031 113788 276065
rect 113822 276031 113856 276065
rect 113890 276031 113924 276065
rect 113958 276031 113992 276065
rect 114026 276031 114060 276065
rect 114094 276031 114128 276065
rect 114162 276031 114196 276065
rect 114230 276031 114266 276065
rect 115852 277544 115970 277576
rect 115852 277442 115860 277544
rect 115962 277442 115970 277544
rect 115852 277410 115970 277442
rect 119005 276093 119031 277669
rect 115939 276065 119031 276093
rect 111174 276003 114266 276031
rect 115939 276031 115975 276065
rect 116009 276031 116043 276065
rect 116077 276031 116111 276065
rect 116145 276031 116179 276065
rect 116213 276031 116247 276065
rect 116281 276031 116315 276065
rect 116349 276031 116383 276065
rect 116417 276031 116451 276065
rect 116485 276031 116519 276065
rect 116553 276031 116587 276065
rect 116621 276031 116655 276065
rect 116689 276031 116723 276065
rect 116757 276031 116791 276065
rect 116825 276031 116859 276065
rect 116893 276031 116927 276065
rect 116961 276031 116995 276065
rect 117029 276031 117063 276065
rect 117097 276031 117131 276065
rect 117165 276031 117199 276065
rect 117233 276031 117267 276065
rect 117301 276031 117335 276065
rect 117369 276031 117403 276065
rect 117437 276031 117471 276065
rect 117505 276031 117539 276065
rect 117573 276031 117607 276065
rect 117641 276031 117675 276065
rect 117709 276031 117743 276065
rect 117777 276031 117811 276065
rect 117845 276031 117879 276065
rect 117913 276031 117947 276065
rect 117981 276031 118015 276065
rect 118049 276031 118083 276065
rect 118117 276031 118151 276065
rect 118185 276031 118219 276065
rect 118253 276031 118287 276065
rect 118321 276031 118355 276065
rect 118389 276031 118423 276065
rect 118457 276031 118491 276065
rect 118525 276031 118559 276065
rect 118593 276031 118627 276065
rect 118661 276031 118695 276065
rect 118729 276031 118763 276065
rect 118797 276031 118831 276065
rect 118865 276031 119031 276065
rect 115939 276003 119031 276031
rect 111174 274427 111200 276003
rect 114235 275878 114353 275910
rect 114235 275776 114243 275878
rect 114345 275776 114353 275878
rect 114235 275744 114353 275776
rect 111174 274399 114266 274427
rect 111174 274365 111340 274399
rect 111374 274365 111408 274399
rect 111442 274365 111476 274399
rect 111510 274365 111544 274399
rect 111578 274365 111612 274399
rect 111646 274365 111680 274399
rect 111714 274365 111748 274399
rect 111782 274365 111816 274399
rect 111850 274365 111884 274399
rect 111918 274365 111952 274399
rect 111986 274365 112020 274399
rect 112054 274365 112088 274399
rect 112122 274365 112156 274399
rect 112190 274365 112224 274399
rect 112258 274365 112292 274399
rect 112326 274365 112360 274399
rect 112394 274365 112428 274399
rect 112462 274365 112496 274399
rect 112530 274365 112564 274399
rect 112598 274365 112632 274399
rect 112666 274365 112700 274399
rect 112734 274365 112768 274399
rect 112802 274365 112836 274399
rect 112870 274365 112904 274399
rect 112938 274365 112972 274399
rect 113006 274365 113040 274399
rect 113074 274365 113108 274399
rect 113142 274365 113176 274399
rect 113210 274365 113244 274399
rect 113278 274365 113312 274399
rect 113346 274365 113380 274399
rect 113414 274365 113448 274399
rect 113482 274365 113516 274399
rect 113550 274365 113584 274399
rect 113618 274365 113652 274399
rect 113686 274365 113720 274399
rect 113754 274365 113788 274399
rect 113822 274365 113856 274399
rect 113890 274365 113924 274399
rect 113958 274365 113992 274399
rect 114026 274365 114060 274399
rect 114094 274365 114128 274399
rect 114162 274365 114196 274399
rect 114230 274365 114266 274399
rect 115852 275878 115970 275910
rect 115852 275776 115860 275878
rect 115962 275776 115970 275878
rect 115852 275744 115970 275776
rect 119005 274427 119031 276003
rect 115939 274399 119031 274427
rect 111174 274337 114266 274365
rect 115939 274365 115975 274399
rect 116009 274365 116043 274399
rect 116077 274365 116111 274399
rect 116145 274365 116179 274399
rect 116213 274365 116247 274399
rect 116281 274365 116315 274399
rect 116349 274365 116383 274399
rect 116417 274365 116451 274399
rect 116485 274365 116519 274399
rect 116553 274365 116587 274399
rect 116621 274365 116655 274399
rect 116689 274365 116723 274399
rect 116757 274365 116791 274399
rect 116825 274365 116859 274399
rect 116893 274365 116927 274399
rect 116961 274365 116995 274399
rect 117029 274365 117063 274399
rect 117097 274365 117131 274399
rect 117165 274365 117199 274399
rect 117233 274365 117267 274399
rect 117301 274365 117335 274399
rect 117369 274365 117403 274399
rect 117437 274365 117471 274399
rect 117505 274365 117539 274399
rect 117573 274365 117607 274399
rect 117641 274365 117675 274399
rect 117709 274365 117743 274399
rect 117777 274365 117811 274399
rect 117845 274365 117879 274399
rect 117913 274365 117947 274399
rect 117981 274365 118015 274399
rect 118049 274365 118083 274399
rect 118117 274365 118151 274399
rect 118185 274365 118219 274399
rect 118253 274365 118287 274399
rect 118321 274365 118355 274399
rect 118389 274365 118423 274399
rect 118457 274365 118491 274399
rect 118525 274365 118559 274399
rect 118593 274365 118627 274399
rect 118661 274365 118695 274399
rect 118729 274365 118763 274399
rect 118797 274365 118831 274399
rect 118865 274365 119031 274399
rect 115939 274337 119031 274365
rect 111174 272761 111200 274337
rect 114235 274212 114353 274244
rect 114235 274110 114243 274212
rect 114345 274110 114353 274212
rect 114235 274078 114353 274110
rect 114143 272761 114266 272766
rect 111174 272733 114266 272761
rect 111174 272704 111340 272733
rect 111046 272699 111340 272704
rect 111374 272699 111408 272733
rect 111442 272699 111476 272733
rect 111510 272699 111544 272733
rect 111578 272699 111612 272733
rect 111646 272699 111680 272733
rect 111714 272699 111748 272733
rect 111782 272699 111816 272733
rect 111850 272699 111884 272733
rect 111918 272699 111952 272733
rect 111986 272699 112020 272733
rect 112054 272699 112088 272733
rect 112122 272699 112156 272733
rect 112190 272699 112224 272733
rect 112258 272699 112292 272733
rect 112326 272699 112360 272733
rect 112394 272699 112428 272733
rect 112462 272699 112496 272733
rect 112530 272699 112564 272733
rect 112598 272699 112632 272733
rect 112666 272699 112700 272733
rect 112734 272699 112768 272733
rect 112802 272699 112836 272733
rect 112870 272699 112904 272733
rect 112938 272699 112972 272733
rect 113006 272699 113040 272733
rect 113074 272699 113108 272733
rect 113142 272699 113176 272733
rect 113210 272699 113244 272733
rect 113278 272699 113312 272733
rect 113346 272699 113380 272733
rect 113414 272699 113448 272733
rect 113482 272699 113516 272733
rect 113550 272699 113584 272733
rect 113618 272699 113652 272733
rect 113686 272699 113720 272733
rect 113754 272699 113788 272733
rect 113822 272699 113856 272733
rect 113890 272699 113924 272733
rect 113958 272699 113992 272733
rect 114026 272699 114060 272733
rect 114094 272699 114128 272733
rect 114162 272699 114196 272733
rect 114230 272699 114266 272733
rect 115852 274212 115970 274244
rect 115852 274110 115860 274212
rect 115962 274110 115970 274212
rect 115852 274078 115970 274110
rect 115939 272761 116062 272766
rect 119005 272761 119031 274337
rect 115939 272733 119031 272761
rect 111046 272671 114266 272699
rect 114143 272551 114266 272671
rect 115939 272699 115975 272733
rect 116009 272699 116043 272733
rect 116077 272699 116111 272733
rect 116145 272699 116179 272733
rect 116213 272699 116247 272733
rect 116281 272699 116315 272733
rect 116349 272699 116383 272733
rect 116417 272699 116451 272733
rect 116485 272699 116519 272733
rect 116553 272699 116587 272733
rect 116621 272699 116655 272733
rect 116689 272699 116723 272733
rect 116757 272699 116791 272733
rect 116825 272699 116859 272733
rect 116893 272699 116927 272733
rect 116961 272699 116995 272733
rect 117029 272699 117063 272733
rect 117097 272699 117131 272733
rect 117165 272699 117199 272733
rect 117233 272699 117267 272733
rect 117301 272699 117335 272733
rect 117369 272699 117403 272733
rect 117437 272699 117471 272733
rect 117505 272699 117539 272733
rect 117573 272699 117607 272733
rect 117641 272699 117675 272733
rect 117709 272699 117743 272733
rect 117777 272699 117811 272733
rect 117845 272699 117879 272733
rect 117913 272699 117947 272733
rect 117981 272699 118015 272733
rect 118049 272699 118083 272733
rect 118117 272699 118151 272733
rect 118185 272699 118219 272733
rect 118253 272699 118287 272733
rect 118321 272699 118355 272733
rect 118389 272699 118423 272733
rect 118457 272699 118491 272733
rect 118525 272699 118559 272733
rect 118593 272699 118627 272733
rect 118661 272699 118695 272733
rect 118729 272699 118763 272733
rect 118797 272699 118831 272733
rect 118865 272704 119031 272733
rect 119133 272704 119159 281102
rect 118865 272699 119159 272704
rect 115939 272671 119159 272699
rect 119938 281139 125172 281165
rect 119938 281059 120256 281139
rect 115939 272551 116062 272671
rect 114143 272460 116062 272551
rect 109951 270204 110259 270212
rect 106281 270169 110259 270204
rect 111939 272249 112069 272273
rect 119021 272249 119151 272273
rect 111939 272247 119151 272249
rect 111939 268677 111953 272247
rect 112055 272238 119035 272247
rect 112055 272136 112178 272238
rect 118944 272136 119035 272238
rect 112055 272125 119035 272136
rect 112055 268826 112069 272125
rect 119021 268826 119035 272125
rect 112055 268815 119035 268826
rect 112055 268713 112171 268815
rect 118937 268713 119035 268815
rect 112055 268702 119035 268713
rect 112055 268677 112069 268702
rect 111939 268651 112069 268677
rect 119021 268677 119035 268702
rect 119137 268677 119151 272247
rect 119938 268785 119970 281059
rect 120072 281037 120256 281059
rect 125118 281037 125172 281139
rect 120072 281012 125172 281037
rect 120072 268861 120104 281012
rect 125047 280856 125171 281012
rect 122027 278588 122144 278643
rect 122027 275562 122034 278588
rect 122136 276212 122144 278588
rect 122136 276205 124321 276212
rect 122136 276103 122531 276205
rect 124265 276103 124321 276205
rect 122136 276097 124321 276103
rect 122136 275562 122144 276097
rect 122027 275507 122144 275562
rect 122792 275002 122891 275036
rect 122925 275002 122959 275036
rect 122993 275002 123027 275036
rect 123061 275002 123095 275036
rect 123129 275002 123163 275036
rect 123197 275002 123231 275036
rect 123265 275002 123299 275036
rect 123333 275002 123367 275036
rect 123401 275002 123435 275036
rect 123469 275002 123503 275036
rect 123537 275002 123571 275036
rect 123605 275002 123639 275036
rect 123673 275002 123707 275036
rect 123741 275002 123775 275036
rect 123809 275002 123843 275036
rect 123877 275002 123911 275036
rect 123945 275002 123979 275036
rect 124013 275002 124112 275036
rect 122792 274915 122826 275002
rect 122792 274847 122826 274881
rect 124078 274915 124112 275002
rect 122792 274779 122826 274813
rect 122792 274711 122826 274745
rect 122792 274643 122826 274677
rect 124078 274847 124112 274881
rect 124078 274779 124112 274813
rect 124078 274711 124112 274745
rect 122792 274562 122826 274609
rect 124078 274643 124112 274677
rect 124078 274582 124112 274609
rect 122060 274541 122826 274562
rect 122060 274507 122110 274541
rect 122144 274507 122178 274541
rect 122212 274507 122246 274541
rect 122280 274507 122314 274541
rect 122348 274507 122382 274541
rect 122416 274507 122450 274541
rect 122484 274507 122518 274541
rect 122552 274507 122586 274541
rect 122620 274507 122654 274541
rect 122688 274522 122826 274541
rect 124078 274552 124848 274582
rect 124078 274522 124232 274552
rect 122688 274507 122891 274522
rect 122060 274488 122891 274507
rect 122925 274488 122959 274522
rect 122993 274488 123027 274522
rect 123061 274488 123095 274522
rect 123129 274488 123163 274522
rect 123197 274488 123231 274522
rect 123265 274488 123299 274522
rect 123333 274488 123367 274522
rect 123401 274488 123435 274522
rect 123469 274488 123503 274522
rect 123537 274488 123571 274522
rect 123605 274488 123639 274522
rect 123673 274488 123707 274522
rect 123741 274488 123775 274522
rect 123809 274488 123843 274522
rect 123877 274488 123911 274522
rect 123945 274488 123979 274522
rect 124013 274518 124232 274522
rect 124266 274518 124300 274552
rect 124334 274518 124368 274552
rect 124402 274518 124436 274552
rect 124470 274518 124504 274552
rect 124538 274518 124572 274552
rect 124606 274518 124640 274552
rect 124674 274518 124708 274552
rect 124742 274518 124776 274552
rect 124810 274518 124848 274552
rect 124013 274488 124848 274518
rect 122060 274486 122807 274488
rect 122060 274384 122150 274486
rect 122062 274281 122150 274384
rect 122062 274247 122089 274281
rect 122123 274247 122150 274281
rect 124726 274297 124814 274488
rect 122062 274213 122150 274247
rect 122062 274179 122089 274213
rect 122123 274179 122150 274213
rect 122062 274145 122150 274179
rect 122062 274111 122089 274145
rect 122123 274111 122150 274145
rect 122062 274077 122150 274111
rect 122062 274043 122089 274077
rect 122123 274043 122150 274077
rect 122062 274009 122150 274043
rect 122062 273975 122089 274009
rect 122123 273975 122150 274009
rect 122062 273941 122150 273975
rect 122062 273907 122089 273941
rect 122123 273907 122150 273941
rect 122062 273873 122150 273907
rect 122062 273839 122089 273873
rect 122123 273839 122150 273873
rect 122062 273805 122150 273839
rect 122062 273771 122089 273805
rect 122123 273771 122150 273805
rect 124726 274263 124753 274297
rect 124787 274263 124814 274297
rect 124726 274229 124814 274263
rect 124726 274195 124753 274229
rect 124787 274195 124814 274229
rect 124726 274161 124814 274195
rect 124726 274127 124753 274161
rect 124787 274127 124814 274161
rect 124726 274093 124814 274127
rect 124726 274059 124753 274093
rect 124787 274059 124814 274093
rect 124726 274025 124814 274059
rect 124726 273991 124753 274025
rect 124787 273991 124814 274025
rect 124726 273957 124814 273991
rect 124726 273923 124753 273957
rect 124787 273923 124814 273957
rect 124726 273889 124814 273923
rect 124726 273855 124753 273889
rect 124787 273855 124814 273889
rect 124726 273821 124814 273855
rect 124726 273787 124753 273821
rect 124787 273787 124814 273821
rect 122062 273737 122150 273771
rect 122062 273703 122089 273737
rect 122123 273703 122150 273737
rect 122062 273669 122150 273703
rect 124726 273753 124814 273787
rect 124726 273719 124753 273753
rect 124787 273719 124814 273753
rect 122062 273635 122089 273669
rect 122123 273635 122150 273669
rect 122062 273618 122150 273635
rect 124726 273685 124814 273719
rect 124726 273651 124753 273685
rect 124787 273651 124814 273685
rect 124726 273618 124814 273651
rect 122062 273598 124814 273618
rect 122062 273564 122243 273598
rect 122277 273564 122311 273598
rect 122345 273564 122379 273598
rect 122413 273564 122447 273598
rect 122481 273564 122515 273598
rect 122549 273564 122583 273598
rect 122617 273564 122651 273598
rect 122685 273564 122719 273598
rect 122753 273564 122787 273598
rect 122821 273564 122855 273598
rect 122889 273564 122923 273598
rect 122957 273564 122991 273598
rect 123025 273564 123059 273598
rect 123093 273564 123127 273598
rect 123161 273564 123195 273598
rect 123229 273564 123263 273598
rect 123297 273564 123331 273598
rect 123365 273564 123399 273598
rect 123433 273564 123467 273598
rect 123501 273564 123535 273598
rect 123569 273564 123603 273598
rect 123637 273564 123671 273598
rect 123705 273564 123739 273598
rect 123773 273564 123807 273598
rect 123841 273564 123875 273598
rect 123909 273564 123943 273598
rect 123977 273564 124011 273598
rect 124045 273564 124079 273598
rect 124113 273564 124147 273598
rect 124181 273564 124215 273598
rect 124249 273564 124283 273598
rect 124317 273564 124351 273598
rect 124385 273564 124419 273598
rect 124453 273564 124487 273598
rect 124521 273564 124555 273598
rect 124589 273564 124814 273598
rect 122062 273545 124814 273564
rect 123978 272750 124880 272777
rect 123978 272716 124065 272750
rect 124099 272716 124133 272750
rect 124167 272716 124201 272750
rect 124235 272716 124269 272750
rect 124303 272716 124337 272750
rect 124371 272716 124405 272750
rect 124439 272716 124473 272750
rect 124507 272716 124541 272750
rect 124575 272716 124609 272750
rect 124643 272716 124677 272750
rect 124711 272716 124880 272750
rect 123978 272689 124880 272716
rect 123978 272592 124029 272689
rect 123978 272558 123986 272592
rect 124020 272558 124029 272592
rect 124811 272687 124880 272689
rect 124811 272653 124828 272687
rect 124862 272653 124880 272687
rect 124811 272619 124880 272653
rect 124811 272585 124828 272619
rect 124862 272585 124880 272619
rect 123978 272524 124029 272558
rect 123978 272490 123986 272524
rect 124020 272490 124029 272524
rect 124811 272551 124880 272585
rect 123978 272456 124029 272490
rect 123978 272422 123986 272456
rect 124020 272422 124029 272456
rect 123978 272388 124029 272422
rect 123978 272354 123986 272388
rect 124020 272354 124029 272388
rect 123978 272320 124029 272354
rect 124811 272517 124828 272551
rect 124862 272517 124880 272551
rect 124811 272483 124880 272517
rect 124811 272449 124828 272483
rect 124862 272449 124880 272483
rect 124811 272415 124880 272449
rect 124811 272381 124828 272415
rect 124862 272381 124880 272415
rect 124811 272347 124880 272381
rect 123978 272286 123986 272320
rect 124020 272286 124029 272320
rect 123978 272252 124029 272286
rect 124811 272313 124828 272347
rect 124862 272313 124880 272347
rect 124811 272279 124880 272313
rect 123978 272218 123986 272252
rect 124020 272218 124029 272252
rect 123978 272184 124029 272218
rect 123978 272150 123986 272184
rect 124020 272150 124029 272184
rect 124811 272245 124828 272279
rect 124862 272245 124880 272279
rect 124811 272211 124880 272245
rect 124811 272177 124828 272211
rect 124862 272177 124880 272211
rect 123978 272116 124029 272150
rect 123978 272082 123986 272116
rect 124020 272082 124029 272116
rect 124811 272143 124880 272177
rect 124811 272109 124828 272143
rect 124862 272109 124880 272143
rect 123978 272048 124029 272082
rect 123978 272014 123986 272048
rect 124020 272014 124029 272048
rect 123978 271980 124029 272014
rect 123978 271946 123986 271980
rect 124020 271946 124029 271980
rect 123978 271912 124029 271946
rect 123978 271878 123986 271912
rect 124020 271878 124029 271912
rect 124811 272075 124880 272109
rect 124811 272041 124828 272075
rect 124862 272041 124880 272075
rect 124811 272007 124880 272041
rect 124811 271973 124828 272007
rect 124862 271973 124880 272007
rect 124811 271939 124880 271973
rect 124811 271905 124828 271939
rect 124862 271905 124880 271939
rect 123978 271844 124029 271878
rect 124811 271871 124880 271905
rect 123978 271810 123986 271844
rect 124020 271810 124029 271844
rect 123978 271776 124029 271810
rect 123978 271742 123986 271776
rect 124020 271742 124029 271776
rect 124811 271837 124828 271871
rect 124862 271837 124880 271871
rect 124811 271803 124880 271837
rect 124811 271769 124828 271803
rect 124862 271769 124880 271803
rect 123978 271708 124029 271742
rect 123978 271674 123986 271708
rect 124020 271674 124029 271708
rect 124811 271735 124880 271769
rect 124811 271701 124828 271735
rect 124862 271701 124880 271735
rect 123978 271640 124029 271674
rect 123978 271606 123986 271640
rect 124020 271606 124029 271640
rect 123978 271572 124029 271606
rect 123978 271538 123986 271572
rect 124020 271538 124029 271572
rect 123978 271504 124029 271538
rect 123978 271470 123986 271504
rect 124020 271470 124029 271504
rect 124811 271667 124880 271701
rect 124811 271633 124828 271667
rect 124862 271633 124880 271667
rect 124811 271599 124880 271633
rect 124811 271565 124828 271599
rect 124862 271565 124880 271599
rect 124811 271531 124880 271565
rect 124811 271497 124828 271531
rect 124862 271497 124880 271531
rect 123978 271436 124029 271470
rect 123978 271402 123986 271436
rect 124020 271402 124029 271436
rect 124811 271463 124880 271497
rect 123978 271368 124029 271402
rect 123978 271334 123986 271368
rect 124020 271334 124029 271368
rect 123978 271300 124029 271334
rect 124811 271429 124828 271463
rect 124862 271429 124880 271463
rect 124811 271395 124880 271429
rect 124811 271361 124828 271395
rect 124862 271361 124880 271395
rect 123978 271266 123986 271300
rect 124020 271266 124029 271300
rect 124811 271327 124880 271361
rect 124811 271293 124828 271327
rect 124862 271293 124880 271327
rect 123978 271232 124029 271266
rect 123978 271198 123986 271232
rect 124020 271198 124029 271232
rect 123978 271164 124029 271198
rect 123978 271130 123986 271164
rect 124020 271130 124029 271164
rect 123978 271096 124029 271130
rect 123978 271062 123986 271096
rect 124020 271062 124029 271096
rect 124811 271259 124880 271293
rect 124811 271225 124828 271259
rect 124862 271225 124880 271259
rect 124811 271191 124880 271225
rect 124811 271157 124828 271191
rect 124862 271157 124880 271191
rect 124811 271123 124880 271157
rect 124811 271089 124828 271123
rect 124862 271089 124880 271123
rect 123978 271028 124029 271062
rect 123978 270994 123986 271028
rect 124020 270994 124029 271028
rect 124811 271055 124880 271089
rect 124811 271021 124828 271055
rect 124862 271021 124880 271055
rect 123978 270960 124029 270994
rect 123978 270926 123986 270960
rect 124020 270926 124029 270960
rect 123978 270892 124029 270926
rect 124811 270987 124880 271021
rect 124811 270953 124828 270987
rect 124862 270953 124880 270987
rect 124811 270919 124880 270953
rect 123978 270858 123986 270892
rect 124020 270858 124029 270892
rect 123978 270824 124029 270858
rect 124811 270885 124828 270919
rect 124862 270885 124880 270919
rect 123978 270790 123986 270824
rect 124020 270790 124029 270824
rect 123978 270756 124029 270790
rect 123978 270722 123986 270756
rect 124020 270722 124029 270756
rect 123978 270688 124029 270722
rect 123978 270654 123986 270688
rect 124020 270654 124029 270688
rect 124811 270851 124880 270885
rect 124811 270817 124828 270851
rect 124862 270817 124880 270851
rect 124811 270783 124880 270817
rect 124811 270749 124828 270783
rect 124862 270749 124880 270783
rect 124811 270715 124880 270749
rect 124811 270681 124828 270715
rect 124862 270681 124880 270715
rect 123978 270620 124029 270654
rect 123978 270586 123986 270620
rect 124020 270586 124029 270620
rect 124811 270647 124880 270681
rect 124811 270613 124828 270647
rect 124862 270613 124880 270647
rect 123978 270552 124029 270586
rect 123978 270518 123986 270552
rect 124020 270518 124029 270552
rect 123978 270484 124029 270518
rect 124811 270579 124880 270613
rect 124811 270545 124828 270579
rect 124862 270545 124880 270579
rect 124811 270511 124880 270545
rect 123978 270450 123986 270484
rect 124020 270450 124029 270484
rect 123978 270416 124029 270450
rect 124811 270477 124828 270511
rect 124862 270477 124880 270511
rect 124811 270443 124880 270477
rect 123978 270382 123986 270416
rect 124020 270382 124029 270416
rect 123978 270348 124029 270382
rect 123978 270314 123986 270348
rect 124020 270314 124029 270348
rect 123978 270280 124029 270314
rect 123978 270246 123986 270280
rect 124020 270246 124029 270280
rect 123978 270212 124029 270246
rect 124811 270409 124828 270443
rect 124862 270409 124880 270443
rect 124811 270375 124880 270409
rect 124811 270341 124828 270375
rect 124862 270341 124880 270375
rect 124811 270307 124880 270341
rect 124811 270273 124828 270307
rect 124862 270273 124880 270307
rect 123978 270178 123986 270212
rect 124020 270178 124029 270212
rect 124811 270239 124880 270273
rect 124811 270205 124828 270239
rect 124862 270205 124880 270239
rect 123978 270144 124029 270178
rect 123978 270110 123986 270144
rect 124020 270110 124029 270144
rect 123978 270076 124029 270110
rect 124811 270171 124880 270205
rect 124811 270137 124828 270171
rect 124862 270137 124880 270171
rect 124811 270103 124880 270137
rect 123978 270042 123986 270076
rect 124020 270042 124029 270076
rect 123978 270008 124029 270042
rect 124811 270069 124828 270103
rect 124862 270069 124880 270103
rect 124811 270035 124880 270069
rect 123978 269974 123986 270008
rect 124020 269974 124029 270008
rect 123978 269940 124029 269974
rect 123978 269906 123986 269940
rect 124020 269906 124029 269940
rect 123978 269872 124029 269906
rect 123978 269838 123986 269872
rect 124020 269838 124029 269872
rect 123978 269804 124029 269838
rect 124811 270001 124828 270035
rect 124862 270001 124880 270035
rect 124811 269967 124880 270001
rect 124811 269933 124828 269967
rect 124862 269933 124880 269967
rect 124811 269899 124880 269933
rect 124811 269865 124828 269899
rect 124862 269865 124880 269899
rect 124811 269831 124880 269865
rect 123978 269770 123986 269804
rect 124020 269770 124029 269804
rect 123978 269736 124029 269770
rect 124811 269797 124828 269831
rect 124862 269797 124880 269831
rect 123978 269702 123986 269736
rect 124020 269702 124029 269736
rect 123978 269668 124029 269702
rect 123978 269634 123986 269668
rect 124020 269634 124029 269668
rect 124811 269763 124880 269797
rect 124811 269729 124828 269763
rect 124862 269729 124880 269763
rect 124811 269695 124880 269729
rect 123978 269600 124029 269634
rect 124811 269661 124828 269695
rect 124862 269661 124880 269695
rect 124811 269627 124880 269661
rect 123978 269566 123986 269600
rect 124020 269566 124029 269600
rect 123978 269532 124029 269566
rect 123978 269498 123986 269532
rect 124020 269498 124029 269532
rect 123978 269464 124029 269498
rect 123978 269430 123986 269464
rect 124020 269430 124029 269464
rect 123978 269396 124029 269430
rect 124811 269593 124828 269627
rect 124862 269593 124880 269627
rect 124811 269559 124880 269593
rect 124811 269525 124828 269559
rect 124862 269525 124880 269559
rect 124811 269491 124880 269525
rect 124811 269457 124828 269491
rect 124862 269457 124880 269491
rect 124811 269423 124880 269457
rect 123978 269362 123986 269396
rect 124020 269362 124029 269396
rect 123978 269281 124029 269362
rect 124811 269389 124828 269423
rect 124862 269389 124880 269423
rect 124811 269355 124880 269389
rect 124811 269321 124828 269355
rect 124862 269321 124880 269355
rect 124811 269281 124880 269321
rect 123978 269254 124880 269281
rect 123978 269220 124049 269254
rect 124083 269220 124117 269254
rect 124151 269220 124185 269254
rect 124219 269220 124253 269254
rect 124287 269220 124321 269254
rect 124355 269220 124389 269254
rect 124423 269220 124457 269254
rect 124491 269220 124525 269254
rect 124559 269220 124593 269254
rect 124627 269220 124661 269254
rect 124695 269220 124880 269254
rect 123978 269193 124880 269220
rect 125047 268990 125058 280856
rect 125160 268990 125171 280856
rect 125047 268861 125171 268990
rect 120072 268835 125199 268861
rect 120072 268785 120283 268835
rect 119938 268733 120283 268785
rect 125145 268733 125199 268835
rect 119938 268708 125199 268733
rect 119021 268651 119151 268677
<< nsubdiff >>
rect 106169 279188 106237 279222
rect 106271 279188 106305 279222
rect 106339 279188 106373 279222
rect 106407 279188 106441 279222
rect 106475 279188 106509 279222
rect 106543 279188 106577 279222
rect 106611 279188 106645 279222
rect 106679 279188 106713 279222
rect 106747 279188 106781 279222
rect 106815 279188 106849 279222
rect 106883 279188 106917 279222
rect 106951 279188 106985 279222
rect 107019 279188 107053 279222
rect 107087 279188 107121 279222
rect 107155 279188 107189 279222
rect 107223 279188 107257 279222
rect 107291 279188 107325 279222
rect 107359 279188 107393 279222
rect 107427 279188 107461 279222
rect 107495 279188 107529 279222
rect 107563 279188 107597 279222
rect 107631 279188 107665 279222
rect 107699 279188 107768 279222
rect 106169 279147 106203 279188
rect 106169 279079 106203 279113
rect 107734 279147 107768 279188
rect 107734 279079 107768 279113
rect 106169 279011 106203 279045
rect 107734 279011 107768 279045
rect 106169 278943 106203 278977
rect 106169 278875 106203 278909
rect 106169 278807 106203 278841
rect 106169 278739 106203 278773
rect 107734 278943 107768 278977
rect 107734 278875 107768 278909
rect 107734 278807 107768 278841
rect 106169 278671 106203 278705
rect 107734 278739 107768 278773
rect 106169 278603 106203 278637
rect 106169 278535 106203 278569
rect 106169 278467 106203 278501
rect 107734 278671 107768 278705
rect 107734 278603 107768 278637
rect 107734 278535 107768 278569
rect 106169 278399 106203 278433
rect 107734 278467 107768 278501
rect 106169 278331 106203 278365
rect 106169 278263 106203 278297
rect 106169 278195 106203 278229
rect 106169 278127 106203 278161
rect 107734 278399 107768 278433
rect 107734 278331 107768 278365
rect 107734 278263 107768 278297
rect 107734 278195 107768 278229
rect 107734 278127 107768 278161
rect 106169 278059 106203 278093
rect 106169 277984 106203 278025
rect 107734 278059 107768 278093
rect 107734 277984 107768 278025
rect 106169 277950 106237 277984
rect 106271 277950 106305 277984
rect 106339 277950 106373 277984
rect 106407 277950 106441 277984
rect 106475 277950 106509 277984
rect 106543 277950 106577 277984
rect 106611 277950 106645 277984
rect 106679 277950 106713 277984
rect 106747 277950 106781 277984
rect 106815 277950 106849 277984
rect 106883 277950 106917 277984
rect 106951 277950 106985 277984
rect 107019 277950 107053 277984
rect 107087 277950 107121 277984
rect 107155 277950 107189 277984
rect 107223 277950 107257 277984
rect 107291 277950 107325 277984
rect 107359 277950 107393 277984
rect 107427 277950 107461 277984
rect 107495 277950 107529 277984
rect 107563 277950 107597 277984
rect 107631 277950 107665 277984
rect 107699 277950 107768 277984
rect 106308 277290 106413 277324
rect 106447 277290 106481 277324
rect 106515 277290 106549 277324
rect 106583 277290 106617 277324
rect 106651 277290 106685 277324
rect 106719 277290 106753 277324
rect 106787 277290 106821 277324
rect 106855 277290 106889 277324
rect 106923 277290 106957 277324
rect 106991 277290 107025 277324
rect 107059 277290 107093 277324
rect 107127 277290 107161 277324
rect 107195 277290 107229 277324
rect 107263 277290 107297 277324
rect 107331 277290 107365 277324
rect 107399 277290 107433 277324
rect 107467 277290 107501 277324
rect 107535 277290 107569 277324
rect 107603 277290 107708 277324
rect 106308 277212 106342 277290
rect 106308 277144 106342 277178
rect 107674 277212 107708 277290
rect 106308 277076 106342 277110
rect 107674 277144 107708 277178
rect 106308 276964 106342 277042
rect 107674 277076 107708 277110
rect 107674 276964 107708 277042
rect 106308 276930 106413 276964
rect 106447 276930 106481 276964
rect 106515 276930 106549 276964
rect 106583 276930 106617 276964
rect 106651 276930 106685 276964
rect 106719 276930 106753 276964
rect 106787 276930 106821 276964
rect 106855 276930 106889 276964
rect 106923 276930 106957 276964
rect 106991 276930 107025 276964
rect 107059 276930 107093 276964
rect 107127 276930 107161 276964
rect 107195 276930 107229 276964
rect 107263 276930 107297 276964
rect 107331 276930 107365 276964
rect 107399 276930 107433 276964
rect 107467 276930 107501 276964
rect 107535 276930 107569 276964
rect 107603 276930 107708 276964
rect 106706 275900 106797 275934
rect 106831 275900 106865 275934
rect 106899 275900 106933 275934
rect 106967 275900 107001 275934
rect 107035 275900 107069 275934
rect 107103 275900 107137 275934
rect 107171 275900 107205 275934
rect 107239 275900 107273 275934
rect 107307 275900 107341 275934
rect 107375 275900 107409 275934
rect 107443 275900 107477 275934
rect 107511 275900 107545 275934
rect 107579 275900 107613 275934
rect 107647 275900 107681 275934
rect 107715 275900 107749 275934
rect 107783 275900 107817 275934
rect 107851 275900 107885 275934
rect 107919 275900 107953 275934
rect 107987 275900 108021 275934
rect 108055 275900 108089 275934
rect 108123 275900 108157 275934
rect 108191 275900 108225 275934
rect 108259 275900 108293 275934
rect 108327 275900 108361 275934
rect 108395 275900 108429 275934
rect 108463 275900 108497 275934
rect 108531 275900 108565 275934
rect 108599 275900 108633 275934
rect 108667 275900 108701 275934
rect 108735 275900 108769 275934
rect 108803 275900 108837 275934
rect 108871 275900 108905 275934
rect 108939 275900 108973 275934
rect 109007 275900 109041 275934
rect 109075 275900 109109 275934
rect 109143 275900 109177 275934
rect 109211 275900 109245 275934
rect 109279 275900 109313 275934
rect 109347 275900 109381 275934
rect 109415 275900 109449 275934
rect 109483 275900 109517 275934
rect 109551 275900 109585 275934
rect 109619 275900 109653 275934
rect 109687 275900 109721 275934
rect 109755 275900 109847 275934
rect 106706 275850 106740 275900
rect 106706 275782 106740 275816
rect 109813 275850 109847 275900
rect 109813 275782 109847 275816
rect 106706 275714 106740 275748
rect 109813 275714 109847 275748
rect 106706 275646 106740 275680
rect 106706 275578 106740 275612
rect 106706 275510 106740 275544
rect 106706 275442 106740 275476
rect 106706 275374 106740 275408
rect 106706 275306 106740 275340
rect 106706 275238 106740 275272
rect 106706 275170 106740 275204
rect 106706 275102 106740 275136
rect 106706 275034 106740 275068
rect 106706 274966 106740 275000
rect 109813 275646 109847 275680
rect 109813 275578 109847 275612
rect 109813 275510 109847 275544
rect 109813 275442 109847 275476
rect 109813 275374 109847 275408
rect 109813 275306 109847 275340
rect 109813 275238 109847 275272
rect 109813 275170 109847 275204
rect 109813 275102 109847 275136
rect 109813 275034 109847 275068
rect 109813 274966 109847 275000
rect 106706 274898 106740 274932
rect 109813 274898 109847 274932
rect 106706 274830 106740 274864
rect 106706 274747 106740 274796
rect 109813 274830 109847 274864
rect 109813 274747 109847 274796
rect 106706 274713 106797 274747
rect 106831 274713 106865 274747
rect 106899 274713 106933 274747
rect 106967 274713 107001 274747
rect 107035 274713 107069 274747
rect 107103 274713 107137 274747
rect 107171 274713 107205 274747
rect 107239 274713 107273 274747
rect 107307 274713 107341 274747
rect 107375 274713 107409 274747
rect 107443 274713 107477 274747
rect 107511 274713 107545 274747
rect 107579 274713 107613 274747
rect 107647 274713 107681 274747
rect 107715 274713 107749 274747
rect 107783 274713 107817 274747
rect 107851 274713 107885 274747
rect 107919 274713 107953 274747
rect 107987 274713 108021 274747
rect 108055 274713 108089 274747
rect 108123 274713 108157 274747
rect 108191 274713 108225 274747
rect 108259 274713 108293 274747
rect 108327 274713 108361 274747
rect 108395 274713 108429 274747
rect 108463 274713 108497 274747
rect 108531 274713 108565 274747
rect 108599 274713 108633 274747
rect 108667 274713 108701 274747
rect 108735 274713 108769 274747
rect 108803 274713 108837 274747
rect 108871 274713 108905 274747
rect 108939 274713 108973 274747
rect 109007 274713 109041 274747
rect 109075 274713 109109 274747
rect 109143 274713 109177 274747
rect 109211 274713 109245 274747
rect 109279 274713 109313 274747
rect 109347 274713 109381 274747
rect 109415 274713 109449 274747
rect 109483 274713 109517 274747
rect 109551 274713 109585 274747
rect 109619 274713 109653 274747
rect 109687 274713 109721 274747
rect 109755 274713 109847 274747
rect 109088 272568 109151 272602
rect 109185 272568 109219 272602
rect 109253 272568 109287 272602
rect 109321 272568 109355 272602
rect 109389 272568 109423 272602
rect 109457 272568 109491 272602
rect 109525 272568 109559 272602
rect 109593 272568 109627 272602
rect 109661 272568 109695 272602
rect 109729 272568 109763 272602
rect 109797 272568 109861 272602
rect 109088 272530 109122 272568
rect 109827 272530 109861 272568
rect 109088 272462 109122 272496
rect 109088 272394 109122 272428
rect 109827 272462 109861 272496
rect 109088 272326 109122 272360
rect 109088 272258 109122 272292
rect 109088 272190 109122 272224
rect 109088 272122 109122 272156
rect 109088 272054 109122 272088
rect 109088 271986 109122 272020
rect 109088 271918 109122 271952
rect 109088 271850 109122 271884
rect 109088 271782 109122 271816
rect 109088 271714 109122 271748
rect 109088 271646 109122 271680
rect 109088 271578 109122 271612
rect 109088 271510 109122 271544
rect 109088 271442 109122 271476
rect 109088 271374 109122 271408
rect 109088 271306 109122 271340
rect 109088 271238 109122 271272
rect 109088 271170 109122 271204
rect 109088 271102 109122 271136
rect 109088 271034 109122 271068
rect 109088 270966 109122 271000
rect 109088 270898 109122 270932
rect 109088 270830 109122 270864
rect 109088 270762 109122 270796
rect 109088 270694 109122 270728
rect 109827 272394 109861 272428
rect 109827 272326 109861 272360
rect 109827 272258 109861 272292
rect 109827 272190 109861 272224
rect 109827 272122 109861 272156
rect 109827 272054 109861 272088
rect 109827 271986 109861 272020
rect 109827 271918 109861 271952
rect 109827 271850 109861 271884
rect 109827 271782 109861 271816
rect 109827 271714 109861 271748
rect 109827 271646 109861 271680
rect 109827 271578 109861 271612
rect 109827 271510 109861 271544
rect 109827 271442 109861 271476
rect 109827 271374 109861 271408
rect 109827 271306 109861 271340
rect 109827 271238 109861 271272
rect 109827 271170 109861 271204
rect 109827 271102 109861 271136
rect 109827 271034 109861 271068
rect 109827 270966 109861 271000
rect 109827 270898 109861 270932
rect 109827 270830 109861 270864
rect 109827 270762 109861 270796
rect 109088 270626 109122 270660
rect 109827 270694 109861 270728
rect 109827 270626 109861 270660
rect 109088 270555 109122 270592
rect 109827 270555 109861 270592
rect 109088 270521 109151 270555
rect 109185 270521 109219 270555
rect 109253 270521 109287 270555
rect 109321 270521 109355 270555
rect 109389 270521 109423 270555
rect 109457 270521 109491 270555
rect 109525 270521 109559 270555
rect 109593 270521 109627 270555
rect 109661 270521 109695 270555
rect 109729 270521 109763 270555
rect 109797 270521 109861 270555
rect 114455 280929 114537 280963
rect 114571 280929 114605 280963
rect 114639 280929 114673 280963
rect 114707 280929 114741 280963
rect 114775 280929 114809 280963
rect 114843 280929 114877 280963
rect 114911 280929 114945 280963
rect 114979 280929 115061 280963
rect 114455 280897 114489 280929
rect 114455 280829 114489 280863
rect 115027 280897 115061 280929
rect 115027 280829 115061 280863
rect 114455 280761 114489 280795
rect 114455 280693 114489 280727
rect 114455 280625 114489 280659
rect 114455 280557 114489 280591
rect 114455 280489 114489 280523
rect 114455 280421 114489 280455
rect 115027 280761 115061 280795
rect 115027 280693 115061 280727
rect 115027 280625 115061 280659
rect 115027 280557 115061 280591
rect 115027 280489 115061 280523
rect 115027 280421 115061 280455
rect 114455 280353 114489 280387
rect 115027 280353 115061 280387
rect 114455 280285 114489 280319
rect 114455 280217 114489 280251
rect 114455 280149 114489 280183
rect 115027 280285 115061 280319
rect 115027 280217 115061 280251
rect 115027 280149 115061 280183
rect 114455 280081 114489 280115
rect 114455 280013 114489 280047
rect 114455 279945 114489 279979
rect 115027 280081 115061 280115
rect 115027 280013 115061 280047
rect 114455 279877 114489 279911
rect 115027 279945 115061 279979
rect 114455 279809 114489 279843
rect 114455 279741 114489 279775
rect 115027 279877 115061 279911
rect 115027 279809 115061 279843
rect 115027 279741 115061 279775
rect 114455 279673 114489 279707
rect 114455 279605 114489 279639
rect 114455 279537 114489 279571
rect 115027 279673 115061 279707
rect 115027 279605 115061 279639
rect 114455 279469 114489 279503
rect 115027 279537 115061 279571
rect 114455 279403 114489 279435
rect 115027 279469 115061 279503
rect 115027 279403 115061 279435
rect 114455 279369 114537 279403
rect 114571 279369 114605 279403
rect 114639 279369 114673 279403
rect 114707 279369 114741 279403
rect 114775 279369 114809 279403
rect 114843 279369 114877 279403
rect 114911 279369 114945 279403
rect 114979 279369 115061 279403
rect 115144 280929 115226 280963
rect 115260 280929 115294 280963
rect 115328 280929 115362 280963
rect 115396 280929 115430 280963
rect 115464 280929 115498 280963
rect 115532 280929 115566 280963
rect 115600 280929 115634 280963
rect 115668 280929 115750 280963
rect 115144 280897 115178 280929
rect 115144 280829 115178 280863
rect 115716 280897 115750 280929
rect 115716 280829 115750 280863
rect 115144 280761 115178 280795
rect 115144 280693 115178 280727
rect 115144 280625 115178 280659
rect 115144 280557 115178 280591
rect 115144 280489 115178 280523
rect 115144 280421 115178 280455
rect 115716 280761 115750 280795
rect 115716 280693 115750 280727
rect 115716 280625 115750 280659
rect 115716 280557 115750 280591
rect 115716 280489 115750 280523
rect 115716 280421 115750 280455
rect 115144 280353 115178 280387
rect 115716 280353 115750 280387
rect 115144 280285 115178 280319
rect 115144 280217 115178 280251
rect 115144 280149 115178 280183
rect 115716 280285 115750 280319
rect 115716 280217 115750 280251
rect 115716 280149 115750 280183
rect 115144 280081 115178 280115
rect 115144 280013 115178 280047
rect 115144 279945 115178 279979
rect 115716 280081 115750 280115
rect 115716 280013 115750 280047
rect 115144 279877 115178 279911
rect 115716 279945 115750 279979
rect 115144 279809 115178 279843
rect 115144 279741 115178 279775
rect 115716 279877 115750 279911
rect 115716 279809 115750 279843
rect 115716 279741 115750 279775
rect 115144 279673 115178 279707
rect 115144 279605 115178 279639
rect 115144 279537 115178 279571
rect 115716 279673 115750 279707
rect 115716 279605 115750 279639
rect 115144 279469 115178 279503
rect 115716 279537 115750 279571
rect 115144 279403 115178 279435
rect 115716 279469 115750 279503
rect 115716 279403 115750 279435
rect 115144 279369 115226 279403
rect 115260 279369 115294 279403
rect 115328 279369 115362 279403
rect 115396 279369 115430 279403
rect 115464 279369 115498 279403
rect 115532 279369 115566 279403
rect 115600 279369 115634 279403
rect 115668 279369 115750 279403
rect 114455 279263 114537 279297
rect 114571 279263 114605 279297
rect 114639 279263 114673 279297
rect 114707 279263 114741 279297
rect 114775 279263 114809 279297
rect 114843 279263 114877 279297
rect 114911 279263 114945 279297
rect 114979 279263 115061 279297
rect 114455 279231 114489 279263
rect 114455 279163 114489 279197
rect 115027 279231 115061 279263
rect 115027 279163 115061 279197
rect 114455 279095 114489 279129
rect 114455 279027 114489 279061
rect 114455 278959 114489 278993
rect 114455 278891 114489 278925
rect 114455 278823 114489 278857
rect 114455 278755 114489 278789
rect 115027 279095 115061 279129
rect 115027 279027 115061 279061
rect 115027 278959 115061 278993
rect 115027 278891 115061 278925
rect 115027 278823 115061 278857
rect 115027 278755 115061 278789
rect 114455 278687 114489 278721
rect 115027 278687 115061 278721
rect 114455 278619 114489 278653
rect 114455 278551 114489 278585
rect 114455 278483 114489 278517
rect 115027 278619 115061 278653
rect 115027 278551 115061 278585
rect 115027 278483 115061 278517
rect 114455 278415 114489 278449
rect 114455 278347 114489 278381
rect 114455 278279 114489 278313
rect 115027 278415 115061 278449
rect 115027 278347 115061 278381
rect 114455 278211 114489 278245
rect 115027 278279 115061 278313
rect 114455 278143 114489 278177
rect 114455 278075 114489 278109
rect 115027 278211 115061 278245
rect 115027 278143 115061 278177
rect 115027 278075 115061 278109
rect 114455 278007 114489 278041
rect 114455 277939 114489 277973
rect 114455 277871 114489 277905
rect 115027 278007 115061 278041
rect 115027 277939 115061 277973
rect 114455 277803 114489 277837
rect 115027 277871 115061 277905
rect 114455 277737 114489 277769
rect 115027 277803 115061 277837
rect 115027 277737 115061 277769
rect 114455 277703 114537 277737
rect 114571 277703 114605 277737
rect 114639 277703 114673 277737
rect 114707 277703 114741 277737
rect 114775 277703 114809 277737
rect 114843 277703 114877 277737
rect 114911 277703 114945 277737
rect 114979 277703 115061 277737
rect 115144 279263 115226 279297
rect 115260 279263 115294 279297
rect 115328 279263 115362 279297
rect 115396 279263 115430 279297
rect 115464 279263 115498 279297
rect 115532 279263 115566 279297
rect 115600 279263 115634 279297
rect 115668 279263 115750 279297
rect 115144 279231 115178 279263
rect 115144 279163 115178 279197
rect 115716 279231 115750 279263
rect 115716 279163 115750 279197
rect 115144 279095 115178 279129
rect 115144 279027 115178 279061
rect 115144 278959 115178 278993
rect 115144 278891 115178 278925
rect 115144 278823 115178 278857
rect 115144 278755 115178 278789
rect 115716 279095 115750 279129
rect 115716 279027 115750 279061
rect 115716 278959 115750 278993
rect 115716 278891 115750 278925
rect 115716 278823 115750 278857
rect 115716 278755 115750 278789
rect 115144 278687 115178 278721
rect 115716 278687 115750 278721
rect 115144 278619 115178 278653
rect 115144 278551 115178 278585
rect 115144 278483 115178 278517
rect 115716 278619 115750 278653
rect 115716 278551 115750 278585
rect 115716 278483 115750 278517
rect 115144 278415 115178 278449
rect 115144 278347 115178 278381
rect 115144 278279 115178 278313
rect 115716 278415 115750 278449
rect 115716 278347 115750 278381
rect 115144 278211 115178 278245
rect 115716 278279 115750 278313
rect 115144 278143 115178 278177
rect 115144 278075 115178 278109
rect 115716 278211 115750 278245
rect 115716 278143 115750 278177
rect 115716 278075 115750 278109
rect 115144 278007 115178 278041
rect 115144 277939 115178 277973
rect 115144 277871 115178 277905
rect 115716 278007 115750 278041
rect 115716 277939 115750 277973
rect 115144 277803 115178 277837
rect 115716 277871 115750 277905
rect 115144 277737 115178 277769
rect 115716 277803 115750 277837
rect 115716 277737 115750 277769
rect 115144 277703 115226 277737
rect 115260 277703 115294 277737
rect 115328 277703 115362 277737
rect 115396 277703 115430 277737
rect 115464 277703 115498 277737
rect 115532 277703 115566 277737
rect 115600 277703 115634 277737
rect 115668 277703 115750 277737
rect 114455 277597 114537 277631
rect 114571 277597 114605 277631
rect 114639 277597 114673 277631
rect 114707 277597 114741 277631
rect 114775 277597 114809 277631
rect 114843 277597 114877 277631
rect 114911 277597 114945 277631
rect 114979 277597 115061 277631
rect 114455 277565 114489 277597
rect 114455 277497 114489 277531
rect 115027 277565 115061 277597
rect 115027 277497 115061 277531
rect 114455 277429 114489 277463
rect 114455 277361 114489 277395
rect 114455 277293 114489 277327
rect 114455 277225 114489 277259
rect 114455 277157 114489 277191
rect 114455 277089 114489 277123
rect 115027 277429 115061 277463
rect 115027 277361 115061 277395
rect 115027 277293 115061 277327
rect 115027 277225 115061 277259
rect 115027 277157 115061 277191
rect 115027 277089 115061 277123
rect 114455 277021 114489 277055
rect 115027 277021 115061 277055
rect 114455 276953 114489 276987
rect 114455 276885 114489 276919
rect 114455 276817 114489 276851
rect 115027 276953 115061 276987
rect 115027 276885 115061 276919
rect 115027 276817 115061 276851
rect 114455 276749 114489 276783
rect 114455 276681 114489 276715
rect 114455 276613 114489 276647
rect 115027 276749 115061 276783
rect 115027 276681 115061 276715
rect 114455 276545 114489 276579
rect 115027 276613 115061 276647
rect 114455 276477 114489 276511
rect 114455 276409 114489 276443
rect 115027 276545 115061 276579
rect 115027 276477 115061 276511
rect 115027 276409 115061 276443
rect 114455 276341 114489 276375
rect 114455 276273 114489 276307
rect 114455 276205 114489 276239
rect 115027 276341 115061 276375
rect 115027 276273 115061 276307
rect 114455 276137 114489 276171
rect 115027 276205 115061 276239
rect 114455 276071 114489 276103
rect 115027 276137 115061 276171
rect 115027 276071 115061 276103
rect 114455 276037 114537 276071
rect 114571 276037 114605 276071
rect 114639 276037 114673 276071
rect 114707 276037 114741 276071
rect 114775 276037 114809 276071
rect 114843 276037 114877 276071
rect 114911 276037 114945 276071
rect 114979 276037 115061 276071
rect 115144 277597 115226 277631
rect 115260 277597 115294 277631
rect 115328 277597 115362 277631
rect 115396 277597 115430 277631
rect 115464 277597 115498 277631
rect 115532 277597 115566 277631
rect 115600 277597 115634 277631
rect 115668 277597 115750 277631
rect 115144 277565 115178 277597
rect 115144 277497 115178 277531
rect 115716 277565 115750 277597
rect 115716 277497 115750 277531
rect 115144 277429 115178 277463
rect 115144 277361 115178 277395
rect 115144 277293 115178 277327
rect 115144 277225 115178 277259
rect 115144 277157 115178 277191
rect 115144 277089 115178 277123
rect 115716 277429 115750 277463
rect 115716 277361 115750 277395
rect 115716 277293 115750 277327
rect 115716 277225 115750 277259
rect 115716 277157 115750 277191
rect 115716 277089 115750 277123
rect 115144 277021 115178 277055
rect 115716 277021 115750 277055
rect 115144 276953 115178 276987
rect 115144 276885 115178 276919
rect 115144 276817 115178 276851
rect 115716 276953 115750 276987
rect 115716 276885 115750 276919
rect 115716 276817 115750 276851
rect 115144 276749 115178 276783
rect 115144 276681 115178 276715
rect 115144 276613 115178 276647
rect 115716 276749 115750 276783
rect 115716 276681 115750 276715
rect 115144 276545 115178 276579
rect 115716 276613 115750 276647
rect 115144 276477 115178 276511
rect 115144 276409 115178 276443
rect 115716 276545 115750 276579
rect 115716 276477 115750 276511
rect 115716 276409 115750 276443
rect 115144 276341 115178 276375
rect 115144 276273 115178 276307
rect 115144 276205 115178 276239
rect 115716 276341 115750 276375
rect 115716 276273 115750 276307
rect 115144 276137 115178 276171
rect 115716 276205 115750 276239
rect 115144 276071 115178 276103
rect 115716 276137 115750 276171
rect 115716 276071 115750 276103
rect 115144 276037 115226 276071
rect 115260 276037 115294 276071
rect 115328 276037 115362 276071
rect 115396 276037 115430 276071
rect 115464 276037 115498 276071
rect 115532 276037 115566 276071
rect 115600 276037 115634 276071
rect 115668 276037 115750 276071
rect 114455 275931 114537 275965
rect 114571 275931 114605 275965
rect 114639 275931 114673 275965
rect 114707 275931 114741 275965
rect 114775 275931 114809 275965
rect 114843 275931 114877 275965
rect 114911 275931 114945 275965
rect 114979 275931 115061 275965
rect 114455 275899 114489 275931
rect 114455 275831 114489 275865
rect 115027 275899 115061 275931
rect 115027 275831 115061 275865
rect 114455 275763 114489 275797
rect 114455 275695 114489 275729
rect 114455 275627 114489 275661
rect 114455 275559 114489 275593
rect 114455 275491 114489 275525
rect 114455 275423 114489 275457
rect 115027 275763 115061 275797
rect 115027 275695 115061 275729
rect 115027 275627 115061 275661
rect 115027 275559 115061 275593
rect 115027 275491 115061 275525
rect 115027 275423 115061 275457
rect 114455 275355 114489 275389
rect 115027 275355 115061 275389
rect 114455 275287 114489 275321
rect 114455 275219 114489 275253
rect 114455 275151 114489 275185
rect 115027 275287 115061 275321
rect 115027 275219 115061 275253
rect 115027 275151 115061 275185
rect 114455 275083 114489 275117
rect 114455 275015 114489 275049
rect 114455 274947 114489 274981
rect 115027 275083 115061 275117
rect 115027 275015 115061 275049
rect 114455 274879 114489 274913
rect 115027 274947 115061 274981
rect 114455 274811 114489 274845
rect 114455 274743 114489 274777
rect 115027 274879 115061 274913
rect 115027 274811 115061 274845
rect 115027 274743 115061 274777
rect 114455 274675 114489 274709
rect 114455 274607 114489 274641
rect 114455 274539 114489 274573
rect 115027 274675 115061 274709
rect 115027 274607 115061 274641
rect 114455 274471 114489 274505
rect 115027 274539 115061 274573
rect 114455 274405 114489 274437
rect 115027 274471 115061 274505
rect 115027 274405 115061 274437
rect 114455 274371 114537 274405
rect 114571 274371 114605 274405
rect 114639 274371 114673 274405
rect 114707 274371 114741 274405
rect 114775 274371 114809 274405
rect 114843 274371 114877 274405
rect 114911 274371 114945 274405
rect 114979 274371 115061 274405
rect 115144 275931 115226 275965
rect 115260 275931 115294 275965
rect 115328 275931 115362 275965
rect 115396 275931 115430 275965
rect 115464 275931 115498 275965
rect 115532 275931 115566 275965
rect 115600 275931 115634 275965
rect 115668 275931 115750 275965
rect 115144 275899 115178 275931
rect 115144 275831 115178 275865
rect 115716 275899 115750 275931
rect 115716 275831 115750 275865
rect 115144 275763 115178 275797
rect 115144 275695 115178 275729
rect 115144 275627 115178 275661
rect 115144 275559 115178 275593
rect 115144 275491 115178 275525
rect 115144 275423 115178 275457
rect 115716 275763 115750 275797
rect 115716 275695 115750 275729
rect 115716 275627 115750 275661
rect 115716 275559 115750 275593
rect 115716 275491 115750 275525
rect 115716 275423 115750 275457
rect 115144 275355 115178 275389
rect 115716 275355 115750 275389
rect 115144 275287 115178 275321
rect 115144 275219 115178 275253
rect 115144 275151 115178 275185
rect 115716 275287 115750 275321
rect 115716 275219 115750 275253
rect 115716 275151 115750 275185
rect 115144 275083 115178 275117
rect 115144 275015 115178 275049
rect 115144 274947 115178 274981
rect 115716 275083 115750 275117
rect 115716 275015 115750 275049
rect 115144 274879 115178 274913
rect 115716 274947 115750 274981
rect 115144 274811 115178 274845
rect 115144 274743 115178 274777
rect 115716 274879 115750 274913
rect 115716 274811 115750 274845
rect 115716 274743 115750 274777
rect 115144 274675 115178 274709
rect 115144 274607 115178 274641
rect 115144 274539 115178 274573
rect 115716 274675 115750 274709
rect 115716 274607 115750 274641
rect 115144 274471 115178 274505
rect 115716 274539 115750 274573
rect 115144 274405 115178 274437
rect 115716 274471 115750 274505
rect 115716 274405 115750 274437
rect 115144 274371 115226 274405
rect 115260 274371 115294 274405
rect 115328 274371 115362 274405
rect 115396 274371 115430 274405
rect 115464 274371 115498 274405
rect 115532 274371 115566 274405
rect 115600 274371 115634 274405
rect 115668 274371 115750 274405
rect 114455 274265 114537 274299
rect 114571 274265 114605 274299
rect 114639 274265 114673 274299
rect 114707 274265 114741 274299
rect 114775 274265 114809 274299
rect 114843 274265 114877 274299
rect 114911 274265 114945 274299
rect 114979 274265 115061 274299
rect 114455 274233 114489 274265
rect 114455 274165 114489 274199
rect 115027 274233 115061 274265
rect 115027 274165 115061 274199
rect 114455 274097 114489 274131
rect 114455 274029 114489 274063
rect 114455 273961 114489 273995
rect 114455 273893 114489 273927
rect 114455 273825 114489 273859
rect 114455 273757 114489 273791
rect 115027 274097 115061 274131
rect 115027 274029 115061 274063
rect 115027 273961 115061 273995
rect 115027 273893 115061 273927
rect 115027 273825 115061 273859
rect 115027 273757 115061 273791
rect 114455 273689 114489 273723
rect 115027 273689 115061 273723
rect 114455 273621 114489 273655
rect 114455 273553 114489 273587
rect 114455 273485 114489 273519
rect 115027 273621 115061 273655
rect 115027 273553 115061 273587
rect 115027 273485 115061 273519
rect 114455 273417 114489 273451
rect 114455 273349 114489 273383
rect 114455 273281 114489 273315
rect 115027 273417 115061 273451
rect 115027 273349 115061 273383
rect 114455 273213 114489 273247
rect 115027 273281 115061 273315
rect 114455 273145 114489 273179
rect 114455 273077 114489 273111
rect 115027 273213 115061 273247
rect 115027 273145 115061 273179
rect 115027 273077 115061 273111
rect 114455 273009 114489 273043
rect 114455 272941 114489 272975
rect 114455 272873 114489 272907
rect 115027 273009 115061 273043
rect 115027 272941 115061 272975
rect 114455 272805 114489 272839
rect 115027 272873 115061 272907
rect 114455 272739 114489 272771
rect 115027 272805 115061 272839
rect 115027 272739 115061 272771
rect 114455 272705 114537 272739
rect 114571 272705 114605 272739
rect 114639 272705 114673 272739
rect 114707 272705 114741 272739
rect 114775 272705 114809 272739
rect 114843 272705 114877 272739
rect 114911 272705 114945 272739
rect 114979 272705 115061 272739
rect 115144 274265 115226 274299
rect 115260 274265 115294 274299
rect 115328 274265 115362 274299
rect 115396 274265 115430 274299
rect 115464 274265 115498 274299
rect 115532 274265 115566 274299
rect 115600 274265 115634 274299
rect 115668 274265 115750 274299
rect 115144 274233 115178 274265
rect 115144 274165 115178 274199
rect 115716 274233 115750 274265
rect 115716 274165 115750 274199
rect 115144 274097 115178 274131
rect 115144 274029 115178 274063
rect 115144 273961 115178 273995
rect 115144 273893 115178 273927
rect 115144 273825 115178 273859
rect 115144 273757 115178 273791
rect 115716 274097 115750 274131
rect 115716 274029 115750 274063
rect 115716 273961 115750 273995
rect 115716 273893 115750 273927
rect 115716 273825 115750 273859
rect 115716 273757 115750 273791
rect 115144 273689 115178 273723
rect 115716 273689 115750 273723
rect 115144 273621 115178 273655
rect 115144 273553 115178 273587
rect 115144 273485 115178 273519
rect 115716 273621 115750 273655
rect 115716 273553 115750 273587
rect 115716 273485 115750 273519
rect 115144 273417 115178 273451
rect 115144 273349 115178 273383
rect 115144 273281 115178 273315
rect 115716 273417 115750 273451
rect 115716 273349 115750 273383
rect 115144 273213 115178 273247
rect 115716 273281 115750 273315
rect 115144 273145 115178 273179
rect 115144 273077 115178 273111
rect 115716 273213 115750 273247
rect 115716 273145 115750 273179
rect 115716 273077 115750 273111
rect 115144 273009 115178 273043
rect 115144 272941 115178 272975
rect 115144 272873 115178 272907
rect 115716 273009 115750 273043
rect 115716 272941 115750 272975
rect 115144 272805 115178 272839
rect 115716 272873 115750 272907
rect 115144 272739 115178 272771
rect 115716 272805 115750 272839
rect 115716 272739 115750 272771
rect 115144 272705 115226 272739
rect 115260 272705 115294 272739
rect 115328 272705 115362 272739
rect 115396 272705 115430 272739
rect 115464 272705 115498 272739
rect 115532 272705 115566 272739
rect 115600 272705 115634 272739
rect 115668 272705 115750 272739
rect 112307 271634 112391 271668
rect 112425 271634 112459 271668
rect 112493 271634 112527 271668
rect 112561 271634 112595 271668
rect 112629 271634 112663 271668
rect 112697 271634 112731 271668
rect 112765 271634 112799 271668
rect 112833 271634 112867 271668
rect 112901 271634 112935 271668
rect 112969 271634 113003 271668
rect 113037 271634 113071 271668
rect 113105 271634 113139 271668
rect 113173 271634 113207 271668
rect 113241 271634 113275 271668
rect 113309 271634 113343 271668
rect 113377 271634 113411 271668
rect 113445 271634 113479 271668
rect 113513 271634 113547 271668
rect 113581 271634 113615 271668
rect 113649 271634 113683 271668
rect 113717 271634 113751 271668
rect 113785 271634 113819 271668
rect 113853 271634 113887 271668
rect 113921 271634 113955 271668
rect 113989 271634 114023 271668
rect 114057 271634 114091 271668
rect 114125 271634 114210 271668
rect 112307 271582 112341 271634
rect 112307 271514 112341 271548
rect 112307 271446 112341 271480
rect 112307 271378 112341 271412
rect 114176 271582 114210 271634
rect 114176 271514 114210 271548
rect 114176 271446 114210 271480
rect 112307 271310 112341 271344
rect 114176 271378 114210 271412
rect 114176 271310 114210 271344
rect 112307 271242 112341 271276
rect 112307 271174 112341 271208
rect 112307 271106 112341 271140
rect 114176 271242 114210 271276
rect 114176 271174 114210 271208
rect 114176 271106 114210 271140
rect 112307 271038 112341 271072
rect 114176 271038 114210 271072
rect 112307 270970 112341 271004
rect 112307 270902 112341 270936
rect 112307 270817 112341 270868
rect 114176 270970 114210 271004
rect 114176 270902 114210 270936
rect 114176 270817 114210 270868
rect 112307 270783 112391 270817
rect 112425 270783 112459 270817
rect 112493 270783 112527 270817
rect 112561 270783 112595 270817
rect 112629 270783 112663 270817
rect 112697 270783 112731 270817
rect 112765 270783 112799 270817
rect 112833 270783 112867 270817
rect 112901 270783 112935 270817
rect 112969 270783 113003 270817
rect 113037 270783 113071 270817
rect 113105 270783 113139 270817
rect 113173 270783 113207 270817
rect 113241 270783 113275 270817
rect 113309 270783 113343 270817
rect 113377 270783 113411 270817
rect 113445 270783 113479 270817
rect 113513 270783 113547 270817
rect 113581 270783 113615 270817
rect 113649 270783 113683 270817
rect 113717 270783 113751 270817
rect 113785 270783 113819 270817
rect 113853 270783 113887 270817
rect 113921 270783 113955 270817
rect 113989 270783 114023 270817
rect 114057 270783 114091 270817
rect 114125 270783 114210 270817
rect 114329 271554 114389 271588
rect 114423 271554 114457 271588
rect 114491 271554 114525 271588
rect 114559 271554 114593 271588
rect 114627 271554 114661 271588
rect 114695 271554 114729 271588
rect 114763 271554 114797 271588
rect 114831 271554 114865 271588
rect 114899 271554 114933 271588
rect 114967 271554 115001 271588
rect 115035 271554 115069 271588
rect 115103 271554 115137 271588
rect 115171 271554 115205 271588
rect 115239 271554 115273 271588
rect 115307 271554 115341 271588
rect 115375 271554 115409 271588
rect 115443 271554 115503 271588
rect 114329 271503 114363 271554
rect 114329 271435 114363 271469
rect 114329 271367 114363 271401
rect 115469 271503 115503 271554
rect 115469 271435 115503 271469
rect 114329 271299 114363 271333
rect 115469 271367 115503 271401
rect 115469 271299 115503 271333
rect 114329 271231 114363 271265
rect 114329 271163 114363 271197
rect 114329 271095 114363 271129
rect 115469 271231 115503 271265
rect 115469 271163 115503 271197
rect 115469 271095 115503 271129
rect 114329 271027 114363 271061
rect 114329 270959 114363 270993
rect 115469 271027 115503 271061
rect 114329 270891 114363 270925
rect 114329 270806 114363 270857
rect 115469 270959 115503 270993
rect 115469 270891 115503 270925
rect 115469 270806 115503 270857
rect 114329 270772 114389 270806
rect 114423 270772 114457 270806
rect 114491 270772 114525 270806
rect 114559 270772 114593 270806
rect 114627 270772 114661 270806
rect 114695 270772 114729 270806
rect 114763 270772 114797 270806
rect 114831 270772 114865 270806
rect 114899 270772 114933 270806
rect 114967 270772 115001 270806
rect 115035 270772 115069 270806
rect 115103 270772 115137 270806
rect 115171 270772 115205 270806
rect 115239 270772 115273 270806
rect 115307 270772 115341 270806
rect 115375 270772 115409 270806
rect 115443 270772 115503 270806
rect 120237 280779 120319 280813
rect 120353 280779 120387 280813
rect 120421 280779 120455 280813
rect 120489 280779 120523 280813
rect 120557 280779 120591 280813
rect 120625 280779 120659 280813
rect 120693 280779 120727 280813
rect 120761 280779 120795 280813
rect 120829 280779 120863 280813
rect 120897 280779 120931 280813
rect 120965 280779 120999 280813
rect 121033 280779 121067 280813
rect 121101 280779 121135 280813
rect 121169 280779 121203 280813
rect 121237 280779 121271 280813
rect 121305 280779 121339 280813
rect 121373 280779 121407 280813
rect 121441 280779 121475 280813
rect 121509 280779 121543 280813
rect 121577 280779 121611 280813
rect 121645 280779 121728 280813
rect 120237 280726 120271 280779
rect 120237 280658 120271 280692
rect 121694 280726 121728 280779
rect 121694 280658 121728 280692
rect 120237 280590 120271 280624
rect 120237 280522 120271 280556
rect 121694 280590 121728 280624
rect 120237 280454 120271 280488
rect 121694 280522 121728 280556
rect 121694 280454 121728 280488
rect 120237 280386 120271 280420
rect 120237 280318 120271 280352
rect 121694 280386 121728 280420
rect 120237 280250 120271 280284
rect 121694 280318 121728 280352
rect 120237 280182 120271 280216
rect 120237 280114 120271 280148
rect 120237 280046 120271 280080
rect 120237 279978 120271 280012
rect 120237 279910 120271 279944
rect 120237 279842 120271 279876
rect 120237 279774 120271 279808
rect 121694 280250 121728 280284
rect 121694 280182 121728 280216
rect 121694 280114 121728 280148
rect 121694 280046 121728 280080
rect 121694 279978 121728 280012
rect 121694 279910 121728 279944
rect 121694 279842 121728 279876
rect 121694 279774 121728 279808
rect 120237 279706 120271 279740
rect 120237 279638 120271 279672
rect 121694 279706 121728 279740
rect 120237 279570 120271 279604
rect 121694 279638 121728 279672
rect 121694 279570 121728 279604
rect 120237 279502 120271 279536
rect 121694 279502 121728 279536
rect 120237 279434 120271 279468
rect 120237 279366 120271 279400
rect 120237 279298 120271 279332
rect 120237 279230 120271 279264
rect 120237 279162 120271 279196
rect 120237 279094 120271 279128
rect 120237 279026 120271 279060
rect 120237 278958 120271 278992
rect 121694 279434 121728 279468
rect 121694 279366 121728 279400
rect 121694 279298 121728 279332
rect 121694 279230 121728 279264
rect 121694 279162 121728 279196
rect 121694 279094 121728 279128
rect 121694 279026 121728 279060
rect 120237 278890 120271 278924
rect 121694 278958 121728 278992
rect 122178 280574 122245 280608
rect 122279 280574 122313 280608
rect 122347 280574 122381 280608
rect 122415 280574 122449 280608
rect 122483 280574 122517 280608
rect 122551 280574 122585 280608
rect 122619 280574 122653 280608
rect 122687 280574 122721 280608
rect 122755 280574 122789 280608
rect 122823 280574 122857 280608
rect 122891 280574 122925 280608
rect 122959 280574 122993 280608
rect 123027 280574 123061 280608
rect 123095 280574 123129 280608
rect 123163 280574 123197 280608
rect 123231 280574 123265 280608
rect 123299 280574 123333 280608
rect 123367 280574 123401 280608
rect 123435 280574 123469 280608
rect 123503 280574 123537 280608
rect 123571 280574 123638 280608
rect 122178 280518 122212 280574
rect 122178 280450 122212 280484
rect 123604 280518 123638 280574
rect 123604 280450 123638 280484
rect 122178 280382 122212 280416
rect 122178 280314 122212 280348
rect 122178 280246 122212 280280
rect 122178 280178 122212 280212
rect 122178 280110 122212 280144
rect 122178 280042 122212 280076
rect 122178 279974 122212 280008
rect 122178 279906 122212 279940
rect 123604 280382 123638 280416
rect 123604 280314 123638 280348
rect 123604 280246 123638 280280
rect 123604 280178 123638 280212
rect 123604 280110 123638 280144
rect 123604 280042 123638 280076
rect 123604 279974 123638 280008
rect 122178 279838 122212 279872
rect 123604 279906 123638 279940
rect 123604 279838 123638 279872
rect 122178 279770 122212 279804
rect 123604 279770 123638 279804
rect 122178 279702 122212 279736
rect 122178 279634 122212 279668
rect 123604 279702 123638 279736
rect 122178 279566 122212 279600
rect 122178 279498 122212 279532
rect 122178 279430 122212 279464
rect 122178 279362 122212 279396
rect 122178 279294 122212 279328
rect 122178 279226 122212 279260
rect 122178 279158 122212 279192
rect 123604 279634 123638 279668
rect 123604 279566 123638 279600
rect 123604 279498 123638 279532
rect 123604 279430 123638 279464
rect 123604 279362 123638 279396
rect 123604 279294 123638 279328
rect 123604 279226 123638 279260
rect 123604 279158 123638 279192
rect 122178 279090 122212 279124
rect 122178 279000 122212 279056
rect 123604 279090 123638 279124
rect 123604 279000 123638 279056
rect 122178 278966 122245 279000
rect 122279 278966 122313 279000
rect 122347 278966 122381 279000
rect 122415 278966 122449 279000
rect 122483 278966 122517 279000
rect 122551 278966 122585 279000
rect 122619 278966 122653 279000
rect 122687 278966 122721 279000
rect 122755 278966 122789 279000
rect 122823 278966 122857 279000
rect 122891 278966 122925 279000
rect 122959 278966 122993 279000
rect 123027 278966 123061 279000
rect 123095 278966 123129 279000
rect 123163 278966 123197 279000
rect 123231 278966 123265 279000
rect 123299 278966 123333 279000
rect 123367 278966 123401 279000
rect 123435 278966 123469 279000
rect 123503 278966 123537 279000
rect 123571 278966 123638 279000
rect 121694 278890 121728 278924
rect 120237 278822 120271 278856
rect 120237 278754 120271 278788
rect 121694 278822 121728 278856
rect 120237 278686 120271 278720
rect 121694 278754 121728 278788
rect 121694 278686 121728 278720
rect 120237 278618 120271 278652
rect 120237 278550 120271 278584
rect 120237 278482 120271 278516
rect 120237 278414 120271 278448
rect 120237 278346 120271 278380
rect 120237 278278 120271 278312
rect 120237 278210 120271 278244
rect 121694 278618 121728 278652
rect 121694 278550 121728 278584
rect 121694 278482 121728 278516
rect 121694 278414 121728 278448
rect 121694 278346 121728 278380
rect 121694 278278 121728 278312
rect 121694 278210 121728 278244
rect 120237 278142 120271 278176
rect 120237 278074 120271 278108
rect 121694 278142 121728 278176
rect 120237 278006 120271 278040
rect 121694 278074 121728 278108
rect 121694 278006 121728 278040
rect 120237 277938 120271 277972
rect 120237 277870 120271 277904
rect 121694 277938 121728 277972
rect 120237 277802 120271 277836
rect 120237 277734 120271 277768
rect 120237 277666 120271 277700
rect 120237 277598 120271 277632
rect 120237 277530 120271 277564
rect 120237 277462 120271 277496
rect 120237 277394 120271 277428
rect 121694 277870 121728 277904
rect 121694 277802 121728 277836
rect 121694 277734 121728 277768
rect 121694 277666 121728 277700
rect 121694 277598 121728 277632
rect 121694 277530 121728 277564
rect 121694 277462 121728 277496
rect 120237 277326 120271 277360
rect 121694 277394 121728 277428
rect 121694 277326 121728 277360
rect 120237 277258 120271 277292
rect 120237 277190 120271 277224
rect 121694 277258 121728 277292
rect 120237 277122 120271 277156
rect 121694 277190 121728 277224
rect 121694 277122 121728 277156
rect 120237 277054 120271 277088
rect 120237 276986 120271 277020
rect 120237 276918 120271 276952
rect 120237 276850 120271 276884
rect 120237 276782 120271 276816
rect 120237 276714 120271 276748
rect 120237 276646 120271 276680
rect 121694 277054 121728 277088
rect 121694 276986 121728 277020
rect 121694 276918 121728 276952
rect 121694 276850 121728 276884
rect 121694 276782 121728 276816
rect 121694 276714 121728 276748
rect 121694 276646 121728 276680
rect 120237 276578 120271 276612
rect 120237 276510 120271 276544
rect 121694 276578 121728 276612
rect 120237 276442 120271 276476
rect 121694 276510 121728 276544
rect 121694 276442 121728 276476
rect 120237 276374 120271 276408
rect 120237 276306 120271 276340
rect 121694 276374 121728 276408
rect 120237 276238 120271 276272
rect 120237 276170 120271 276204
rect 120237 276102 120271 276136
rect 120237 276034 120271 276068
rect 120237 275966 120271 276000
rect 120237 275898 120271 275932
rect 120237 275830 120271 275864
rect 121694 276306 121728 276340
rect 121694 276238 121728 276272
rect 121694 276170 121728 276204
rect 121694 276102 121728 276136
rect 121694 276034 121728 276068
rect 121694 275966 121728 276000
rect 121694 275898 121728 275932
rect 120237 275762 120271 275796
rect 121694 275830 121728 275864
rect 121694 275762 121728 275796
rect 120237 275694 120271 275728
rect 120237 275626 120271 275660
rect 121694 275694 121728 275728
rect 120237 275558 120271 275592
rect 121694 275626 121728 275660
rect 121694 275558 121728 275592
rect 120237 275490 120271 275524
rect 120237 275422 120271 275456
rect 120237 275354 120271 275388
rect 120237 275286 120271 275320
rect 120237 275218 120271 275252
rect 120237 275150 120271 275184
rect 120237 275082 120271 275116
rect 121694 275490 121728 275524
rect 122254 278448 122343 278482
rect 122377 278448 122411 278482
rect 122445 278448 122479 278482
rect 122513 278448 122547 278482
rect 122581 278448 122615 278482
rect 122649 278448 122683 278482
rect 122717 278448 122751 278482
rect 122785 278448 122819 278482
rect 122853 278448 122887 278482
rect 122921 278448 122955 278482
rect 122989 278448 123023 278482
rect 123057 278448 123091 278482
rect 123125 278448 123159 278482
rect 123193 278448 123227 278482
rect 123261 278448 123295 278482
rect 123329 278448 123363 278482
rect 123397 278448 123431 278482
rect 123465 278448 123499 278482
rect 123533 278448 123567 278482
rect 123601 278448 123635 278482
rect 123669 278448 123703 278482
rect 123737 278448 123771 278482
rect 123805 278448 123839 278482
rect 123873 278448 123907 278482
rect 123941 278448 123975 278482
rect 124009 278448 124043 278482
rect 124077 278448 124111 278482
rect 124145 278448 124179 278482
rect 124213 278448 124247 278482
rect 124281 278448 124370 278482
rect 122254 278395 122288 278448
rect 124336 278395 124370 278448
rect 122254 278327 122288 278361
rect 122254 278259 122288 278293
rect 124336 278327 124370 278361
rect 122254 278191 122288 278225
rect 122254 278123 122288 278157
rect 122254 278055 122288 278089
rect 122254 277987 122288 278021
rect 122254 277919 122288 277953
rect 122254 277851 122288 277885
rect 122254 277783 122288 277817
rect 124336 278259 124370 278293
rect 124336 278191 124370 278225
rect 124336 278123 124370 278157
rect 122254 277715 122288 277749
rect 122254 277647 122288 277681
rect 122254 277579 122288 277613
rect 122254 277511 122288 277545
rect 122254 277443 122288 277477
rect 122254 277375 122288 277409
rect 122254 277307 122288 277341
rect 124336 278055 124370 278089
rect 124336 277987 124370 278021
rect 124336 277919 124370 277953
rect 124336 277851 124370 277885
rect 124336 277783 124370 277817
rect 124336 277715 124370 277749
rect 124336 277647 124370 277681
rect 124336 277579 124370 277613
rect 124336 277511 124370 277545
rect 124336 277443 124370 277477
rect 124336 277375 124370 277409
rect 124336 277307 124370 277341
rect 122254 277221 122288 277273
rect 124336 277221 124370 277273
rect 122254 277187 122343 277221
rect 122377 277187 122411 277221
rect 122445 277187 122479 277221
rect 122513 277187 122547 277221
rect 122581 277187 122615 277221
rect 122649 277187 122683 277221
rect 122717 277187 122751 277221
rect 122785 277187 122819 277221
rect 122853 277187 122887 277221
rect 122921 277187 122955 277221
rect 122989 277187 123023 277221
rect 123057 277187 123091 277221
rect 123125 277187 123159 277221
rect 123193 277187 123227 277221
rect 123261 277187 123295 277221
rect 123329 277187 123363 277221
rect 123397 277187 123431 277221
rect 123465 277187 123499 277221
rect 123533 277187 123567 277221
rect 123601 277187 123635 277221
rect 123669 277187 123703 277221
rect 123737 277187 123771 277221
rect 123805 277187 123839 277221
rect 123873 277187 123907 277221
rect 123941 277187 123975 277221
rect 124009 277187 124043 277221
rect 124077 277187 124111 277221
rect 124145 277187 124179 277221
rect 124213 277187 124247 277221
rect 124281 277187 124370 277221
rect 122278 276817 122404 276851
rect 122438 276817 122472 276851
rect 122506 276817 122540 276851
rect 122574 276817 122608 276851
rect 122642 276817 122676 276851
rect 122710 276817 122744 276851
rect 122778 276817 122812 276851
rect 122846 276817 122880 276851
rect 122914 276817 122948 276851
rect 122982 276817 123016 276851
rect 123050 276817 123084 276851
rect 123118 276817 123152 276851
rect 123186 276817 123220 276851
rect 123254 276817 123288 276851
rect 123322 276817 123356 276851
rect 123390 276817 123424 276851
rect 123458 276817 123492 276851
rect 123526 276817 123560 276851
rect 123594 276817 123628 276851
rect 123662 276817 123696 276851
rect 123730 276817 123764 276851
rect 123798 276817 123832 276851
rect 123866 276817 123992 276851
rect 122278 276733 122312 276817
rect 122278 276665 122312 276699
rect 123958 276733 123992 276817
rect 122278 276597 122312 276631
rect 122278 276529 122312 276563
rect 122278 276461 122312 276495
rect 123958 276665 123992 276699
rect 123958 276597 123992 276631
rect 123958 276529 123992 276563
rect 122278 276343 122312 276427
rect 123958 276461 123992 276495
rect 123958 276343 123992 276427
rect 122278 276309 122404 276343
rect 122438 276309 122472 276343
rect 122506 276309 122540 276343
rect 122574 276309 122608 276343
rect 122642 276309 122676 276343
rect 122710 276309 122744 276343
rect 122778 276309 122812 276343
rect 122846 276309 122880 276343
rect 122914 276309 122948 276343
rect 122982 276309 123016 276343
rect 123050 276309 123084 276343
rect 123118 276309 123152 276343
rect 123186 276309 123220 276343
rect 123254 276309 123288 276343
rect 123322 276309 123356 276343
rect 123390 276309 123424 276343
rect 123458 276309 123492 276343
rect 123526 276309 123560 276343
rect 123594 276309 123628 276343
rect 123662 276309 123696 276343
rect 123730 276309 123764 276343
rect 123798 276309 123832 276343
rect 123866 276309 123992 276343
rect 122283 275937 122379 275971
rect 122413 275937 122447 275971
rect 122481 275937 122515 275971
rect 122549 275937 122583 275971
rect 122617 275937 122651 275971
rect 122685 275937 122719 275971
rect 122753 275937 122787 275971
rect 122821 275937 122855 275971
rect 122889 275937 122923 275971
rect 122957 275937 122991 275971
rect 123025 275937 123059 275971
rect 123093 275937 123127 275971
rect 123161 275937 123195 275971
rect 123229 275937 123263 275971
rect 123297 275937 123331 275971
rect 123365 275937 123399 275971
rect 123433 275937 123467 275971
rect 123501 275937 123535 275971
rect 123569 275937 123603 275971
rect 123637 275937 123671 275971
rect 123705 275937 123739 275971
rect 123773 275937 123807 275971
rect 123841 275937 123875 275971
rect 123909 275937 123943 275971
rect 123977 275937 124011 275971
rect 124045 275937 124079 275971
rect 124113 275937 124147 275971
rect 124181 275937 124215 275971
rect 124249 275937 124283 275971
rect 124317 275937 124351 275971
rect 124385 275937 124419 275971
rect 124453 275937 124487 275971
rect 124521 275937 124555 275971
rect 124589 275937 124623 275971
rect 124657 275937 124691 275971
rect 124725 275937 124759 275971
rect 124793 275937 124827 275971
rect 124861 275937 124957 275971
rect 122283 275846 122317 275937
rect 122283 275778 122317 275812
rect 124923 275846 124957 275937
rect 122283 275710 122317 275744
rect 124923 275778 124957 275812
rect 122283 275585 122317 275676
rect 124923 275710 124957 275744
rect 124923 275585 124957 275676
rect 122283 275551 122379 275585
rect 122413 275551 122447 275585
rect 122481 275551 122515 275585
rect 122549 275551 122583 275585
rect 122617 275551 122651 275585
rect 122685 275551 122719 275585
rect 122753 275551 122787 275585
rect 122821 275551 122855 275585
rect 122889 275551 122923 275585
rect 122957 275551 122991 275585
rect 123025 275551 123059 275585
rect 123093 275551 123127 275585
rect 123161 275551 123195 275585
rect 123229 275551 123263 275585
rect 123297 275551 123331 275585
rect 123365 275551 123399 275585
rect 123433 275551 123467 275585
rect 123501 275551 123535 275585
rect 123569 275551 123603 275585
rect 123637 275551 123671 275585
rect 123705 275551 123739 275585
rect 123773 275551 123807 275585
rect 123841 275551 123875 275585
rect 123909 275551 123943 275585
rect 123977 275551 124011 275585
rect 124045 275551 124079 275585
rect 124113 275551 124147 275585
rect 124181 275551 124215 275585
rect 124249 275551 124283 275585
rect 124317 275551 124351 275585
rect 124385 275551 124419 275585
rect 124453 275551 124487 275585
rect 124521 275551 124555 275585
rect 124589 275551 124623 275585
rect 124657 275551 124691 275585
rect 124725 275551 124759 275585
rect 124793 275551 124827 275585
rect 124861 275551 124957 275585
rect 121694 275422 121728 275456
rect 121694 275354 121728 275388
rect 121694 275286 121728 275320
rect 121694 275218 121728 275252
rect 121694 275150 121728 275184
rect 121694 275082 121728 275116
rect 120237 275014 120271 275048
rect 120237 274946 120271 274980
rect 121694 275014 121728 275048
rect 120237 274878 120271 274912
rect 121694 274946 121728 274980
rect 121694 274878 121728 274912
rect 120237 274810 120271 274844
rect 120237 274742 120271 274776
rect 121694 274810 121728 274844
rect 120237 274674 120271 274708
rect 120237 274606 120271 274640
rect 120237 274538 120271 274572
rect 120237 274470 120271 274504
rect 120237 274402 120271 274436
rect 120237 274334 120271 274368
rect 120237 274266 120271 274300
rect 121694 274742 121728 274776
rect 121694 274674 121728 274708
rect 121694 274606 121728 274640
rect 121694 274538 121728 274572
rect 121694 274470 121728 274504
rect 121694 274402 121728 274436
rect 121694 274334 121728 274368
rect 121694 274266 121728 274300
rect 120237 274198 120271 274232
rect 121694 274198 121728 274232
rect 120237 274130 120271 274164
rect 120237 274062 120271 274096
rect 121694 274130 121728 274164
rect 120237 273994 120271 274028
rect 121694 274062 121728 274096
rect 121694 273994 121728 274028
rect 120237 273926 120271 273960
rect 120237 273858 120271 273892
rect 120237 273790 120271 273824
rect 120237 273722 120271 273756
rect 120237 273654 120271 273688
rect 120237 273586 120271 273620
rect 120237 273518 120271 273552
rect 120237 273450 120271 273484
rect 121694 273926 121728 273960
rect 121694 273858 121728 273892
rect 121694 273790 121728 273824
rect 121694 273722 121728 273756
rect 121694 273654 121728 273688
rect 121694 273586 121728 273620
rect 121694 273518 121728 273552
rect 120237 273382 120271 273416
rect 121694 273450 121728 273484
rect 120237 273314 120271 273348
rect 121694 273382 121728 273416
rect 121694 273314 121728 273348
rect 120237 273246 120271 273280
rect 120237 273178 120271 273212
rect 121694 273246 121728 273280
rect 120237 273110 120271 273144
rect 120237 273042 120271 273076
rect 120237 272974 120271 273008
rect 120237 272906 120271 272940
rect 120237 272838 120271 272872
rect 120237 272770 120271 272804
rect 120237 272702 120271 272736
rect 121694 273178 121728 273212
rect 121694 273110 121728 273144
rect 121694 273042 121728 273076
rect 121694 272974 121728 273008
rect 121694 272906 121728 272940
rect 121694 272838 121728 272872
rect 121694 272770 121728 272804
rect 121694 272702 121728 272736
rect 120237 272634 120271 272668
rect 121694 272634 121728 272668
rect 120237 272566 120271 272600
rect 120237 272498 120271 272532
rect 121694 272566 121728 272600
rect 120237 272430 120271 272464
rect 121694 272498 121728 272532
rect 121694 272430 121728 272464
rect 120237 272362 120271 272396
rect 120237 272294 120271 272328
rect 120237 272226 120271 272260
rect 120237 272158 120271 272192
rect 120237 272090 120271 272124
rect 120237 272022 120271 272056
rect 120237 271954 120271 271988
rect 120237 271886 120271 271920
rect 121694 272362 121728 272396
rect 121694 272294 121728 272328
rect 121694 272226 121728 272260
rect 121694 272158 121728 272192
rect 121694 272090 121728 272124
rect 121694 272022 121728 272056
rect 121694 271954 121728 271988
rect 120237 271818 120271 271852
rect 121694 271886 121728 271920
rect 121694 271818 121728 271852
rect 120237 271750 120271 271784
rect 121694 271750 121728 271784
rect 120237 271682 120271 271716
rect 120237 271614 120271 271648
rect 121694 271682 121728 271716
rect 120237 271546 120271 271580
rect 120237 271478 120271 271512
rect 120237 271410 120271 271444
rect 120237 271342 120271 271376
rect 120237 271274 120271 271308
rect 120237 271206 120271 271240
rect 120237 271138 120271 271172
rect 121694 271614 121728 271648
rect 121694 271546 121728 271580
rect 121694 271478 121728 271512
rect 121694 271410 121728 271444
rect 121694 271342 121728 271376
rect 121694 271274 121728 271308
rect 121694 271206 121728 271240
rect 121694 271138 121728 271172
rect 120237 271070 120271 271104
rect 120237 271002 120271 271036
rect 121694 271070 121728 271104
rect 120237 270934 120271 270968
rect 121694 271002 121728 271036
rect 120237 270866 120271 270900
rect 121694 270934 121728 270968
rect 121694 270866 121728 270900
rect 120237 270798 120271 270832
rect 120237 270730 120271 270764
rect 120237 270662 120271 270696
rect 120237 270594 120271 270628
rect 120237 270526 120271 270560
rect 120237 270458 120271 270492
rect 120237 270390 120271 270424
rect 120237 270322 120271 270356
rect 121694 270798 121728 270832
rect 121694 270730 121728 270764
rect 121694 270662 121728 270696
rect 121694 270594 121728 270628
rect 121694 270526 121728 270560
rect 121694 270458 121728 270492
rect 121694 270390 121728 270424
rect 120237 270254 120271 270288
rect 121694 270322 121728 270356
rect 121694 270254 121728 270288
rect 120237 270186 120271 270220
rect 121694 270186 121728 270220
rect 120237 270118 120271 270152
rect 120237 270050 120271 270084
rect 121694 270118 121728 270152
rect 120237 269982 120271 270016
rect 120237 269914 120271 269948
rect 120237 269846 120271 269880
rect 120237 269778 120271 269812
rect 120237 269710 120271 269744
rect 120237 269642 120271 269676
rect 120237 269574 120271 269608
rect 121694 270050 121728 270084
rect 121694 269982 121728 270016
rect 121694 269914 121728 269948
rect 121694 269846 121728 269880
rect 121694 269778 121728 269812
rect 121694 269710 121728 269744
rect 121694 269642 121728 269676
rect 121694 269574 121728 269608
rect 120237 269506 120271 269540
rect 120237 269438 120271 269472
rect 121694 269506 121728 269540
rect 120237 269370 120271 269404
rect 121694 269438 121728 269472
rect 120237 269302 120271 269336
rect 121694 269370 121728 269404
rect 121694 269302 121728 269336
rect 120237 269234 120271 269268
rect 120237 269166 120271 269200
rect 121694 269234 121728 269268
rect 120237 269098 120271 269132
rect 121694 269166 121728 269200
rect 121694 269098 121728 269132
rect 120237 269012 120271 269064
rect 121694 269012 121728 269064
rect 120237 268978 120319 269012
rect 120353 268978 120387 269012
rect 120421 268978 120455 269012
rect 120489 268978 120523 269012
rect 120557 268978 120591 269012
rect 120625 268978 120659 269012
rect 120693 268978 120727 269012
rect 120761 268978 120795 269012
rect 120829 268978 120863 269012
rect 120897 268978 120931 269012
rect 120965 268978 120999 269012
rect 121033 268978 121067 269012
rect 121101 268978 121135 269012
rect 121169 268978 121203 269012
rect 121237 268978 121271 269012
rect 121305 268978 121339 269012
rect 121373 268978 121407 269012
rect 121441 268978 121475 269012
rect 121509 268978 121543 269012
rect 121577 268978 121611 269012
rect 121645 268978 121728 269012
rect 121920 272964 122006 272998
rect 122040 272964 122074 272998
rect 122108 272964 122142 272998
rect 122176 272964 122210 272998
rect 122244 272964 122278 272998
rect 122312 272964 122346 272998
rect 122380 272964 122414 272998
rect 122448 272964 122482 272998
rect 122516 272964 122550 272998
rect 122584 272964 122618 272998
rect 122652 272964 122686 272998
rect 122720 272964 122754 272998
rect 122788 272964 122822 272998
rect 122856 272964 122890 272998
rect 122924 272964 122958 272998
rect 122992 272964 123026 272998
rect 123060 272964 123094 272998
rect 123128 272964 123162 272998
rect 123196 272964 123230 272998
rect 123264 272964 123298 272998
rect 123332 272964 123366 272998
rect 123400 272964 123434 272998
rect 123468 272964 123554 272998
rect 121920 272917 121954 272964
rect 123520 272917 123554 272964
rect 121920 272849 121954 272883
rect 121920 272781 121954 272815
rect 123520 272849 123554 272883
rect 121920 272713 121954 272747
rect 123520 272781 123554 272815
rect 123520 272713 123554 272747
rect 121920 272645 121954 272679
rect 123520 272645 123554 272679
rect 121920 272577 121954 272611
rect 121920 272509 121954 272543
rect 123520 272577 123554 272611
rect 121920 272441 121954 272475
rect 123520 272509 123554 272543
rect 123520 272441 123554 272475
rect 121920 272373 121954 272407
rect 121920 272305 121954 272339
rect 121920 272237 121954 272271
rect 121920 272169 121954 272203
rect 121920 272101 121954 272135
rect 121920 272033 121954 272067
rect 121920 271965 121954 271999
rect 121920 271897 121954 271931
rect 123520 272373 123554 272407
rect 123520 272305 123554 272339
rect 123520 272237 123554 272271
rect 123520 272169 123554 272203
rect 123520 272101 123554 272135
rect 123520 272033 123554 272067
rect 123520 271965 123554 271999
rect 121920 271829 121954 271863
rect 123520 271897 123554 271931
rect 121920 271761 121954 271795
rect 123520 271829 123554 271863
rect 123520 271761 123554 271795
rect 121920 271693 121954 271727
rect 121920 271625 121954 271659
rect 123520 271693 123554 271727
rect 121920 271557 121954 271591
rect 121920 271489 121954 271523
rect 121920 271421 121954 271455
rect 121920 271353 121954 271387
rect 121920 271285 121954 271319
rect 121920 271217 121954 271251
rect 121920 271149 121954 271183
rect 123520 271625 123554 271659
rect 123520 271557 123554 271591
rect 123520 271489 123554 271523
rect 123520 271421 123554 271455
rect 123520 271353 123554 271387
rect 123520 271285 123554 271319
rect 123520 271217 123554 271251
rect 123520 271149 123554 271183
rect 121920 271081 121954 271115
rect 123520 271081 123554 271115
rect 121920 271013 121954 271047
rect 121920 270945 121954 270979
rect 123520 271013 123554 271047
rect 121920 270877 121954 270911
rect 123520 270945 123554 270979
rect 123520 270877 123554 270911
rect 121920 270809 121954 270843
rect 121920 270741 121954 270775
rect 121920 270673 121954 270707
rect 121920 270605 121954 270639
rect 121920 270537 121954 270571
rect 121920 270469 121954 270503
rect 121920 270401 121954 270435
rect 121920 270333 121954 270367
rect 123520 270809 123554 270843
rect 123520 270741 123554 270775
rect 123520 270673 123554 270707
rect 123520 270605 123554 270639
rect 123520 270537 123554 270571
rect 123520 270469 123554 270503
rect 123520 270401 123554 270435
rect 121920 270265 121954 270299
rect 123520 270333 123554 270367
rect 123520 270265 123554 270299
rect 121920 270197 121954 270231
rect 123520 270197 123554 270231
rect 121920 270129 121954 270163
rect 121920 270061 121954 270095
rect 123520 270129 123554 270163
rect 121920 269993 121954 270027
rect 121920 269925 121954 269959
rect 121920 269857 121954 269891
rect 121920 269789 121954 269823
rect 121920 269721 121954 269755
rect 121920 269653 121954 269687
rect 121920 269585 121954 269619
rect 123520 270061 123554 270095
rect 123520 269993 123554 270027
rect 123520 269925 123554 269959
rect 123520 269857 123554 269891
rect 123520 269789 123554 269823
rect 123520 269721 123554 269755
rect 123520 269653 123554 269687
rect 123520 269585 123554 269619
rect 121920 269517 121954 269551
rect 121920 269449 121954 269483
rect 123520 269517 123554 269551
rect 121920 269381 121954 269415
rect 123520 269449 123554 269483
rect 121920 269313 121954 269347
rect 123520 269381 123554 269415
rect 123520 269313 123554 269347
rect 121920 269245 121954 269279
rect 121920 269177 121954 269211
rect 123520 269245 123554 269279
rect 121920 269109 121954 269143
rect 123520 269177 123554 269211
rect 123520 269109 123554 269143
rect 121920 269028 121954 269075
rect 123520 269028 123554 269075
rect 121920 268994 122006 269028
rect 122040 268994 122074 269028
rect 122108 268994 122142 269028
rect 122176 268994 122210 269028
rect 122244 268994 122278 269028
rect 122312 268994 122346 269028
rect 122380 268994 122414 269028
rect 122448 268994 122482 269028
rect 122516 268994 122550 269028
rect 122584 268994 122618 269028
rect 122652 268994 122686 269028
rect 122720 268994 122754 269028
rect 122788 268994 122822 269028
rect 122856 268994 122890 269028
rect 122924 268994 122958 269028
rect 122992 268994 123026 269028
rect 123060 268994 123094 269028
rect 123128 268994 123162 269028
rect 123196 268994 123230 269028
rect 123264 268994 123298 269028
rect 123332 268994 123366 269028
rect 123400 268994 123434 269028
rect 123468 268994 123554 269028
<< psubdiffcont >>
rect 111264 281122 111298 281156
rect 111332 281122 111366 281156
rect 111400 281122 111434 281156
rect 111468 281122 111502 281156
rect 111536 281122 111570 281156
rect 111604 281122 111638 281156
rect 111672 281122 111706 281156
rect 111740 281122 111774 281156
rect 111808 281122 111842 281156
rect 111876 281122 111910 281156
rect 111944 281122 111978 281156
rect 112012 281122 112046 281156
rect 112080 281122 112114 281156
rect 112148 281122 112182 281156
rect 112216 281122 112250 281156
rect 112284 281122 112318 281156
rect 112352 281122 112386 281156
rect 112420 281122 112454 281156
rect 112488 281122 112522 281156
rect 112556 281122 112590 281156
rect 112624 281122 112658 281156
rect 112692 281122 112726 281156
rect 112760 281122 112794 281156
rect 112828 281122 112862 281156
rect 112896 281122 112930 281156
rect 112964 281122 112998 281156
rect 113032 281122 113066 281156
rect 113100 281122 113134 281156
rect 113168 281122 113202 281156
rect 113236 281122 113270 281156
rect 113304 281122 113338 281156
rect 113372 281122 113406 281156
rect 113440 281122 113474 281156
rect 113508 281122 113542 281156
rect 113576 281122 113610 281156
rect 113644 281122 113678 281156
rect 113712 281122 113746 281156
rect 113780 281122 113814 281156
rect 113848 281122 113882 281156
rect 113916 281122 113950 281156
rect 113984 281122 114018 281156
rect 114052 281122 114086 281156
rect 114120 281122 114154 281156
rect 114188 281122 114222 281156
rect 114256 281122 114290 281156
rect 114324 281122 114358 281156
rect 114392 281122 114426 281156
rect 114460 281122 114494 281156
rect 114528 281122 114562 281156
rect 114596 281122 114630 281156
rect 114664 281122 114698 281156
rect 114732 281122 114766 281156
rect 114800 281122 114834 281156
rect 114868 281122 114902 281156
rect 114936 281122 114970 281156
rect 115004 281122 115038 281156
rect 115072 281122 115106 281156
rect 115140 281122 115174 281156
rect 115208 281122 115242 281156
rect 115276 281122 115310 281156
rect 115344 281122 115378 281156
rect 115412 281122 115446 281156
rect 115480 281122 115514 281156
rect 115548 281122 115582 281156
rect 115616 281122 115650 281156
rect 115684 281122 115718 281156
rect 115752 281122 115786 281156
rect 115820 281122 115854 281156
rect 115888 281122 115922 281156
rect 115956 281122 115990 281156
rect 116024 281122 116058 281156
rect 116092 281122 116126 281156
rect 116160 281122 116194 281156
rect 116228 281122 116262 281156
rect 116296 281122 116330 281156
rect 116364 281122 116398 281156
rect 116432 281122 116466 281156
rect 116500 281122 116534 281156
rect 116568 281122 116602 281156
rect 116636 281122 116670 281156
rect 116704 281122 116738 281156
rect 116772 281122 116806 281156
rect 116840 281122 116874 281156
rect 116908 281122 116942 281156
rect 116976 281122 117010 281156
rect 117044 281122 117078 281156
rect 117112 281122 117146 281156
rect 117180 281122 117214 281156
rect 117248 281122 117282 281156
rect 117316 281122 117350 281156
rect 117384 281122 117418 281156
rect 117452 281122 117486 281156
rect 117520 281122 117554 281156
rect 117588 281122 117622 281156
rect 117656 281122 117690 281156
rect 117724 281122 117758 281156
rect 117792 281122 117826 281156
rect 117860 281122 117894 281156
rect 117928 281122 117962 281156
rect 117996 281122 118030 281156
rect 118064 281122 118098 281156
rect 118132 281122 118166 281156
rect 118200 281122 118234 281156
rect 118268 281122 118302 281156
rect 118336 281122 118370 281156
rect 118404 281122 118438 281156
rect 118472 281122 118506 281156
rect 118540 281122 118574 281156
rect 118608 281122 118642 281156
rect 118676 281122 118710 281156
rect 118744 281122 118778 281156
rect 118812 281122 118846 281156
rect 106000 280983 106034 281017
rect 106176 280986 106210 281020
rect 106244 280986 106278 281020
rect 106312 280986 106346 281020
rect 106380 280986 106414 281020
rect 106448 280986 106482 281020
rect 106516 280986 106550 281020
rect 106584 280986 106618 281020
rect 106652 280986 106686 281020
rect 106720 280986 106754 281020
rect 106788 280986 106822 281020
rect 106856 280986 106890 281020
rect 106924 280986 106958 281020
rect 106992 280986 107026 281020
rect 107060 280986 107094 281020
rect 107128 280986 107162 281020
rect 107196 280986 107230 281020
rect 107264 280986 107298 281020
rect 107332 280986 107366 281020
rect 107400 280986 107434 281020
rect 107468 280986 107502 281020
rect 107536 280986 107570 281020
rect 107604 280986 107638 281020
rect 107672 280986 107706 281020
rect 107740 280986 107774 281020
rect 107808 280986 107842 281020
rect 107876 280986 107910 281020
rect 107944 280986 107978 281020
rect 108012 280986 108046 281020
rect 108080 280986 108114 281020
rect 108148 280986 108182 281020
rect 108216 280986 108250 281020
rect 108284 280986 108318 281020
rect 108352 280986 108386 281020
rect 108420 280986 108454 281020
rect 108488 280986 108522 281020
rect 108556 280986 108590 281020
rect 108624 280986 108658 281020
rect 108692 280986 108726 281020
rect 108760 280986 108794 281020
rect 108828 280986 108862 281020
rect 108896 280986 108930 281020
rect 108964 280986 108998 281020
rect 109032 280986 109066 281020
rect 109100 280986 109134 281020
rect 109168 280986 109202 281020
rect 109236 280986 109270 281020
rect 109304 280986 109338 281020
rect 109372 280986 109406 281020
rect 109440 280986 109474 281020
rect 109508 280986 109542 281020
rect 109576 280986 109610 281020
rect 109644 280986 109678 281020
rect 109712 280986 109746 281020
rect 109780 280986 109814 281020
rect 109848 280986 109882 281020
rect 109916 280986 109950 281020
rect 109984 280986 110018 281020
rect 110052 280986 110086 281020
rect 110120 280986 110154 281020
rect 110188 280986 110222 281020
rect 106000 280915 106034 280949
rect 106000 280847 106034 280881
rect 106149 280825 106183 280859
rect 106000 280779 106034 280813
rect 106149 280757 106183 280791
rect 106000 280711 106034 280745
rect 106149 280689 106183 280723
rect 106000 280643 106034 280677
rect 106149 280621 106183 280655
rect 106000 280575 106034 280609
rect 106149 280553 106183 280587
rect 106000 280507 106034 280541
rect 106149 280485 106183 280519
rect 106000 280439 106034 280473
rect 106149 280417 106183 280451
rect 106000 280371 106034 280405
rect 106149 280349 106183 280383
rect 106000 280303 106034 280337
rect 106149 280281 106183 280315
rect 106000 280235 106034 280269
rect 106149 280213 106183 280247
rect 106000 280167 106034 280201
rect 106149 280145 106183 280179
rect 106000 280099 106034 280133
rect 106149 280077 106183 280111
rect 106000 280031 106034 280065
rect 106149 280009 106183 280043
rect 106000 279963 106034 279997
rect 106149 279941 106183 279975
rect 106000 279895 106034 279929
rect 106149 279873 106183 279907
rect 106000 279827 106034 279861
rect 106149 279805 106183 279839
rect 110255 280807 110289 280841
rect 110255 280739 110289 280773
rect 110255 280671 110289 280705
rect 110255 280603 110289 280637
rect 110255 280535 110289 280569
rect 110255 280467 110289 280501
rect 110255 280399 110289 280433
rect 110255 280331 110289 280365
rect 110255 280263 110289 280297
rect 110255 280195 110289 280229
rect 110255 280127 110289 280161
rect 110255 280059 110289 280093
rect 110255 279991 110289 280025
rect 110255 279923 110289 279957
rect 110255 279855 110289 279889
rect 106000 279759 106034 279793
rect 106149 279737 106183 279771
rect 106000 279691 106034 279725
rect 110255 279787 110289 279821
rect 110255 279719 110289 279753
rect 106000 279623 106034 279657
rect 106000 279555 106034 279589
rect 106176 279566 106210 279600
rect 106244 279566 106278 279600
rect 106312 279566 106346 279600
rect 106380 279566 106414 279600
rect 106448 279566 106482 279600
rect 106516 279566 106550 279600
rect 106584 279566 106618 279600
rect 106652 279566 106686 279600
rect 106720 279566 106754 279600
rect 106788 279566 106822 279600
rect 106856 279566 106890 279600
rect 106924 279566 106958 279600
rect 106992 279566 107026 279600
rect 107060 279566 107094 279600
rect 107128 279566 107162 279600
rect 107196 279566 107230 279600
rect 107264 279566 107298 279600
rect 107332 279566 107366 279600
rect 107400 279566 107434 279600
rect 107468 279566 107502 279600
rect 107536 279566 107570 279600
rect 107604 279566 107638 279600
rect 107672 279566 107706 279600
rect 107740 279566 107774 279600
rect 107808 279566 107842 279600
rect 107876 279566 107910 279600
rect 107944 279566 107978 279600
rect 108012 279566 108046 279600
rect 108080 279566 108114 279600
rect 108148 279566 108182 279600
rect 108216 279566 108250 279600
rect 108284 279566 108318 279600
rect 108352 279566 108386 279600
rect 108420 279566 108454 279600
rect 108488 279566 108522 279600
rect 108556 279566 108590 279600
rect 108624 279566 108658 279600
rect 108692 279566 108726 279600
rect 108760 279566 108794 279600
rect 108828 279566 108862 279600
rect 108896 279566 108930 279600
rect 108964 279566 108998 279600
rect 109032 279566 109066 279600
rect 109100 279566 109134 279600
rect 109168 279566 109202 279600
rect 109236 279566 109270 279600
rect 109304 279566 109338 279600
rect 109372 279566 109406 279600
rect 109440 279566 109474 279600
rect 109508 279566 109542 279600
rect 109576 279566 109610 279600
rect 109644 279566 109678 279600
rect 109712 279566 109746 279600
rect 109780 279566 109814 279600
rect 109848 279566 109882 279600
rect 109916 279566 109950 279600
rect 109984 279566 110018 279600
rect 110052 279566 110086 279600
rect 110120 279566 110154 279600
rect 110188 279566 110222 279600
rect 106000 279487 106034 279521
rect 106000 279419 106034 279453
rect 106000 279351 106034 279385
rect 106000 279283 106034 279317
rect 106000 279215 106034 279249
rect 106000 279147 106034 279181
rect 106000 279079 106034 279113
rect 106000 279011 106034 279045
rect 106000 278943 106034 278977
rect 106000 278875 106034 278909
rect 106000 278807 106034 278841
rect 106000 278739 106034 278773
rect 106000 278671 106034 278705
rect 106000 278603 106034 278637
rect 106000 278535 106034 278569
rect 106000 278467 106034 278501
rect 106000 278399 106034 278433
rect 106000 278331 106034 278365
rect 106000 278263 106034 278297
rect 106000 278195 106034 278229
rect 106000 278127 106034 278161
rect 106000 278059 106034 278093
rect 106000 277991 106034 278025
rect 106000 277923 106034 277957
rect 109733 279151 109767 279185
rect 109801 279151 109835 279185
rect 109869 279151 109903 279185
rect 109937 279151 109971 279185
rect 110005 279151 110039 279185
rect 110073 279151 110107 279185
rect 109617 279037 109651 279071
rect 110189 279037 110223 279071
rect 109617 278969 109651 279003
rect 109617 278901 109651 278935
rect 109617 278833 109651 278867
rect 109617 278765 109651 278799
rect 109617 278697 109651 278731
rect 109617 278629 109651 278663
rect 109617 278561 109651 278595
rect 109617 278493 109651 278527
rect 109617 278425 109651 278459
rect 109617 278357 109651 278391
rect 109617 278289 109651 278323
rect 109617 278221 109651 278255
rect 109617 278153 109651 278187
rect 109617 278085 109651 278119
rect 109617 278017 109651 278051
rect 106000 277855 106034 277889
rect 106000 277787 106034 277821
rect 106000 277719 106034 277753
rect 106000 277651 106034 277685
rect 106000 277583 106034 277617
rect 106000 277515 106034 277549
rect 106000 277447 106034 277481
rect 106000 277379 106034 277413
rect 106000 277311 106034 277345
rect 109617 277949 109651 277983
rect 110189 278969 110223 279003
rect 110189 278901 110223 278935
rect 110189 278833 110223 278867
rect 110189 278765 110223 278799
rect 110189 278697 110223 278731
rect 110189 278629 110223 278663
rect 110189 278561 110223 278595
rect 110189 278493 110223 278527
rect 110189 278425 110223 278459
rect 110189 278357 110223 278391
rect 110189 278289 110223 278323
rect 110189 278221 110223 278255
rect 110189 278153 110223 278187
rect 110189 278085 110223 278119
rect 110189 278017 110223 278051
rect 109617 277881 109651 277915
rect 110189 277949 110223 277983
rect 109617 277813 109651 277847
rect 110189 277881 110223 277915
rect 109617 277745 109651 277779
rect 110189 277813 110223 277847
rect 109617 277677 109651 277711
rect 109617 277609 109651 277643
rect 109617 277541 109651 277575
rect 109617 277473 109651 277507
rect 109617 277405 109651 277439
rect 109617 277337 109651 277371
rect 106000 277243 106034 277277
rect 106000 277175 106034 277209
rect 106000 277107 106034 277141
rect 106000 277039 106034 277073
rect 106000 276971 106034 277005
rect 106000 276903 106034 276937
rect 109617 277269 109651 277303
rect 109617 277201 109651 277235
rect 109617 277133 109651 277167
rect 109617 277065 109651 277099
rect 109617 276997 109651 277031
rect 106000 276835 106034 276869
rect 106000 276767 106034 276801
rect 106000 276699 106034 276733
rect 106000 276631 106034 276665
rect 106000 276563 106034 276597
rect 109617 276929 109651 276963
rect 109617 276861 109651 276895
rect 109617 276793 109651 276827
rect 109617 276725 109651 276759
rect 110189 277745 110223 277779
rect 110189 277677 110223 277711
rect 110189 277609 110223 277643
rect 110189 277541 110223 277575
rect 110189 277473 110223 277507
rect 110189 277405 110223 277439
rect 110189 277337 110223 277371
rect 110189 277269 110223 277303
rect 110189 277201 110223 277235
rect 110189 277133 110223 277167
rect 110189 277065 110223 277099
rect 110189 276997 110223 277031
rect 110189 276929 110223 276963
rect 110189 276861 110223 276895
rect 110189 276793 110223 276827
rect 110189 276725 110223 276759
rect 109617 276657 109651 276691
rect 110189 276657 110223 276691
rect 109733 276543 109767 276577
rect 109801 276543 109835 276577
rect 109869 276543 109903 276577
rect 109937 276543 109971 276577
rect 110005 276543 110039 276577
rect 110073 276543 110107 276577
rect 106000 276495 106034 276529
rect 106000 276427 106034 276461
rect 106000 276359 106034 276393
rect 106000 276291 106034 276325
rect 106000 276223 106034 276257
rect 106000 276155 106034 276189
rect 106000 276087 106034 276121
rect 106000 276019 106034 276053
rect 106000 275951 106034 275985
rect 110167 275991 110201 276025
rect 106000 275883 106034 275917
rect 106000 275815 106034 275849
rect 106000 275747 106034 275781
rect 106000 275679 106034 275713
rect 106000 275611 106034 275645
rect 106000 275543 106034 275577
rect 106000 275475 106034 275509
rect 106000 275407 106034 275441
rect 106000 275339 106034 275373
rect 106000 275271 106034 275305
rect 106000 275203 106034 275237
rect 106000 275135 106034 275169
rect 106000 275067 106034 275101
rect 106000 274999 106034 275033
rect 106000 274931 106034 274965
rect 106000 274863 106034 274897
rect 106000 274795 106034 274829
rect 106000 274727 106034 274761
rect 110167 275923 110201 275957
rect 110167 275855 110201 275889
rect 110167 275787 110201 275821
rect 110167 275719 110201 275753
rect 110167 275651 110201 275685
rect 110167 275583 110201 275617
rect 110167 275515 110201 275549
rect 110167 275447 110201 275481
rect 110167 275379 110201 275413
rect 110167 275311 110201 275345
rect 110167 275243 110201 275277
rect 110167 275175 110201 275209
rect 110167 275107 110201 275141
rect 110167 275039 110201 275073
rect 110167 274971 110201 275005
rect 110167 274903 110201 274937
rect 110167 274835 110201 274869
rect 110167 274767 110201 274801
rect 106000 274659 106034 274693
rect 110167 274699 110201 274733
rect 106117 274556 106151 274590
rect 106185 274556 106219 274590
rect 106253 274556 106287 274590
rect 106321 274556 106355 274590
rect 106389 274556 106423 274590
rect 106457 274556 106491 274590
rect 106525 274556 106559 274590
rect 106593 274556 106627 274590
rect 106661 274556 106695 274590
rect 106729 274556 106763 274590
rect 106797 274556 106831 274590
rect 106865 274556 106899 274590
rect 106933 274556 106967 274590
rect 107001 274556 107035 274590
rect 107069 274556 107103 274590
rect 107137 274556 107171 274590
rect 107205 274556 107239 274590
rect 107273 274556 107307 274590
rect 107341 274556 107375 274590
rect 107409 274556 107443 274590
rect 107477 274556 107511 274590
rect 107545 274556 107579 274590
rect 107613 274556 107647 274590
rect 107681 274556 107715 274590
rect 107749 274556 107783 274590
rect 107817 274556 107851 274590
rect 107885 274556 107919 274590
rect 107953 274556 107987 274590
rect 108021 274556 108055 274590
rect 108089 274556 108123 274590
rect 108157 274556 108191 274590
rect 108225 274556 108259 274590
rect 108293 274556 108327 274590
rect 108361 274556 108395 274590
rect 108429 274556 108463 274590
rect 108497 274556 108531 274590
rect 108565 274556 108599 274590
rect 108633 274556 108667 274590
rect 108701 274556 108735 274590
rect 108769 274556 108803 274590
rect 108837 274556 108871 274590
rect 108905 274556 108939 274590
rect 108973 274556 109007 274590
rect 109041 274556 109075 274590
rect 109109 274556 109143 274590
rect 109177 274556 109211 274590
rect 109245 274556 109279 274590
rect 109313 274556 109347 274590
rect 109381 274556 109415 274590
rect 109449 274556 109483 274590
rect 109517 274556 109551 274590
rect 109585 274556 109619 274590
rect 109653 274556 109687 274590
rect 109721 274556 109755 274590
rect 109789 274556 109823 274590
rect 109857 274556 109891 274590
rect 109925 274556 109959 274590
rect 109993 274556 110027 274590
rect 110061 274556 110095 274590
rect 110129 274556 110163 274590
rect 106285 270212 106455 272898
rect 106595 272821 109961 272923
rect 106735 272287 106769 272321
rect 106848 272316 106882 272350
rect 106977 272316 107011 272350
rect 107045 272316 107079 272350
rect 107113 272316 107147 272350
rect 107181 272316 107215 272350
rect 107249 272316 107283 272350
rect 107317 272316 107351 272350
rect 107385 272316 107419 272350
rect 107453 272316 107487 272350
rect 107521 272316 107555 272350
rect 107589 272316 107623 272350
rect 107657 272316 107691 272350
rect 107725 272316 107759 272350
rect 107793 272316 107827 272350
rect 107861 272316 107895 272350
rect 107929 272316 107963 272350
rect 107997 272316 108031 272350
rect 108065 272316 108099 272350
rect 108133 272316 108167 272350
rect 108201 272316 108235 272350
rect 108269 272316 108303 272350
rect 108337 272316 108371 272350
rect 108405 272316 108439 272350
rect 108473 272316 108507 272350
rect 108541 272316 108575 272350
rect 108609 272316 108643 272350
rect 106735 272219 106769 272253
rect 106735 272151 106769 272185
rect 108749 272287 108783 272321
rect 108749 272219 108783 272253
rect 106735 272083 106769 272117
rect 108749 272151 108783 272185
rect 108749 272083 108783 272117
rect 106735 272015 106769 272049
rect 106735 271947 106769 271981
rect 106735 271879 106769 271913
rect 106735 271811 106769 271845
rect 106735 271743 106769 271777
rect 108749 272015 108783 272049
rect 108749 271947 108783 271981
rect 108749 271879 108783 271913
rect 108749 271811 108783 271845
rect 108749 271743 108783 271777
rect 106735 271675 106769 271709
rect 108749 271675 108783 271709
rect 106735 271607 106769 271641
rect 106735 271539 106769 271573
rect 108749 271607 108783 271641
rect 106735 271471 106769 271505
rect 108749 271539 108783 271573
rect 106735 271403 106769 271437
rect 106735 271335 106769 271369
rect 108749 271471 108783 271505
rect 108749 271403 108783 271437
rect 108749 271335 108783 271369
rect 106735 271267 106769 271301
rect 108749 271267 108783 271301
rect 106735 271199 106769 271233
rect 108749 271199 108783 271233
rect 106735 271131 106769 271165
rect 108749 271131 108783 271165
rect 106735 271063 106769 271097
rect 106735 270995 106769 271029
rect 106735 270927 106769 270961
rect 108749 271063 108783 271097
rect 108749 270995 108783 271029
rect 106735 270859 106769 270893
rect 108749 270927 108783 270961
rect 106735 270791 106769 270825
rect 108749 270859 108783 270893
rect 108749 270791 108783 270825
rect 106875 270750 106909 270784
rect 106943 270750 106977 270784
rect 107011 270750 107045 270784
rect 107079 270750 107113 270784
rect 107147 270750 107181 270784
rect 107215 270750 107249 270784
rect 107283 270750 107317 270784
rect 107351 270750 107385 270784
rect 107419 270750 107453 270784
rect 107487 270750 107521 270784
rect 107555 270750 107589 270784
rect 107623 270750 107657 270784
rect 107691 270750 107725 270784
rect 107759 270750 107793 270784
rect 107827 270750 107861 270784
rect 107895 270750 107929 270784
rect 107963 270750 107997 270784
rect 108031 270750 108065 270784
rect 108099 270750 108133 270784
rect 108167 270750 108201 270784
rect 108235 270750 108269 270784
rect 108303 270750 108337 270784
rect 108371 270750 108405 270784
rect 108439 270750 108473 270784
rect 108507 270750 108541 270784
rect 108575 270750 108609 270784
rect 108643 270750 108677 270784
rect 106585 270204 109951 270306
rect 110085 270212 110255 272898
rect 111072 272704 111174 281102
rect 114243 280774 114345 280876
rect 111340 279363 111374 279397
rect 111408 279363 111442 279397
rect 111476 279363 111510 279397
rect 111544 279363 111578 279397
rect 111612 279363 111646 279397
rect 111680 279363 111714 279397
rect 111748 279363 111782 279397
rect 111816 279363 111850 279397
rect 111884 279363 111918 279397
rect 111952 279363 111986 279397
rect 112020 279363 112054 279397
rect 112088 279363 112122 279397
rect 112156 279363 112190 279397
rect 112224 279363 112258 279397
rect 112292 279363 112326 279397
rect 112360 279363 112394 279397
rect 112428 279363 112462 279397
rect 112496 279363 112530 279397
rect 112564 279363 112598 279397
rect 112632 279363 112666 279397
rect 112700 279363 112734 279397
rect 112768 279363 112802 279397
rect 112836 279363 112870 279397
rect 112904 279363 112938 279397
rect 112972 279363 113006 279397
rect 113040 279363 113074 279397
rect 113108 279363 113142 279397
rect 113176 279363 113210 279397
rect 113244 279363 113278 279397
rect 113312 279363 113346 279397
rect 113380 279363 113414 279397
rect 113448 279363 113482 279397
rect 113516 279363 113550 279397
rect 113584 279363 113618 279397
rect 113652 279363 113686 279397
rect 113720 279363 113754 279397
rect 113788 279363 113822 279397
rect 113856 279363 113890 279397
rect 113924 279363 113958 279397
rect 113992 279363 114026 279397
rect 114060 279363 114094 279397
rect 114128 279363 114162 279397
rect 114196 279363 114230 279397
rect 115860 280774 115962 280876
rect 115975 279363 116009 279397
rect 116043 279363 116077 279397
rect 116111 279363 116145 279397
rect 116179 279363 116213 279397
rect 116247 279363 116281 279397
rect 116315 279363 116349 279397
rect 116383 279363 116417 279397
rect 116451 279363 116485 279397
rect 116519 279363 116553 279397
rect 116587 279363 116621 279397
rect 116655 279363 116689 279397
rect 116723 279363 116757 279397
rect 116791 279363 116825 279397
rect 116859 279363 116893 279397
rect 116927 279363 116961 279397
rect 116995 279363 117029 279397
rect 117063 279363 117097 279397
rect 117131 279363 117165 279397
rect 117199 279363 117233 279397
rect 117267 279363 117301 279397
rect 117335 279363 117369 279397
rect 117403 279363 117437 279397
rect 117471 279363 117505 279397
rect 117539 279363 117573 279397
rect 117607 279363 117641 279397
rect 117675 279363 117709 279397
rect 117743 279363 117777 279397
rect 117811 279363 117845 279397
rect 117879 279363 117913 279397
rect 117947 279363 117981 279397
rect 118015 279363 118049 279397
rect 118083 279363 118117 279397
rect 118151 279363 118185 279397
rect 118219 279363 118253 279397
rect 118287 279363 118321 279397
rect 118355 279363 118389 279397
rect 118423 279363 118457 279397
rect 118491 279363 118525 279397
rect 118559 279363 118593 279397
rect 118627 279363 118661 279397
rect 118695 279363 118729 279397
rect 118763 279363 118797 279397
rect 118831 279363 118865 279397
rect 114243 279108 114345 279210
rect 111340 277697 111374 277731
rect 111408 277697 111442 277731
rect 111476 277697 111510 277731
rect 111544 277697 111578 277731
rect 111612 277697 111646 277731
rect 111680 277697 111714 277731
rect 111748 277697 111782 277731
rect 111816 277697 111850 277731
rect 111884 277697 111918 277731
rect 111952 277697 111986 277731
rect 112020 277697 112054 277731
rect 112088 277697 112122 277731
rect 112156 277697 112190 277731
rect 112224 277697 112258 277731
rect 112292 277697 112326 277731
rect 112360 277697 112394 277731
rect 112428 277697 112462 277731
rect 112496 277697 112530 277731
rect 112564 277697 112598 277731
rect 112632 277697 112666 277731
rect 112700 277697 112734 277731
rect 112768 277697 112802 277731
rect 112836 277697 112870 277731
rect 112904 277697 112938 277731
rect 112972 277697 113006 277731
rect 113040 277697 113074 277731
rect 113108 277697 113142 277731
rect 113176 277697 113210 277731
rect 113244 277697 113278 277731
rect 113312 277697 113346 277731
rect 113380 277697 113414 277731
rect 113448 277697 113482 277731
rect 113516 277697 113550 277731
rect 113584 277697 113618 277731
rect 113652 277697 113686 277731
rect 113720 277697 113754 277731
rect 113788 277697 113822 277731
rect 113856 277697 113890 277731
rect 113924 277697 113958 277731
rect 113992 277697 114026 277731
rect 114060 277697 114094 277731
rect 114128 277697 114162 277731
rect 114196 277697 114230 277731
rect 115860 279108 115962 279210
rect 115975 277697 116009 277731
rect 116043 277697 116077 277731
rect 116111 277697 116145 277731
rect 116179 277697 116213 277731
rect 116247 277697 116281 277731
rect 116315 277697 116349 277731
rect 116383 277697 116417 277731
rect 116451 277697 116485 277731
rect 116519 277697 116553 277731
rect 116587 277697 116621 277731
rect 116655 277697 116689 277731
rect 116723 277697 116757 277731
rect 116791 277697 116825 277731
rect 116859 277697 116893 277731
rect 116927 277697 116961 277731
rect 116995 277697 117029 277731
rect 117063 277697 117097 277731
rect 117131 277697 117165 277731
rect 117199 277697 117233 277731
rect 117267 277697 117301 277731
rect 117335 277697 117369 277731
rect 117403 277697 117437 277731
rect 117471 277697 117505 277731
rect 117539 277697 117573 277731
rect 117607 277697 117641 277731
rect 117675 277697 117709 277731
rect 117743 277697 117777 277731
rect 117811 277697 117845 277731
rect 117879 277697 117913 277731
rect 117947 277697 117981 277731
rect 118015 277697 118049 277731
rect 118083 277697 118117 277731
rect 118151 277697 118185 277731
rect 118219 277697 118253 277731
rect 118287 277697 118321 277731
rect 118355 277697 118389 277731
rect 118423 277697 118457 277731
rect 118491 277697 118525 277731
rect 118559 277697 118593 277731
rect 118627 277697 118661 277731
rect 118695 277697 118729 277731
rect 118763 277697 118797 277731
rect 118831 277697 118865 277731
rect 114243 277442 114345 277544
rect 111340 276031 111374 276065
rect 111408 276031 111442 276065
rect 111476 276031 111510 276065
rect 111544 276031 111578 276065
rect 111612 276031 111646 276065
rect 111680 276031 111714 276065
rect 111748 276031 111782 276065
rect 111816 276031 111850 276065
rect 111884 276031 111918 276065
rect 111952 276031 111986 276065
rect 112020 276031 112054 276065
rect 112088 276031 112122 276065
rect 112156 276031 112190 276065
rect 112224 276031 112258 276065
rect 112292 276031 112326 276065
rect 112360 276031 112394 276065
rect 112428 276031 112462 276065
rect 112496 276031 112530 276065
rect 112564 276031 112598 276065
rect 112632 276031 112666 276065
rect 112700 276031 112734 276065
rect 112768 276031 112802 276065
rect 112836 276031 112870 276065
rect 112904 276031 112938 276065
rect 112972 276031 113006 276065
rect 113040 276031 113074 276065
rect 113108 276031 113142 276065
rect 113176 276031 113210 276065
rect 113244 276031 113278 276065
rect 113312 276031 113346 276065
rect 113380 276031 113414 276065
rect 113448 276031 113482 276065
rect 113516 276031 113550 276065
rect 113584 276031 113618 276065
rect 113652 276031 113686 276065
rect 113720 276031 113754 276065
rect 113788 276031 113822 276065
rect 113856 276031 113890 276065
rect 113924 276031 113958 276065
rect 113992 276031 114026 276065
rect 114060 276031 114094 276065
rect 114128 276031 114162 276065
rect 114196 276031 114230 276065
rect 115860 277442 115962 277544
rect 115975 276031 116009 276065
rect 116043 276031 116077 276065
rect 116111 276031 116145 276065
rect 116179 276031 116213 276065
rect 116247 276031 116281 276065
rect 116315 276031 116349 276065
rect 116383 276031 116417 276065
rect 116451 276031 116485 276065
rect 116519 276031 116553 276065
rect 116587 276031 116621 276065
rect 116655 276031 116689 276065
rect 116723 276031 116757 276065
rect 116791 276031 116825 276065
rect 116859 276031 116893 276065
rect 116927 276031 116961 276065
rect 116995 276031 117029 276065
rect 117063 276031 117097 276065
rect 117131 276031 117165 276065
rect 117199 276031 117233 276065
rect 117267 276031 117301 276065
rect 117335 276031 117369 276065
rect 117403 276031 117437 276065
rect 117471 276031 117505 276065
rect 117539 276031 117573 276065
rect 117607 276031 117641 276065
rect 117675 276031 117709 276065
rect 117743 276031 117777 276065
rect 117811 276031 117845 276065
rect 117879 276031 117913 276065
rect 117947 276031 117981 276065
rect 118015 276031 118049 276065
rect 118083 276031 118117 276065
rect 118151 276031 118185 276065
rect 118219 276031 118253 276065
rect 118287 276031 118321 276065
rect 118355 276031 118389 276065
rect 118423 276031 118457 276065
rect 118491 276031 118525 276065
rect 118559 276031 118593 276065
rect 118627 276031 118661 276065
rect 118695 276031 118729 276065
rect 118763 276031 118797 276065
rect 118831 276031 118865 276065
rect 114243 275776 114345 275878
rect 111340 274365 111374 274399
rect 111408 274365 111442 274399
rect 111476 274365 111510 274399
rect 111544 274365 111578 274399
rect 111612 274365 111646 274399
rect 111680 274365 111714 274399
rect 111748 274365 111782 274399
rect 111816 274365 111850 274399
rect 111884 274365 111918 274399
rect 111952 274365 111986 274399
rect 112020 274365 112054 274399
rect 112088 274365 112122 274399
rect 112156 274365 112190 274399
rect 112224 274365 112258 274399
rect 112292 274365 112326 274399
rect 112360 274365 112394 274399
rect 112428 274365 112462 274399
rect 112496 274365 112530 274399
rect 112564 274365 112598 274399
rect 112632 274365 112666 274399
rect 112700 274365 112734 274399
rect 112768 274365 112802 274399
rect 112836 274365 112870 274399
rect 112904 274365 112938 274399
rect 112972 274365 113006 274399
rect 113040 274365 113074 274399
rect 113108 274365 113142 274399
rect 113176 274365 113210 274399
rect 113244 274365 113278 274399
rect 113312 274365 113346 274399
rect 113380 274365 113414 274399
rect 113448 274365 113482 274399
rect 113516 274365 113550 274399
rect 113584 274365 113618 274399
rect 113652 274365 113686 274399
rect 113720 274365 113754 274399
rect 113788 274365 113822 274399
rect 113856 274365 113890 274399
rect 113924 274365 113958 274399
rect 113992 274365 114026 274399
rect 114060 274365 114094 274399
rect 114128 274365 114162 274399
rect 114196 274365 114230 274399
rect 115860 275776 115962 275878
rect 115975 274365 116009 274399
rect 116043 274365 116077 274399
rect 116111 274365 116145 274399
rect 116179 274365 116213 274399
rect 116247 274365 116281 274399
rect 116315 274365 116349 274399
rect 116383 274365 116417 274399
rect 116451 274365 116485 274399
rect 116519 274365 116553 274399
rect 116587 274365 116621 274399
rect 116655 274365 116689 274399
rect 116723 274365 116757 274399
rect 116791 274365 116825 274399
rect 116859 274365 116893 274399
rect 116927 274365 116961 274399
rect 116995 274365 117029 274399
rect 117063 274365 117097 274399
rect 117131 274365 117165 274399
rect 117199 274365 117233 274399
rect 117267 274365 117301 274399
rect 117335 274365 117369 274399
rect 117403 274365 117437 274399
rect 117471 274365 117505 274399
rect 117539 274365 117573 274399
rect 117607 274365 117641 274399
rect 117675 274365 117709 274399
rect 117743 274365 117777 274399
rect 117811 274365 117845 274399
rect 117879 274365 117913 274399
rect 117947 274365 117981 274399
rect 118015 274365 118049 274399
rect 118083 274365 118117 274399
rect 118151 274365 118185 274399
rect 118219 274365 118253 274399
rect 118287 274365 118321 274399
rect 118355 274365 118389 274399
rect 118423 274365 118457 274399
rect 118491 274365 118525 274399
rect 118559 274365 118593 274399
rect 118627 274365 118661 274399
rect 118695 274365 118729 274399
rect 118763 274365 118797 274399
rect 118831 274365 118865 274399
rect 114243 274110 114345 274212
rect 111340 272699 111374 272733
rect 111408 272699 111442 272733
rect 111476 272699 111510 272733
rect 111544 272699 111578 272733
rect 111612 272699 111646 272733
rect 111680 272699 111714 272733
rect 111748 272699 111782 272733
rect 111816 272699 111850 272733
rect 111884 272699 111918 272733
rect 111952 272699 111986 272733
rect 112020 272699 112054 272733
rect 112088 272699 112122 272733
rect 112156 272699 112190 272733
rect 112224 272699 112258 272733
rect 112292 272699 112326 272733
rect 112360 272699 112394 272733
rect 112428 272699 112462 272733
rect 112496 272699 112530 272733
rect 112564 272699 112598 272733
rect 112632 272699 112666 272733
rect 112700 272699 112734 272733
rect 112768 272699 112802 272733
rect 112836 272699 112870 272733
rect 112904 272699 112938 272733
rect 112972 272699 113006 272733
rect 113040 272699 113074 272733
rect 113108 272699 113142 272733
rect 113176 272699 113210 272733
rect 113244 272699 113278 272733
rect 113312 272699 113346 272733
rect 113380 272699 113414 272733
rect 113448 272699 113482 272733
rect 113516 272699 113550 272733
rect 113584 272699 113618 272733
rect 113652 272699 113686 272733
rect 113720 272699 113754 272733
rect 113788 272699 113822 272733
rect 113856 272699 113890 272733
rect 113924 272699 113958 272733
rect 113992 272699 114026 272733
rect 114060 272699 114094 272733
rect 114128 272699 114162 272733
rect 114196 272699 114230 272733
rect 115860 274110 115962 274212
rect 115975 272699 116009 272733
rect 116043 272699 116077 272733
rect 116111 272699 116145 272733
rect 116179 272699 116213 272733
rect 116247 272699 116281 272733
rect 116315 272699 116349 272733
rect 116383 272699 116417 272733
rect 116451 272699 116485 272733
rect 116519 272699 116553 272733
rect 116587 272699 116621 272733
rect 116655 272699 116689 272733
rect 116723 272699 116757 272733
rect 116791 272699 116825 272733
rect 116859 272699 116893 272733
rect 116927 272699 116961 272733
rect 116995 272699 117029 272733
rect 117063 272699 117097 272733
rect 117131 272699 117165 272733
rect 117199 272699 117233 272733
rect 117267 272699 117301 272733
rect 117335 272699 117369 272733
rect 117403 272699 117437 272733
rect 117471 272699 117505 272733
rect 117539 272699 117573 272733
rect 117607 272699 117641 272733
rect 117675 272699 117709 272733
rect 117743 272699 117777 272733
rect 117811 272699 117845 272733
rect 117879 272699 117913 272733
rect 117947 272699 117981 272733
rect 118015 272699 118049 272733
rect 118083 272699 118117 272733
rect 118151 272699 118185 272733
rect 118219 272699 118253 272733
rect 118287 272699 118321 272733
rect 118355 272699 118389 272733
rect 118423 272699 118457 272733
rect 118491 272699 118525 272733
rect 118559 272699 118593 272733
rect 118627 272699 118661 272733
rect 118695 272699 118729 272733
rect 118763 272699 118797 272733
rect 118831 272699 118865 272733
rect 119031 272704 119133 281102
rect 111953 268677 112055 272247
rect 112178 272136 118944 272238
rect 112171 268713 118937 268815
rect 119035 268677 119137 272247
rect 119970 268785 120072 281059
rect 120256 281037 125118 281139
rect 122034 275562 122136 278588
rect 122531 276103 124265 276205
rect 122891 275002 122925 275036
rect 122959 275002 122993 275036
rect 123027 275002 123061 275036
rect 123095 275002 123129 275036
rect 123163 275002 123197 275036
rect 123231 275002 123265 275036
rect 123299 275002 123333 275036
rect 123367 275002 123401 275036
rect 123435 275002 123469 275036
rect 123503 275002 123537 275036
rect 123571 275002 123605 275036
rect 123639 275002 123673 275036
rect 123707 275002 123741 275036
rect 123775 275002 123809 275036
rect 123843 275002 123877 275036
rect 123911 275002 123945 275036
rect 123979 275002 124013 275036
rect 122792 274881 122826 274915
rect 124078 274881 124112 274915
rect 122792 274813 122826 274847
rect 122792 274745 122826 274779
rect 122792 274677 122826 274711
rect 124078 274813 124112 274847
rect 124078 274745 124112 274779
rect 124078 274677 124112 274711
rect 122792 274609 122826 274643
rect 124078 274609 124112 274643
rect 122110 274507 122144 274541
rect 122178 274507 122212 274541
rect 122246 274507 122280 274541
rect 122314 274507 122348 274541
rect 122382 274507 122416 274541
rect 122450 274507 122484 274541
rect 122518 274507 122552 274541
rect 122586 274507 122620 274541
rect 122654 274507 122688 274541
rect 122891 274488 122925 274522
rect 122959 274488 122993 274522
rect 123027 274488 123061 274522
rect 123095 274488 123129 274522
rect 123163 274488 123197 274522
rect 123231 274488 123265 274522
rect 123299 274488 123333 274522
rect 123367 274488 123401 274522
rect 123435 274488 123469 274522
rect 123503 274488 123537 274522
rect 123571 274488 123605 274522
rect 123639 274488 123673 274522
rect 123707 274488 123741 274522
rect 123775 274488 123809 274522
rect 123843 274488 123877 274522
rect 123911 274488 123945 274522
rect 123979 274488 124013 274522
rect 124232 274518 124266 274552
rect 124300 274518 124334 274552
rect 124368 274518 124402 274552
rect 124436 274518 124470 274552
rect 124504 274518 124538 274552
rect 124572 274518 124606 274552
rect 124640 274518 124674 274552
rect 124708 274518 124742 274552
rect 124776 274518 124810 274552
rect 122089 274247 122123 274281
rect 122089 274179 122123 274213
rect 122089 274111 122123 274145
rect 122089 274043 122123 274077
rect 122089 273975 122123 274009
rect 122089 273907 122123 273941
rect 122089 273839 122123 273873
rect 122089 273771 122123 273805
rect 124753 274263 124787 274297
rect 124753 274195 124787 274229
rect 124753 274127 124787 274161
rect 124753 274059 124787 274093
rect 124753 273991 124787 274025
rect 124753 273923 124787 273957
rect 124753 273855 124787 273889
rect 124753 273787 124787 273821
rect 122089 273703 122123 273737
rect 124753 273719 124787 273753
rect 122089 273635 122123 273669
rect 124753 273651 124787 273685
rect 122243 273564 122277 273598
rect 122311 273564 122345 273598
rect 122379 273564 122413 273598
rect 122447 273564 122481 273598
rect 122515 273564 122549 273598
rect 122583 273564 122617 273598
rect 122651 273564 122685 273598
rect 122719 273564 122753 273598
rect 122787 273564 122821 273598
rect 122855 273564 122889 273598
rect 122923 273564 122957 273598
rect 122991 273564 123025 273598
rect 123059 273564 123093 273598
rect 123127 273564 123161 273598
rect 123195 273564 123229 273598
rect 123263 273564 123297 273598
rect 123331 273564 123365 273598
rect 123399 273564 123433 273598
rect 123467 273564 123501 273598
rect 123535 273564 123569 273598
rect 123603 273564 123637 273598
rect 123671 273564 123705 273598
rect 123739 273564 123773 273598
rect 123807 273564 123841 273598
rect 123875 273564 123909 273598
rect 123943 273564 123977 273598
rect 124011 273564 124045 273598
rect 124079 273564 124113 273598
rect 124147 273564 124181 273598
rect 124215 273564 124249 273598
rect 124283 273564 124317 273598
rect 124351 273564 124385 273598
rect 124419 273564 124453 273598
rect 124487 273564 124521 273598
rect 124555 273564 124589 273598
rect 124065 272716 124099 272750
rect 124133 272716 124167 272750
rect 124201 272716 124235 272750
rect 124269 272716 124303 272750
rect 124337 272716 124371 272750
rect 124405 272716 124439 272750
rect 124473 272716 124507 272750
rect 124541 272716 124575 272750
rect 124609 272716 124643 272750
rect 124677 272716 124711 272750
rect 123986 272558 124020 272592
rect 124828 272653 124862 272687
rect 124828 272585 124862 272619
rect 123986 272490 124020 272524
rect 123986 272422 124020 272456
rect 123986 272354 124020 272388
rect 124828 272517 124862 272551
rect 124828 272449 124862 272483
rect 124828 272381 124862 272415
rect 123986 272286 124020 272320
rect 124828 272313 124862 272347
rect 123986 272218 124020 272252
rect 123986 272150 124020 272184
rect 124828 272245 124862 272279
rect 124828 272177 124862 272211
rect 123986 272082 124020 272116
rect 124828 272109 124862 272143
rect 123986 272014 124020 272048
rect 123986 271946 124020 271980
rect 123986 271878 124020 271912
rect 124828 272041 124862 272075
rect 124828 271973 124862 272007
rect 124828 271905 124862 271939
rect 123986 271810 124020 271844
rect 123986 271742 124020 271776
rect 124828 271837 124862 271871
rect 124828 271769 124862 271803
rect 123986 271674 124020 271708
rect 124828 271701 124862 271735
rect 123986 271606 124020 271640
rect 123986 271538 124020 271572
rect 123986 271470 124020 271504
rect 124828 271633 124862 271667
rect 124828 271565 124862 271599
rect 124828 271497 124862 271531
rect 123986 271402 124020 271436
rect 123986 271334 124020 271368
rect 124828 271429 124862 271463
rect 124828 271361 124862 271395
rect 123986 271266 124020 271300
rect 124828 271293 124862 271327
rect 123986 271198 124020 271232
rect 123986 271130 124020 271164
rect 123986 271062 124020 271096
rect 124828 271225 124862 271259
rect 124828 271157 124862 271191
rect 124828 271089 124862 271123
rect 123986 270994 124020 271028
rect 124828 271021 124862 271055
rect 123986 270926 124020 270960
rect 124828 270953 124862 270987
rect 123986 270858 124020 270892
rect 124828 270885 124862 270919
rect 123986 270790 124020 270824
rect 123986 270722 124020 270756
rect 123986 270654 124020 270688
rect 124828 270817 124862 270851
rect 124828 270749 124862 270783
rect 124828 270681 124862 270715
rect 123986 270586 124020 270620
rect 124828 270613 124862 270647
rect 123986 270518 124020 270552
rect 124828 270545 124862 270579
rect 123986 270450 124020 270484
rect 124828 270477 124862 270511
rect 123986 270382 124020 270416
rect 123986 270314 124020 270348
rect 123986 270246 124020 270280
rect 124828 270409 124862 270443
rect 124828 270341 124862 270375
rect 124828 270273 124862 270307
rect 123986 270178 124020 270212
rect 124828 270205 124862 270239
rect 123986 270110 124020 270144
rect 124828 270137 124862 270171
rect 123986 270042 124020 270076
rect 124828 270069 124862 270103
rect 123986 269974 124020 270008
rect 123986 269906 124020 269940
rect 123986 269838 124020 269872
rect 124828 270001 124862 270035
rect 124828 269933 124862 269967
rect 124828 269865 124862 269899
rect 123986 269770 124020 269804
rect 124828 269797 124862 269831
rect 123986 269702 124020 269736
rect 123986 269634 124020 269668
rect 124828 269729 124862 269763
rect 124828 269661 124862 269695
rect 123986 269566 124020 269600
rect 123986 269498 124020 269532
rect 123986 269430 124020 269464
rect 124828 269593 124862 269627
rect 124828 269525 124862 269559
rect 124828 269457 124862 269491
rect 123986 269362 124020 269396
rect 124828 269389 124862 269423
rect 124828 269321 124862 269355
rect 124049 269220 124083 269254
rect 124117 269220 124151 269254
rect 124185 269220 124219 269254
rect 124253 269220 124287 269254
rect 124321 269220 124355 269254
rect 124389 269220 124423 269254
rect 124457 269220 124491 269254
rect 124525 269220 124559 269254
rect 124593 269220 124627 269254
rect 124661 269220 124695 269254
rect 125058 268990 125160 280856
rect 120283 268733 125145 268835
<< nsubdiffcont >>
rect 106237 279188 106271 279222
rect 106305 279188 106339 279222
rect 106373 279188 106407 279222
rect 106441 279188 106475 279222
rect 106509 279188 106543 279222
rect 106577 279188 106611 279222
rect 106645 279188 106679 279222
rect 106713 279188 106747 279222
rect 106781 279188 106815 279222
rect 106849 279188 106883 279222
rect 106917 279188 106951 279222
rect 106985 279188 107019 279222
rect 107053 279188 107087 279222
rect 107121 279188 107155 279222
rect 107189 279188 107223 279222
rect 107257 279188 107291 279222
rect 107325 279188 107359 279222
rect 107393 279188 107427 279222
rect 107461 279188 107495 279222
rect 107529 279188 107563 279222
rect 107597 279188 107631 279222
rect 107665 279188 107699 279222
rect 106169 279113 106203 279147
rect 106169 279045 106203 279079
rect 107734 279113 107768 279147
rect 107734 279045 107768 279079
rect 106169 278977 106203 279011
rect 106169 278909 106203 278943
rect 106169 278841 106203 278875
rect 106169 278773 106203 278807
rect 107734 278977 107768 279011
rect 107734 278909 107768 278943
rect 107734 278841 107768 278875
rect 107734 278773 107768 278807
rect 106169 278705 106203 278739
rect 107734 278705 107768 278739
rect 106169 278637 106203 278671
rect 106169 278569 106203 278603
rect 106169 278501 106203 278535
rect 107734 278637 107768 278671
rect 107734 278569 107768 278603
rect 107734 278501 107768 278535
rect 106169 278433 106203 278467
rect 107734 278433 107768 278467
rect 106169 278365 106203 278399
rect 106169 278297 106203 278331
rect 106169 278229 106203 278263
rect 106169 278161 106203 278195
rect 107734 278365 107768 278399
rect 107734 278297 107768 278331
rect 107734 278229 107768 278263
rect 107734 278161 107768 278195
rect 106169 278093 106203 278127
rect 106169 278025 106203 278059
rect 107734 278093 107768 278127
rect 107734 278025 107768 278059
rect 106237 277950 106271 277984
rect 106305 277950 106339 277984
rect 106373 277950 106407 277984
rect 106441 277950 106475 277984
rect 106509 277950 106543 277984
rect 106577 277950 106611 277984
rect 106645 277950 106679 277984
rect 106713 277950 106747 277984
rect 106781 277950 106815 277984
rect 106849 277950 106883 277984
rect 106917 277950 106951 277984
rect 106985 277950 107019 277984
rect 107053 277950 107087 277984
rect 107121 277950 107155 277984
rect 107189 277950 107223 277984
rect 107257 277950 107291 277984
rect 107325 277950 107359 277984
rect 107393 277950 107427 277984
rect 107461 277950 107495 277984
rect 107529 277950 107563 277984
rect 107597 277950 107631 277984
rect 107665 277950 107699 277984
rect 106413 277290 106447 277324
rect 106481 277290 106515 277324
rect 106549 277290 106583 277324
rect 106617 277290 106651 277324
rect 106685 277290 106719 277324
rect 106753 277290 106787 277324
rect 106821 277290 106855 277324
rect 106889 277290 106923 277324
rect 106957 277290 106991 277324
rect 107025 277290 107059 277324
rect 107093 277290 107127 277324
rect 107161 277290 107195 277324
rect 107229 277290 107263 277324
rect 107297 277290 107331 277324
rect 107365 277290 107399 277324
rect 107433 277290 107467 277324
rect 107501 277290 107535 277324
rect 107569 277290 107603 277324
rect 106308 277178 106342 277212
rect 107674 277178 107708 277212
rect 106308 277110 106342 277144
rect 107674 277110 107708 277144
rect 106308 277042 106342 277076
rect 107674 277042 107708 277076
rect 106413 276930 106447 276964
rect 106481 276930 106515 276964
rect 106549 276930 106583 276964
rect 106617 276930 106651 276964
rect 106685 276930 106719 276964
rect 106753 276930 106787 276964
rect 106821 276930 106855 276964
rect 106889 276930 106923 276964
rect 106957 276930 106991 276964
rect 107025 276930 107059 276964
rect 107093 276930 107127 276964
rect 107161 276930 107195 276964
rect 107229 276930 107263 276964
rect 107297 276930 107331 276964
rect 107365 276930 107399 276964
rect 107433 276930 107467 276964
rect 107501 276930 107535 276964
rect 107569 276930 107603 276964
rect 106797 275900 106831 275934
rect 106865 275900 106899 275934
rect 106933 275900 106967 275934
rect 107001 275900 107035 275934
rect 107069 275900 107103 275934
rect 107137 275900 107171 275934
rect 107205 275900 107239 275934
rect 107273 275900 107307 275934
rect 107341 275900 107375 275934
rect 107409 275900 107443 275934
rect 107477 275900 107511 275934
rect 107545 275900 107579 275934
rect 107613 275900 107647 275934
rect 107681 275900 107715 275934
rect 107749 275900 107783 275934
rect 107817 275900 107851 275934
rect 107885 275900 107919 275934
rect 107953 275900 107987 275934
rect 108021 275900 108055 275934
rect 108089 275900 108123 275934
rect 108157 275900 108191 275934
rect 108225 275900 108259 275934
rect 108293 275900 108327 275934
rect 108361 275900 108395 275934
rect 108429 275900 108463 275934
rect 108497 275900 108531 275934
rect 108565 275900 108599 275934
rect 108633 275900 108667 275934
rect 108701 275900 108735 275934
rect 108769 275900 108803 275934
rect 108837 275900 108871 275934
rect 108905 275900 108939 275934
rect 108973 275900 109007 275934
rect 109041 275900 109075 275934
rect 109109 275900 109143 275934
rect 109177 275900 109211 275934
rect 109245 275900 109279 275934
rect 109313 275900 109347 275934
rect 109381 275900 109415 275934
rect 109449 275900 109483 275934
rect 109517 275900 109551 275934
rect 109585 275900 109619 275934
rect 109653 275900 109687 275934
rect 109721 275900 109755 275934
rect 106706 275816 106740 275850
rect 106706 275748 106740 275782
rect 109813 275816 109847 275850
rect 106706 275680 106740 275714
rect 109813 275748 109847 275782
rect 106706 275612 106740 275646
rect 106706 275544 106740 275578
rect 106706 275476 106740 275510
rect 106706 275408 106740 275442
rect 106706 275340 106740 275374
rect 106706 275272 106740 275306
rect 106706 275204 106740 275238
rect 106706 275136 106740 275170
rect 106706 275068 106740 275102
rect 106706 275000 106740 275034
rect 106706 274932 106740 274966
rect 109813 275680 109847 275714
rect 109813 275612 109847 275646
rect 109813 275544 109847 275578
rect 109813 275476 109847 275510
rect 109813 275408 109847 275442
rect 109813 275340 109847 275374
rect 109813 275272 109847 275306
rect 109813 275204 109847 275238
rect 109813 275136 109847 275170
rect 109813 275068 109847 275102
rect 109813 275000 109847 275034
rect 106706 274864 106740 274898
rect 109813 274932 109847 274966
rect 106706 274796 106740 274830
rect 109813 274864 109847 274898
rect 109813 274796 109847 274830
rect 106797 274713 106831 274747
rect 106865 274713 106899 274747
rect 106933 274713 106967 274747
rect 107001 274713 107035 274747
rect 107069 274713 107103 274747
rect 107137 274713 107171 274747
rect 107205 274713 107239 274747
rect 107273 274713 107307 274747
rect 107341 274713 107375 274747
rect 107409 274713 107443 274747
rect 107477 274713 107511 274747
rect 107545 274713 107579 274747
rect 107613 274713 107647 274747
rect 107681 274713 107715 274747
rect 107749 274713 107783 274747
rect 107817 274713 107851 274747
rect 107885 274713 107919 274747
rect 107953 274713 107987 274747
rect 108021 274713 108055 274747
rect 108089 274713 108123 274747
rect 108157 274713 108191 274747
rect 108225 274713 108259 274747
rect 108293 274713 108327 274747
rect 108361 274713 108395 274747
rect 108429 274713 108463 274747
rect 108497 274713 108531 274747
rect 108565 274713 108599 274747
rect 108633 274713 108667 274747
rect 108701 274713 108735 274747
rect 108769 274713 108803 274747
rect 108837 274713 108871 274747
rect 108905 274713 108939 274747
rect 108973 274713 109007 274747
rect 109041 274713 109075 274747
rect 109109 274713 109143 274747
rect 109177 274713 109211 274747
rect 109245 274713 109279 274747
rect 109313 274713 109347 274747
rect 109381 274713 109415 274747
rect 109449 274713 109483 274747
rect 109517 274713 109551 274747
rect 109585 274713 109619 274747
rect 109653 274713 109687 274747
rect 109721 274713 109755 274747
rect 109151 272568 109185 272602
rect 109219 272568 109253 272602
rect 109287 272568 109321 272602
rect 109355 272568 109389 272602
rect 109423 272568 109457 272602
rect 109491 272568 109525 272602
rect 109559 272568 109593 272602
rect 109627 272568 109661 272602
rect 109695 272568 109729 272602
rect 109763 272568 109797 272602
rect 109088 272496 109122 272530
rect 109088 272428 109122 272462
rect 109827 272496 109861 272530
rect 109827 272428 109861 272462
rect 109088 272360 109122 272394
rect 109088 272292 109122 272326
rect 109088 272224 109122 272258
rect 109088 272156 109122 272190
rect 109088 272088 109122 272122
rect 109088 272020 109122 272054
rect 109088 271952 109122 271986
rect 109088 271884 109122 271918
rect 109088 271816 109122 271850
rect 109088 271748 109122 271782
rect 109088 271680 109122 271714
rect 109088 271612 109122 271646
rect 109088 271544 109122 271578
rect 109088 271476 109122 271510
rect 109088 271408 109122 271442
rect 109088 271340 109122 271374
rect 109088 271272 109122 271306
rect 109088 271204 109122 271238
rect 109088 271136 109122 271170
rect 109088 271068 109122 271102
rect 109088 271000 109122 271034
rect 109088 270932 109122 270966
rect 109088 270864 109122 270898
rect 109088 270796 109122 270830
rect 109088 270728 109122 270762
rect 109827 272360 109861 272394
rect 109827 272292 109861 272326
rect 109827 272224 109861 272258
rect 109827 272156 109861 272190
rect 109827 272088 109861 272122
rect 109827 272020 109861 272054
rect 109827 271952 109861 271986
rect 109827 271884 109861 271918
rect 109827 271816 109861 271850
rect 109827 271748 109861 271782
rect 109827 271680 109861 271714
rect 109827 271612 109861 271646
rect 109827 271544 109861 271578
rect 109827 271476 109861 271510
rect 109827 271408 109861 271442
rect 109827 271340 109861 271374
rect 109827 271272 109861 271306
rect 109827 271204 109861 271238
rect 109827 271136 109861 271170
rect 109827 271068 109861 271102
rect 109827 271000 109861 271034
rect 109827 270932 109861 270966
rect 109827 270864 109861 270898
rect 109827 270796 109861 270830
rect 109827 270728 109861 270762
rect 109088 270660 109122 270694
rect 109088 270592 109122 270626
rect 109827 270660 109861 270694
rect 109827 270592 109861 270626
rect 109151 270521 109185 270555
rect 109219 270521 109253 270555
rect 109287 270521 109321 270555
rect 109355 270521 109389 270555
rect 109423 270521 109457 270555
rect 109491 270521 109525 270555
rect 109559 270521 109593 270555
rect 109627 270521 109661 270555
rect 109695 270521 109729 270555
rect 109763 270521 109797 270555
rect 114537 280929 114571 280963
rect 114605 280929 114639 280963
rect 114673 280929 114707 280963
rect 114741 280929 114775 280963
rect 114809 280929 114843 280963
rect 114877 280929 114911 280963
rect 114945 280929 114979 280963
rect 114455 280863 114489 280897
rect 115027 280863 115061 280897
rect 114455 280795 114489 280829
rect 114455 280727 114489 280761
rect 114455 280659 114489 280693
rect 114455 280591 114489 280625
rect 114455 280523 114489 280557
rect 114455 280455 114489 280489
rect 114455 280387 114489 280421
rect 115027 280795 115061 280829
rect 115027 280727 115061 280761
rect 115027 280659 115061 280693
rect 115027 280591 115061 280625
rect 115027 280523 115061 280557
rect 115027 280455 115061 280489
rect 114455 280319 114489 280353
rect 115027 280387 115061 280421
rect 114455 280251 114489 280285
rect 114455 280183 114489 280217
rect 115027 280319 115061 280353
rect 115027 280251 115061 280285
rect 115027 280183 115061 280217
rect 114455 280115 114489 280149
rect 114455 280047 114489 280081
rect 114455 279979 114489 280013
rect 115027 280115 115061 280149
rect 115027 280047 115061 280081
rect 115027 279979 115061 280013
rect 114455 279911 114489 279945
rect 115027 279911 115061 279945
rect 114455 279843 114489 279877
rect 114455 279775 114489 279809
rect 115027 279843 115061 279877
rect 115027 279775 115061 279809
rect 114455 279707 114489 279741
rect 114455 279639 114489 279673
rect 114455 279571 114489 279605
rect 115027 279707 115061 279741
rect 115027 279639 115061 279673
rect 115027 279571 115061 279605
rect 114455 279503 114489 279537
rect 115027 279503 115061 279537
rect 114455 279435 114489 279469
rect 115027 279435 115061 279469
rect 114537 279369 114571 279403
rect 114605 279369 114639 279403
rect 114673 279369 114707 279403
rect 114741 279369 114775 279403
rect 114809 279369 114843 279403
rect 114877 279369 114911 279403
rect 114945 279369 114979 279403
rect 115226 280929 115260 280963
rect 115294 280929 115328 280963
rect 115362 280929 115396 280963
rect 115430 280929 115464 280963
rect 115498 280929 115532 280963
rect 115566 280929 115600 280963
rect 115634 280929 115668 280963
rect 115144 280863 115178 280897
rect 115716 280863 115750 280897
rect 115144 280795 115178 280829
rect 115144 280727 115178 280761
rect 115144 280659 115178 280693
rect 115144 280591 115178 280625
rect 115144 280523 115178 280557
rect 115144 280455 115178 280489
rect 115144 280387 115178 280421
rect 115716 280795 115750 280829
rect 115716 280727 115750 280761
rect 115716 280659 115750 280693
rect 115716 280591 115750 280625
rect 115716 280523 115750 280557
rect 115716 280455 115750 280489
rect 115144 280319 115178 280353
rect 115716 280387 115750 280421
rect 115144 280251 115178 280285
rect 115144 280183 115178 280217
rect 115716 280319 115750 280353
rect 115716 280251 115750 280285
rect 115716 280183 115750 280217
rect 115144 280115 115178 280149
rect 115144 280047 115178 280081
rect 115144 279979 115178 280013
rect 115716 280115 115750 280149
rect 115716 280047 115750 280081
rect 115716 279979 115750 280013
rect 115144 279911 115178 279945
rect 115716 279911 115750 279945
rect 115144 279843 115178 279877
rect 115144 279775 115178 279809
rect 115716 279843 115750 279877
rect 115716 279775 115750 279809
rect 115144 279707 115178 279741
rect 115144 279639 115178 279673
rect 115144 279571 115178 279605
rect 115716 279707 115750 279741
rect 115716 279639 115750 279673
rect 115716 279571 115750 279605
rect 115144 279503 115178 279537
rect 115716 279503 115750 279537
rect 115144 279435 115178 279469
rect 115716 279435 115750 279469
rect 115226 279369 115260 279403
rect 115294 279369 115328 279403
rect 115362 279369 115396 279403
rect 115430 279369 115464 279403
rect 115498 279369 115532 279403
rect 115566 279369 115600 279403
rect 115634 279369 115668 279403
rect 114537 279263 114571 279297
rect 114605 279263 114639 279297
rect 114673 279263 114707 279297
rect 114741 279263 114775 279297
rect 114809 279263 114843 279297
rect 114877 279263 114911 279297
rect 114945 279263 114979 279297
rect 114455 279197 114489 279231
rect 115027 279197 115061 279231
rect 114455 279129 114489 279163
rect 114455 279061 114489 279095
rect 114455 278993 114489 279027
rect 114455 278925 114489 278959
rect 114455 278857 114489 278891
rect 114455 278789 114489 278823
rect 114455 278721 114489 278755
rect 115027 279129 115061 279163
rect 115027 279061 115061 279095
rect 115027 278993 115061 279027
rect 115027 278925 115061 278959
rect 115027 278857 115061 278891
rect 115027 278789 115061 278823
rect 114455 278653 114489 278687
rect 115027 278721 115061 278755
rect 114455 278585 114489 278619
rect 114455 278517 114489 278551
rect 115027 278653 115061 278687
rect 115027 278585 115061 278619
rect 115027 278517 115061 278551
rect 114455 278449 114489 278483
rect 114455 278381 114489 278415
rect 114455 278313 114489 278347
rect 115027 278449 115061 278483
rect 115027 278381 115061 278415
rect 115027 278313 115061 278347
rect 114455 278245 114489 278279
rect 115027 278245 115061 278279
rect 114455 278177 114489 278211
rect 114455 278109 114489 278143
rect 115027 278177 115061 278211
rect 115027 278109 115061 278143
rect 114455 278041 114489 278075
rect 114455 277973 114489 278007
rect 114455 277905 114489 277939
rect 115027 278041 115061 278075
rect 115027 277973 115061 278007
rect 115027 277905 115061 277939
rect 114455 277837 114489 277871
rect 115027 277837 115061 277871
rect 114455 277769 114489 277803
rect 115027 277769 115061 277803
rect 114537 277703 114571 277737
rect 114605 277703 114639 277737
rect 114673 277703 114707 277737
rect 114741 277703 114775 277737
rect 114809 277703 114843 277737
rect 114877 277703 114911 277737
rect 114945 277703 114979 277737
rect 115226 279263 115260 279297
rect 115294 279263 115328 279297
rect 115362 279263 115396 279297
rect 115430 279263 115464 279297
rect 115498 279263 115532 279297
rect 115566 279263 115600 279297
rect 115634 279263 115668 279297
rect 115144 279197 115178 279231
rect 115716 279197 115750 279231
rect 115144 279129 115178 279163
rect 115144 279061 115178 279095
rect 115144 278993 115178 279027
rect 115144 278925 115178 278959
rect 115144 278857 115178 278891
rect 115144 278789 115178 278823
rect 115144 278721 115178 278755
rect 115716 279129 115750 279163
rect 115716 279061 115750 279095
rect 115716 278993 115750 279027
rect 115716 278925 115750 278959
rect 115716 278857 115750 278891
rect 115716 278789 115750 278823
rect 115144 278653 115178 278687
rect 115716 278721 115750 278755
rect 115144 278585 115178 278619
rect 115144 278517 115178 278551
rect 115716 278653 115750 278687
rect 115716 278585 115750 278619
rect 115716 278517 115750 278551
rect 115144 278449 115178 278483
rect 115144 278381 115178 278415
rect 115144 278313 115178 278347
rect 115716 278449 115750 278483
rect 115716 278381 115750 278415
rect 115716 278313 115750 278347
rect 115144 278245 115178 278279
rect 115716 278245 115750 278279
rect 115144 278177 115178 278211
rect 115144 278109 115178 278143
rect 115716 278177 115750 278211
rect 115716 278109 115750 278143
rect 115144 278041 115178 278075
rect 115144 277973 115178 278007
rect 115144 277905 115178 277939
rect 115716 278041 115750 278075
rect 115716 277973 115750 278007
rect 115716 277905 115750 277939
rect 115144 277837 115178 277871
rect 115716 277837 115750 277871
rect 115144 277769 115178 277803
rect 115716 277769 115750 277803
rect 115226 277703 115260 277737
rect 115294 277703 115328 277737
rect 115362 277703 115396 277737
rect 115430 277703 115464 277737
rect 115498 277703 115532 277737
rect 115566 277703 115600 277737
rect 115634 277703 115668 277737
rect 114537 277597 114571 277631
rect 114605 277597 114639 277631
rect 114673 277597 114707 277631
rect 114741 277597 114775 277631
rect 114809 277597 114843 277631
rect 114877 277597 114911 277631
rect 114945 277597 114979 277631
rect 114455 277531 114489 277565
rect 115027 277531 115061 277565
rect 114455 277463 114489 277497
rect 114455 277395 114489 277429
rect 114455 277327 114489 277361
rect 114455 277259 114489 277293
rect 114455 277191 114489 277225
rect 114455 277123 114489 277157
rect 114455 277055 114489 277089
rect 115027 277463 115061 277497
rect 115027 277395 115061 277429
rect 115027 277327 115061 277361
rect 115027 277259 115061 277293
rect 115027 277191 115061 277225
rect 115027 277123 115061 277157
rect 114455 276987 114489 277021
rect 115027 277055 115061 277089
rect 114455 276919 114489 276953
rect 114455 276851 114489 276885
rect 115027 276987 115061 277021
rect 115027 276919 115061 276953
rect 115027 276851 115061 276885
rect 114455 276783 114489 276817
rect 114455 276715 114489 276749
rect 114455 276647 114489 276681
rect 115027 276783 115061 276817
rect 115027 276715 115061 276749
rect 115027 276647 115061 276681
rect 114455 276579 114489 276613
rect 115027 276579 115061 276613
rect 114455 276511 114489 276545
rect 114455 276443 114489 276477
rect 115027 276511 115061 276545
rect 115027 276443 115061 276477
rect 114455 276375 114489 276409
rect 114455 276307 114489 276341
rect 114455 276239 114489 276273
rect 115027 276375 115061 276409
rect 115027 276307 115061 276341
rect 115027 276239 115061 276273
rect 114455 276171 114489 276205
rect 115027 276171 115061 276205
rect 114455 276103 114489 276137
rect 115027 276103 115061 276137
rect 114537 276037 114571 276071
rect 114605 276037 114639 276071
rect 114673 276037 114707 276071
rect 114741 276037 114775 276071
rect 114809 276037 114843 276071
rect 114877 276037 114911 276071
rect 114945 276037 114979 276071
rect 115226 277597 115260 277631
rect 115294 277597 115328 277631
rect 115362 277597 115396 277631
rect 115430 277597 115464 277631
rect 115498 277597 115532 277631
rect 115566 277597 115600 277631
rect 115634 277597 115668 277631
rect 115144 277531 115178 277565
rect 115716 277531 115750 277565
rect 115144 277463 115178 277497
rect 115144 277395 115178 277429
rect 115144 277327 115178 277361
rect 115144 277259 115178 277293
rect 115144 277191 115178 277225
rect 115144 277123 115178 277157
rect 115144 277055 115178 277089
rect 115716 277463 115750 277497
rect 115716 277395 115750 277429
rect 115716 277327 115750 277361
rect 115716 277259 115750 277293
rect 115716 277191 115750 277225
rect 115716 277123 115750 277157
rect 115144 276987 115178 277021
rect 115716 277055 115750 277089
rect 115144 276919 115178 276953
rect 115144 276851 115178 276885
rect 115716 276987 115750 277021
rect 115716 276919 115750 276953
rect 115716 276851 115750 276885
rect 115144 276783 115178 276817
rect 115144 276715 115178 276749
rect 115144 276647 115178 276681
rect 115716 276783 115750 276817
rect 115716 276715 115750 276749
rect 115716 276647 115750 276681
rect 115144 276579 115178 276613
rect 115716 276579 115750 276613
rect 115144 276511 115178 276545
rect 115144 276443 115178 276477
rect 115716 276511 115750 276545
rect 115716 276443 115750 276477
rect 115144 276375 115178 276409
rect 115144 276307 115178 276341
rect 115144 276239 115178 276273
rect 115716 276375 115750 276409
rect 115716 276307 115750 276341
rect 115716 276239 115750 276273
rect 115144 276171 115178 276205
rect 115716 276171 115750 276205
rect 115144 276103 115178 276137
rect 115716 276103 115750 276137
rect 115226 276037 115260 276071
rect 115294 276037 115328 276071
rect 115362 276037 115396 276071
rect 115430 276037 115464 276071
rect 115498 276037 115532 276071
rect 115566 276037 115600 276071
rect 115634 276037 115668 276071
rect 114537 275931 114571 275965
rect 114605 275931 114639 275965
rect 114673 275931 114707 275965
rect 114741 275931 114775 275965
rect 114809 275931 114843 275965
rect 114877 275931 114911 275965
rect 114945 275931 114979 275965
rect 114455 275865 114489 275899
rect 115027 275865 115061 275899
rect 114455 275797 114489 275831
rect 114455 275729 114489 275763
rect 114455 275661 114489 275695
rect 114455 275593 114489 275627
rect 114455 275525 114489 275559
rect 114455 275457 114489 275491
rect 114455 275389 114489 275423
rect 115027 275797 115061 275831
rect 115027 275729 115061 275763
rect 115027 275661 115061 275695
rect 115027 275593 115061 275627
rect 115027 275525 115061 275559
rect 115027 275457 115061 275491
rect 114455 275321 114489 275355
rect 115027 275389 115061 275423
rect 114455 275253 114489 275287
rect 114455 275185 114489 275219
rect 115027 275321 115061 275355
rect 115027 275253 115061 275287
rect 115027 275185 115061 275219
rect 114455 275117 114489 275151
rect 114455 275049 114489 275083
rect 114455 274981 114489 275015
rect 115027 275117 115061 275151
rect 115027 275049 115061 275083
rect 115027 274981 115061 275015
rect 114455 274913 114489 274947
rect 115027 274913 115061 274947
rect 114455 274845 114489 274879
rect 114455 274777 114489 274811
rect 115027 274845 115061 274879
rect 115027 274777 115061 274811
rect 114455 274709 114489 274743
rect 114455 274641 114489 274675
rect 114455 274573 114489 274607
rect 115027 274709 115061 274743
rect 115027 274641 115061 274675
rect 115027 274573 115061 274607
rect 114455 274505 114489 274539
rect 115027 274505 115061 274539
rect 114455 274437 114489 274471
rect 115027 274437 115061 274471
rect 114537 274371 114571 274405
rect 114605 274371 114639 274405
rect 114673 274371 114707 274405
rect 114741 274371 114775 274405
rect 114809 274371 114843 274405
rect 114877 274371 114911 274405
rect 114945 274371 114979 274405
rect 115226 275931 115260 275965
rect 115294 275931 115328 275965
rect 115362 275931 115396 275965
rect 115430 275931 115464 275965
rect 115498 275931 115532 275965
rect 115566 275931 115600 275965
rect 115634 275931 115668 275965
rect 115144 275865 115178 275899
rect 115716 275865 115750 275899
rect 115144 275797 115178 275831
rect 115144 275729 115178 275763
rect 115144 275661 115178 275695
rect 115144 275593 115178 275627
rect 115144 275525 115178 275559
rect 115144 275457 115178 275491
rect 115144 275389 115178 275423
rect 115716 275797 115750 275831
rect 115716 275729 115750 275763
rect 115716 275661 115750 275695
rect 115716 275593 115750 275627
rect 115716 275525 115750 275559
rect 115716 275457 115750 275491
rect 115144 275321 115178 275355
rect 115716 275389 115750 275423
rect 115144 275253 115178 275287
rect 115144 275185 115178 275219
rect 115716 275321 115750 275355
rect 115716 275253 115750 275287
rect 115716 275185 115750 275219
rect 115144 275117 115178 275151
rect 115144 275049 115178 275083
rect 115144 274981 115178 275015
rect 115716 275117 115750 275151
rect 115716 275049 115750 275083
rect 115716 274981 115750 275015
rect 115144 274913 115178 274947
rect 115716 274913 115750 274947
rect 115144 274845 115178 274879
rect 115144 274777 115178 274811
rect 115716 274845 115750 274879
rect 115716 274777 115750 274811
rect 115144 274709 115178 274743
rect 115144 274641 115178 274675
rect 115144 274573 115178 274607
rect 115716 274709 115750 274743
rect 115716 274641 115750 274675
rect 115716 274573 115750 274607
rect 115144 274505 115178 274539
rect 115716 274505 115750 274539
rect 115144 274437 115178 274471
rect 115716 274437 115750 274471
rect 115226 274371 115260 274405
rect 115294 274371 115328 274405
rect 115362 274371 115396 274405
rect 115430 274371 115464 274405
rect 115498 274371 115532 274405
rect 115566 274371 115600 274405
rect 115634 274371 115668 274405
rect 114537 274265 114571 274299
rect 114605 274265 114639 274299
rect 114673 274265 114707 274299
rect 114741 274265 114775 274299
rect 114809 274265 114843 274299
rect 114877 274265 114911 274299
rect 114945 274265 114979 274299
rect 114455 274199 114489 274233
rect 115027 274199 115061 274233
rect 114455 274131 114489 274165
rect 114455 274063 114489 274097
rect 114455 273995 114489 274029
rect 114455 273927 114489 273961
rect 114455 273859 114489 273893
rect 114455 273791 114489 273825
rect 114455 273723 114489 273757
rect 115027 274131 115061 274165
rect 115027 274063 115061 274097
rect 115027 273995 115061 274029
rect 115027 273927 115061 273961
rect 115027 273859 115061 273893
rect 115027 273791 115061 273825
rect 114455 273655 114489 273689
rect 115027 273723 115061 273757
rect 114455 273587 114489 273621
rect 114455 273519 114489 273553
rect 115027 273655 115061 273689
rect 115027 273587 115061 273621
rect 115027 273519 115061 273553
rect 114455 273451 114489 273485
rect 114455 273383 114489 273417
rect 114455 273315 114489 273349
rect 115027 273451 115061 273485
rect 115027 273383 115061 273417
rect 115027 273315 115061 273349
rect 114455 273247 114489 273281
rect 115027 273247 115061 273281
rect 114455 273179 114489 273213
rect 114455 273111 114489 273145
rect 115027 273179 115061 273213
rect 115027 273111 115061 273145
rect 114455 273043 114489 273077
rect 114455 272975 114489 273009
rect 114455 272907 114489 272941
rect 115027 273043 115061 273077
rect 115027 272975 115061 273009
rect 115027 272907 115061 272941
rect 114455 272839 114489 272873
rect 115027 272839 115061 272873
rect 114455 272771 114489 272805
rect 115027 272771 115061 272805
rect 114537 272705 114571 272739
rect 114605 272705 114639 272739
rect 114673 272705 114707 272739
rect 114741 272705 114775 272739
rect 114809 272705 114843 272739
rect 114877 272705 114911 272739
rect 114945 272705 114979 272739
rect 115226 274265 115260 274299
rect 115294 274265 115328 274299
rect 115362 274265 115396 274299
rect 115430 274265 115464 274299
rect 115498 274265 115532 274299
rect 115566 274265 115600 274299
rect 115634 274265 115668 274299
rect 115144 274199 115178 274233
rect 115716 274199 115750 274233
rect 115144 274131 115178 274165
rect 115144 274063 115178 274097
rect 115144 273995 115178 274029
rect 115144 273927 115178 273961
rect 115144 273859 115178 273893
rect 115144 273791 115178 273825
rect 115144 273723 115178 273757
rect 115716 274131 115750 274165
rect 115716 274063 115750 274097
rect 115716 273995 115750 274029
rect 115716 273927 115750 273961
rect 115716 273859 115750 273893
rect 115716 273791 115750 273825
rect 115144 273655 115178 273689
rect 115716 273723 115750 273757
rect 115144 273587 115178 273621
rect 115144 273519 115178 273553
rect 115716 273655 115750 273689
rect 115716 273587 115750 273621
rect 115716 273519 115750 273553
rect 115144 273451 115178 273485
rect 115144 273383 115178 273417
rect 115144 273315 115178 273349
rect 115716 273451 115750 273485
rect 115716 273383 115750 273417
rect 115716 273315 115750 273349
rect 115144 273247 115178 273281
rect 115716 273247 115750 273281
rect 115144 273179 115178 273213
rect 115144 273111 115178 273145
rect 115716 273179 115750 273213
rect 115716 273111 115750 273145
rect 115144 273043 115178 273077
rect 115144 272975 115178 273009
rect 115144 272907 115178 272941
rect 115716 273043 115750 273077
rect 115716 272975 115750 273009
rect 115716 272907 115750 272941
rect 115144 272839 115178 272873
rect 115716 272839 115750 272873
rect 115144 272771 115178 272805
rect 115716 272771 115750 272805
rect 115226 272705 115260 272739
rect 115294 272705 115328 272739
rect 115362 272705 115396 272739
rect 115430 272705 115464 272739
rect 115498 272705 115532 272739
rect 115566 272705 115600 272739
rect 115634 272705 115668 272739
rect 112391 271634 112425 271668
rect 112459 271634 112493 271668
rect 112527 271634 112561 271668
rect 112595 271634 112629 271668
rect 112663 271634 112697 271668
rect 112731 271634 112765 271668
rect 112799 271634 112833 271668
rect 112867 271634 112901 271668
rect 112935 271634 112969 271668
rect 113003 271634 113037 271668
rect 113071 271634 113105 271668
rect 113139 271634 113173 271668
rect 113207 271634 113241 271668
rect 113275 271634 113309 271668
rect 113343 271634 113377 271668
rect 113411 271634 113445 271668
rect 113479 271634 113513 271668
rect 113547 271634 113581 271668
rect 113615 271634 113649 271668
rect 113683 271634 113717 271668
rect 113751 271634 113785 271668
rect 113819 271634 113853 271668
rect 113887 271634 113921 271668
rect 113955 271634 113989 271668
rect 114023 271634 114057 271668
rect 114091 271634 114125 271668
rect 112307 271548 112341 271582
rect 112307 271480 112341 271514
rect 112307 271412 112341 271446
rect 114176 271548 114210 271582
rect 114176 271480 114210 271514
rect 114176 271412 114210 271446
rect 112307 271344 112341 271378
rect 112307 271276 112341 271310
rect 114176 271344 114210 271378
rect 112307 271208 112341 271242
rect 112307 271140 112341 271174
rect 114176 271276 114210 271310
rect 114176 271208 114210 271242
rect 114176 271140 114210 271174
rect 112307 271072 112341 271106
rect 112307 271004 112341 271038
rect 114176 271072 114210 271106
rect 112307 270936 112341 270970
rect 112307 270868 112341 270902
rect 114176 271004 114210 271038
rect 114176 270936 114210 270970
rect 114176 270868 114210 270902
rect 112391 270783 112425 270817
rect 112459 270783 112493 270817
rect 112527 270783 112561 270817
rect 112595 270783 112629 270817
rect 112663 270783 112697 270817
rect 112731 270783 112765 270817
rect 112799 270783 112833 270817
rect 112867 270783 112901 270817
rect 112935 270783 112969 270817
rect 113003 270783 113037 270817
rect 113071 270783 113105 270817
rect 113139 270783 113173 270817
rect 113207 270783 113241 270817
rect 113275 270783 113309 270817
rect 113343 270783 113377 270817
rect 113411 270783 113445 270817
rect 113479 270783 113513 270817
rect 113547 270783 113581 270817
rect 113615 270783 113649 270817
rect 113683 270783 113717 270817
rect 113751 270783 113785 270817
rect 113819 270783 113853 270817
rect 113887 270783 113921 270817
rect 113955 270783 113989 270817
rect 114023 270783 114057 270817
rect 114091 270783 114125 270817
rect 114389 271554 114423 271588
rect 114457 271554 114491 271588
rect 114525 271554 114559 271588
rect 114593 271554 114627 271588
rect 114661 271554 114695 271588
rect 114729 271554 114763 271588
rect 114797 271554 114831 271588
rect 114865 271554 114899 271588
rect 114933 271554 114967 271588
rect 115001 271554 115035 271588
rect 115069 271554 115103 271588
rect 115137 271554 115171 271588
rect 115205 271554 115239 271588
rect 115273 271554 115307 271588
rect 115341 271554 115375 271588
rect 115409 271554 115443 271588
rect 114329 271469 114363 271503
rect 114329 271401 114363 271435
rect 115469 271469 115503 271503
rect 115469 271401 115503 271435
rect 114329 271333 114363 271367
rect 114329 271265 114363 271299
rect 115469 271333 115503 271367
rect 114329 271197 114363 271231
rect 114329 271129 114363 271163
rect 114329 271061 114363 271095
rect 115469 271265 115503 271299
rect 115469 271197 115503 271231
rect 115469 271129 115503 271163
rect 114329 270993 114363 271027
rect 115469 271061 115503 271095
rect 115469 270993 115503 271027
rect 114329 270925 114363 270959
rect 114329 270857 114363 270891
rect 115469 270925 115503 270959
rect 115469 270857 115503 270891
rect 114389 270772 114423 270806
rect 114457 270772 114491 270806
rect 114525 270772 114559 270806
rect 114593 270772 114627 270806
rect 114661 270772 114695 270806
rect 114729 270772 114763 270806
rect 114797 270772 114831 270806
rect 114865 270772 114899 270806
rect 114933 270772 114967 270806
rect 115001 270772 115035 270806
rect 115069 270772 115103 270806
rect 115137 270772 115171 270806
rect 115205 270772 115239 270806
rect 115273 270772 115307 270806
rect 115341 270772 115375 270806
rect 115409 270772 115443 270806
rect 120319 280779 120353 280813
rect 120387 280779 120421 280813
rect 120455 280779 120489 280813
rect 120523 280779 120557 280813
rect 120591 280779 120625 280813
rect 120659 280779 120693 280813
rect 120727 280779 120761 280813
rect 120795 280779 120829 280813
rect 120863 280779 120897 280813
rect 120931 280779 120965 280813
rect 120999 280779 121033 280813
rect 121067 280779 121101 280813
rect 121135 280779 121169 280813
rect 121203 280779 121237 280813
rect 121271 280779 121305 280813
rect 121339 280779 121373 280813
rect 121407 280779 121441 280813
rect 121475 280779 121509 280813
rect 121543 280779 121577 280813
rect 121611 280779 121645 280813
rect 120237 280692 120271 280726
rect 120237 280624 120271 280658
rect 121694 280692 121728 280726
rect 120237 280556 120271 280590
rect 121694 280624 121728 280658
rect 121694 280556 121728 280590
rect 120237 280488 120271 280522
rect 120237 280420 120271 280454
rect 121694 280488 121728 280522
rect 120237 280352 120271 280386
rect 121694 280420 121728 280454
rect 121694 280352 121728 280386
rect 120237 280284 120271 280318
rect 121694 280284 121728 280318
rect 120237 280216 120271 280250
rect 120237 280148 120271 280182
rect 120237 280080 120271 280114
rect 120237 280012 120271 280046
rect 120237 279944 120271 279978
rect 120237 279876 120271 279910
rect 120237 279808 120271 279842
rect 120237 279740 120271 279774
rect 121694 280216 121728 280250
rect 121694 280148 121728 280182
rect 121694 280080 121728 280114
rect 121694 280012 121728 280046
rect 121694 279944 121728 279978
rect 121694 279876 121728 279910
rect 121694 279808 121728 279842
rect 120237 279672 120271 279706
rect 121694 279740 121728 279774
rect 121694 279672 121728 279706
rect 120237 279604 120271 279638
rect 120237 279536 120271 279570
rect 121694 279604 121728 279638
rect 120237 279468 120271 279502
rect 121694 279536 121728 279570
rect 120237 279400 120271 279434
rect 120237 279332 120271 279366
rect 120237 279264 120271 279298
rect 120237 279196 120271 279230
rect 120237 279128 120271 279162
rect 120237 279060 120271 279094
rect 120237 278992 120271 279026
rect 121694 279468 121728 279502
rect 121694 279400 121728 279434
rect 121694 279332 121728 279366
rect 121694 279264 121728 279298
rect 121694 279196 121728 279230
rect 121694 279128 121728 279162
rect 121694 279060 121728 279094
rect 121694 278992 121728 279026
rect 120237 278924 120271 278958
rect 120237 278856 120271 278890
rect 122245 280574 122279 280608
rect 122313 280574 122347 280608
rect 122381 280574 122415 280608
rect 122449 280574 122483 280608
rect 122517 280574 122551 280608
rect 122585 280574 122619 280608
rect 122653 280574 122687 280608
rect 122721 280574 122755 280608
rect 122789 280574 122823 280608
rect 122857 280574 122891 280608
rect 122925 280574 122959 280608
rect 122993 280574 123027 280608
rect 123061 280574 123095 280608
rect 123129 280574 123163 280608
rect 123197 280574 123231 280608
rect 123265 280574 123299 280608
rect 123333 280574 123367 280608
rect 123401 280574 123435 280608
rect 123469 280574 123503 280608
rect 123537 280574 123571 280608
rect 122178 280484 122212 280518
rect 122178 280416 122212 280450
rect 123604 280484 123638 280518
rect 122178 280348 122212 280382
rect 122178 280280 122212 280314
rect 122178 280212 122212 280246
rect 122178 280144 122212 280178
rect 122178 280076 122212 280110
rect 122178 280008 122212 280042
rect 122178 279940 122212 279974
rect 123604 280416 123638 280450
rect 123604 280348 123638 280382
rect 123604 280280 123638 280314
rect 123604 280212 123638 280246
rect 123604 280144 123638 280178
rect 123604 280076 123638 280110
rect 123604 280008 123638 280042
rect 123604 279940 123638 279974
rect 122178 279872 122212 279906
rect 122178 279804 122212 279838
rect 123604 279872 123638 279906
rect 122178 279736 122212 279770
rect 123604 279804 123638 279838
rect 123604 279736 123638 279770
rect 122178 279668 122212 279702
rect 123604 279668 123638 279702
rect 122178 279600 122212 279634
rect 122178 279532 122212 279566
rect 122178 279464 122212 279498
rect 122178 279396 122212 279430
rect 122178 279328 122212 279362
rect 122178 279260 122212 279294
rect 122178 279192 122212 279226
rect 122178 279124 122212 279158
rect 123604 279600 123638 279634
rect 123604 279532 123638 279566
rect 123604 279464 123638 279498
rect 123604 279396 123638 279430
rect 123604 279328 123638 279362
rect 123604 279260 123638 279294
rect 123604 279192 123638 279226
rect 122178 279056 122212 279090
rect 123604 279124 123638 279158
rect 123604 279056 123638 279090
rect 122245 278966 122279 279000
rect 122313 278966 122347 279000
rect 122381 278966 122415 279000
rect 122449 278966 122483 279000
rect 122517 278966 122551 279000
rect 122585 278966 122619 279000
rect 122653 278966 122687 279000
rect 122721 278966 122755 279000
rect 122789 278966 122823 279000
rect 122857 278966 122891 279000
rect 122925 278966 122959 279000
rect 122993 278966 123027 279000
rect 123061 278966 123095 279000
rect 123129 278966 123163 279000
rect 123197 278966 123231 279000
rect 123265 278966 123299 279000
rect 123333 278966 123367 279000
rect 123401 278966 123435 279000
rect 123469 278966 123503 279000
rect 123537 278966 123571 279000
rect 121694 278924 121728 278958
rect 120237 278788 120271 278822
rect 121694 278856 121728 278890
rect 121694 278788 121728 278822
rect 120237 278720 120271 278754
rect 120237 278652 120271 278686
rect 121694 278720 121728 278754
rect 120237 278584 120271 278618
rect 120237 278516 120271 278550
rect 120237 278448 120271 278482
rect 120237 278380 120271 278414
rect 120237 278312 120271 278346
rect 120237 278244 120271 278278
rect 120237 278176 120271 278210
rect 121694 278652 121728 278686
rect 121694 278584 121728 278618
rect 121694 278516 121728 278550
rect 121694 278448 121728 278482
rect 121694 278380 121728 278414
rect 121694 278312 121728 278346
rect 121694 278244 121728 278278
rect 120237 278108 120271 278142
rect 121694 278176 121728 278210
rect 121694 278108 121728 278142
rect 120237 278040 120271 278074
rect 120237 277972 120271 278006
rect 121694 278040 121728 278074
rect 120237 277904 120271 277938
rect 121694 277972 121728 278006
rect 121694 277904 121728 277938
rect 120237 277836 120271 277870
rect 120237 277768 120271 277802
rect 120237 277700 120271 277734
rect 120237 277632 120271 277666
rect 120237 277564 120271 277598
rect 120237 277496 120271 277530
rect 120237 277428 120271 277462
rect 121694 277836 121728 277870
rect 121694 277768 121728 277802
rect 121694 277700 121728 277734
rect 121694 277632 121728 277666
rect 121694 277564 121728 277598
rect 121694 277496 121728 277530
rect 121694 277428 121728 277462
rect 120237 277360 120271 277394
rect 120237 277292 120271 277326
rect 121694 277360 121728 277394
rect 120237 277224 120271 277258
rect 121694 277292 121728 277326
rect 121694 277224 121728 277258
rect 120237 277156 120271 277190
rect 120237 277088 120271 277122
rect 121694 277156 121728 277190
rect 120237 277020 120271 277054
rect 120237 276952 120271 276986
rect 120237 276884 120271 276918
rect 120237 276816 120271 276850
rect 120237 276748 120271 276782
rect 120237 276680 120271 276714
rect 120237 276612 120271 276646
rect 121694 277088 121728 277122
rect 121694 277020 121728 277054
rect 121694 276952 121728 276986
rect 121694 276884 121728 276918
rect 121694 276816 121728 276850
rect 121694 276748 121728 276782
rect 121694 276680 121728 276714
rect 120237 276544 120271 276578
rect 121694 276612 121728 276646
rect 121694 276544 121728 276578
rect 120237 276476 120271 276510
rect 120237 276408 120271 276442
rect 121694 276476 121728 276510
rect 120237 276340 120271 276374
rect 121694 276408 121728 276442
rect 121694 276340 121728 276374
rect 120237 276272 120271 276306
rect 120237 276204 120271 276238
rect 120237 276136 120271 276170
rect 120237 276068 120271 276102
rect 120237 276000 120271 276034
rect 120237 275932 120271 275966
rect 120237 275864 120271 275898
rect 121694 276272 121728 276306
rect 121694 276204 121728 276238
rect 121694 276136 121728 276170
rect 121694 276068 121728 276102
rect 121694 276000 121728 276034
rect 121694 275932 121728 275966
rect 121694 275864 121728 275898
rect 120237 275796 120271 275830
rect 120237 275728 120271 275762
rect 121694 275796 121728 275830
rect 120237 275660 120271 275694
rect 121694 275728 121728 275762
rect 121694 275660 121728 275694
rect 120237 275592 120271 275626
rect 120237 275524 120271 275558
rect 121694 275592 121728 275626
rect 120237 275456 120271 275490
rect 120237 275388 120271 275422
rect 120237 275320 120271 275354
rect 120237 275252 120271 275286
rect 120237 275184 120271 275218
rect 120237 275116 120271 275150
rect 120237 275048 120271 275082
rect 121694 275524 121728 275558
rect 122343 278448 122377 278482
rect 122411 278448 122445 278482
rect 122479 278448 122513 278482
rect 122547 278448 122581 278482
rect 122615 278448 122649 278482
rect 122683 278448 122717 278482
rect 122751 278448 122785 278482
rect 122819 278448 122853 278482
rect 122887 278448 122921 278482
rect 122955 278448 122989 278482
rect 123023 278448 123057 278482
rect 123091 278448 123125 278482
rect 123159 278448 123193 278482
rect 123227 278448 123261 278482
rect 123295 278448 123329 278482
rect 123363 278448 123397 278482
rect 123431 278448 123465 278482
rect 123499 278448 123533 278482
rect 123567 278448 123601 278482
rect 123635 278448 123669 278482
rect 123703 278448 123737 278482
rect 123771 278448 123805 278482
rect 123839 278448 123873 278482
rect 123907 278448 123941 278482
rect 123975 278448 124009 278482
rect 124043 278448 124077 278482
rect 124111 278448 124145 278482
rect 124179 278448 124213 278482
rect 124247 278448 124281 278482
rect 122254 278361 122288 278395
rect 122254 278293 122288 278327
rect 124336 278361 124370 278395
rect 124336 278293 124370 278327
rect 122254 278225 122288 278259
rect 122254 278157 122288 278191
rect 122254 278089 122288 278123
rect 122254 278021 122288 278055
rect 122254 277953 122288 277987
rect 122254 277885 122288 277919
rect 122254 277817 122288 277851
rect 124336 278225 124370 278259
rect 124336 278157 124370 278191
rect 124336 278089 124370 278123
rect 122254 277749 122288 277783
rect 122254 277681 122288 277715
rect 122254 277613 122288 277647
rect 122254 277545 122288 277579
rect 122254 277477 122288 277511
rect 122254 277409 122288 277443
rect 122254 277341 122288 277375
rect 122254 277273 122288 277307
rect 124336 278021 124370 278055
rect 124336 277953 124370 277987
rect 124336 277885 124370 277919
rect 124336 277817 124370 277851
rect 124336 277749 124370 277783
rect 124336 277681 124370 277715
rect 124336 277613 124370 277647
rect 124336 277545 124370 277579
rect 124336 277477 124370 277511
rect 124336 277409 124370 277443
rect 124336 277341 124370 277375
rect 124336 277273 124370 277307
rect 122343 277187 122377 277221
rect 122411 277187 122445 277221
rect 122479 277187 122513 277221
rect 122547 277187 122581 277221
rect 122615 277187 122649 277221
rect 122683 277187 122717 277221
rect 122751 277187 122785 277221
rect 122819 277187 122853 277221
rect 122887 277187 122921 277221
rect 122955 277187 122989 277221
rect 123023 277187 123057 277221
rect 123091 277187 123125 277221
rect 123159 277187 123193 277221
rect 123227 277187 123261 277221
rect 123295 277187 123329 277221
rect 123363 277187 123397 277221
rect 123431 277187 123465 277221
rect 123499 277187 123533 277221
rect 123567 277187 123601 277221
rect 123635 277187 123669 277221
rect 123703 277187 123737 277221
rect 123771 277187 123805 277221
rect 123839 277187 123873 277221
rect 123907 277187 123941 277221
rect 123975 277187 124009 277221
rect 124043 277187 124077 277221
rect 124111 277187 124145 277221
rect 124179 277187 124213 277221
rect 124247 277187 124281 277221
rect 122404 276817 122438 276851
rect 122472 276817 122506 276851
rect 122540 276817 122574 276851
rect 122608 276817 122642 276851
rect 122676 276817 122710 276851
rect 122744 276817 122778 276851
rect 122812 276817 122846 276851
rect 122880 276817 122914 276851
rect 122948 276817 122982 276851
rect 123016 276817 123050 276851
rect 123084 276817 123118 276851
rect 123152 276817 123186 276851
rect 123220 276817 123254 276851
rect 123288 276817 123322 276851
rect 123356 276817 123390 276851
rect 123424 276817 123458 276851
rect 123492 276817 123526 276851
rect 123560 276817 123594 276851
rect 123628 276817 123662 276851
rect 123696 276817 123730 276851
rect 123764 276817 123798 276851
rect 123832 276817 123866 276851
rect 122278 276699 122312 276733
rect 123958 276699 123992 276733
rect 122278 276631 122312 276665
rect 122278 276563 122312 276597
rect 122278 276495 122312 276529
rect 123958 276631 123992 276665
rect 123958 276563 123992 276597
rect 123958 276495 123992 276529
rect 122278 276427 122312 276461
rect 123958 276427 123992 276461
rect 122404 276309 122438 276343
rect 122472 276309 122506 276343
rect 122540 276309 122574 276343
rect 122608 276309 122642 276343
rect 122676 276309 122710 276343
rect 122744 276309 122778 276343
rect 122812 276309 122846 276343
rect 122880 276309 122914 276343
rect 122948 276309 122982 276343
rect 123016 276309 123050 276343
rect 123084 276309 123118 276343
rect 123152 276309 123186 276343
rect 123220 276309 123254 276343
rect 123288 276309 123322 276343
rect 123356 276309 123390 276343
rect 123424 276309 123458 276343
rect 123492 276309 123526 276343
rect 123560 276309 123594 276343
rect 123628 276309 123662 276343
rect 123696 276309 123730 276343
rect 123764 276309 123798 276343
rect 123832 276309 123866 276343
rect 122379 275937 122413 275971
rect 122447 275937 122481 275971
rect 122515 275937 122549 275971
rect 122583 275937 122617 275971
rect 122651 275937 122685 275971
rect 122719 275937 122753 275971
rect 122787 275937 122821 275971
rect 122855 275937 122889 275971
rect 122923 275937 122957 275971
rect 122991 275937 123025 275971
rect 123059 275937 123093 275971
rect 123127 275937 123161 275971
rect 123195 275937 123229 275971
rect 123263 275937 123297 275971
rect 123331 275937 123365 275971
rect 123399 275937 123433 275971
rect 123467 275937 123501 275971
rect 123535 275937 123569 275971
rect 123603 275937 123637 275971
rect 123671 275937 123705 275971
rect 123739 275937 123773 275971
rect 123807 275937 123841 275971
rect 123875 275937 123909 275971
rect 123943 275937 123977 275971
rect 124011 275937 124045 275971
rect 124079 275937 124113 275971
rect 124147 275937 124181 275971
rect 124215 275937 124249 275971
rect 124283 275937 124317 275971
rect 124351 275937 124385 275971
rect 124419 275937 124453 275971
rect 124487 275937 124521 275971
rect 124555 275937 124589 275971
rect 124623 275937 124657 275971
rect 124691 275937 124725 275971
rect 124759 275937 124793 275971
rect 124827 275937 124861 275971
rect 122283 275812 122317 275846
rect 124923 275812 124957 275846
rect 122283 275744 122317 275778
rect 124923 275744 124957 275778
rect 122283 275676 122317 275710
rect 124923 275676 124957 275710
rect 122379 275551 122413 275585
rect 122447 275551 122481 275585
rect 122515 275551 122549 275585
rect 122583 275551 122617 275585
rect 122651 275551 122685 275585
rect 122719 275551 122753 275585
rect 122787 275551 122821 275585
rect 122855 275551 122889 275585
rect 122923 275551 122957 275585
rect 122991 275551 123025 275585
rect 123059 275551 123093 275585
rect 123127 275551 123161 275585
rect 123195 275551 123229 275585
rect 123263 275551 123297 275585
rect 123331 275551 123365 275585
rect 123399 275551 123433 275585
rect 123467 275551 123501 275585
rect 123535 275551 123569 275585
rect 123603 275551 123637 275585
rect 123671 275551 123705 275585
rect 123739 275551 123773 275585
rect 123807 275551 123841 275585
rect 123875 275551 123909 275585
rect 123943 275551 123977 275585
rect 124011 275551 124045 275585
rect 124079 275551 124113 275585
rect 124147 275551 124181 275585
rect 124215 275551 124249 275585
rect 124283 275551 124317 275585
rect 124351 275551 124385 275585
rect 124419 275551 124453 275585
rect 124487 275551 124521 275585
rect 124555 275551 124589 275585
rect 124623 275551 124657 275585
rect 124691 275551 124725 275585
rect 124759 275551 124793 275585
rect 124827 275551 124861 275585
rect 121694 275456 121728 275490
rect 121694 275388 121728 275422
rect 121694 275320 121728 275354
rect 121694 275252 121728 275286
rect 121694 275184 121728 275218
rect 121694 275116 121728 275150
rect 120237 274980 120271 275014
rect 121694 275048 121728 275082
rect 121694 274980 121728 275014
rect 120237 274912 120271 274946
rect 120237 274844 120271 274878
rect 121694 274912 121728 274946
rect 120237 274776 120271 274810
rect 121694 274844 121728 274878
rect 121694 274776 121728 274810
rect 120237 274708 120271 274742
rect 120237 274640 120271 274674
rect 120237 274572 120271 274606
rect 120237 274504 120271 274538
rect 120237 274436 120271 274470
rect 120237 274368 120271 274402
rect 120237 274300 120271 274334
rect 120237 274232 120271 274266
rect 121694 274708 121728 274742
rect 121694 274640 121728 274674
rect 121694 274572 121728 274606
rect 121694 274504 121728 274538
rect 121694 274436 121728 274470
rect 121694 274368 121728 274402
rect 121694 274300 121728 274334
rect 120237 274164 120271 274198
rect 121694 274232 121728 274266
rect 120237 274096 120271 274130
rect 121694 274164 121728 274198
rect 121694 274096 121728 274130
rect 120237 274028 120271 274062
rect 120237 273960 120271 273994
rect 121694 274028 121728 274062
rect 120237 273892 120271 273926
rect 120237 273824 120271 273858
rect 120237 273756 120271 273790
rect 120237 273688 120271 273722
rect 120237 273620 120271 273654
rect 120237 273552 120271 273586
rect 120237 273484 120271 273518
rect 121694 273960 121728 273994
rect 121694 273892 121728 273926
rect 121694 273824 121728 273858
rect 121694 273756 121728 273790
rect 121694 273688 121728 273722
rect 121694 273620 121728 273654
rect 121694 273552 121728 273586
rect 121694 273484 121728 273518
rect 120237 273416 120271 273450
rect 121694 273416 121728 273450
rect 120237 273348 120271 273382
rect 120237 273280 120271 273314
rect 121694 273348 121728 273382
rect 120237 273212 120271 273246
rect 121694 273280 121728 273314
rect 121694 273212 121728 273246
rect 120237 273144 120271 273178
rect 120237 273076 120271 273110
rect 120237 273008 120271 273042
rect 120237 272940 120271 272974
rect 120237 272872 120271 272906
rect 120237 272804 120271 272838
rect 120237 272736 120271 272770
rect 120237 272668 120271 272702
rect 121694 273144 121728 273178
rect 121694 273076 121728 273110
rect 121694 273008 121728 273042
rect 121694 272940 121728 272974
rect 121694 272872 121728 272906
rect 121694 272804 121728 272838
rect 121694 272736 121728 272770
rect 120237 272600 120271 272634
rect 121694 272668 121728 272702
rect 121694 272600 121728 272634
rect 120237 272532 120271 272566
rect 121694 272532 121728 272566
rect 120237 272464 120271 272498
rect 120237 272396 120271 272430
rect 121694 272464 121728 272498
rect 120237 272328 120271 272362
rect 120237 272260 120271 272294
rect 120237 272192 120271 272226
rect 120237 272124 120271 272158
rect 120237 272056 120271 272090
rect 120237 271988 120271 272022
rect 120237 271920 120271 271954
rect 121694 272396 121728 272430
rect 121694 272328 121728 272362
rect 121694 272260 121728 272294
rect 121694 272192 121728 272226
rect 121694 272124 121728 272158
rect 121694 272056 121728 272090
rect 121694 271988 121728 272022
rect 121694 271920 121728 271954
rect 120237 271852 120271 271886
rect 120237 271784 120271 271818
rect 121694 271852 121728 271886
rect 120237 271716 120271 271750
rect 121694 271784 121728 271818
rect 120237 271648 120271 271682
rect 121694 271716 121728 271750
rect 121694 271648 121728 271682
rect 120237 271580 120271 271614
rect 120237 271512 120271 271546
rect 120237 271444 120271 271478
rect 120237 271376 120271 271410
rect 120237 271308 120271 271342
rect 120237 271240 120271 271274
rect 120237 271172 120271 271206
rect 120237 271104 120271 271138
rect 121694 271580 121728 271614
rect 121694 271512 121728 271546
rect 121694 271444 121728 271478
rect 121694 271376 121728 271410
rect 121694 271308 121728 271342
rect 121694 271240 121728 271274
rect 121694 271172 121728 271206
rect 120237 271036 120271 271070
rect 121694 271104 121728 271138
rect 121694 271036 121728 271070
rect 120237 270968 120271 271002
rect 121694 270968 121728 271002
rect 120237 270900 120271 270934
rect 120237 270832 120271 270866
rect 121694 270900 121728 270934
rect 120237 270764 120271 270798
rect 120237 270696 120271 270730
rect 120237 270628 120271 270662
rect 120237 270560 120271 270594
rect 120237 270492 120271 270526
rect 120237 270424 120271 270458
rect 120237 270356 120271 270390
rect 121694 270832 121728 270866
rect 121694 270764 121728 270798
rect 121694 270696 121728 270730
rect 121694 270628 121728 270662
rect 121694 270560 121728 270594
rect 121694 270492 121728 270526
rect 121694 270424 121728 270458
rect 121694 270356 121728 270390
rect 120237 270288 120271 270322
rect 120237 270220 120271 270254
rect 121694 270288 121728 270322
rect 120237 270152 120271 270186
rect 121694 270220 121728 270254
rect 120237 270084 120271 270118
rect 121694 270152 121728 270186
rect 121694 270084 121728 270118
rect 120237 270016 120271 270050
rect 120237 269948 120271 269982
rect 120237 269880 120271 269914
rect 120237 269812 120271 269846
rect 120237 269744 120271 269778
rect 120237 269676 120271 269710
rect 120237 269608 120271 269642
rect 120237 269540 120271 269574
rect 121694 270016 121728 270050
rect 121694 269948 121728 269982
rect 121694 269880 121728 269914
rect 121694 269812 121728 269846
rect 121694 269744 121728 269778
rect 121694 269676 121728 269710
rect 121694 269608 121728 269642
rect 120237 269472 120271 269506
rect 121694 269540 121728 269574
rect 121694 269472 121728 269506
rect 120237 269404 120271 269438
rect 121694 269404 121728 269438
rect 120237 269336 120271 269370
rect 120237 269268 120271 269302
rect 121694 269336 121728 269370
rect 120237 269200 120271 269234
rect 121694 269268 121728 269302
rect 121694 269200 121728 269234
rect 120237 269132 120271 269166
rect 120237 269064 120271 269098
rect 121694 269132 121728 269166
rect 121694 269064 121728 269098
rect 120319 268978 120353 269012
rect 120387 268978 120421 269012
rect 120455 268978 120489 269012
rect 120523 268978 120557 269012
rect 120591 268978 120625 269012
rect 120659 268978 120693 269012
rect 120727 268978 120761 269012
rect 120795 268978 120829 269012
rect 120863 268978 120897 269012
rect 120931 268978 120965 269012
rect 120999 268978 121033 269012
rect 121067 268978 121101 269012
rect 121135 268978 121169 269012
rect 121203 268978 121237 269012
rect 121271 268978 121305 269012
rect 121339 268978 121373 269012
rect 121407 268978 121441 269012
rect 121475 268978 121509 269012
rect 121543 268978 121577 269012
rect 121611 268978 121645 269012
rect 122006 272964 122040 272998
rect 122074 272964 122108 272998
rect 122142 272964 122176 272998
rect 122210 272964 122244 272998
rect 122278 272964 122312 272998
rect 122346 272964 122380 272998
rect 122414 272964 122448 272998
rect 122482 272964 122516 272998
rect 122550 272964 122584 272998
rect 122618 272964 122652 272998
rect 122686 272964 122720 272998
rect 122754 272964 122788 272998
rect 122822 272964 122856 272998
rect 122890 272964 122924 272998
rect 122958 272964 122992 272998
rect 123026 272964 123060 272998
rect 123094 272964 123128 272998
rect 123162 272964 123196 272998
rect 123230 272964 123264 272998
rect 123298 272964 123332 272998
rect 123366 272964 123400 272998
rect 123434 272964 123468 272998
rect 121920 272883 121954 272917
rect 121920 272815 121954 272849
rect 123520 272883 123554 272917
rect 123520 272815 123554 272849
rect 121920 272747 121954 272781
rect 123520 272747 123554 272781
rect 121920 272679 121954 272713
rect 121920 272611 121954 272645
rect 123520 272679 123554 272713
rect 121920 272543 121954 272577
rect 123520 272611 123554 272645
rect 123520 272543 123554 272577
rect 121920 272475 121954 272509
rect 121920 272407 121954 272441
rect 123520 272475 123554 272509
rect 121920 272339 121954 272373
rect 121920 272271 121954 272305
rect 121920 272203 121954 272237
rect 121920 272135 121954 272169
rect 121920 272067 121954 272101
rect 121920 271999 121954 272033
rect 121920 271931 121954 271965
rect 123520 272407 123554 272441
rect 123520 272339 123554 272373
rect 123520 272271 123554 272305
rect 123520 272203 123554 272237
rect 123520 272135 123554 272169
rect 123520 272067 123554 272101
rect 123520 271999 123554 272033
rect 123520 271931 123554 271965
rect 121920 271863 121954 271897
rect 123520 271863 123554 271897
rect 121920 271795 121954 271829
rect 121920 271727 121954 271761
rect 123520 271795 123554 271829
rect 121920 271659 121954 271693
rect 123520 271727 123554 271761
rect 123520 271659 123554 271693
rect 121920 271591 121954 271625
rect 121920 271523 121954 271557
rect 121920 271455 121954 271489
rect 121920 271387 121954 271421
rect 121920 271319 121954 271353
rect 121920 271251 121954 271285
rect 121920 271183 121954 271217
rect 121920 271115 121954 271149
rect 123520 271591 123554 271625
rect 123520 271523 123554 271557
rect 123520 271455 123554 271489
rect 123520 271387 123554 271421
rect 123520 271319 123554 271353
rect 123520 271251 123554 271285
rect 123520 271183 123554 271217
rect 121920 271047 121954 271081
rect 123520 271115 123554 271149
rect 121920 270979 121954 271013
rect 123520 271047 123554 271081
rect 123520 270979 123554 271013
rect 121920 270911 121954 270945
rect 121920 270843 121954 270877
rect 123520 270911 123554 270945
rect 121920 270775 121954 270809
rect 121920 270707 121954 270741
rect 121920 270639 121954 270673
rect 121920 270571 121954 270605
rect 121920 270503 121954 270537
rect 121920 270435 121954 270469
rect 121920 270367 121954 270401
rect 123520 270843 123554 270877
rect 123520 270775 123554 270809
rect 123520 270707 123554 270741
rect 123520 270639 123554 270673
rect 123520 270571 123554 270605
rect 123520 270503 123554 270537
rect 123520 270435 123554 270469
rect 123520 270367 123554 270401
rect 121920 270299 121954 270333
rect 121920 270231 121954 270265
rect 123520 270299 123554 270333
rect 121920 270163 121954 270197
rect 123520 270231 123554 270265
rect 121920 270095 121954 270129
rect 123520 270163 123554 270197
rect 123520 270095 123554 270129
rect 121920 270027 121954 270061
rect 121920 269959 121954 269993
rect 121920 269891 121954 269925
rect 121920 269823 121954 269857
rect 121920 269755 121954 269789
rect 121920 269687 121954 269721
rect 121920 269619 121954 269653
rect 121920 269551 121954 269585
rect 123520 270027 123554 270061
rect 123520 269959 123554 269993
rect 123520 269891 123554 269925
rect 123520 269823 123554 269857
rect 123520 269755 123554 269789
rect 123520 269687 123554 269721
rect 123520 269619 123554 269653
rect 121920 269483 121954 269517
rect 123520 269551 123554 269585
rect 123520 269483 123554 269517
rect 121920 269415 121954 269449
rect 123520 269415 123554 269449
rect 121920 269347 121954 269381
rect 121920 269279 121954 269313
rect 123520 269347 123554 269381
rect 121920 269211 121954 269245
rect 123520 269279 123554 269313
rect 123520 269211 123554 269245
rect 121920 269143 121954 269177
rect 121920 269075 121954 269109
rect 123520 269143 123554 269177
rect 123520 269075 123554 269109
rect 122006 268994 122040 269028
rect 122074 268994 122108 269028
rect 122142 268994 122176 269028
rect 122210 268994 122244 269028
rect 122278 268994 122312 269028
rect 122346 268994 122380 269028
rect 122414 268994 122448 269028
rect 122482 268994 122516 269028
rect 122550 268994 122584 269028
rect 122618 268994 122652 269028
rect 122686 268994 122720 269028
rect 122754 268994 122788 269028
rect 122822 268994 122856 269028
rect 122890 268994 122924 269028
rect 122958 268994 122992 269028
rect 123026 268994 123060 269028
rect 123094 268994 123128 269028
rect 123162 268994 123196 269028
rect 123230 268994 123264 269028
rect 123298 268994 123332 269028
rect 123366 268994 123400 269028
rect 123434 268994 123468 269028
<< poly >>
rect 106357 280885 106489 280901
rect 106357 280851 106406 280885
rect 106440 280851 106489 280885
rect 106357 280813 106489 280851
rect 106757 280885 106889 280901
rect 106757 280851 106806 280885
rect 106840 280851 106889 280885
rect 106757 280813 106889 280851
rect 107157 280885 107289 280901
rect 107157 280851 107206 280885
rect 107240 280851 107289 280885
rect 107157 280813 107289 280851
rect 107557 280885 107689 280901
rect 107557 280851 107606 280885
rect 107640 280851 107689 280885
rect 107557 280813 107689 280851
rect 107957 280885 108089 280901
rect 107957 280851 108006 280885
rect 108040 280851 108089 280885
rect 107957 280813 108089 280851
rect 108357 280885 108489 280901
rect 108357 280851 108406 280885
rect 108440 280851 108489 280885
rect 108357 280813 108489 280851
rect 108757 280885 108889 280901
rect 108757 280851 108806 280885
rect 108840 280851 108889 280885
rect 108757 280813 108889 280851
rect 109157 280885 109289 280901
rect 109157 280851 109206 280885
rect 109240 280851 109289 280885
rect 109157 280813 109289 280851
rect 109557 280885 109689 280901
rect 109557 280851 109606 280885
rect 109640 280851 109689 280885
rect 109557 280813 109689 280851
rect 109957 280885 110089 280901
rect 109957 280851 110006 280885
rect 110040 280851 110089 280885
rect 109957 280813 110089 280851
rect 106357 279755 106489 279793
rect 106357 279721 106406 279755
rect 106440 279721 106489 279755
rect 106357 279705 106489 279721
rect 106757 279755 106889 279793
rect 106757 279721 106806 279755
rect 106840 279721 106889 279755
rect 106757 279705 106889 279721
rect 107157 279755 107289 279793
rect 107157 279721 107206 279755
rect 107240 279721 107289 279755
rect 107157 279705 107289 279721
rect 107557 279755 107689 279793
rect 107557 279721 107606 279755
rect 107640 279721 107689 279755
rect 107557 279705 107689 279721
rect 107957 279755 108089 279793
rect 107957 279721 108006 279755
rect 108040 279721 108089 279755
rect 107957 279705 108089 279721
rect 108357 279755 108489 279793
rect 108357 279721 108406 279755
rect 108440 279721 108489 279755
rect 108357 279705 108489 279721
rect 108757 279755 108889 279793
rect 108757 279721 108806 279755
rect 108840 279721 108889 279755
rect 108757 279705 108889 279721
rect 109157 279755 109289 279793
rect 109157 279721 109206 279755
rect 109240 279721 109289 279755
rect 109157 279705 109289 279721
rect 109557 279755 109689 279793
rect 109557 279721 109606 279755
rect 109640 279721 109689 279755
rect 109557 279705 109689 279721
rect 109957 279755 110089 279793
rect 109957 279721 110006 279755
rect 110040 279721 110089 279755
rect 109957 279705 110089 279721
rect 106271 278969 106368 279011
rect 106271 278935 106287 278969
rect 106321 278935 106368 278969
rect 106271 278901 106368 278935
rect 106271 278867 106287 278901
rect 106321 278867 106368 278901
rect 106271 278833 106368 278867
rect 106271 278799 106287 278833
rect 106321 278799 106368 278833
rect 106271 278757 106368 278799
rect 107582 278969 107679 279011
rect 107582 278935 107629 278969
rect 107663 278935 107679 278969
rect 107582 278901 107679 278935
rect 107582 278867 107629 278901
rect 107663 278867 107679 278901
rect 107582 278833 107679 278867
rect 107582 278799 107629 278833
rect 107663 278799 107679 278833
rect 107582 278757 107679 278799
rect 106271 278369 106368 278411
rect 106271 278335 106287 278369
rect 106321 278335 106368 278369
rect 106271 278301 106368 278335
rect 106271 278267 106287 278301
rect 106321 278267 106368 278301
rect 106271 278233 106368 278267
rect 106271 278199 106287 278233
rect 106321 278199 106368 278233
rect 106271 278157 106368 278199
rect 107582 278369 107679 278411
rect 107582 278335 107629 278369
rect 107663 278335 107679 278369
rect 107582 278301 107679 278335
rect 107582 278267 107629 278301
rect 107663 278267 107679 278301
rect 107582 278233 107679 278267
rect 107582 278199 107629 278233
rect 107663 278199 107679 278233
rect 107582 278157 107679 278199
rect 109777 279083 110063 279099
rect 109777 279049 109801 279083
rect 109835 279049 109869 279083
rect 109903 279049 109937 279083
rect 109971 279049 110005 279083
rect 110039 279049 110063 279083
rect 109777 279011 110063 279049
rect 109777 277935 110063 277973
rect 109777 277901 109801 277935
rect 109835 277901 109869 277935
rect 109903 277901 109937 277935
rect 109971 277901 110005 277935
rect 110039 277901 110063 277935
rect 109777 277885 110063 277901
rect 109777 277827 110063 277843
rect 109777 277793 109801 277827
rect 109835 277793 109869 277827
rect 109903 277793 109937 277827
rect 109971 277793 110005 277827
rect 110039 277793 110063 277827
rect 109777 277755 110063 277793
rect 106394 277144 106491 277164
rect 106394 277110 106410 277144
rect 106444 277110 106491 277144
rect 106394 277090 106491 277110
rect 107525 277144 107622 277164
rect 107525 277110 107572 277144
rect 107606 277110 107622 277144
rect 107525 277090 107622 277110
rect 109777 276679 110063 276717
rect 109777 276645 109801 276679
rect 109835 276645 109869 276679
rect 109903 276645 109937 276679
rect 109971 276645 110005 276679
rect 110039 276645 110063 276679
rect 109777 276629 110063 276645
rect 106854 275681 106951 275713
rect 106854 275647 106870 275681
rect 106904 275647 106951 275681
rect 106854 275613 106951 275647
rect 106854 275579 106870 275613
rect 106904 275579 106951 275613
rect 106854 275545 106951 275579
rect 106854 275511 106870 275545
rect 106904 275511 106951 275545
rect 106854 275477 106951 275511
rect 106854 275443 106870 275477
rect 106904 275443 106951 275477
rect 106854 275409 106951 275443
rect 106854 275375 106870 275409
rect 106904 275375 106951 275409
rect 106854 275341 106951 275375
rect 106854 275307 106870 275341
rect 106904 275307 106951 275341
rect 106854 275273 106951 275307
rect 106854 275239 106870 275273
rect 106904 275239 106951 275273
rect 106854 275205 106951 275239
rect 106854 275171 106870 275205
rect 106904 275171 106951 275205
rect 106854 275137 106951 275171
rect 106854 275103 106870 275137
rect 106904 275103 106951 275137
rect 106854 275069 106951 275103
rect 106854 275035 106870 275069
rect 106904 275035 106951 275069
rect 106854 275001 106951 275035
rect 106854 274967 106870 275001
rect 106904 274967 106951 275001
rect 106854 274935 106951 274967
rect 107129 275681 107226 275713
rect 107129 275647 107176 275681
rect 107210 275647 107226 275681
rect 107129 275613 107226 275647
rect 107129 275579 107176 275613
rect 107210 275579 107226 275613
rect 107129 275545 107226 275579
rect 107129 275511 107176 275545
rect 107210 275511 107226 275545
rect 107129 275477 107226 275511
rect 107129 275443 107176 275477
rect 107210 275443 107226 275477
rect 107129 275409 107226 275443
rect 107129 275375 107176 275409
rect 107210 275375 107226 275409
rect 107129 275341 107226 275375
rect 107129 275307 107176 275341
rect 107210 275307 107226 275341
rect 107129 275273 107226 275307
rect 107129 275239 107176 275273
rect 107210 275239 107226 275273
rect 107129 275205 107226 275239
rect 107129 275171 107176 275205
rect 107210 275171 107226 275205
rect 107129 275137 107226 275171
rect 107129 275103 107176 275137
rect 107210 275103 107226 275137
rect 107129 275069 107226 275103
rect 107129 275035 107176 275069
rect 107210 275035 107226 275069
rect 107129 275001 107226 275035
rect 107129 274967 107176 275001
rect 107210 274967 107226 275001
rect 107129 274935 107226 274967
rect 107354 275681 107451 275713
rect 107354 275647 107370 275681
rect 107404 275647 107451 275681
rect 107354 275613 107451 275647
rect 107354 275579 107370 275613
rect 107404 275579 107451 275613
rect 107354 275545 107451 275579
rect 107354 275511 107370 275545
rect 107404 275511 107451 275545
rect 107354 275477 107451 275511
rect 107354 275443 107370 275477
rect 107404 275443 107451 275477
rect 107354 275409 107451 275443
rect 107354 275375 107370 275409
rect 107404 275375 107451 275409
rect 107354 275341 107451 275375
rect 107354 275307 107370 275341
rect 107404 275307 107451 275341
rect 107354 275273 107451 275307
rect 107354 275239 107370 275273
rect 107404 275239 107451 275273
rect 107354 275205 107451 275239
rect 107354 275171 107370 275205
rect 107404 275171 107451 275205
rect 107354 275137 107451 275171
rect 107354 275103 107370 275137
rect 107404 275103 107451 275137
rect 107354 275069 107451 275103
rect 107354 275035 107370 275069
rect 107404 275035 107451 275069
rect 107354 275001 107451 275035
rect 107354 274967 107370 275001
rect 107404 274967 107451 275001
rect 107354 274935 107451 274967
rect 107629 275681 107726 275713
rect 107629 275647 107676 275681
rect 107710 275647 107726 275681
rect 107629 275613 107726 275647
rect 107629 275579 107676 275613
rect 107710 275579 107726 275613
rect 107629 275545 107726 275579
rect 107629 275511 107676 275545
rect 107710 275511 107726 275545
rect 107629 275477 107726 275511
rect 107629 275443 107676 275477
rect 107710 275443 107726 275477
rect 107629 275409 107726 275443
rect 107629 275375 107676 275409
rect 107710 275375 107726 275409
rect 107629 275341 107726 275375
rect 107629 275307 107676 275341
rect 107710 275307 107726 275341
rect 107629 275273 107726 275307
rect 107629 275239 107676 275273
rect 107710 275239 107726 275273
rect 107629 275205 107726 275239
rect 107629 275171 107676 275205
rect 107710 275171 107726 275205
rect 107629 275137 107726 275171
rect 107629 275103 107676 275137
rect 107710 275103 107726 275137
rect 107629 275069 107726 275103
rect 107629 275035 107676 275069
rect 107710 275035 107726 275069
rect 107629 275001 107726 275035
rect 107629 274967 107676 275001
rect 107710 274967 107726 275001
rect 107629 274935 107726 274967
rect 107854 275681 107951 275713
rect 107854 275647 107870 275681
rect 107904 275647 107951 275681
rect 107854 275613 107951 275647
rect 107854 275579 107870 275613
rect 107904 275579 107951 275613
rect 107854 275545 107951 275579
rect 107854 275511 107870 275545
rect 107904 275511 107951 275545
rect 107854 275477 107951 275511
rect 107854 275443 107870 275477
rect 107904 275443 107951 275477
rect 107854 275409 107951 275443
rect 107854 275375 107870 275409
rect 107904 275375 107951 275409
rect 107854 275341 107951 275375
rect 107854 275307 107870 275341
rect 107904 275307 107951 275341
rect 107854 275273 107951 275307
rect 107854 275239 107870 275273
rect 107904 275239 107951 275273
rect 107854 275205 107951 275239
rect 107854 275171 107870 275205
rect 107904 275171 107951 275205
rect 107854 275137 107951 275171
rect 107854 275103 107870 275137
rect 107904 275103 107951 275137
rect 107854 275069 107951 275103
rect 107854 275035 107870 275069
rect 107904 275035 107951 275069
rect 107854 275001 107951 275035
rect 107854 274967 107870 275001
rect 107904 274967 107951 275001
rect 107854 274935 107951 274967
rect 108129 275681 108226 275713
rect 108129 275647 108176 275681
rect 108210 275647 108226 275681
rect 108129 275613 108226 275647
rect 108129 275579 108176 275613
rect 108210 275579 108226 275613
rect 108129 275545 108226 275579
rect 108129 275511 108176 275545
rect 108210 275511 108226 275545
rect 108129 275477 108226 275511
rect 108129 275443 108176 275477
rect 108210 275443 108226 275477
rect 108129 275409 108226 275443
rect 108129 275375 108176 275409
rect 108210 275375 108226 275409
rect 108129 275341 108226 275375
rect 108129 275307 108176 275341
rect 108210 275307 108226 275341
rect 108129 275273 108226 275307
rect 108129 275239 108176 275273
rect 108210 275239 108226 275273
rect 108129 275205 108226 275239
rect 108129 275171 108176 275205
rect 108210 275171 108226 275205
rect 108129 275137 108226 275171
rect 108129 275103 108176 275137
rect 108210 275103 108226 275137
rect 108129 275069 108226 275103
rect 108129 275035 108176 275069
rect 108210 275035 108226 275069
rect 108129 275001 108226 275035
rect 108129 274967 108176 275001
rect 108210 274967 108226 275001
rect 108129 274935 108226 274967
rect 108354 275681 108451 275713
rect 108354 275647 108370 275681
rect 108404 275647 108451 275681
rect 108354 275613 108451 275647
rect 108354 275579 108370 275613
rect 108404 275579 108451 275613
rect 108354 275545 108451 275579
rect 108354 275511 108370 275545
rect 108404 275511 108451 275545
rect 108354 275477 108451 275511
rect 108354 275443 108370 275477
rect 108404 275443 108451 275477
rect 108354 275409 108451 275443
rect 108354 275375 108370 275409
rect 108404 275375 108451 275409
rect 108354 275341 108451 275375
rect 108354 275307 108370 275341
rect 108404 275307 108451 275341
rect 108354 275273 108451 275307
rect 108354 275239 108370 275273
rect 108404 275239 108451 275273
rect 108354 275205 108451 275239
rect 108354 275171 108370 275205
rect 108404 275171 108451 275205
rect 108354 275137 108451 275171
rect 108354 275103 108370 275137
rect 108404 275103 108451 275137
rect 108354 275069 108451 275103
rect 108354 275035 108370 275069
rect 108404 275035 108451 275069
rect 108354 275001 108451 275035
rect 108354 274967 108370 275001
rect 108404 274967 108451 275001
rect 108354 274935 108451 274967
rect 108629 275681 108726 275713
rect 108629 275647 108676 275681
rect 108710 275647 108726 275681
rect 108629 275613 108726 275647
rect 108629 275579 108676 275613
rect 108710 275579 108726 275613
rect 108629 275545 108726 275579
rect 108629 275511 108676 275545
rect 108710 275511 108726 275545
rect 108629 275477 108726 275511
rect 108629 275443 108676 275477
rect 108710 275443 108726 275477
rect 108629 275409 108726 275443
rect 108629 275375 108676 275409
rect 108710 275375 108726 275409
rect 108629 275341 108726 275375
rect 108629 275307 108676 275341
rect 108710 275307 108726 275341
rect 108629 275273 108726 275307
rect 108629 275239 108676 275273
rect 108710 275239 108726 275273
rect 108629 275205 108726 275239
rect 108629 275171 108676 275205
rect 108710 275171 108726 275205
rect 108629 275137 108726 275171
rect 108629 275103 108676 275137
rect 108710 275103 108726 275137
rect 108629 275069 108726 275103
rect 108629 275035 108676 275069
rect 108710 275035 108726 275069
rect 108629 275001 108726 275035
rect 108629 274967 108676 275001
rect 108710 274967 108726 275001
rect 108629 274935 108726 274967
rect 108854 275681 108951 275713
rect 108854 275647 108870 275681
rect 108904 275647 108951 275681
rect 108854 275613 108951 275647
rect 108854 275579 108870 275613
rect 108904 275579 108951 275613
rect 108854 275545 108951 275579
rect 108854 275511 108870 275545
rect 108904 275511 108951 275545
rect 108854 275477 108951 275511
rect 108854 275443 108870 275477
rect 108904 275443 108951 275477
rect 108854 275409 108951 275443
rect 108854 275375 108870 275409
rect 108904 275375 108951 275409
rect 108854 275341 108951 275375
rect 108854 275307 108870 275341
rect 108904 275307 108951 275341
rect 108854 275273 108951 275307
rect 108854 275239 108870 275273
rect 108904 275239 108951 275273
rect 108854 275205 108951 275239
rect 108854 275171 108870 275205
rect 108904 275171 108951 275205
rect 108854 275137 108951 275171
rect 108854 275103 108870 275137
rect 108904 275103 108951 275137
rect 108854 275069 108951 275103
rect 108854 275035 108870 275069
rect 108904 275035 108951 275069
rect 108854 275001 108951 275035
rect 108854 274967 108870 275001
rect 108904 274967 108951 275001
rect 108854 274935 108951 274967
rect 109129 275681 109226 275713
rect 109129 275647 109176 275681
rect 109210 275647 109226 275681
rect 109129 275613 109226 275647
rect 109129 275579 109176 275613
rect 109210 275579 109226 275613
rect 109129 275545 109226 275579
rect 109129 275511 109176 275545
rect 109210 275511 109226 275545
rect 109129 275477 109226 275511
rect 109129 275443 109176 275477
rect 109210 275443 109226 275477
rect 109129 275409 109226 275443
rect 109129 275375 109176 275409
rect 109210 275375 109226 275409
rect 109129 275341 109226 275375
rect 109129 275307 109176 275341
rect 109210 275307 109226 275341
rect 109129 275273 109226 275307
rect 109129 275239 109176 275273
rect 109210 275239 109226 275273
rect 109129 275205 109226 275239
rect 109129 275171 109176 275205
rect 109210 275171 109226 275205
rect 109129 275137 109226 275171
rect 109129 275103 109176 275137
rect 109210 275103 109226 275137
rect 109129 275069 109226 275103
rect 109129 275035 109176 275069
rect 109210 275035 109226 275069
rect 109129 275001 109226 275035
rect 109129 274967 109176 275001
rect 109210 274967 109226 275001
rect 109129 274935 109226 274967
rect 109354 275681 109451 275713
rect 109354 275647 109370 275681
rect 109404 275647 109451 275681
rect 109354 275613 109451 275647
rect 109354 275579 109370 275613
rect 109404 275579 109451 275613
rect 109354 275545 109451 275579
rect 109354 275511 109370 275545
rect 109404 275511 109451 275545
rect 109354 275477 109451 275511
rect 109354 275443 109370 275477
rect 109404 275443 109451 275477
rect 109354 275409 109451 275443
rect 109354 275375 109370 275409
rect 109404 275375 109451 275409
rect 109354 275341 109451 275375
rect 109354 275307 109370 275341
rect 109404 275307 109451 275341
rect 109354 275273 109451 275307
rect 109354 275239 109370 275273
rect 109404 275239 109451 275273
rect 109354 275205 109451 275239
rect 109354 275171 109370 275205
rect 109404 275171 109451 275205
rect 109354 275137 109451 275171
rect 109354 275103 109370 275137
rect 109404 275103 109451 275137
rect 109354 275069 109451 275103
rect 109354 275035 109370 275069
rect 109404 275035 109451 275069
rect 109354 275001 109451 275035
rect 109354 274967 109370 275001
rect 109404 274967 109451 275001
rect 109354 274935 109451 274967
rect 109629 275681 109726 275713
rect 109629 275647 109676 275681
rect 109710 275647 109726 275681
rect 109629 275613 109726 275647
rect 109629 275579 109676 275613
rect 109710 275579 109726 275613
rect 109629 275545 109726 275579
rect 109629 275511 109676 275545
rect 109710 275511 109726 275545
rect 109629 275477 109726 275511
rect 109629 275443 109676 275477
rect 109710 275443 109726 275477
rect 109629 275409 109726 275443
rect 109629 275375 109676 275409
rect 109710 275375 109726 275409
rect 109629 275341 109726 275375
rect 109629 275307 109676 275341
rect 109710 275307 109726 275341
rect 109629 275273 109726 275307
rect 109629 275239 109676 275273
rect 109710 275239 109726 275273
rect 109629 275205 109726 275239
rect 109629 275171 109676 275205
rect 109710 275171 109726 275205
rect 109629 275137 109726 275171
rect 109629 275103 109676 275137
rect 109710 275103 109726 275137
rect 109629 275069 109726 275103
rect 109629 275035 109676 275069
rect 109710 275035 109726 275069
rect 109629 275001 109726 275035
rect 109629 274967 109676 275001
rect 109710 274967 109726 275001
rect 109629 274935 109726 274967
rect 109440 272507 109510 272523
rect 109440 272473 109458 272507
rect 109492 272473 109510 272507
rect 109440 272426 109510 272473
rect 107459 272151 108079 272167
rect 107459 272117 107480 272151
rect 107514 272117 107548 272151
rect 107582 272117 107616 272151
rect 107650 272117 107684 272151
rect 107718 272117 107752 272151
rect 107786 272117 107820 272151
rect 107854 272117 107888 272151
rect 107922 272117 107956 272151
rect 107990 272117 108024 272151
rect 108058 272117 108079 272151
rect 107459 272079 108079 272117
rect 106981 272043 107191 272059
rect 106981 272009 107001 272043
rect 107035 272009 107069 272043
rect 107103 272009 107137 272043
rect 107171 272009 107191 272043
rect 106981 271971 107191 272009
rect 106981 271769 107191 271807
rect 106981 271735 107001 271769
rect 107035 271735 107069 271769
rect 107103 271735 107137 271769
rect 107171 271735 107191 271769
rect 106981 271719 107191 271735
rect 107459 271697 108079 271735
rect 107459 271663 107480 271697
rect 107514 271663 107548 271697
rect 107582 271663 107616 271697
rect 107650 271663 107684 271697
rect 107718 271663 107752 271697
rect 107786 271663 107820 271697
rect 107854 271663 107888 271697
rect 107922 271663 107956 271697
rect 107990 271663 108024 271697
rect 108058 271663 108079 271697
rect 107459 271647 108079 271663
rect 107085 271451 107173 271489
rect 107085 271417 107101 271451
rect 107135 271417 107173 271451
rect 107085 271383 107173 271417
rect 107085 271349 107101 271383
rect 107135 271349 107173 271383
rect 107085 271311 107173 271349
rect 108373 271451 108461 271489
rect 108373 271417 108411 271451
rect 108445 271417 108461 271451
rect 108373 271383 108461 271417
rect 108373 271349 108411 271383
rect 108445 271349 108461 271383
rect 108373 271311 108461 271349
rect 107085 271081 107173 271119
rect 107085 271047 107101 271081
rect 107135 271047 107173 271081
rect 107085 271013 107173 271047
rect 107085 270979 107101 271013
rect 107135 270979 107173 271013
rect 107085 270941 107173 270979
rect 108373 271081 108461 271119
rect 108373 271047 108411 271081
rect 108445 271047 108461 271081
rect 108373 271013 108461 271047
rect 108373 270979 108411 271013
rect 108445 270979 108461 271013
rect 108373 270941 108461 270979
rect 109440 270659 109510 270706
rect 109440 270625 109458 270659
rect 109492 270625 109510 270659
rect 109440 270609 109510 270625
rect 111436 280791 111524 280820
rect 111436 280757 111452 280791
rect 111486 280757 111524 280791
rect 111436 280723 111524 280757
rect 111436 280689 111452 280723
rect 111486 280689 111524 280723
rect 111436 280660 111524 280689
rect 112624 280791 112712 280820
rect 112624 280757 112662 280791
rect 112696 280757 112712 280791
rect 112624 280723 112712 280757
rect 112624 280689 112662 280723
rect 112696 280689 112712 280723
rect 112624 280660 112712 280689
rect 112882 280779 112970 280828
rect 112882 280745 112898 280779
rect 112932 280745 112970 280779
rect 112882 280711 112970 280745
rect 112882 280677 112898 280711
rect 112932 280677 112970 280711
rect 112882 280628 112970 280677
rect 114070 280779 114158 280828
rect 114070 280745 114108 280779
rect 114142 280745 114158 280779
rect 114070 280711 114158 280745
rect 114070 280677 114108 280711
rect 114142 280677 114158 280711
rect 114070 280628 114158 280677
rect 111436 280431 111524 280460
rect 111436 280397 111452 280431
rect 111486 280397 111524 280431
rect 111436 280363 111524 280397
rect 111436 280329 111452 280363
rect 111486 280329 111524 280363
rect 111436 280300 111524 280329
rect 112624 280431 112712 280460
rect 112624 280397 112662 280431
rect 112696 280397 112712 280431
rect 112624 280363 112712 280397
rect 112624 280329 112662 280363
rect 112696 280329 112712 280363
rect 112624 280300 112712 280329
rect 112882 280355 112970 280404
rect 112882 280321 112898 280355
rect 112932 280321 112970 280355
rect 112882 280287 112970 280321
rect 112882 280253 112898 280287
rect 112932 280253 112970 280287
rect 112882 280204 112970 280253
rect 114070 280355 114158 280404
rect 114070 280321 114108 280355
rect 114142 280321 114158 280355
rect 114070 280287 114158 280321
rect 114070 280253 114108 280287
rect 114142 280253 114158 280287
rect 114070 280204 114158 280253
rect 114560 280756 114657 280803
rect 114560 280722 114576 280756
rect 114610 280722 114657 280756
rect 114560 280688 114657 280722
rect 114560 280654 114576 280688
rect 114610 280654 114657 280688
rect 114560 280620 114657 280654
rect 114560 280586 114576 280620
rect 114610 280586 114657 280620
rect 114560 280552 114657 280586
rect 114560 280518 114576 280552
rect 114610 280518 114657 280552
rect 114560 280484 114657 280518
rect 114560 280450 114576 280484
rect 114610 280450 114657 280484
rect 114560 280403 114657 280450
rect 114857 280756 114954 280803
rect 114857 280722 114904 280756
rect 114938 280722 114954 280756
rect 114857 280688 114954 280722
rect 114857 280654 114904 280688
rect 114938 280654 114954 280688
rect 114857 280620 114954 280654
rect 114857 280586 114904 280620
rect 114938 280586 114954 280620
rect 114857 280552 114954 280586
rect 114857 280518 114904 280552
rect 114938 280518 114954 280552
rect 114857 280484 114954 280518
rect 114857 280450 114904 280484
rect 114938 280450 114954 280484
rect 114857 280403 114954 280450
rect 111436 280071 111524 280100
rect 111436 280037 111452 280071
rect 111486 280037 111524 280071
rect 111436 280003 111524 280037
rect 111436 279969 111452 280003
rect 111486 279969 111524 280003
rect 111436 279940 111524 279969
rect 112624 280071 112712 280100
rect 112624 280037 112662 280071
rect 112696 280037 112712 280071
rect 112624 280003 112712 280037
rect 112624 279969 112662 280003
rect 112696 279969 112712 280003
rect 112624 279940 112712 279969
rect 112912 279979 113000 280002
rect 112912 279945 112928 279979
rect 112962 279945 113000 279979
rect 112912 279922 113000 279945
rect 114100 279979 114188 280002
rect 114100 279945 114138 279979
rect 114172 279945 114188 279979
rect 114100 279922 114188 279945
rect 114560 280088 114657 280117
rect 114560 280054 114576 280088
rect 114610 280054 114657 280088
rect 114560 280020 114657 280054
rect 114560 279986 114576 280020
rect 114610 279986 114657 280020
rect 114560 279957 114657 279986
rect 114857 280088 114954 280117
rect 114857 280054 114904 280088
rect 114938 280054 114954 280088
rect 114857 280020 114954 280054
rect 114857 279986 114904 280020
rect 114938 279986 114954 280020
rect 114857 279957 114954 279986
rect 111436 279711 111524 279740
rect 111436 279677 111452 279711
rect 111486 279677 111524 279711
rect 111436 279643 111524 279677
rect 111436 279609 111452 279643
rect 111486 279609 111524 279643
rect 111436 279580 111524 279609
rect 112624 279711 112712 279740
rect 112624 279677 112662 279711
rect 112696 279677 112712 279711
rect 112624 279643 112712 279677
rect 112624 279609 112662 279643
rect 112696 279609 112712 279643
rect 112912 279681 113000 279704
rect 112912 279647 112928 279681
rect 112962 279647 113000 279681
rect 112912 279624 113000 279647
rect 114100 279681 114188 279704
rect 114100 279647 114138 279681
rect 114172 279647 114188 279681
rect 114100 279624 114188 279647
rect 112624 279580 112712 279609
rect 114560 279680 114657 279709
rect 114560 279646 114576 279680
rect 114610 279646 114657 279680
rect 114560 279612 114657 279646
rect 114560 279578 114576 279612
rect 114610 279578 114657 279612
rect 114560 279549 114657 279578
rect 114857 279680 114954 279709
rect 114857 279646 114904 279680
rect 114938 279646 114954 279680
rect 114857 279612 114954 279646
rect 114857 279578 114904 279612
rect 114938 279578 114954 279612
rect 114857 279549 114954 279578
rect 115251 280756 115348 280803
rect 115251 280722 115267 280756
rect 115301 280722 115348 280756
rect 115251 280688 115348 280722
rect 115251 280654 115267 280688
rect 115301 280654 115348 280688
rect 115251 280620 115348 280654
rect 115251 280586 115267 280620
rect 115301 280586 115348 280620
rect 115251 280552 115348 280586
rect 115251 280518 115267 280552
rect 115301 280518 115348 280552
rect 115251 280484 115348 280518
rect 115251 280450 115267 280484
rect 115301 280450 115348 280484
rect 115251 280403 115348 280450
rect 115548 280756 115645 280803
rect 115548 280722 115595 280756
rect 115629 280722 115645 280756
rect 115548 280688 115645 280722
rect 115548 280654 115595 280688
rect 115629 280654 115645 280688
rect 115548 280620 115645 280654
rect 115548 280586 115595 280620
rect 115629 280586 115645 280620
rect 115548 280552 115645 280586
rect 115548 280518 115595 280552
rect 115629 280518 115645 280552
rect 115548 280484 115645 280518
rect 115548 280450 115595 280484
rect 115629 280450 115645 280484
rect 115548 280403 115645 280450
rect 116047 280779 116135 280828
rect 116047 280745 116063 280779
rect 116097 280745 116135 280779
rect 116047 280711 116135 280745
rect 116047 280677 116063 280711
rect 116097 280677 116135 280711
rect 116047 280628 116135 280677
rect 117235 280779 117323 280828
rect 117235 280745 117273 280779
rect 117307 280745 117323 280779
rect 117235 280711 117323 280745
rect 117235 280677 117273 280711
rect 117307 280677 117323 280711
rect 117235 280628 117323 280677
rect 117493 280791 117581 280820
rect 117493 280757 117509 280791
rect 117543 280757 117581 280791
rect 117493 280723 117581 280757
rect 117493 280689 117509 280723
rect 117543 280689 117581 280723
rect 117493 280660 117581 280689
rect 118681 280791 118769 280820
rect 118681 280757 118719 280791
rect 118753 280757 118769 280791
rect 118681 280723 118769 280757
rect 118681 280689 118719 280723
rect 118753 280689 118769 280723
rect 118681 280660 118769 280689
rect 117493 280431 117581 280460
rect 116047 280355 116135 280404
rect 116047 280321 116063 280355
rect 116097 280321 116135 280355
rect 116047 280287 116135 280321
rect 116047 280253 116063 280287
rect 116097 280253 116135 280287
rect 116047 280204 116135 280253
rect 117235 280355 117323 280404
rect 117235 280321 117273 280355
rect 117307 280321 117323 280355
rect 117235 280287 117323 280321
rect 117493 280397 117509 280431
rect 117543 280397 117581 280431
rect 117493 280363 117581 280397
rect 117493 280329 117509 280363
rect 117543 280329 117581 280363
rect 117493 280300 117581 280329
rect 118681 280431 118769 280460
rect 118681 280397 118719 280431
rect 118753 280397 118769 280431
rect 118681 280363 118769 280397
rect 118681 280329 118719 280363
rect 118753 280329 118769 280363
rect 118681 280300 118769 280329
rect 117235 280253 117273 280287
rect 117307 280253 117323 280287
rect 117235 280204 117323 280253
rect 115251 280088 115348 280117
rect 115251 280054 115267 280088
rect 115301 280054 115348 280088
rect 115251 280020 115348 280054
rect 115251 279986 115267 280020
rect 115301 279986 115348 280020
rect 115251 279957 115348 279986
rect 115548 280088 115645 280117
rect 115548 280054 115595 280088
rect 115629 280054 115645 280088
rect 115548 280020 115645 280054
rect 115548 279986 115595 280020
rect 115629 279986 115645 280020
rect 115548 279957 115645 279986
rect 117493 280071 117581 280100
rect 117493 280037 117509 280071
rect 117543 280037 117581 280071
rect 117493 280003 117581 280037
rect 116017 279979 116105 280002
rect 116017 279945 116033 279979
rect 116067 279945 116105 279979
rect 116017 279922 116105 279945
rect 117205 279979 117293 280002
rect 117205 279945 117243 279979
rect 117277 279945 117293 279979
rect 117205 279922 117293 279945
rect 117493 279969 117509 280003
rect 117543 279969 117581 280003
rect 117493 279940 117581 279969
rect 118681 280071 118769 280100
rect 118681 280037 118719 280071
rect 118753 280037 118769 280071
rect 118681 280003 118769 280037
rect 118681 279969 118719 280003
rect 118753 279969 118769 280003
rect 118681 279940 118769 279969
rect 115251 279680 115348 279709
rect 115251 279646 115267 279680
rect 115301 279646 115348 279680
rect 115251 279612 115348 279646
rect 115251 279578 115267 279612
rect 115301 279578 115348 279612
rect 115251 279549 115348 279578
rect 115548 279680 115645 279709
rect 115548 279646 115595 279680
rect 115629 279646 115645 279680
rect 115548 279612 115645 279646
rect 115548 279578 115595 279612
rect 115629 279578 115645 279612
rect 115548 279549 115645 279578
rect 117493 279711 117581 279740
rect 116017 279681 116105 279704
rect 116017 279647 116033 279681
rect 116067 279647 116105 279681
rect 116017 279624 116105 279647
rect 117205 279681 117293 279704
rect 117205 279647 117243 279681
rect 117277 279647 117293 279681
rect 117205 279624 117293 279647
rect 117493 279677 117509 279711
rect 117543 279677 117581 279711
rect 117493 279643 117581 279677
rect 117493 279609 117509 279643
rect 117543 279609 117581 279643
rect 117493 279580 117581 279609
rect 118681 279711 118769 279740
rect 118681 279677 118719 279711
rect 118753 279677 118769 279711
rect 118681 279643 118769 279677
rect 118681 279609 118719 279643
rect 118753 279609 118769 279643
rect 118681 279580 118769 279609
rect 111436 279125 111524 279154
rect 111436 279091 111452 279125
rect 111486 279091 111524 279125
rect 111436 279057 111524 279091
rect 111436 279023 111452 279057
rect 111486 279023 111524 279057
rect 111436 278994 111524 279023
rect 112624 279125 112712 279154
rect 112624 279091 112662 279125
rect 112696 279091 112712 279125
rect 112624 279057 112712 279091
rect 112624 279023 112662 279057
rect 112696 279023 112712 279057
rect 112624 278994 112712 279023
rect 112882 279113 112970 279162
rect 112882 279079 112898 279113
rect 112932 279079 112970 279113
rect 112882 279045 112970 279079
rect 112882 279011 112898 279045
rect 112932 279011 112970 279045
rect 112882 278962 112970 279011
rect 114070 279113 114158 279162
rect 114070 279079 114108 279113
rect 114142 279079 114158 279113
rect 114070 279045 114158 279079
rect 114070 279011 114108 279045
rect 114142 279011 114158 279045
rect 114070 278962 114158 279011
rect 111436 278765 111524 278794
rect 111436 278731 111452 278765
rect 111486 278731 111524 278765
rect 111436 278697 111524 278731
rect 111436 278663 111452 278697
rect 111486 278663 111524 278697
rect 111436 278634 111524 278663
rect 112624 278765 112712 278794
rect 112624 278731 112662 278765
rect 112696 278731 112712 278765
rect 112624 278697 112712 278731
rect 112624 278663 112662 278697
rect 112696 278663 112712 278697
rect 112624 278634 112712 278663
rect 112882 278689 112970 278738
rect 112882 278655 112898 278689
rect 112932 278655 112970 278689
rect 112882 278621 112970 278655
rect 112882 278587 112898 278621
rect 112932 278587 112970 278621
rect 112882 278538 112970 278587
rect 114070 278689 114158 278738
rect 114070 278655 114108 278689
rect 114142 278655 114158 278689
rect 114070 278621 114158 278655
rect 114070 278587 114108 278621
rect 114142 278587 114158 278621
rect 114070 278538 114158 278587
rect 114560 279090 114657 279137
rect 114560 279056 114576 279090
rect 114610 279056 114657 279090
rect 114560 279022 114657 279056
rect 114560 278988 114576 279022
rect 114610 278988 114657 279022
rect 114560 278954 114657 278988
rect 114560 278920 114576 278954
rect 114610 278920 114657 278954
rect 114560 278886 114657 278920
rect 114560 278852 114576 278886
rect 114610 278852 114657 278886
rect 114560 278818 114657 278852
rect 114560 278784 114576 278818
rect 114610 278784 114657 278818
rect 114560 278737 114657 278784
rect 114857 279090 114954 279137
rect 114857 279056 114904 279090
rect 114938 279056 114954 279090
rect 114857 279022 114954 279056
rect 114857 278988 114904 279022
rect 114938 278988 114954 279022
rect 114857 278954 114954 278988
rect 114857 278920 114904 278954
rect 114938 278920 114954 278954
rect 114857 278886 114954 278920
rect 114857 278852 114904 278886
rect 114938 278852 114954 278886
rect 114857 278818 114954 278852
rect 114857 278784 114904 278818
rect 114938 278784 114954 278818
rect 114857 278737 114954 278784
rect 111436 278405 111524 278434
rect 111436 278371 111452 278405
rect 111486 278371 111524 278405
rect 111436 278337 111524 278371
rect 111436 278303 111452 278337
rect 111486 278303 111524 278337
rect 111436 278274 111524 278303
rect 112624 278405 112712 278434
rect 112624 278371 112662 278405
rect 112696 278371 112712 278405
rect 112624 278337 112712 278371
rect 112624 278303 112662 278337
rect 112696 278303 112712 278337
rect 112624 278274 112712 278303
rect 112912 278313 113000 278336
rect 112912 278279 112928 278313
rect 112962 278279 113000 278313
rect 112912 278256 113000 278279
rect 114100 278313 114188 278336
rect 114100 278279 114138 278313
rect 114172 278279 114188 278313
rect 114100 278256 114188 278279
rect 114560 278422 114657 278451
rect 114560 278388 114576 278422
rect 114610 278388 114657 278422
rect 114560 278354 114657 278388
rect 114560 278320 114576 278354
rect 114610 278320 114657 278354
rect 114560 278291 114657 278320
rect 114857 278422 114954 278451
rect 114857 278388 114904 278422
rect 114938 278388 114954 278422
rect 114857 278354 114954 278388
rect 114857 278320 114904 278354
rect 114938 278320 114954 278354
rect 114857 278291 114954 278320
rect 111436 278045 111524 278074
rect 111436 278011 111452 278045
rect 111486 278011 111524 278045
rect 111436 277977 111524 278011
rect 111436 277943 111452 277977
rect 111486 277943 111524 277977
rect 111436 277914 111524 277943
rect 112624 278045 112712 278074
rect 112624 278011 112662 278045
rect 112696 278011 112712 278045
rect 112624 277977 112712 278011
rect 112624 277943 112662 277977
rect 112696 277943 112712 277977
rect 112912 278015 113000 278038
rect 112912 277981 112928 278015
rect 112962 277981 113000 278015
rect 112912 277958 113000 277981
rect 114100 278015 114188 278038
rect 114100 277981 114138 278015
rect 114172 277981 114188 278015
rect 114100 277958 114188 277981
rect 112624 277914 112712 277943
rect 114560 278014 114657 278043
rect 114560 277980 114576 278014
rect 114610 277980 114657 278014
rect 114560 277946 114657 277980
rect 114560 277912 114576 277946
rect 114610 277912 114657 277946
rect 114560 277883 114657 277912
rect 114857 278014 114954 278043
rect 114857 277980 114904 278014
rect 114938 277980 114954 278014
rect 114857 277946 114954 277980
rect 114857 277912 114904 277946
rect 114938 277912 114954 277946
rect 114857 277883 114954 277912
rect 115251 279090 115348 279137
rect 115251 279056 115267 279090
rect 115301 279056 115348 279090
rect 115251 279022 115348 279056
rect 115251 278988 115267 279022
rect 115301 278988 115348 279022
rect 115251 278954 115348 278988
rect 115251 278920 115267 278954
rect 115301 278920 115348 278954
rect 115251 278886 115348 278920
rect 115251 278852 115267 278886
rect 115301 278852 115348 278886
rect 115251 278818 115348 278852
rect 115251 278784 115267 278818
rect 115301 278784 115348 278818
rect 115251 278737 115348 278784
rect 115548 279090 115645 279137
rect 115548 279056 115595 279090
rect 115629 279056 115645 279090
rect 115548 279022 115645 279056
rect 115548 278988 115595 279022
rect 115629 278988 115645 279022
rect 115548 278954 115645 278988
rect 115548 278920 115595 278954
rect 115629 278920 115645 278954
rect 115548 278886 115645 278920
rect 115548 278852 115595 278886
rect 115629 278852 115645 278886
rect 115548 278818 115645 278852
rect 115548 278784 115595 278818
rect 115629 278784 115645 278818
rect 115548 278737 115645 278784
rect 116047 279113 116135 279162
rect 116047 279079 116063 279113
rect 116097 279079 116135 279113
rect 116047 279045 116135 279079
rect 116047 279011 116063 279045
rect 116097 279011 116135 279045
rect 116047 278962 116135 279011
rect 117235 279113 117323 279162
rect 117235 279079 117273 279113
rect 117307 279079 117323 279113
rect 117235 279045 117323 279079
rect 117235 279011 117273 279045
rect 117307 279011 117323 279045
rect 117235 278962 117323 279011
rect 117493 279125 117581 279154
rect 117493 279091 117509 279125
rect 117543 279091 117581 279125
rect 117493 279057 117581 279091
rect 117493 279023 117509 279057
rect 117543 279023 117581 279057
rect 117493 278994 117581 279023
rect 118681 279125 118769 279154
rect 118681 279091 118719 279125
rect 118753 279091 118769 279125
rect 118681 279057 118769 279091
rect 118681 279023 118719 279057
rect 118753 279023 118769 279057
rect 118681 278994 118769 279023
rect 117493 278765 117581 278794
rect 116047 278689 116135 278738
rect 116047 278655 116063 278689
rect 116097 278655 116135 278689
rect 116047 278621 116135 278655
rect 116047 278587 116063 278621
rect 116097 278587 116135 278621
rect 116047 278538 116135 278587
rect 117235 278689 117323 278738
rect 117235 278655 117273 278689
rect 117307 278655 117323 278689
rect 117235 278621 117323 278655
rect 117493 278731 117509 278765
rect 117543 278731 117581 278765
rect 117493 278697 117581 278731
rect 117493 278663 117509 278697
rect 117543 278663 117581 278697
rect 117493 278634 117581 278663
rect 118681 278765 118769 278794
rect 118681 278731 118719 278765
rect 118753 278731 118769 278765
rect 118681 278697 118769 278731
rect 118681 278663 118719 278697
rect 118753 278663 118769 278697
rect 118681 278634 118769 278663
rect 117235 278587 117273 278621
rect 117307 278587 117323 278621
rect 117235 278538 117323 278587
rect 115251 278422 115348 278451
rect 115251 278388 115267 278422
rect 115301 278388 115348 278422
rect 115251 278354 115348 278388
rect 115251 278320 115267 278354
rect 115301 278320 115348 278354
rect 115251 278291 115348 278320
rect 115548 278422 115645 278451
rect 115548 278388 115595 278422
rect 115629 278388 115645 278422
rect 115548 278354 115645 278388
rect 115548 278320 115595 278354
rect 115629 278320 115645 278354
rect 115548 278291 115645 278320
rect 117493 278405 117581 278434
rect 117493 278371 117509 278405
rect 117543 278371 117581 278405
rect 117493 278337 117581 278371
rect 116017 278313 116105 278336
rect 116017 278279 116033 278313
rect 116067 278279 116105 278313
rect 116017 278256 116105 278279
rect 117205 278313 117293 278336
rect 117205 278279 117243 278313
rect 117277 278279 117293 278313
rect 117205 278256 117293 278279
rect 117493 278303 117509 278337
rect 117543 278303 117581 278337
rect 117493 278274 117581 278303
rect 118681 278405 118769 278434
rect 118681 278371 118719 278405
rect 118753 278371 118769 278405
rect 118681 278337 118769 278371
rect 118681 278303 118719 278337
rect 118753 278303 118769 278337
rect 118681 278274 118769 278303
rect 115251 278014 115348 278043
rect 115251 277980 115267 278014
rect 115301 277980 115348 278014
rect 115251 277946 115348 277980
rect 115251 277912 115267 277946
rect 115301 277912 115348 277946
rect 115251 277883 115348 277912
rect 115548 278014 115645 278043
rect 115548 277980 115595 278014
rect 115629 277980 115645 278014
rect 115548 277946 115645 277980
rect 115548 277912 115595 277946
rect 115629 277912 115645 277946
rect 115548 277883 115645 277912
rect 117493 278045 117581 278074
rect 116017 278015 116105 278038
rect 116017 277981 116033 278015
rect 116067 277981 116105 278015
rect 116017 277958 116105 277981
rect 117205 278015 117293 278038
rect 117205 277981 117243 278015
rect 117277 277981 117293 278015
rect 117205 277958 117293 277981
rect 117493 278011 117509 278045
rect 117543 278011 117581 278045
rect 117493 277977 117581 278011
rect 117493 277943 117509 277977
rect 117543 277943 117581 277977
rect 117493 277914 117581 277943
rect 118681 278045 118769 278074
rect 118681 278011 118719 278045
rect 118753 278011 118769 278045
rect 118681 277977 118769 278011
rect 118681 277943 118719 277977
rect 118753 277943 118769 277977
rect 118681 277914 118769 277943
rect 111436 277459 111524 277488
rect 111436 277425 111452 277459
rect 111486 277425 111524 277459
rect 111436 277391 111524 277425
rect 111436 277357 111452 277391
rect 111486 277357 111524 277391
rect 111436 277328 111524 277357
rect 112624 277459 112712 277488
rect 112624 277425 112662 277459
rect 112696 277425 112712 277459
rect 112624 277391 112712 277425
rect 112624 277357 112662 277391
rect 112696 277357 112712 277391
rect 112624 277328 112712 277357
rect 112882 277447 112970 277496
rect 112882 277413 112898 277447
rect 112932 277413 112970 277447
rect 112882 277379 112970 277413
rect 112882 277345 112898 277379
rect 112932 277345 112970 277379
rect 112882 277296 112970 277345
rect 114070 277447 114158 277496
rect 114070 277413 114108 277447
rect 114142 277413 114158 277447
rect 114070 277379 114158 277413
rect 114070 277345 114108 277379
rect 114142 277345 114158 277379
rect 114070 277296 114158 277345
rect 111436 277099 111524 277128
rect 111436 277065 111452 277099
rect 111486 277065 111524 277099
rect 111436 277031 111524 277065
rect 111436 276997 111452 277031
rect 111486 276997 111524 277031
rect 111436 276968 111524 276997
rect 112624 277099 112712 277128
rect 112624 277065 112662 277099
rect 112696 277065 112712 277099
rect 112624 277031 112712 277065
rect 112624 276997 112662 277031
rect 112696 276997 112712 277031
rect 112624 276968 112712 276997
rect 112882 277023 112970 277072
rect 112882 276989 112898 277023
rect 112932 276989 112970 277023
rect 112882 276955 112970 276989
rect 112882 276921 112898 276955
rect 112932 276921 112970 276955
rect 112882 276872 112970 276921
rect 114070 277023 114158 277072
rect 114070 276989 114108 277023
rect 114142 276989 114158 277023
rect 114070 276955 114158 276989
rect 114070 276921 114108 276955
rect 114142 276921 114158 276955
rect 114070 276872 114158 276921
rect 114560 277424 114657 277471
rect 114560 277390 114576 277424
rect 114610 277390 114657 277424
rect 114560 277356 114657 277390
rect 114560 277322 114576 277356
rect 114610 277322 114657 277356
rect 114560 277288 114657 277322
rect 114560 277254 114576 277288
rect 114610 277254 114657 277288
rect 114560 277220 114657 277254
rect 114560 277186 114576 277220
rect 114610 277186 114657 277220
rect 114560 277152 114657 277186
rect 114560 277118 114576 277152
rect 114610 277118 114657 277152
rect 114560 277071 114657 277118
rect 114857 277424 114954 277471
rect 114857 277390 114904 277424
rect 114938 277390 114954 277424
rect 114857 277356 114954 277390
rect 114857 277322 114904 277356
rect 114938 277322 114954 277356
rect 114857 277288 114954 277322
rect 114857 277254 114904 277288
rect 114938 277254 114954 277288
rect 114857 277220 114954 277254
rect 114857 277186 114904 277220
rect 114938 277186 114954 277220
rect 114857 277152 114954 277186
rect 114857 277118 114904 277152
rect 114938 277118 114954 277152
rect 114857 277071 114954 277118
rect 111436 276739 111524 276768
rect 111436 276705 111452 276739
rect 111486 276705 111524 276739
rect 111436 276671 111524 276705
rect 111436 276637 111452 276671
rect 111486 276637 111524 276671
rect 111436 276608 111524 276637
rect 112624 276739 112712 276768
rect 112624 276705 112662 276739
rect 112696 276705 112712 276739
rect 112624 276671 112712 276705
rect 112624 276637 112662 276671
rect 112696 276637 112712 276671
rect 112624 276608 112712 276637
rect 112912 276647 113000 276670
rect 112912 276613 112928 276647
rect 112962 276613 113000 276647
rect 112912 276590 113000 276613
rect 114100 276647 114188 276670
rect 114100 276613 114138 276647
rect 114172 276613 114188 276647
rect 114100 276590 114188 276613
rect 114560 276756 114657 276785
rect 114560 276722 114576 276756
rect 114610 276722 114657 276756
rect 114560 276688 114657 276722
rect 114560 276654 114576 276688
rect 114610 276654 114657 276688
rect 114560 276625 114657 276654
rect 114857 276756 114954 276785
rect 114857 276722 114904 276756
rect 114938 276722 114954 276756
rect 114857 276688 114954 276722
rect 114857 276654 114904 276688
rect 114938 276654 114954 276688
rect 114857 276625 114954 276654
rect 111436 276379 111524 276408
rect 111436 276345 111452 276379
rect 111486 276345 111524 276379
rect 111436 276311 111524 276345
rect 111436 276277 111452 276311
rect 111486 276277 111524 276311
rect 111436 276248 111524 276277
rect 112624 276379 112712 276408
rect 112624 276345 112662 276379
rect 112696 276345 112712 276379
rect 112624 276311 112712 276345
rect 112624 276277 112662 276311
rect 112696 276277 112712 276311
rect 112912 276349 113000 276372
rect 112912 276315 112928 276349
rect 112962 276315 113000 276349
rect 112912 276292 113000 276315
rect 114100 276349 114188 276372
rect 114100 276315 114138 276349
rect 114172 276315 114188 276349
rect 114100 276292 114188 276315
rect 112624 276248 112712 276277
rect 114560 276348 114657 276377
rect 114560 276314 114576 276348
rect 114610 276314 114657 276348
rect 114560 276280 114657 276314
rect 114560 276246 114576 276280
rect 114610 276246 114657 276280
rect 114560 276217 114657 276246
rect 114857 276348 114954 276377
rect 114857 276314 114904 276348
rect 114938 276314 114954 276348
rect 114857 276280 114954 276314
rect 114857 276246 114904 276280
rect 114938 276246 114954 276280
rect 114857 276217 114954 276246
rect 115251 277424 115348 277471
rect 115251 277390 115267 277424
rect 115301 277390 115348 277424
rect 115251 277356 115348 277390
rect 115251 277322 115267 277356
rect 115301 277322 115348 277356
rect 115251 277288 115348 277322
rect 115251 277254 115267 277288
rect 115301 277254 115348 277288
rect 115251 277220 115348 277254
rect 115251 277186 115267 277220
rect 115301 277186 115348 277220
rect 115251 277152 115348 277186
rect 115251 277118 115267 277152
rect 115301 277118 115348 277152
rect 115251 277071 115348 277118
rect 115548 277424 115645 277471
rect 115548 277390 115595 277424
rect 115629 277390 115645 277424
rect 115548 277356 115645 277390
rect 115548 277322 115595 277356
rect 115629 277322 115645 277356
rect 115548 277288 115645 277322
rect 115548 277254 115595 277288
rect 115629 277254 115645 277288
rect 115548 277220 115645 277254
rect 115548 277186 115595 277220
rect 115629 277186 115645 277220
rect 115548 277152 115645 277186
rect 115548 277118 115595 277152
rect 115629 277118 115645 277152
rect 115548 277071 115645 277118
rect 116047 277447 116135 277496
rect 116047 277413 116063 277447
rect 116097 277413 116135 277447
rect 116047 277379 116135 277413
rect 116047 277345 116063 277379
rect 116097 277345 116135 277379
rect 116047 277296 116135 277345
rect 117235 277447 117323 277496
rect 117235 277413 117273 277447
rect 117307 277413 117323 277447
rect 117235 277379 117323 277413
rect 117235 277345 117273 277379
rect 117307 277345 117323 277379
rect 117235 277296 117323 277345
rect 117493 277459 117581 277488
rect 117493 277425 117509 277459
rect 117543 277425 117581 277459
rect 117493 277391 117581 277425
rect 117493 277357 117509 277391
rect 117543 277357 117581 277391
rect 117493 277328 117581 277357
rect 118681 277459 118769 277488
rect 118681 277425 118719 277459
rect 118753 277425 118769 277459
rect 118681 277391 118769 277425
rect 118681 277357 118719 277391
rect 118753 277357 118769 277391
rect 118681 277328 118769 277357
rect 117493 277099 117581 277128
rect 116047 277023 116135 277072
rect 116047 276989 116063 277023
rect 116097 276989 116135 277023
rect 116047 276955 116135 276989
rect 116047 276921 116063 276955
rect 116097 276921 116135 276955
rect 116047 276872 116135 276921
rect 117235 277023 117323 277072
rect 117235 276989 117273 277023
rect 117307 276989 117323 277023
rect 117235 276955 117323 276989
rect 117493 277065 117509 277099
rect 117543 277065 117581 277099
rect 117493 277031 117581 277065
rect 117493 276997 117509 277031
rect 117543 276997 117581 277031
rect 117493 276968 117581 276997
rect 118681 277099 118769 277128
rect 118681 277065 118719 277099
rect 118753 277065 118769 277099
rect 118681 277031 118769 277065
rect 118681 276997 118719 277031
rect 118753 276997 118769 277031
rect 118681 276968 118769 276997
rect 117235 276921 117273 276955
rect 117307 276921 117323 276955
rect 117235 276872 117323 276921
rect 115251 276756 115348 276785
rect 115251 276722 115267 276756
rect 115301 276722 115348 276756
rect 115251 276688 115348 276722
rect 115251 276654 115267 276688
rect 115301 276654 115348 276688
rect 115251 276625 115348 276654
rect 115548 276756 115645 276785
rect 115548 276722 115595 276756
rect 115629 276722 115645 276756
rect 115548 276688 115645 276722
rect 115548 276654 115595 276688
rect 115629 276654 115645 276688
rect 115548 276625 115645 276654
rect 117493 276739 117581 276768
rect 117493 276705 117509 276739
rect 117543 276705 117581 276739
rect 117493 276671 117581 276705
rect 116017 276647 116105 276670
rect 116017 276613 116033 276647
rect 116067 276613 116105 276647
rect 116017 276590 116105 276613
rect 117205 276647 117293 276670
rect 117205 276613 117243 276647
rect 117277 276613 117293 276647
rect 117205 276590 117293 276613
rect 117493 276637 117509 276671
rect 117543 276637 117581 276671
rect 117493 276608 117581 276637
rect 118681 276739 118769 276768
rect 118681 276705 118719 276739
rect 118753 276705 118769 276739
rect 118681 276671 118769 276705
rect 118681 276637 118719 276671
rect 118753 276637 118769 276671
rect 118681 276608 118769 276637
rect 115251 276348 115348 276377
rect 115251 276314 115267 276348
rect 115301 276314 115348 276348
rect 115251 276280 115348 276314
rect 115251 276246 115267 276280
rect 115301 276246 115348 276280
rect 115251 276217 115348 276246
rect 115548 276348 115645 276377
rect 115548 276314 115595 276348
rect 115629 276314 115645 276348
rect 115548 276280 115645 276314
rect 115548 276246 115595 276280
rect 115629 276246 115645 276280
rect 115548 276217 115645 276246
rect 117493 276379 117581 276408
rect 116017 276349 116105 276372
rect 116017 276315 116033 276349
rect 116067 276315 116105 276349
rect 116017 276292 116105 276315
rect 117205 276349 117293 276372
rect 117205 276315 117243 276349
rect 117277 276315 117293 276349
rect 117205 276292 117293 276315
rect 117493 276345 117509 276379
rect 117543 276345 117581 276379
rect 117493 276311 117581 276345
rect 117493 276277 117509 276311
rect 117543 276277 117581 276311
rect 117493 276248 117581 276277
rect 118681 276379 118769 276408
rect 118681 276345 118719 276379
rect 118753 276345 118769 276379
rect 118681 276311 118769 276345
rect 118681 276277 118719 276311
rect 118753 276277 118769 276311
rect 118681 276248 118769 276277
rect 111436 275793 111524 275822
rect 111436 275759 111452 275793
rect 111486 275759 111524 275793
rect 111436 275725 111524 275759
rect 111436 275691 111452 275725
rect 111486 275691 111524 275725
rect 111436 275662 111524 275691
rect 112624 275793 112712 275822
rect 112624 275759 112662 275793
rect 112696 275759 112712 275793
rect 112624 275725 112712 275759
rect 112624 275691 112662 275725
rect 112696 275691 112712 275725
rect 112624 275662 112712 275691
rect 112882 275781 112970 275830
rect 112882 275747 112898 275781
rect 112932 275747 112970 275781
rect 112882 275713 112970 275747
rect 112882 275679 112898 275713
rect 112932 275679 112970 275713
rect 112882 275630 112970 275679
rect 114070 275781 114158 275830
rect 114070 275747 114108 275781
rect 114142 275747 114158 275781
rect 114070 275713 114158 275747
rect 114070 275679 114108 275713
rect 114142 275679 114158 275713
rect 114070 275630 114158 275679
rect 111436 275433 111524 275462
rect 111436 275399 111452 275433
rect 111486 275399 111524 275433
rect 111436 275365 111524 275399
rect 111436 275331 111452 275365
rect 111486 275331 111524 275365
rect 111436 275302 111524 275331
rect 112624 275433 112712 275462
rect 112624 275399 112662 275433
rect 112696 275399 112712 275433
rect 112624 275365 112712 275399
rect 112624 275331 112662 275365
rect 112696 275331 112712 275365
rect 112624 275302 112712 275331
rect 112882 275357 112970 275406
rect 112882 275323 112898 275357
rect 112932 275323 112970 275357
rect 112882 275289 112970 275323
rect 112882 275255 112898 275289
rect 112932 275255 112970 275289
rect 112882 275206 112970 275255
rect 114070 275357 114158 275406
rect 114070 275323 114108 275357
rect 114142 275323 114158 275357
rect 114070 275289 114158 275323
rect 114070 275255 114108 275289
rect 114142 275255 114158 275289
rect 114070 275206 114158 275255
rect 114560 275758 114657 275805
rect 114560 275724 114576 275758
rect 114610 275724 114657 275758
rect 114560 275690 114657 275724
rect 114560 275656 114576 275690
rect 114610 275656 114657 275690
rect 114560 275622 114657 275656
rect 114560 275588 114576 275622
rect 114610 275588 114657 275622
rect 114560 275554 114657 275588
rect 114560 275520 114576 275554
rect 114610 275520 114657 275554
rect 114560 275486 114657 275520
rect 114560 275452 114576 275486
rect 114610 275452 114657 275486
rect 114560 275405 114657 275452
rect 114857 275758 114954 275805
rect 114857 275724 114904 275758
rect 114938 275724 114954 275758
rect 114857 275690 114954 275724
rect 114857 275656 114904 275690
rect 114938 275656 114954 275690
rect 114857 275622 114954 275656
rect 114857 275588 114904 275622
rect 114938 275588 114954 275622
rect 114857 275554 114954 275588
rect 114857 275520 114904 275554
rect 114938 275520 114954 275554
rect 114857 275486 114954 275520
rect 114857 275452 114904 275486
rect 114938 275452 114954 275486
rect 114857 275405 114954 275452
rect 111436 275073 111524 275102
rect 111436 275039 111452 275073
rect 111486 275039 111524 275073
rect 111436 275005 111524 275039
rect 111436 274971 111452 275005
rect 111486 274971 111524 275005
rect 111436 274942 111524 274971
rect 112624 275073 112712 275102
rect 112624 275039 112662 275073
rect 112696 275039 112712 275073
rect 112624 275005 112712 275039
rect 112624 274971 112662 275005
rect 112696 274971 112712 275005
rect 112624 274942 112712 274971
rect 112912 274981 113000 275004
rect 112912 274947 112928 274981
rect 112962 274947 113000 274981
rect 112912 274924 113000 274947
rect 114100 274981 114188 275004
rect 114100 274947 114138 274981
rect 114172 274947 114188 274981
rect 114100 274924 114188 274947
rect 114560 275090 114657 275119
rect 114560 275056 114576 275090
rect 114610 275056 114657 275090
rect 114560 275022 114657 275056
rect 114560 274988 114576 275022
rect 114610 274988 114657 275022
rect 114560 274959 114657 274988
rect 114857 275090 114954 275119
rect 114857 275056 114904 275090
rect 114938 275056 114954 275090
rect 114857 275022 114954 275056
rect 114857 274988 114904 275022
rect 114938 274988 114954 275022
rect 114857 274959 114954 274988
rect 111436 274713 111524 274742
rect 111436 274679 111452 274713
rect 111486 274679 111524 274713
rect 111436 274645 111524 274679
rect 111436 274611 111452 274645
rect 111486 274611 111524 274645
rect 111436 274582 111524 274611
rect 112624 274713 112712 274742
rect 112624 274679 112662 274713
rect 112696 274679 112712 274713
rect 112624 274645 112712 274679
rect 112624 274611 112662 274645
rect 112696 274611 112712 274645
rect 112912 274683 113000 274706
rect 112912 274649 112928 274683
rect 112962 274649 113000 274683
rect 112912 274626 113000 274649
rect 114100 274683 114188 274706
rect 114100 274649 114138 274683
rect 114172 274649 114188 274683
rect 114100 274626 114188 274649
rect 112624 274582 112712 274611
rect 114560 274682 114657 274711
rect 114560 274648 114576 274682
rect 114610 274648 114657 274682
rect 114560 274614 114657 274648
rect 114560 274580 114576 274614
rect 114610 274580 114657 274614
rect 114560 274551 114657 274580
rect 114857 274682 114954 274711
rect 114857 274648 114904 274682
rect 114938 274648 114954 274682
rect 114857 274614 114954 274648
rect 114857 274580 114904 274614
rect 114938 274580 114954 274614
rect 114857 274551 114954 274580
rect 115251 275758 115348 275805
rect 115251 275724 115267 275758
rect 115301 275724 115348 275758
rect 115251 275690 115348 275724
rect 115251 275656 115267 275690
rect 115301 275656 115348 275690
rect 115251 275622 115348 275656
rect 115251 275588 115267 275622
rect 115301 275588 115348 275622
rect 115251 275554 115348 275588
rect 115251 275520 115267 275554
rect 115301 275520 115348 275554
rect 115251 275486 115348 275520
rect 115251 275452 115267 275486
rect 115301 275452 115348 275486
rect 115251 275405 115348 275452
rect 115548 275758 115645 275805
rect 115548 275724 115595 275758
rect 115629 275724 115645 275758
rect 115548 275690 115645 275724
rect 115548 275656 115595 275690
rect 115629 275656 115645 275690
rect 115548 275622 115645 275656
rect 115548 275588 115595 275622
rect 115629 275588 115645 275622
rect 115548 275554 115645 275588
rect 115548 275520 115595 275554
rect 115629 275520 115645 275554
rect 115548 275486 115645 275520
rect 115548 275452 115595 275486
rect 115629 275452 115645 275486
rect 115548 275405 115645 275452
rect 116047 275781 116135 275830
rect 116047 275747 116063 275781
rect 116097 275747 116135 275781
rect 116047 275713 116135 275747
rect 116047 275679 116063 275713
rect 116097 275679 116135 275713
rect 116047 275630 116135 275679
rect 117235 275781 117323 275830
rect 117235 275747 117273 275781
rect 117307 275747 117323 275781
rect 117235 275713 117323 275747
rect 117235 275679 117273 275713
rect 117307 275679 117323 275713
rect 117235 275630 117323 275679
rect 117493 275793 117581 275822
rect 117493 275759 117509 275793
rect 117543 275759 117581 275793
rect 117493 275725 117581 275759
rect 117493 275691 117509 275725
rect 117543 275691 117581 275725
rect 117493 275662 117581 275691
rect 118681 275793 118769 275822
rect 118681 275759 118719 275793
rect 118753 275759 118769 275793
rect 118681 275725 118769 275759
rect 118681 275691 118719 275725
rect 118753 275691 118769 275725
rect 118681 275662 118769 275691
rect 117493 275433 117581 275462
rect 116047 275357 116135 275406
rect 116047 275323 116063 275357
rect 116097 275323 116135 275357
rect 116047 275289 116135 275323
rect 116047 275255 116063 275289
rect 116097 275255 116135 275289
rect 116047 275206 116135 275255
rect 117235 275357 117323 275406
rect 117235 275323 117273 275357
rect 117307 275323 117323 275357
rect 117235 275289 117323 275323
rect 117493 275399 117509 275433
rect 117543 275399 117581 275433
rect 117493 275365 117581 275399
rect 117493 275331 117509 275365
rect 117543 275331 117581 275365
rect 117493 275302 117581 275331
rect 118681 275433 118769 275462
rect 118681 275399 118719 275433
rect 118753 275399 118769 275433
rect 118681 275365 118769 275399
rect 118681 275331 118719 275365
rect 118753 275331 118769 275365
rect 118681 275302 118769 275331
rect 117235 275255 117273 275289
rect 117307 275255 117323 275289
rect 117235 275206 117323 275255
rect 115251 275090 115348 275119
rect 115251 275056 115267 275090
rect 115301 275056 115348 275090
rect 115251 275022 115348 275056
rect 115251 274988 115267 275022
rect 115301 274988 115348 275022
rect 115251 274959 115348 274988
rect 115548 275090 115645 275119
rect 115548 275056 115595 275090
rect 115629 275056 115645 275090
rect 115548 275022 115645 275056
rect 115548 274988 115595 275022
rect 115629 274988 115645 275022
rect 115548 274959 115645 274988
rect 117493 275073 117581 275102
rect 117493 275039 117509 275073
rect 117543 275039 117581 275073
rect 117493 275005 117581 275039
rect 116017 274981 116105 275004
rect 116017 274947 116033 274981
rect 116067 274947 116105 274981
rect 116017 274924 116105 274947
rect 117205 274981 117293 275004
rect 117205 274947 117243 274981
rect 117277 274947 117293 274981
rect 117205 274924 117293 274947
rect 117493 274971 117509 275005
rect 117543 274971 117581 275005
rect 117493 274942 117581 274971
rect 118681 275073 118769 275102
rect 118681 275039 118719 275073
rect 118753 275039 118769 275073
rect 118681 275005 118769 275039
rect 118681 274971 118719 275005
rect 118753 274971 118769 275005
rect 118681 274942 118769 274971
rect 115251 274682 115348 274711
rect 115251 274648 115267 274682
rect 115301 274648 115348 274682
rect 115251 274614 115348 274648
rect 115251 274580 115267 274614
rect 115301 274580 115348 274614
rect 115251 274551 115348 274580
rect 115548 274682 115645 274711
rect 115548 274648 115595 274682
rect 115629 274648 115645 274682
rect 115548 274614 115645 274648
rect 115548 274580 115595 274614
rect 115629 274580 115645 274614
rect 115548 274551 115645 274580
rect 117493 274713 117581 274742
rect 116017 274683 116105 274706
rect 116017 274649 116033 274683
rect 116067 274649 116105 274683
rect 116017 274626 116105 274649
rect 117205 274683 117293 274706
rect 117205 274649 117243 274683
rect 117277 274649 117293 274683
rect 117205 274626 117293 274649
rect 117493 274679 117509 274713
rect 117543 274679 117581 274713
rect 117493 274645 117581 274679
rect 117493 274611 117509 274645
rect 117543 274611 117581 274645
rect 117493 274582 117581 274611
rect 118681 274713 118769 274742
rect 118681 274679 118719 274713
rect 118753 274679 118769 274713
rect 118681 274645 118769 274679
rect 118681 274611 118719 274645
rect 118753 274611 118769 274645
rect 118681 274582 118769 274611
rect 111436 274127 111524 274156
rect 111436 274093 111452 274127
rect 111486 274093 111524 274127
rect 111436 274059 111524 274093
rect 111436 274025 111452 274059
rect 111486 274025 111524 274059
rect 111436 273996 111524 274025
rect 112624 274127 112712 274156
rect 112624 274093 112662 274127
rect 112696 274093 112712 274127
rect 112624 274059 112712 274093
rect 112624 274025 112662 274059
rect 112696 274025 112712 274059
rect 112624 273996 112712 274025
rect 112882 274115 112970 274164
rect 112882 274081 112898 274115
rect 112932 274081 112970 274115
rect 112882 274047 112970 274081
rect 112882 274013 112898 274047
rect 112932 274013 112970 274047
rect 112882 273964 112970 274013
rect 114070 274115 114158 274164
rect 114070 274081 114108 274115
rect 114142 274081 114158 274115
rect 114070 274047 114158 274081
rect 114070 274013 114108 274047
rect 114142 274013 114158 274047
rect 114070 273964 114158 274013
rect 111436 273767 111524 273796
rect 111436 273733 111452 273767
rect 111486 273733 111524 273767
rect 111436 273699 111524 273733
rect 111436 273665 111452 273699
rect 111486 273665 111524 273699
rect 111436 273636 111524 273665
rect 112624 273767 112712 273796
rect 112624 273733 112662 273767
rect 112696 273733 112712 273767
rect 112624 273699 112712 273733
rect 112624 273665 112662 273699
rect 112696 273665 112712 273699
rect 112624 273636 112712 273665
rect 112882 273691 112970 273740
rect 112882 273657 112898 273691
rect 112932 273657 112970 273691
rect 112882 273623 112970 273657
rect 112882 273589 112898 273623
rect 112932 273589 112970 273623
rect 112882 273540 112970 273589
rect 114070 273691 114158 273740
rect 114070 273657 114108 273691
rect 114142 273657 114158 273691
rect 114070 273623 114158 273657
rect 114070 273589 114108 273623
rect 114142 273589 114158 273623
rect 114070 273540 114158 273589
rect 114560 274092 114657 274139
rect 114560 274058 114576 274092
rect 114610 274058 114657 274092
rect 114560 274024 114657 274058
rect 114560 273990 114576 274024
rect 114610 273990 114657 274024
rect 114560 273956 114657 273990
rect 114560 273922 114576 273956
rect 114610 273922 114657 273956
rect 114560 273888 114657 273922
rect 114560 273854 114576 273888
rect 114610 273854 114657 273888
rect 114560 273820 114657 273854
rect 114560 273786 114576 273820
rect 114610 273786 114657 273820
rect 114560 273739 114657 273786
rect 114857 274092 114954 274139
rect 114857 274058 114904 274092
rect 114938 274058 114954 274092
rect 114857 274024 114954 274058
rect 114857 273990 114904 274024
rect 114938 273990 114954 274024
rect 114857 273956 114954 273990
rect 114857 273922 114904 273956
rect 114938 273922 114954 273956
rect 114857 273888 114954 273922
rect 114857 273854 114904 273888
rect 114938 273854 114954 273888
rect 114857 273820 114954 273854
rect 114857 273786 114904 273820
rect 114938 273786 114954 273820
rect 114857 273739 114954 273786
rect 111436 273407 111524 273436
rect 111436 273373 111452 273407
rect 111486 273373 111524 273407
rect 111436 273339 111524 273373
rect 111436 273305 111452 273339
rect 111486 273305 111524 273339
rect 111436 273276 111524 273305
rect 112624 273407 112712 273436
rect 112624 273373 112662 273407
rect 112696 273373 112712 273407
rect 112624 273339 112712 273373
rect 112624 273305 112662 273339
rect 112696 273305 112712 273339
rect 112624 273276 112712 273305
rect 112912 273315 113000 273338
rect 112912 273281 112928 273315
rect 112962 273281 113000 273315
rect 112912 273258 113000 273281
rect 114100 273315 114188 273338
rect 114100 273281 114138 273315
rect 114172 273281 114188 273315
rect 114100 273258 114188 273281
rect 114560 273424 114657 273453
rect 114560 273390 114576 273424
rect 114610 273390 114657 273424
rect 114560 273356 114657 273390
rect 114560 273322 114576 273356
rect 114610 273322 114657 273356
rect 114560 273293 114657 273322
rect 114857 273424 114954 273453
rect 114857 273390 114904 273424
rect 114938 273390 114954 273424
rect 114857 273356 114954 273390
rect 114857 273322 114904 273356
rect 114938 273322 114954 273356
rect 114857 273293 114954 273322
rect 111436 273047 111524 273076
rect 111436 273013 111452 273047
rect 111486 273013 111524 273047
rect 111436 272979 111524 273013
rect 111436 272945 111452 272979
rect 111486 272945 111524 272979
rect 111436 272916 111524 272945
rect 112624 273047 112712 273076
rect 112624 273013 112662 273047
rect 112696 273013 112712 273047
rect 112624 272979 112712 273013
rect 112624 272945 112662 272979
rect 112696 272945 112712 272979
rect 112912 273017 113000 273040
rect 112912 272983 112928 273017
rect 112962 272983 113000 273017
rect 112912 272960 113000 272983
rect 114100 273017 114188 273040
rect 114100 272983 114138 273017
rect 114172 272983 114188 273017
rect 114100 272960 114188 272983
rect 112624 272916 112712 272945
rect 114560 273016 114657 273045
rect 114560 272982 114576 273016
rect 114610 272982 114657 273016
rect 114560 272948 114657 272982
rect 114560 272914 114576 272948
rect 114610 272914 114657 272948
rect 114560 272885 114657 272914
rect 114857 273016 114954 273045
rect 114857 272982 114904 273016
rect 114938 272982 114954 273016
rect 114857 272948 114954 272982
rect 114857 272914 114904 272948
rect 114938 272914 114954 272948
rect 114857 272885 114954 272914
rect 115251 274092 115348 274139
rect 115251 274058 115267 274092
rect 115301 274058 115348 274092
rect 115251 274024 115348 274058
rect 115251 273990 115267 274024
rect 115301 273990 115348 274024
rect 115251 273956 115348 273990
rect 115251 273922 115267 273956
rect 115301 273922 115348 273956
rect 115251 273888 115348 273922
rect 115251 273854 115267 273888
rect 115301 273854 115348 273888
rect 115251 273820 115348 273854
rect 115251 273786 115267 273820
rect 115301 273786 115348 273820
rect 115251 273739 115348 273786
rect 115548 274092 115645 274139
rect 115548 274058 115595 274092
rect 115629 274058 115645 274092
rect 115548 274024 115645 274058
rect 115548 273990 115595 274024
rect 115629 273990 115645 274024
rect 115548 273956 115645 273990
rect 115548 273922 115595 273956
rect 115629 273922 115645 273956
rect 115548 273888 115645 273922
rect 115548 273854 115595 273888
rect 115629 273854 115645 273888
rect 115548 273820 115645 273854
rect 115548 273786 115595 273820
rect 115629 273786 115645 273820
rect 115548 273739 115645 273786
rect 116047 274115 116135 274164
rect 116047 274081 116063 274115
rect 116097 274081 116135 274115
rect 116047 274047 116135 274081
rect 116047 274013 116063 274047
rect 116097 274013 116135 274047
rect 116047 273964 116135 274013
rect 117235 274115 117323 274164
rect 117235 274081 117273 274115
rect 117307 274081 117323 274115
rect 117235 274047 117323 274081
rect 117235 274013 117273 274047
rect 117307 274013 117323 274047
rect 117235 273964 117323 274013
rect 117493 274127 117581 274156
rect 117493 274093 117509 274127
rect 117543 274093 117581 274127
rect 117493 274059 117581 274093
rect 117493 274025 117509 274059
rect 117543 274025 117581 274059
rect 117493 273996 117581 274025
rect 118681 274127 118769 274156
rect 118681 274093 118719 274127
rect 118753 274093 118769 274127
rect 118681 274059 118769 274093
rect 118681 274025 118719 274059
rect 118753 274025 118769 274059
rect 118681 273996 118769 274025
rect 117493 273767 117581 273796
rect 116047 273691 116135 273740
rect 116047 273657 116063 273691
rect 116097 273657 116135 273691
rect 116047 273623 116135 273657
rect 116047 273589 116063 273623
rect 116097 273589 116135 273623
rect 116047 273540 116135 273589
rect 117235 273691 117323 273740
rect 117235 273657 117273 273691
rect 117307 273657 117323 273691
rect 117235 273623 117323 273657
rect 117493 273733 117509 273767
rect 117543 273733 117581 273767
rect 117493 273699 117581 273733
rect 117493 273665 117509 273699
rect 117543 273665 117581 273699
rect 117493 273636 117581 273665
rect 118681 273767 118769 273796
rect 118681 273733 118719 273767
rect 118753 273733 118769 273767
rect 118681 273699 118769 273733
rect 118681 273665 118719 273699
rect 118753 273665 118769 273699
rect 118681 273636 118769 273665
rect 117235 273589 117273 273623
rect 117307 273589 117323 273623
rect 117235 273540 117323 273589
rect 115251 273424 115348 273453
rect 115251 273390 115267 273424
rect 115301 273390 115348 273424
rect 115251 273356 115348 273390
rect 115251 273322 115267 273356
rect 115301 273322 115348 273356
rect 115251 273293 115348 273322
rect 115548 273424 115645 273453
rect 115548 273390 115595 273424
rect 115629 273390 115645 273424
rect 115548 273356 115645 273390
rect 115548 273322 115595 273356
rect 115629 273322 115645 273356
rect 115548 273293 115645 273322
rect 117493 273407 117581 273436
rect 117493 273373 117509 273407
rect 117543 273373 117581 273407
rect 117493 273339 117581 273373
rect 116017 273315 116105 273338
rect 116017 273281 116033 273315
rect 116067 273281 116105 273315
rect 116017 273258 116105 273281
rect 117205 273315 117293 273338
rect 117205 273281 117243 273315
rect 117277 273281 117293 273315
rect 117205 273258 117293 273281
rect 117493 273305 117509 273339
rect 117543 273305 117581 273339
rect 117493 273276 117581 273305
rect 118681 273407 118769 273436
rect 118681 273373 118719 273407
rect 118753 273373 118769 273407
rect 118681 273339 118769 273373
rect 118681 273305 118719 273339
rect 118753 273305 118769 273339
rect 118681 273276 118769 273305
rect 115251 273016 115348 273045
rect 115251 272982 115267 273016
rect 115301 272982 115348 273016
rect 115251 272948 115348 272982
rect 115251 272914 115267 272948
rect 115301 272914 115348 272948
rect 115251 272885 115348 272914
rect 115548 273016 115645 273045
rect 115548 272982 115595 273016
rect 115629 272982 115645 273016
rect 115548 272948 115645 272982
rect 115548 272914 115595 272948
rect 115629 272914 115645 272948
rect 115548 272885 115645 272914
rect 117493 273047 117581 273076
rect 116017 273017 116105 273040
rect 116017 272983 116033 273017
rect 116067 272983 116105 273017
rect 116017 272960 116105 272983
rect 117205 273017 117293 273040
rect 117205 272983 117243 273017
rect 117277 272983 117293 273017
rect 117205 272960 117293 272983
rect 117493 273013 117509 273047
rect 117543 273013 117581 273047
rect 117493 272979 117581 273013
rect 117493 272945 117509 272979
rect 117543 272945 117581 272979
rect 117493 272916 117581 272945
rect 118681 273047 118769 273076
rect 118681 273013 118719 273047
rect 118753 273013 118769 273047
rect 118681 272979 118769 273013
rect 118681 272945 118719 272979
rect 118753 272945 118769 272979
rect 118681 272916 118769 272945
rect 115881 271996 116041 272012
rect 115881 271962 115910 271996
rect 115944 271962 115978 271996
rect 116012 271962 116041 271996
rect 115881 271924 116041 271962
rect 116281 271996 116441 272012
rect 116281 271962 116310 271996
rect 116344 271962 116378 271996
rect 116412 271962 116441 271996
rect 116281 271924 116441 271962
rect 116681 271996 116841 272012
rect 116681 271962 116710 271996
rect 116744 271962 116778 271996
rect 116812 271962 116841 271996
rect 116681 271924 116841 271962
rect 117081 271996 117241 272012
rect 117081 271962 117110 271996
rect 117144 271962 117178 271996
rect 117212 271962 117241 271996
rect 117081 271924 117241 271962
rect 117481 271996 117641 272012
rect 117481 271962 117510 271996
rect 117544 271962 117578 271996
rect 117612 271962 117641 271996
rect 117481 271924 117641 271962
rect 117881 271996 118041 272012
rect 117881 271962 117910 271996
rect 117944 271962 117978 271996
rect 118012 271962 118041 271996
rect 117881 271924 118041 271962
rect 118281 271996 118441 272012
rect 118281 271962 118310 271996
rect 118344 271962 118378 271996
rect 118412 271962 118441 271996
rect 118281 271924 118441 271962
rect 118681 271996 118841 272012
rect 118681 271962 118710 271996
rect 118744 271962 118778 271996
rect 118812 271962 118841 271996
rect 118681 271924 118841 271962
rect 112578 271387 112738 271403
rect 112578 271353 112607 271387
rect 112641 271353 112675 271387
rect 112709 271353 112738 271387
rect 112578 271306 112738 271353
rect 112978 271387 113138 271403
rect 112978 271353 113007 271387
rect 113041 271353 113075 271387
rect 113109 271353 113138 271387
rect 112978 271306 113138 271353
rect 113378 271387 113538 271403
rect 113378 271353 113407 271387
rect 113441 271353 113475 271387
rect 113509 271353 113538 271387
rect 113378 271306 113538 271353
rect 113778 271387 113938 271403
rect 113778 271353 113807 271387
rect 113841 271353 113875 271387
rect 113909 271353 113938 271387
rect 113778 271306 113938 271353
rect 112578 271059 112738 271106
rect 112578 271025 112607 271059
rect 112641 271025 112675 271059
rect 112709 271025 112738 271059
rect 112578 271009 112738 271025
rect 112978 271059 113138 271106
rect 112978 271025 113007 271059
rect 113041 271025 113075 271059
rect 113109 271025 113138 271059
rect 112978 271009 113138 271025
rect 113378 271059 113538 271106
rect 113378 271025 113407 271059
rect 113441 271025 113475 271059
rect 113509 271025 113538 271059
rect 113378 271009 113538 271025
rect 113778 271059 113938 271106
rect 113778 271025 113807 271059
rect 113841 271025 113875 271059
rect 113909 271025 113938 271059
rect 113778 271009 113938 271025
rect 114637 271358 114797 271374
rect 114637 271324 114666 271358
rect 114700 271324 114734 271358
rect 114768 271324 114797 271358
rect 114637 271277 114797 271324
rect 115037 271358 115197 271374
rect 115037 271324 115066 271358
rect 115100 271324 115134 271358
rect 115168 271324 115197 271358
rect 115037 271277 115197 271324
rect 114637 271030 114797 271077
rect 114637 270996 114666 271030
rect 114700 270996 114734 271030
rect 114768 270996 114797 271030
rect 114637 270980 114797 270996
rect 115037 271030 115197 271077
rect 115037 270996 115066 271030
rect 115100 270996 115134 271030
rect 115168 270996 115197 271030
rect 115037 270980 115197 270996
rect 115881 270786 116041 270824
rect 115881 270752 115910 270786
rect 115944 270752 115978 270786
rect 116012 270752 116041 270786
rect 115881 270736 116041 270752
rect 116281 270786 116441 270824
rect 116281 270752 116310 270786
rect 116344 270752 116378 270786
rect 116412 270752 116441 270786
rect 116281 270736 116441 270752
rect 116681 270786 116841 270824
rect 116681 270752 116710 270786
rect 116744 270752 116778 270786
rect 116812 270752 116841 270786
rect 116681 270736 116841 270752
rect 117081 270786 117241 270824
rect 117081 270752 117110 270786
rect 117144 270752 117178 270786
rect 117212 270752 117241 270786
rect 117081 270736 117241 270752
rect 117481 270786 117641 270824
rect 117481 270752 117510 270786
rect 117544 270752 117578 270786
rect 117612 270752 117641 270786
rect 117481 270736 117641 270752
rect 117881 270786 118041 270824
rect 117881 270752 117910 270786
rect 117944 270752 117978 270786
rect 118012 270752 118041 270786
rect 117881 270736 118041 270752
rect 118281 270786 118441 270824
rect 118281 270752 118310 270786
rect 118344 270752 118378 270786
rect 118412 270752 118441 270786
rect 118281 270736 118441 270752
rect 118681 270786 118841 270824
rect 118681 270752 118710 270786
rect 118744 270752 118778 270786
rect 118812 270752 118841 270786
rect 118681 270736 118841 270752
rect 112560 270296 112720 270312
rect 112560 270262 112589 270296
rect 112623 270262 112657 270296
rect 112691 270262 112720 270296
rect 112560 270224 112720 270262
rect 112960 270296 113120 270312
rect 112960 270262 112989 270296
rect 113023 270262 113057 270296
rect 113091 270262 113120 270296
rect 112960 270224 113120 270262
rect 113360 270296 113520 270312
rect 113360 270262 113389 270296
rect 113423 270262 113457 270296
rect 113491 270262 113520 270296
rect 113360 270224 113520 270262
rect 113760 270296 113920 270312
rect 113760 270262 113789 270296
rect 113823 270262 113857 270296
rect 113891 270262 113920 270296
rect 113760 270224 113920 270262
rect 114160 270296 114320 270312
rect 114160 270262 114189 270296
rect 114223 270262 114257 270296
rect 114291 270262 114320 270296
rect 114160 270224 114320 270262
rect 114560 270296 114720 270312
rect 114560 270262 114589 270296
rect 114623 270262 114657 270296
rect 114691 270262 114720 270296
rect 114560 270224 114720 270262
rect 114960 270296 115120 270312
rect 114960 270262 114989 270296
rect 115023 270262 115057 270296
rect 115091 270262 115120 270296
rect 114960 270224 115120 270262
rect 115360 270296 115520 270312
rect 115360 270262 115389 270296
rect 115423 270262 115457 270296
rect 115491 270262 115520 270296
rect 115360 270224 115520 270262
rect 115760 270296 115920 270312
rect 115760 270262 115789 270296
rect 115823 270262 115857 270296
rect 115891 270262 115920 270296
rect 115760 270224 115920 270262
rect 116160 270296 116320 270312
rect 116160 270262 116189 270296
rect 116223 270262 116257 270296
rect 116291 270262 116320 270296
rect 116160 270224 116320 270262
rect 116560 270296 116720 270312
rect 116560 270262 116589 270296
rect 116623 270262 116657 270296
rect 116691 270262 116720 270296
rect 116560 270224 116720 270262
rect 116960 270296 117120 270312
rect 116960 270262 116989 270296
rect 117023 270262 117057 270296
rect 117091 270262 117120 270296
rect 116960 270224 117120 270262
rect 117360 270296 117520 270312
rect 117360 270262 117389 270296
rect 117423 270262 117457 270296
rect 117491 270262 117520 270296
rect 117360 270224 117520 270262
rect 117760 270296 117920 270312
rect 117760 270262 117789 270296
rect 117823 270262 117857 270296
rect 117891 270262 117920 270296
rect 117760 270224 117920 270262
rect 118160 270296 118320 270312
rect 118160 270262 118189 270296
rect 118223 270262 118257 270296
rect 118291 270262 118320 270296
rect 118160 270224 118320 270262
rect 118560 270296 118720 270312
rect 118560 270262 118589 270296
rect 118623 270262 118657 270296
rect 118691 270262 118720 270296
rect 118560 270224 118720 270262
rect 112560 269086 112720 269124
rect 112560 269052 112589 269086
rect 112623 269052 112657 269086
rect 112691 269052 112720 269086
rect 112560 269036 112720 269052
rect 112960 269086 113120 269124
rect 112960 269052 112989 269086
rect 113023 269052 113057 269086
rect 113091 269052 113120 269086
rect 112960 269036 113120 269052
rect 113360 269086 113520 269124
rect 113360 269052 113389 269086
rect 113423 269052 113457 269086
rect 113491 269052 113520 269086
rect 113360 269036 113520 269052
rect 113760 269086 113920 269124
rect 113760 269052 113789 269086
rect 113823 269052 113857 269086
rect 113891 269052 113920 269086
rect 113760 269036 113920 269052
rect 114160 269086 114320 269124
rect 114160 269052 114189 269086
rect 114223 269052 114257 269086
rect 114291 269052 114320 269086
rect 114160 269036 114320 269052
rect 114560 269086 114720 269124
rect 114560 269052 114589 269086
rect 114623 269052 114657 269086
rect 114691 269052 114720 269086
rect 114560 269036 114720 269052
rect 114960 269086 115120 269124
rect 114960 269052 114989 269086
rect 115023 269052 115057 269086
rect 115091 269052 115120 269086
rect 114960 269036 115120 269052
rect 115360 269086 115520 269124
rect 115360 269052 115389 269086
rect 115423 269052 115457 269086
rect 115491 269052 115520 269086
rect 115360 269036 115520 269052
rect 115760 269086 115920 269124
rect 115760 269052 115789 269086
rect 115823 269052 115857 269086
rect 115891 269052 115920 269086
rect 115760 269036 115920 269052
rect 116160 269086 116320 269124
rect 116160 269052 116189 269086
rect 116223 269052 116257 269086
rect 116291 269052 116320 269086
rect 116160 269036 116320 269052
rect 116560 269086 116720 269124
rect 116560 269052 116589 269086
rect 116623 269052 116657 269086
rect 116691 269052 116720 269086
rect 116560 269036 116720 269052
rect 116960 269086 117120 269124
rect 116960 269052 116989 269086
rect 117023 269052 117057 269086
rect 117091 269052 117120 269086
rect 116960 269036 117120 269052
rect 117360 269086 117520 269124
rect 117360 269052 117389 269086
rect 117423 269052 117457 269086
rect 117491 269052 117520 269086
rect 117360 269036 117520 269052
rect 117760 269086 117920 269124
rect 117760 269052 117789 269086
rect 117823 269052 117857 269086
rect 117891 269052 117920 269086
rect 117760 269036 117920 269052
rect 118160 269086 118320 269124
rect 118160 269052 118189 269086
rect 118223 269052 118257 269086
rect 118291 269052 118320 269086
rect 118160 269036 118320 269052
rect 118560 269086 118720 269124
rect 118560 269052 118589 269086
rect 118623 269052 118657 269086
rect 118691 269052 118720 269086
rect 118560 269036 118720 269052
rect 120429 280718 120829 280734
rect 120429 280684 120476 280718
rect 120510 280684 120544 280718
rect 120578 280684 120612 280718
rect 120646 280684 120680 280718
rect 120714 280684 120748 280718
rect 120782 280684 120829 280718
rect 120429 280637 120829 280684
rect 121129 280718 121529 280734
rect 121129 280684 121176 280718
rect 121210 280684 121244 280718
rect 121278 280684 121312 280718
rect 121346 280684 121380 280718
rect 121414 280684 121448 280718
rect 121482 280684 121529 280718
rect 121129 280637 121529 280684
rect 120429 280490 120829 280537
rect 120429 280456 120476 280490
rect 120510 280456 120544 280490
rect 120578 280456 120612 280490
rect 120646 280456 120680 280490
rect 120714 280456 120748 280490
rect 120782 280456 120829 280490
rect 120429 280440 120829 280456
rect 121129 280490 121529 280537
rect 121129 280456 121176 280490
rect 121210 280456 121244 280490
rect 121278 280456 121312 280490
rect 121346 280456 121380 280490
rect 121414 280456 121448 280490
rect 121482 280456 121529 280490
rect 121129 280440 121529 280456
rect 120429 280334 120829 280350
rect 120429 280300 120476 280334
rect 120510 280300 120544 280334
rect 120578 280300 120612 280334
rect 120646 280300 120680 280334
rect 120714 280300 120748 280334
rect 120782 280300 120829 280334
rect 120429 280253 120829 280300
rect 121129 280334 121529 280350
rect 121129 280300 121176 280334
rect 121210 280300 121244 280334
rect 121278 280300 121312 280334
rect 121346 280300 121380 280334
rect 121414 280300 121448 280334
rect 121482 280300 121529 280334
rect 121129 280253 121529 280300
rect 120429 279706 120829 279753
rect 120429 279672 120476 279706
rect 120510 279672 120544 279706
rect 120578 279672 120612 279706
rect 120646 279672 120680 279706
rect 120714 279672 120748 279706
rect 120782 279672 120829 279706
rect 120429 279656 120829 279672
rect 121129 279706 121529 279753
rect 121129 279672 121176 279706
rect 121210 279672 121244 279706
rect 121278 279672 121312 279706
rect 121346 279672 121380 279706
rect 121414 279672 121448 279706
rect 121482 279672 121529 279706
rect 121129 279656 121529 279672
rect 120429 279550 120829 279566
rect 120429 279516 120476 279550
rect 120510 279516 120544 279550
rect 120578 279516 120612 279550
rect 120646 279516 120680 279550
rect 120714 279516 120748 279550
rect 120782 279516 120829 279550
rect 120429 279469 120829 279516
rect 121129 279550 121529 279566
rect 121129 279516 121176 279550
rect 121210 279516 121244 279550
rect 121278 279516 121312 279550
rect 121346 279516 121380 279550
rect 121414 279516 121448 279550
rect 121482 279516 121529 279550
rect 121129 279469 121529 279516
rect 120429 278922 120829 278969
rect 120429 278888 120476 278922
rect 120510 278888 120544 278922
rect 120578 278888 120612 278922
rect 120646 278888 120680 278922
rect 120714 278888 120748 278922
rect 120782 278888 120829 278922
rect 120429 278872 120829 278888
rect 121129 278922 121529 278969
rect 121129 278888 121176 278922
rect 121210 278888 121244 278922
rect 121278 278888 121312 278922
rect 121346 278888 121380 278922
rect 121414 278888 121448 278922
rect 121482 278888 121529 278922
rect 121129 278872 121529 278888
rect 122356 280504 122756 280520
rect 122356 280470 122403 280504
rect 122437 280470 122471 280504
rect 122505 280470 122539 280504
rect 122573 280470 122607 280504
rect 122641 280470 122675 280504
rect 122709 280470 122756 280504
rect 122356 280423 122756 280470
rect 123056 280504 123456 280520
rect 123056 280470 123103 280504
rect 123137 280470 123171 280504
rect 123205 280470 123239 280504
rect 123273 280470 123307 280504
rect 123341 280470 123375 280504
rect 123409 280470 123456 280504
rect 123056 280423 123456 280470
rect 122356 279876 122756 279923
rect 122356 279842 122403 279876
rect 122437 279842 122471 279876
rect 122505 279842 122539 279876
rect 122573 279842 122607 279876
rect 122641 279842 122675 279876
rect 122709 279842 122756 279876
rect 122356 279826 122756 279842
rect 123056 279876 123456 279923
rect 123056 279842 123103 279876
rect 123137 279842 123171 279876
rect 123205 279842 123239 279876
rect 123273 279842 123307 279876
rect 123341 279842 123375 279876
rect 123409 279842 123456 279876
rect 123056 279826 123456 279842
rect 122356 279720 122756 279736
rect 122356 279686 122403 279720
rect 122437 279686 122471 279720
rect 122505 279686 122539 279720
rect 122573 279686 122607 279720
rect 122641 279686 122675 279720
rect 122709 279686 122756 279720
rect 122356 279639 122756 279686
rect 123056 279720 123456 279736
rect 123056 279686 123103 279720
rect 123137 279686 123171 279720
rect 123205 279686 123239 279720
rect 123273 279686 123307 279720
rect 123341 279686 123375 279720
rect 123409 279686 123456 279720
rect 123056 279639 123456 279686
rect 122356 279092 122756 279139
rect 122356 279058 122403 279092
rect 122437 279058 122471 279092
rect 122505 279058 122539 279092
rect 122573 279058 122607 279092
rect 122641 279058 122675 279092
rect 122709 279058 122756 279092
rect 122356 279042 122756 279058
rect 123056 279092 123456 279139
rect 123056 279058 123103 279092
rect 123137 279058 123171 279092
rect 123205 279058 123239 279092
rect 123273 279058 123307 279092
rect 123341 279058 123375 279092
rect 123409 279058 123456 279092
rect 123056 279042 123456 279058
rect 120429 278766 120829 278782
rect 120429 278732 120476 278766
rect 120510 278732 120544 278766
rect 120578 278732 120612 278766
rect 120646 278732 120680 278766
rect 120714 278732 120748 278766
rect 120782 278732 120829 278766
rect 120429 278685 120829 278732
rect 121129 278766 121529 278782
rect 121129 278732 121176 278766
rect 121210 278732 121244 278766
rect 121278 278732 121312 278766
rect 121346 278732 121380 278766
rect 121414 278732 121448 278766
rect 121482 278732 121529 278766
rect 121129 278685 121529 278732
rect 120429 278138 120829 278185
rect 120429 278104 120476 278138
rect 120510 278104 120544 278138
rect 120578 278104 120612 278138
rect 120646 278104 120680 278138
rect 120714 278104 120748 278138
rect 120782 278104 120829 278138
rect 120429 278088 120829 278104
rect 121129 278138 121529 278185
rect 121129 278104 121176 278138
rect 121210 278104 121244 278138
rect 121278 278104 121312 278138
rect 121346 278104 121380 278138
rect 121414 278104 121448 278138
rect 121482 278104 121529 278138
rect 121129 278088 121529 278104
rect 120429 277982 120829 277998
rect 120429 277948 120476 277982
rect 120510 277948 120544 277982
rect 120578 277948 120612 277982
rect 120646 277948 120680 277982
rect 120714 277948 120748 277982
rect 120782 277948 120829 277982
rect 120429 277901 120829 277948
rect 121129 277982 121529 277998
rect 121129 277948 121176 277982
rect 121210 277948 121244 277982
rect 121278 277948 121312 277982
rect 121346 277948 121380 277982
rect 121414 277948 121448 277982
rect 121482 277948 121529 277982
rect 121129 277901 121529 277948
rect 120429 277354 120829 277401
rect 120429 277320 120476 277354
rect 120510 277320 120544 277354
rect 120578 277320 120612 277354
rect 120646 277320 120680 277354
rect 120714 277320 120748 277354
rect 120782 277320 120829 277354
rect 120429 277304 120829 277320
rect 121129 277354 121529 277401
rect 121129 277320 121176 277354
rect 121210 277320 121244 277354
rect 121278 277320 121312 277354
rect 121346 277320 121380 277354
rect 121414 277320 121448 277354
rect 121482 277320 121529 277354
rect 121129 277304 121529 277320
rect 120429 277198 120829 277214
rect 120429 277164 120476 277198
rect 120510 277164 120544 277198
rect 120578 277164 120612 277198
rect 120646 277164 120680 277198
rect 120714 277164 120748 277198
rect 120782 277164 120829 277198
rect 120429 277117 120829 277164
rect 121129 277198 121529 277214
rect 121129 277164 121176 277198
rect 121210 277164 121244 277198
rect 121278 277164 121312 277198
rect 121346 277164 121380 277198
rect 121414 277164 121448 277198
rect 121482 277164 121529 277198
rect 121129 277117 121529 277164
rect 120429 276570 120829 276617
rect 120429 276536 120476 276570
rect 120510 276536 120544 276570
rect 120578 276536 120612 276570
rect 120646 276536 120680 276570
rect 120714 276536 120748 276570
rect 120782 276536 120829 276570
rect 120429 276520 120829 276536
rect 121129 276570 121529 276617
rect 121129 276536 121176 276570
rect 121210 276536 121244 276570
rect 121278 276536 121312 276570
rect 121346 276536 121380 276570
rect 121414 276536 121448 276570
rect 121482 276536 121529 276570
rect 121129 276520 121529 276536
rect 120429 276414 120829 276430
rect 120429 276380 120476 276414
rect 120510 276380 120544 276414
rect 120578 276380 120612 276414
rect 120646 276380 120680 276414
rect 120714 276380 120748 276414
rect 120782 276380 120829 276414
rect 120429 276333 120829 276380
rect 121129 276414 121529 276430
rect 121129 276380 121176 276414
rect 121210 276380 121244 276414
rect 121278 276380 121312 276414
rect 121346 276380 121380 276414
rect 121414 276380 121448 276414
rect 121482 276380 121529 276414
rect 121129 276333 121529 276380
rect 120429 275786 120829 275833
rect 120429 275752 120476 275786
rect 120510 275752 120544 275786
rect 120578 275752 120612 275786
rect 120646 275752 120680 275786
rect 120714 275752 120748 275786
rect 120782 275752 120829 275786
rect 120429 275736 120829 275752
rect 121129 275786 121529 275833
rect 121129 275752 121176 275786
rect 121210 275752 121244 275786
rect 121278 275752 121312 275786
rect 121346 275752 121380 275786
rect 121414 275752 121448 275786
rect 121482 275752 121529 275786
rect 121129 275736 121529 275752
rect 120429 275630 120829 275646
rect 120429 275596 120476 275630
rect 120510 275596 120544 275630
rect 120578 275596 120612 275630
rect 120646 275596 120680 275630
rect 120714 275596 120748 275630
rect 120782 275596 120829 275630
rect 120429 275549 120829 275596
rect 121129 275630 121529 275646
rect 121129 275596 121176 275630
rect 121210 275596 121244 275630
rect 121278 275596 121312 275630
rect 121346 275596 121380 275630
rect 121414 275596 121448 275630
rect 121482 275596 121529 275630
rect 121129 275549 121529 275596
rect 122414 278347 123290 278363
rect 122414 278313 122461 278347
rect 122495 278313 122529 278347
rect 122563 278313 122597 278347
rect 122631 278313 122665 278347
rect 122699 278313 122733 278347
rect 122767 278313 122801 278347
rect 122835 278313 122869 278347
rect 122903 278313 122937 278347
rect 122971 278313 123005 278347
rect 123039 278313 123073 278347
rect 123107 278313 123141 278347
rect 123175 278313 123209 278347
rect 123243 278313 123290 278347
rect 122414 278266 123290 278313
rect 123656 278161 124210 278177
rect 123656 278127 123678 278161
rect 123712 278127 123746 278161
rect 123780 278127 123814 278161
rect 123848 278127 123882 278161
rect 123916 278127 123950 278161
rect 123984 278127 124018 278161
rect 124052 278127 124086 278161
rect 124120 278127 124154 278161
rect 124188 278127 124210 278161
rect 123656 278080 124210 278127
rect 122414 277745 123290 277792
rect 122414 277711 122461 277745
rect 122495 277711 122529 277745
rect 122563 277711 122597 277745
rect 122631 277711 122665 277745
rect 122699 277711 122733 277745
rect 122767 277711 122801 277745
rect 122835 277711 122869 277745
rect 122903 277711 122937 277745
rect 122971 277711 123005 277745
rect 123039 277711 123073 277745
rect 123107 277711 123141 277745
rect 123175 277711 123209 277745
rect 123243 277711 123290 277745
rect 122414 277695 123290 277711
rect 122416 277581 123216 277597
rect 122416 277547 122459 277581
rect 122493 277547 122527 277581
rect 122561 277547 122595 277581
rect 122629 277547 122663 277581
rect 122697 277547 122731 277581
rect 122765 277547 122799 277581
rect 122833 277547 122867 277581
rect 122901 277547 122935 277581
rect 122969 277547 123003 277581
rect 123037 277547 123071 277581
rect 123105 277547 123139 277581
rect 123173 277547 123216 277581
rect 122416 277500 123216 277547
rect 122416 277353 123216 277400
rect 122416 277319 122459 277353
rect 122493 277319 122527 277353
rect 122561 277319 122595 277353
rect 122629 277319 122663 277353
rect 122697 277319 122731 277353
rect 122765 277319 122799 277353
rect 122833 277319 122867 277353
rect 122901 277319 122935 277353
rect 122969 277319 123003 277353
rect 123037 277319 123071 277353
rect 123105 277319 123139 277353
rect 123173 277319 123216 277353
rect 122416 277303 123216 277319
rect 123656 277347 124210 277394
rect 123656 277313 123678 277347
rect 123712 277313 123746 277347
rect 123780 277313 123814 277347
rect 123848 277313 123882 277347
rect 123916 277313 123950 277347
rect 123984 277313 124018 277347
rect 124052 277313 124086 277347
rect 124120 277313 124154 277347
rect 124188 277313 124210 277347
rect 123656 277297 124210 277313
rect 122438 276749 123832 276765
rect 122438 276715 122472 276749
rect 122506 276715 122540 276749
rect 122574 276715 122608 276749
rect 122642 276715 122676 276749
rect 122710 276715 122744 276749
rect 122778 276715 122812 276749
rect 122846 276715 122880 276749
rect 122914 276715 122948 276749
rect 122982 276715 123016 276749
rect 123050 276715 123084 276749
rect 123118 276715 123152 276749
rect 123186 276715 123220 276749
rect 123254 276715 123288 276749
rect 123322 276715 123356 276749
rect 123390 276715 123424 276749
rect 123458 276715 123492 276749
rect 123526 276715 123560 276749
rect 123594 276715 123628 276749
rect 123662 276715 123696 276749
rect 123730 276715 123764 276749
rect 123798 276715 123832 276749
rect 122438 276668 123832 276715
rect 122438 276445 123832 276492
rect 122438 276411 122472 276445
rect 122506 276411 122540 276445
rect 122574 276411 122608 276445
rect 122642 276411 122676 276445
rect 122710 276411 122744 276445
rect 122778 276411 122812 276445
rect 122846 276411 122880 276445
rect 122914 276411 122948 276445
rect 122982 276411 123016 276445
rect 123050 276411 123084 276445
rect 123118 276411 123152 276445
rect 123186 276411 123220 276445
rect 123254 276411 123288 276445
rect 123322 276411 123356 276445
rect 123390 276411 123424 276445
rect 123458 276411 123492 276445
rect 123526 276411 123560 276445
rect 123594 276411 123628 276445
rect 123662 276411 123696 276445
rect 123730 276411 123764 276445
rect 123798 276411 123832 276445
rect 122438 276395 123832 276411
rect 122369 275778 122466 275811
rect 122369 275744 122385 275778
rect 122419 275744 122466 275778
rect 122369 275711 122466 275744
rect 122866 275778 122963 275811
rect 122866 275744 122913 275778
rect 122947 275744 122963 275778
rect 122866 275711 122963 275744
rect 123005 275778 123102 275811
rect 123005 275744 123021 275778
rect 123055 275744 123102 275778
rect 123005 275711 123102 275744
rect 123502 275778 123599 275811
rect 123502 275744 123549 275778
rect 123583 275744 123599 275778
rect 123502 275711 123599 275744
rect 123641 275778 123738 275811
rect 123641 275744 123657 275778
rect 123691 275744 123738 275778
rect 123641 275711 123738 275744
rect 124138 275778 124235 275811
rect 124138 275744 124185 275778
rect 124219 275744 124235 275778
rect 124138 275711 124235 275744
rect 124277 275778 124374 275811
rect 124277 275744 124293 275778
rect 124327 275744 124374 275778
rect 124277 275711 124374 275744
rect 124774 275778 124871 275811
rect 124774 275744 124821 275778
rect 124855 275744 124871 275778
rect 124774 275711 124871 275744
rect 120429 275002 120829 275049
rect 120429 274968 120476 275002
rect 120510 274968 120544 275002
rect 120578 274968 120612 275002
rect 120646 274968 120680 275002
rect 120714 274968 120748 275002
rect 120782 274968 120829 275002
rect 120429 274952 120829 274968
rect 121129 275002 121529 275049
rect 121129 274968 121176 275002
rect 121210 274968 121244 275002
rect 121278 274968 121312 275002
rect 121346 274968 121380 275002
rect 121414 274968 121448 275002
rect 121482 274968 121529 275002
rect 121129 274952 121529 274968
rect 120429 274846 120829 274862
rect 120429 274812 120476 274846
rect 120510 274812 120544 274846
rect 120578 274812 120612 274846
rect 120646 274812 120680 274846
rect 120714 274812 120748 274846
rect 120782 274812 120829 274846
rect 120429 274765 120829 274812
rect 121129 274846 121529 274862
rect 121129 274812 121176 274846
rect 121210 274812 121244 274846
rect 121278 274812 121312 274846
rect 121346 274812 121380 274846
rect 121414 274812 121448 274846
rect 121482 274812 121529 274846
rect 121129 274765 121529 274812
rect 122952 274934 123952 274950
rect 122952 274900 122993 274934
rect 123027 274900 123061 274934
rect 123095 274900 123129 274934
rect 123163 274900 123197 274934
rect 123231 274900 123265 274934
rect 123299 274900 123333 274934
rect 123367 274900 123401 274934
rect 123435 274900 123469 274934
rect 123503 274900 123537 274934
rect 123571 274900 123605 274934
rect 123639 274900 123673 274934
rect 123707 274900 123741 274934
rect 123775 274900 123809 274934
rect 123843 274900 123877 274934
rect 123911 274900 123952 274934
rect 122952 274862 123952 274900
rect 122952 274624 123952 274662
rect 122952 274590 122993 274624
rect 123027 274590 123061 274624
rect 123095 274590 123129 274624
rect 123163 274590 123197 274624
rect 123231 274590 123265 274624
rect 123299 274590 123333 274624
rect 123367 274590 123401 274624
rect 123435 274590 123469 274624
rect 123503 274590 123537 274624
rect 123571 274590 123605 274624
rect 123639 274590 123673 274624
rect 123707 274590 123741 274624
rect 123775 274590 123809 274624
rect 123843 274590 123877 274624
rect 123911 274590 123952 274624
rect 122952 274574 123952 274590
rect 120429 274218 120829 274265
rect 120429 274184 120476 274218
rect 120510 274184 120544 274218
rect 120578 274184 120612 274218
rect 120646 274184 120680 274218
rect 120714 274184 120748 274218
rect 120782 274184 120829 274218
rect 120429 274168 120829 274184
rect 121129 274218 121529 274265
rect 121129 274184 121176 274218
rect 121210 274184 121244 274218
rect 121278 274184 121312 274218
rect 121346 274184 121380 274218
rect 121414 274184 121448 274218
rect 121482 274184 121529 274218
rect 121129 274168 121529 274184
rect 120429 274062 120829 274078
rect 120429 274028 120476 274062
rect 120510 274028 120544 274062
rect 120578 274028 120612 274062
rect 120646 274028 120680 274062
rect 120714 274028 120748 274062
rect 120782 274028 120829 274062
rect 120429 273981 120829 274028
rect 121129 274062 121529 274078
rect 121129 274028 121176 274062
rect 121210 274028 121244 274062
rect 121278 274028 121312 274062
rect 121346 274028 121380 274062
rect 121414 274028 121448 274062
rect 121482 274028 121529 274062
rect 121129 273981 121529 274028
rect 122277 274350 122477 274366
rect 122277 274316 122326 274350
rect 122360 274316 122394 274350
rect 122428 274316 122477 274350
rect 122277 274278 122477 274316
rect 122693 274350 122893 274366
rect 122693 274316 122742 274350
rect 122776 274316 122810 274350
rect 122844 274316 122893 274350
rect 122693 274278 122893 274316
rect 123109 274350 123309 274366
rect 123109 274316 123158 274350
rect 123192 274316 123226 274350
rect 123260 274316 123309 274350
rect 123109 274278 123309 274316
rect 123525 274350 123725 274366
rect 123525 274316 123574 274350
rect 123608 274316 123642 274350
rect 123676 274316 123725 274350
rect 123525 274278 123725 274316
rect 123941 274350 124141 274366
rect 123941 274316 123990 274350
rect 124024 274316 124058 274350
rect 124092 274316 124141 274350
rect 123941 274278 124141 274316
rect 124357 274350 124557 274366
rect 124357 274316 124406 274350
rect 124440 274316 124474 274350
rect 124508 274316 124557 274350
rect 124357 274278 124557 274316
rect 122277 273740 122477 273778
rect 122277 273706 122326 273740
rect 122360 273706 122394 273740
rect 122428 273706 122477 273740
rect 122277 273690 122477 273706
rect 122693 273740 122893 273778
rect 122693 273706 122742 273740
rect 122776 273706 122810 273740
rect 122844 273706 122893 273740
rect 122693 273690 122893 273706
rect 123109 273740 123309 273778
rect 123109 273706 123158 273740
rect 123192 273706 123226 273740
rect 123260 273706 123309 273740
rect 123109 273690 123309 273706
rect 123525 273740 123725 273778
rect 123525 273706 123574 273740
rect 123608 273706 123642 273740
rect 123676 273706 123725 273740
rect 123525 273690 123725 273706
rect 123941 273740 124141 273778
rect 123941 273706 123990 273740
rect 124024 273706 124058 273740
rect 124092 273706 124141 273740
rect 123941 273690 124141 273706
rect 124357 273740 124557 273778
rect 124357 273706 124406 273740
rect 124440 273706 124474 273740
rect 124508 273706 124557 273740
rect 124357 273690 124557 273706
rect 120429 273434 120829 273481
rect 120429 273400 120476 273434
rect 120510 273400 120544 273434
rect 120578 273400 120612 273434
rect 120646 273400 120680 273434
rect 120714 273400 120748 273434
rect 120782 273400 120829 273434
rect 120429 273384 120829 273400
rect 121129 273434 121529 273481
rect 121129 273400 121176 273434
rect 121210 273400 121244 273434
rect 121278 273400 121312 273434
rect 121346 273400 121380 273434
rect 121414 273400 121448 273434
rect 121482 273400 121529 273434
rect 121129 273384 121529 273400
rect 120429 273278 120829 273294
rect 120429 273244 120476 273278
rect 120510 273244 120544 273278
rect 120578 273244 120612 273278
rect 120646 273244 120680 273278
rect 120714 273244 120748 273278
rect 120782 273244 120829 273278
rect 120429 273197 120829 273244
rect 121129 273278 121529 273294
rect 121129 273244 121176 273278
rect 121210 273244 121244 273278
rect 121278 273244 121312 273278
rect 121346 273244 121380 273278
rect 121414 273244 121448 273278
rect 121482 273244 121529 273278
rect 121129 273197 121529 273244
rect 120429 272650 120829 272697
rect 120429 272616 120476 272650
rect 120510 272616 120544 272650
rect 120578 272616 120612 272650
rect 120646 272616 120680 272650
rect 120714 272616 120748 272650
rect 120782 272616 120829 272650
rect 120429 272600 120829 272616
rect 121129 272650 121529 272697
rect 121129 272616 121176 272650
rect 121210 272616 121244 272650
rect 121278 272616 121312 272650
rect 121346 272616 121380 272650
rect 121414 272616 121448 272650
rect 121482 272616 121529 272650
rect 121129 272600 121529 272616
rect 120429 272494 120829 272510
rect 120429 272460 120476 272494
rect 120510 272460 120544 272494
rect 120578 272460 120612 272494
rect 120646 272460 120680 272494
rect 120714 272460 120748 272494
rect 120782 272460 120829 272494
rect 120429 272413 120829 272460
rect 121129 272494 121529 272510
rect 121129 272460 121176 272494
rect 121210 272460 121244 272494
rect 121278 272460 121312 272494
rect 121346 272460 121380 272494
rect 121414 272460 121448 272494
rect 121482 272460 121529 272494
rect 121129 272413 121529 272460
rect 120429 271866 120829 271913
rect 120429 271832 120476 271866
rect 120510 271832 120544 271866
rect 120578 271832 120612 271866
rect 120646 271832 120680 271866
rect 120714 271832 120748 271866
rect 120782 271832 120829 271866
rect 120429 271816 120829 271832
rect 121129 271866 121529 271913
rect 121129 271832 121176 271866
rect 121210 271832 121244 271866
rect 121278 271832 121312 271866
rect 121346 271832 121380 271866
rect 121414 271832 121448 271866
rect 121482 271832 121529 271866
rect 121129 271816 121529 271832
rect 120429 271710 120829 271726
rect 120429 271676 120476 271710
rect 120510 271676 120544 271710
rect 120578 271676 120612 271710
rect 120646 271676 120680 271710
rect 120714 271676 120748 271710
rect 120782 271676 120829 271710
rect 120429 271629 120829 271676
rect 121129 271710 121529 271726
rect 121129 271676 121176 271710
rect 121210 271676 121244 271710
rect 121278 271676 121312 271710
rect 121346 271676 121380 271710
rect 121414 271676 121448 271710
rect 121482 271676 121529 271710
rect 121129 271629 121529 271676
rect 120429 271082 120829 271129
rect 120429 271048 120476 271082
rect 120510 271048 120544 271082
rect 120578 271048 120612 271082
rect 120646 271048 120680 271082
rect 120714 271048 120748 271082
rect 120782 271048 120829 271082
rect 120429 271032 120829 271048
rect 121129 271082 121529 271129
rect 121129 271048 121176 271082
rect 121210 271048 121244 271082
rect 121278 271048 121312 271082
rect 121346 271048 121380 271082
rect 121414 271048 121448 271082
rect 121482 271048 121529 271082
rect 121129 271032 121529 271048
rect 120429 270926 120829 270942
rect 120429 270892 120476 270926
rect 120510 270892 120544 270926
rect 120578 270892 120612 270926
rect 120646 270892 120680 270926
rect 120714 270892 120748 270926
rect 120782 270892 120829 270926
rect 120429 270845 120829 270892
rect 121129 270926 121529 270942
rect 121129 270892 121176 270926
rect 121210 270892 121244 270926
rect 121278 270892 121312 270926
rect 121346 270892 121380 270926
rect 121414 270892 121448 270926
rect 121482 270892 121529 270926
rect 121129 270845 121529 270892
rect 120429 270298 120829 270345
rect 120429 270264 120476 270298
rect 120510 270264 120544 270298
rect 120578 270264 120612 270298
rect 120646 270264 120680 270298
rect 120714 270264 120748 270298
rect 120782 270264 120829 270298
rect 120429 270248 120829 270264
rect 121129 270298 121529 270345
rect 121129 270264 121176 270298
rect 121210 270264 121244 270298
rect 121278 270264 121312 270298
rect 121346 270264 121380 270298
rect 121414 270264 121448 270298
rect 121482 270264 121529 270298
rect 121129 270248 121529 270264
rect 120429 270142 120829 270158
rect 120429 270108 120476 270142
rect 120510 270108 120544 270142
rect 120578 270108 120612 270142
rect 120646 270108 120680 270142
rect 120714 270108 120748 270142
rect 120782 270108 120829 270142
rect 120429 270061 120829 270108
rect 121129 270142 121529 270158
rect 121129 270108 121176 270142
rect 121210 270108 121244 270142
rect 121278 270108 121312 270142
rect 121346 270108 121380 270142
rect 121414 270108 121448 270142
rect 121482 270108 121529 270142
rect 121129 270061 121529 270108
rect 120429 269514 120829 269561
rect 120429 269480 120476 269514
rect 120510 269480 120544 269514
rect 120578 269480 120612 269514
rect 120646 269480 120680 269514
rect 120714 269480 120748 269514
rect 120782 269480 120829 269514
rect 120429 269464 120829 269480
rect 121129 269514 121529 269561
rect 121129 269480 121176 269514
rect 121210 269480 121244 269514
rect 121278 269480 121312 269514
rect 121346 269480 121380 269514
rect 121414 269480 121448 269514
rect 121482 269480 121529 269514
rect 121129 269464 121529 269480
rect 120429 269358 120829 269374
rect 120429 269324 120476 269358
rect 120510 269324 120544 269358
rect 120578 269324 120612 269358
rect 120646 269324 120680 269358
rect 120714 269324 120748 269358
rect 120782 269324 120829 269358
rect 120429 269277 120829 269324
rect 121129 269358 121529 269374
rect 121129 269324 121176 269358
rect 121210 269324 121244 269358
rect 121278 269324 121312 269358
rect 121346 269324 121380 269358
rect 121414 269324 121448 269358
rect 121482 269324 121529 269358
rect 121129 269277 121529 269324
rect 120429 269130 120829 269177
rect 120429 269096 120476 269130
rect 120510 269096 120544 269130
rect 120578 269096 120612 269130
rect 120646 269096 120680 269130
rect 120714 269096 120748 269130
rect 120782 269096 120829 269130
rect 120429 269080 120829 269096
rect 121129 269130 121529 269177
rect 121129 269096 121176 269130
rect 121210 269096 121244 269130
rect 121278 269096 121312 269130
rect 121346 269096 121380 269130
rect 121414 269096 121448 269130
rect 121482 269096 121529 269130
rect 121129 269080 121529 269096
rect 122125 272894 122525 272910
rect 122125 272860 122172 272894
rect 122206 272860 122240 272894
rect 122274 272860 122308 272894
rect 122342 272860 122376 272894
rect 122410 272860 122444 272894
rect 122478 272860 122525 272894
rect 122125 272813 122525 272860
rect 122825 272894 123225 272910
rect 122825 272860 122872 272894
rect 122906 272860 122940 272894
rect 122974 272860 123008 272894
rect 123042 272860 123076 272894
rect 123110 272860 123144 272894
rect 123178 272860 123225 272894
rect 122825 272813 123225 272860
rect 122125 272666 122525 272713
rect 122125 272632 122172 272666
rect 122206 272632 122240 272666
rect 122274 272632 122308 272666
rect 122342 272632 122376 272666
rect 122410 272632 122444 272666
rect 122478 272632 122525 272666
rect 122125 272616 122525 272632
rect 122825 272666 123225 272713
rect 122825 272632 122872 272666
rect 122906 272632 122940 272666
rect 122974 272632 123008 272666
rect 123042 272632 123076 272666
rect 123110 272632 123144 272666
rect 123178 272632 123225 272666
rect 122825 272616 123225 272632
rect 122125 272510 122525 272526
rect 122125 272476 122172 272510
rect 122206 272476 122240 272510
rect 122274 272476 122308 272510
rect 122342 272476 122376 272510
rect 122410 272476 122444 272510
rect 122478 272476 122525 272510
rect 122125 272429 122525 272476
rect 122825 272510 123225 272526
rect 122825 272476 122872 272510
rect 122906 272476 122940 272510
rect 122974 272476 123008 272510
rect 123042 272476 123076 272510
rect 123110 272476 123144 272510
rect 123178 272476 123225 272510
rect 122825 272429 123225 272476
rect 122125 271882 122525 271929
rect 122125 271848 122172 271882
rect 122206 271848 122240 271882
rect 122274 271848 122308 271882
rect 122342 271848 122376 271882
rect 122410 271848 122444 271882
rect 122478 271848 122525 271882
rect 122125 271832 122525 271848
rect 122825 271882 123225 271929
rect 122825 271848 122872 271882
rect 122906 271848 122940 271882
rect 122974 271848 123008 271882
rect 123042 271848 123076 271882
rect 123110 271848 123144 271882
rect 123178 271848 123225 271882
rect 122825 271832 123225 271848
rect 122125 271726 122525 271742
rect 122125 271692 122172 271726
rect 122206 271692 122240 271726
rect 122274 271692 122308 271726
rect 122342 271692 122376 271726
rect 122410 271692 122444 271726
rect 122478 271692 122525 271726
rect 122125 271645 122525 271692
rect 122825 271726 123225 271742
rect 122825 271692 122872 271726
rect 122906 271692 122940 271726
rect 122974 271692 123008 271726
rect 123042 271692 123076 271726
rect 123110 271692 123144 271726
rect 123178 271692 123225 271726
rect 122825 271645 123225 271692
rect 122125 271098 122525 271145
rect 122125 271064 122172 271098
rect 122206 271064 122240 271098
rect 122274 271064 122308 271098
rect 122342 271064 122376 271098
rect 122410 271064 122444 271098
rect 122478 271064 122525 271098
rect 122125 271048 122525 271064
rect 122825 271098 123225 271145
rect 122825 271064 122872 271098
rect 122906 271064 122940 271098
rect 122974 271064 123008 271098
rect 123042 271064 123076 271098
rect 123110 271064 123144 271098
rect 123178 271064 123225 271098
rect 122825 271048 123225 271064
rect 122125 270942 122525 270958
rect 122125 270908 122172 270942
rect 122206 270908 122240 270942
rect 122274 270908 122308 270942
rect 122342 270908 122376 270942
rect 122410 270908 122444 270942
rect 122478 270908 122525 270942
rect 122125 270861 122525 270908
rect 122825 270942 123225 270958
rect 122825 270908 122872 270942
rect 122906 270908 122940 270942
rect 122974 270908 123008 270942
rect 123042 270908 123076 270942
rect 123110 270908 123144 270942
rect 123178 270908 123225 270942
rect 122825 270861 123225 270908
rect 122125 270314 122525 270361
rect 122125 270280 122172 270314
rect 122206 270280 122240 270314
rect 122274 270280 122308 270314
rect 122342 270280 122376 270314
rect 122410 270280 122444 270314
rect 122478 270280 122525 270314
rect 122125 270264 122525 270280
rect 122825 270314 123225 270361
rect 122825 270280 122872 270314
rect 122906 270280 122940 270314
rect 122974 270280 123008 270314
rect 123042 270280 123076 270314
rect 123110 270280 123144 270314
rect 123178 270280 123225 270314
rect 122825 270264 123225 270280
rect 122125 270158 122525 270174
rect 122125 270124 122172 270158
rect 122206 270124 122240 270158
rect 122274 270124 122308 270158
rect 122342 270124 122376 270158
rect 122410 270124 122444 270158
rect 122478 270124 122525 270158
rect 122125 270077 122525 270124
rect 122825 270158 123225 270174
rect 122825 270124 122872 270158
rect 122906 270124 122940 270158
rect 122974 270124 123008 270158
rect 123042 270124 123076 270158
rect 123110 270124 123144 270158
rect 123178 270124 123225 270158
rect 122825 270077 123225 270124
rect 122125 269530 122525 269577
rect 122125 269496 122172 269530
rect 122206 269496 122240 269530
rect 122274 269496 122308 269530
rect 122342 269496 122376 269530
rect 122410 269496 122444 269530
rect 122478 269496 122525 269530
rect 122125 269480 122525 269496
rect 122825 269530 123225 269577
rect 122825 269496 122872 269530
rect 122906 269496 122940 269530
rect 122974 269496 123008 269530
rect 123042 269496 123076 269530
rect 123110 269496 123144 269530
rect 123178 269496 123225 269530
rect 122825 269480 123225 269496
rect 122125 269374 122525 269390
rect 122125 269340 122172 269374
rect 122206 269340 122240 269374
rect 122274 269340 122308 269374
rect 122342 269340 122376 269374
rect 122410 269340 122444 269374
rect 122478 269340 122525 269374
rect 122125 269293 122525 269340
rect 122825 269374 123225 269390
rect 122825 269340 122872 269374
rect 122906 269340 122940 269374
rect 122974 269340 123008 269374
rect 123042 269340 123076 269374
rect 123110 269340 123144 269374
rect 123178 269340 123225 269374
rect 122825 269293 123225 269340
rect 122125 269146 122525 269193
rect 122125 269112 122172 269146
rect 122206 269112 122240 269146
rect 122274 269112 122308 269146
rect 122342 269112 122376 269146
rect 122410 269112 122444 269146
rect 122478 269112 122525 269146
rect 122125 269096 122525 269112
rect 122825 269146 123225 269193
rect 122825 269112 122872 269146
rect 122906 269112 122940 269146
rect 122974 269112 123008 269146
rect 123042 269112 123076 269146
rect 123110 269112 123144 269146
rect 123178 269112 123225 269146
rect 122825 269096 123225 269112
rect 124104 272471 124192 272520
rect 124104 272437 124120 272471
rect 124154 272437 124192 272471
rect 124104 272403 124192 272437
rect 124104 272369 124120 272403
rect 124154 272369 124192 272403
rect 124104 272320 124192 272369
rect 124692 272471 124780 272520
rect 124692 272437 124730 272471
rect 124764 272437 124780 272471
rect 124692 272403 124780 272437
rect 124692 272369 124730 272403
rect 124764 272369 124780 272403
rect 124692 272320 124780 272369
rect 124104 272055 124192 272104
rect 124104 272021 124120 272055
rect 124154 272021 124192 272055
rect 124104 271987 124192 272021
rect 124104 271953 124120 271987
rect 124154 271953 124192 271987
rect 124104 271904 124192 271953
rect 124692 272055 124780 272104
rect 124692 272021 124730 272055
rect 124764 272021 124780 272055
rect 124692 271987 124780 272021
rect 124692 271953 124730 271987
rect 124764 271953 124780 271987
rect 124692 271904 124780 271953
rect 124104 271639 124192 271688
rect 124104 271605 124120 271639
rect 124154 271605 124192 271639
rect 124104 271571 124192 271605
rect 124104 271537 124120 271571
rect 124154 271537 124192 271571
rect 124104 271488 124192 271537
rect 124692 271639 124780 271688
rect 124692 271605 124730 271639
rect 124764 271605 124780 271639
rect 124692 271571 124780 271605
rect 124692 271537 124730 271571
rect 124764 271537 124780 271571
rect 124692 271488 124780 271537
rect 124104 271223 124192 271272
rect 124104 271189 124120 271223
rect 124154 271189 124192 271223
rect 124104 271155 124192 271189
rect 124104 271121 124120 271155
rect 124154 271121 124192 271155
rect 124104 271072 124192 271121
rect 124692 271223 124780 271272
rect 124692 271189 124730 271223
rect 124764 271189 124780 271223
rect 124692 271155 124780 271189
rect 124692 271121 124730 271155
rect 124764 271121 124780 271155
rect 124692 271072 124780 271121
rect 124104 270807 124192 270856
rect 124104 270773 124120 270807
rect 124154 270773 124192 270807
rect 124104 270739 124192 270773
rect 124104 270705 124120 270739
rect 124154 270705 124192 270739
rect 124104 270656 124192 270705
rect 124692 270807 124780 270856
rect 124692 270773 124730 270807
rect 124764 270773 124780 270807
rect 124692 270739 124780 270773
rect 124692 270705 124730 270739
rect 124764 270705 124780 270739
rect 124692 270656 124780 270705
rect 124104 270391 124192 270440
rect 124104 270357 124120 270391
rect 124154 270357 124192 270391
rect 124104 270323 124192 270357
rect 124104 270289 124120 270323
rect 124154 270289 124192 270323
rect 124104 270240 124192 270289
rect 124692 270391 124780 270440
rect 124692 270357 124730 270391
rect 124764 270357 124780 270391
rect 124692 270323 124780 270357
rect 124692 270289 124730 270323
rect 124764 270289 124780 270323
rect 124692 270240 124780 270289
rect 124104 269975 124192 270024
rect 124104 269941 124120 269975
rect 124154 269941 124192 269975
rect 124104 269907 124192 269941
rect 124104 269873 124120 269907
rect 124154 269873 124192 269907
rect 124104 269824 124192 269873
rect 124692 269975 124780 270024
rect 124692 269941 124730 269975
rect 124764 269941 124780 269975
rect 124692 269907 124780 269941
rect 124692 269873 124730 269907
rect 124764 269873 124780 269907
rect 124692 269824 124780 269873
rect 124104 269559 124192 269608
rect 124104 269525 124120 269559
rect 124154 269525 124192 269559
rect 124104 269491 124192 269525
rect 124104 269457 124120 269491
rect 124154 269457 124192 269491
rect 124104 269408 124192 269457
rect 124692 269559 124780 269608
rect 124692 269525 124730 269559
rect 124764 269525 124780 269559
rect 124692 269491 124780 269525
rect 124692 269457 124730 269491
rect 124764 269457 124780 269491
rect 124692 269408 124780 269457
<< polycont >>
rect 106406 280851 106440 280885
rect 106806 280851 106840 280885
rect 107206 280851 107240 280885
rect 107606 280851 107640 280885
rect 108006 280851 108040 280885
rect 108406 280851 108440 280885
rect 108806 280851 108840 280885
rect 109206 280851 109240 280885
rect 109606 280851 109640 280885
rect 110006 280851 110040 280885
rect 106406 279721 106440 279755
rect 106806 279721 106840 279755
rect 107206 279721 107240 279755
rect 107606 279721 107640 279755
rect 108006 279721 108040 279755
rect 108406 279721 108440 279755
rect 108806 279721 108840 279755
rect 109206 279721 109240 279755
rect 109606 279721 109640 279755
rect 110006 279721 110040 279755
rect 106287 278935 106321 278969
rect 106287 278867 106321 278901
rect 106287 278799 106321 278833
rect 107629 278935 107663 278969
rect 107629 278867 107663 278901
rect 107629 278799 107663 278833
rect 106287 278335 106321 278369
rect 106287 278267 106321 278301
rect 106287 278199 106321 278233
rect 107629 278335 107663 278369
rect 107629 278267 107663 278301
rect 107629 278199 107663 278233
rect 109801 279049 109835 279083
rect 109869 279049 109903 279083
rect 109937 279049 109971 279083
rect 110005 279049 110039 279083
rect 109801 277901 109835 277935
rect 109869 277901 109903 277935
rect 109937 277901 109971 277935
rect 110005 277901 110039 277935
rect 109801 277793 109835 277827
rect 109869 277793 109903 277827
rect 109937 277793 109971 277827
rect 110005 277793 110039 277827
rect 106410 277110 106444 277144
rect 107572 277110 107606 277144
rect 109801 276645 109835 276679
rect 109869 276645 109903 276679
rect 109937 276645 109971 276679
rect 110005 276645 110039 276679
rect 106870 275647 106904 275681
rect 106870 275579 106904 275613
rect 106870 275511 106904 275545
rect 106870 275443 106904 275477
rect 106870 275375 106904 275409
rect 106870 275307 106904 275341
rect 106870 275239 106904 275273
rect 106870 275171 106904 275205
rect 106870 275103 106904 275137
rect 106870 275035 106904 275069
rect 106870 274967 106904 275001
rect 107176 275647 107210 275681
rect 107176 275579 107210 275613
rect 107176 275511 107210 275545
rect 107176 275443 107210 275477
rect 107176 275375 107210 275409
rect 107176 275307 107210 275341
rect 107176 275239 107210 275273
rect 107176 275171 107210 275205
rect 107176 275103 107210 275137
rect 107176 275035 107210 275069
rect 107176 274967 107210 275001
rect 107370 275647 107404 275681
rect 107370 275579 107404 275613
rect 107370 275511 107404 275545
rect 107370 275443 107404 275477
rect 107370 275375 107404 275409
rect 107370 275307 107404 275341
rect 107370 275239 107404 275273
rect 107370 275171 107404 275205
rect 107370 275103 107404 275137
rect 107370 275035 107404 275069
rect 107370 274967 107404 275001
rect 107676 275647 107710 275681
rect 107676 275579 107710 275613
rect 107676 275511 107710 275545
rect 107676 275443 107710 275477
rect 107676 275375 107710 275409
rect 107676 275307 107710 275341
rect 107676 275239 107710 275273
rect 107676 275171 107710 275205
rect 107676 275103 107710 275137
rect 107676 275035 107710 275069
rect 107676 274967 107710 275001
rect 107870 275647 107904 275681
rect 107870 275579 107904 275613
rect 107870 275511 107904 275545
rect 107870 275443 107904 275477
rect 107870 275375 107904 275409
rect 107870 275307 107904 275341
rect 107870 275239 107904 275273
rect 107870 275171 107904 275205
rect 107870 275103 107904 275137
rect 107870 275035 107904 275069
rect 107870 274967 107904 275001
rect 108176 275647 108210 275681
rect 108176 275579 108210 275613
rect 108176 275511 108210 275545
rect 108176 275443 108210 275477
rect 108176 275375 108210 275409
rect 108176 275307 108210 275341
rect 108176 275239 108210 275273
rect 108176 275171 108210 275205
rect 108176 275103 108210 275137
rect 108176 275035 108210 275069
rect 108176 274967 108210 275001
rect 108370 275647 108404 275681
rect 108370 275579 108404 275613
rect 108370 275511 108404 275545
rect 108370 275443 108404 275477
rect 108370 275375 108404 275409
rect 108370 275307 108404 275341
rect 108370 275239 108404 275273
rect 108370 275171 108404 275205
rect 108370 275103 108404 275137
rect 108370 275035 108404 275069
rect 108370 274967 108404 275001
rect 108676 275647 108710 275681
rect 108676 275579 108710 275613
rect 108676 275511 108710 275545
rect 108676 275443 108710 275477
rect 108676 275375 108710 275409
rect 108676 275307 108710 275341
rect 108676 275239 108710 275273
rect 108676 275171 108710 275205
rect 108676 275103 108710 275137
rect 108676 275035 108710 275069
rect 108676 274967 108710 275001
rect 108870 275647 108904 275681
rect 108870 275579 108904 275613
rect 108870 275511 108904 275545
rect 108870 275443 108904 275477
rect 108870 275375 108904 275409
rect 108870 275307 108904 275341
rect 108870 275239 108904 275273
rect 108870 275171 108904 275205
rect 108870 275103 108904 275137
rect 108870 275035 108904 275069
rect 108870 274967 108904 275001
rect 109176 275647 109210 275681
rect 109176 275579 109210 275613
rect 109176 275511 109210 275545
rect 109176 275443 109210 275477
rect 109176 275375 109210 275409
rect 109176 275307 109210 275341
rect 109176 275239 109210 275273
rect 109176 275171 109210 275205
rect 109176 275103 109210 275137
rect 109176 275035 109210 275069
rect 109176 274967 109210 275001
rect 109370 275647 109404 275681
rect 109370 275579 109404 275613
rect 109370 275511 109404 275545
rect 109370 275443 109404 275477
rect 109370 275375 109404 275409
rect 109370 275307 109404 275341
rect 109370 275239 109404 275273
rect 109370 275171 109404 275205
rect 109370 275103 109404 275137
rect 109370 275035 109404 275069
rect 109370 274967 109404 275001
rect 109676 275647 109710 275681
rect 109676 275579 109710 275613
rect 109676 275511 109710 275545
rect 109676 275443 109710 275477
rect 109676 275375 109710 275409
rect 109676 275307 109710 275341
rect 109676 275239 109710 275273
rect 109676 275171 109710 275205
rect 109676 275103 109710 275137
rect 109676 275035 109710 275069
rect 109676 274967 109710 275001
rect 109458 272473 109492 272507
rect 107480 272117 107514 272151
rect 107548 272117 107582 272151
rect 107616 272117 107650 272151
rect 107684 272117 107718 272151
rect 107752 272117 107786 272151
rect 107820 272117 107854 272151
rect 107888 272117 107922 272151
rect 107956 272117 107990 272151
rect 108024 272117 108058 272151
rect 107001 272009 107035 272043
rect 107069 272009 107103 272043
rect 107137 272009 107171 272043
rect 107001 271735 107035 271769
rect 107069 271735 107103 271769
rect 107137 271735 107171 271769
rect 107480 271663 107514 271697
rect 107548 271663 107582 271697
rect 107616 271663 107650 271697
rect 107684 271663 107718 271697
rect 107752 271663 107786 271697
rect 107820 271663 107854 271697
rect 107888 271663 107922 271697
rect 107956 271663 107990 271697
rect 108024 271663 108058 271697
rect 107101 271417 107135 271451
rect 107101 271349 107135 271383
rect 108411 271417 108445 271451
rect 108411 271349 108445 271383
rect 107101 271047 107135 271081
rect 107101 270979 107135 271013
rect 108411 271047 108445 271081
rect 108411 270979 108445 271013
rect 109458 270625 109492 270659
rect 111452 280757 111486 280791
rect 111452 280689 111486 280723
rect 112662 280757 112696 280791
rect 112662 280689 112696 280723
rect 112898 280745 112932 280779
rect 112898 280677 112932 280711
rect 114108 280745 114142 280779
rect 114108 280677 114142 280711
rect 111452 280397 111486 280431
rect 111452 280329 111486 280363
rect 112662 280397 112696 280431
rect 112662 280329 112696 280363
rect 112898 280321 112932 280355
rect 112898 280253 112932 280287
rect 114108 280321 114142 280355
rect 114108 280253 114142 280287
rect 114576 280722 114610 280756
rect 114576 280654 114610 280688
rect 114576 280586 114610 280620
rect 114576 280518 114610 280552
rect 114576 280450 114610 280484
rect 114904 280722 114938 280756
rect 114904 280654 114938 280688
rect 114904 280586 114938 280620
rect 114904 280518 114938 280552
rect 114904 280450 114938 280484
rect 111452 280037 111486 280071
rect 111452 279969 111486 280003
rect 112662 280037 112696 280071
rect 112662 279969 112696 280003
rect 112928 279945 112962 279979
rect 114138 279945 114172 279979
rect 114576 280054 114610 280088
rect 114576 279986 114610 280020
rect 114904 280054 114938 280088
rect 114904 279986 114938 280020
rect 111452 279677 111486 279711
rect 111452 279609 111486 279643
rect 112662 279677 112696 279711
rect 112662 279609 112696 279643
rect 112928 279647 112962 279681
rect 114138 279647 114172 279681
rect 114576 279646 114610 279680
rect 114576 279578 114610 279612
rect 114904 279646 114938 279680
rect 114904 279578 114938 279612
rect 115267 280722 115301 280756
rect 115267 280654 115301 280688
rect 115267 280586 115301 280620
rect 115267 280518 115301 280552
rect 115267 280450 115301 280484
rect 115595 280722 115629 280756
rect 115595 280654 115629 280688
rect 115595 280586 115629 280620
rect 115595 280518 115629 280552
rect 115595 280450 115629 280484
rect 116063 280745 116097 280779
rect 116063 280677 116097 280711
rect 117273 280745 117307 280779
rect 117273 280677 117307 280711
rect 117509 280757 117543 280791
rect 117509 280689 117543 280723
rect 118719 280757 118753 280791
rect 118719 280689 118753 280723
rect 116063 280321 116097 280355
rect 116063 280253 116097 280287
rect 117273 280321 117307 280355
rect 117509 280397 117543 280431
rect 117509 280329 117543 280363
rect 118719 280397 118753 280431
rect 118719 280329 118753 280363
rect 117273 280253 117307 280287
rect 115267 280054 115301 280088
rect 115267 279986 115301 280020
rect 115595 280054 115629 280088
rect 115595 279986 115629 280020
rect 117509 280037 117543 280071
rect 116033 279945 116067 279979
rect 117243 279945 117277 279979
rect 117509 279969 117543 280003
rect 118719 280037 118753 280071
rect 118719 279969 118753 280003
rect 115267 279646 115301 279680
rect 115267 279578 115301 279612
rect 115595 279646 115629 279680
rect 115595 279578 115629 279612
rect 116033 279647 116067 279681
rect 117243 279647 117277 279681
rect 117509 279677 117543 279711
rect 117509 279609 117543 279643
rect 118719 279677 118753 279711
rect 118719 279609 118753 279643
rect 111452 279091 111486 279125
rect 111452 279023 111486 279057
rect 112662 279091 112696 279125
rect 112662 279023 112696 279057
rect 112898 279079 112932 279113
rect 112898 279011 112932 279045
rect 114108 279079 114142 279113
rect 114108 279011 114142 279045
rect 111452 278731 111486 278765
rect 111452 278663 111486 278697
rect 112662 278731 112696 278765
rect 112662 278663 112696 278697
rect 112898 278655 112932 278689
rect 112898 278587 112932 278621
rect 114108 278655 114142 278689
rect 114108 278587 114142 278621
rect 114576 279056 114610 279090
rect 114576 278988 114610 279022
rect 114576 278920 114610 278954
rect 114576 278852 114610 278886
rect 114576 278784 114610 278818
rect 114904 279056 114938 279090
rect 114904 278988 114938 279022
rect 114904 278920 114938 278954
rect 114904 278852 114938 278886
rect 114904 278784 114938 278818
rect 111452 278371 111486 278405
rect 111452 278303 111486 278337
rect 112662 278371 112696 278405
rect 112662 278303 112696 278337
rect 112928 278279 112962 278313
rect 114138 278279 114172 278313
rect 114576 278388 114610 278422
rect 114576 278320 114610 278354
rect 114904 278388 114938 278422
rect 114904 278320 114938 278354
rect 111452 278011 111486 278045
rect 111452 277943 111486 277977
rect 112662 278011 112696 278045
rect 112662 277943 112696 277977
rect 112928 277981 112962 278015
rect 114138 277981 114172 278015
rect 114576 277980 114610 278014
rect 114576 277912 114610 277946
rect 114904 277980 114938 278014
rect 114904 277912 114938 277946
rect 115267 279056 115301 279090
rect 115267 278988 115301 279022
rect 115267 278920 115301 278954
rect 115267 278852 115301 278886
rect 115267 278784 115301 278818
rect 115595 279056 115629 279090
rect 115595 278988 115629 279022
rect 115595 278920 115629 278954
rect 115595 278852 115629 278886
rect 115595 278784 115629 278818
rect 116063 279079 116097 279113
rect 116063 279011 116097 279045
rect 117273 279079 117307 279113
rect 117273 279011 117307 279045
rect 117509 279091 117543 279125
rect 117509 279023 117543 279057
rect 118719 279091 118753 279125
rect 118719 279023 118753 279057
rect 116063 278655 116097 278689
rect 116063 278587 116097 278621
rect 117273 278655 117307 278689
rect 117509 278731 117543 278765
rect 117509 278663 117543 278697
rect 118719 278731 118753 278765
rect 118719 278663 118753 278697
rect 117273 278587 117307 278621
rect 115267 278388 115301 278422
rect 115267 278320 115301 278354
rect 115595 278388 115629 278422
rect 115595 278320 115629 278354
rect 117509 278371 117543 278405
rect 116033 278279 116067 278313
rect 117243 278279 117277 278313
rect 117509 278303 117543 278337
rect 118719 278371 118753 278405
rect 118719 278303 118753 278337
rect 115267 277980 115301 278014
rect 115267 277912 115301 277946
rect 115595 277980 115629 278014
rect 115595 277912 115629 277946
rect 116033 277981 116067 278015
rect 117243 277981 117277 278015
rect 117509 278011 117543 278045
rect 117509 277943 117543 277977
rect 118719 278011 118753 278045
rect 118719 277943 118753 277977
rect 111452 277425 111486 277459
rect 111452 277357 111486 277391
rect 112662 277425 112696 277459
rect 112662 277357 112696 277391
rect 112898 277413 112932 277447
rect 112898 277345 112932 277379
rect 114108 277413 114142 277447
rect 114108 277345 114142 277379
rect 111452 277065 111486 277099
rect 111452 276997 111486 277031
rect 112662 277065 112696 277099
rect 112662 276997 112696 277031
rect 112898 276989 112932 277023
rect 112898 276921 112932 276955
rect 114108 276989 114142 277023
rect 114108 276921 114142 276955
rect 114576 277390 114610 277424
rect 114576 277322 114610 277356
rect 114576 277254 114610 277288
rect 114576 277186 114610 277220
rect 114576 277118 114610 277152
rect 114904 277390 114938 277424
rect 114904 277322 114938 277356
rect 114904 277254 114938 277288
rect 114904 277186 114938 277220
rect 114904 277118 114938 277152
rect 111452 276705 111486 276739
rect 111452 276637 111486 276671
rect 112662 276705 112696 276739
rect 112662 276637 112696 276671
rect 112928 276613 112962 276647
rect 114138 276613 114172 276647
rect 114576 276722 114610 276756
rect 114576 276654 114610 276688
rect 114904 276722 114938 276756
rect 114904 276654 114938 276688
rect 111452 276345 111486 276379
rect 111452 276277 111486 276311
rect 112662 276345 112696 276379
rect 112662 276277 112696 276311
rect 112928 276315 112962 276349
rect 114138 276315 114172 276349
rect 114576 276314 114610 276348
rect 114576 276246 114610 276280
rect 114904 276314 114938 276348
rect 114904 276246 114938 276280
rect 115267 277390 115301 277424
rect 115267 277322 115301 277356
rect 115267 277254 115301 277288
rect 115267 277186 115301 277220
rect 115267 277118 115301 277152
rect 115595 277390 115629 277424
rect 115595 277322 115629 277356
rect 115595 277254 115629 277288
rect 115595 277186 115629 277220
rect 115595 277118 115629 277152
rect 116063 277413 116097 277447
rect 116063 277345 116097 277379
rect 117273 277413 117307 277447
rect 117273 277345 117307 277379
rect 117509 277425 117543 277459
rect 117509 277357 117543 277391
rect 118719 277425 118753 277459
rect 118719 277357 118753 277391
rect 116063 276989 116097 277023
rect 116063 276921 116097 276955
rect 117273 276989 117307 277023
rect 117509 277065 117543 277099
rect 117509 276997 117543 277031
rect 118719 277065 118753 277099
rect 118719 276997 118753 277031
rect 117273 276921 117307 276955
rect 115267 276722 115301 276756
rect 115267 276654 115301 276688
rect 115595 276722 115629 276756
rect 115595 276654 115629 276688
rect 117509 276705 117543 276739
rect 116033 276613 116067 276647
rect 117243 276613 117277 276647
rect 117509 276637 117543 276671
rect 118719 276705 118753 276739
rect 118719 276637 118753 276671
rect 115267 276314 115301 276348
rect 115267 276246 115301 276280
rect 115595 276314 115629 276348
rect 115595 276246 115629 276280
rect 116033 276315 116067 276349
rect 117243 276315 117277 276349
rect 117509 276345 117543 276379
rect 117509 276277 117543 276311
rect 118719 276345 118753 276379
rect 118719 276277 118753 276311
rect 111452 275759 111486 275793
rect 111452 275691 111486 275725
rect 112662 275759 112696 275793
rect 112662 275691 112696 275725
rect 112898 275747 112932 275781
rect 112898 275679 112932 275713
rect 114108 275747 114142 275781
rect 114108 275679 114142 275713
rect 111452 275399 111486 275433
rect 111452 275331 111486 275365
rect 112662 275399 112696 275433
rect 112662 275331 112696 275365
rect 112898 275323 112932 275357
rect 112898 275255 112932 275289
rect 114108 275323 114142 275357
rect 114108 275255 114142 275289
rect 114576 275724 114610 275758
rect 114576 275656 114610 275690
rect 114576 275588 114610 275622
rect 114576 275520 114610 275554
rect 114576 275452 114610 275486
rect 114904 275724 114938 275758
rect 114904 275656 114938 275690
rect 114904 275588 114938 275622
rect 114904 275520 114938 275554
rect 114904 275452 114938 275486
rect 111452 275039 111486 275073
rect 111452 274971 111486 275005
rect 112662 275039 112696 275073
rect 112662 274971 112696 275005
rect 112928 274947 112962 274981
rect 114138 274947 114172 274981
rect 114576 275056 114610 275090
rect 114576 274988 114610 275022
rect 114904 275056 114938 275090
rect 114904 274988 114938 275022
rect 111452 274679 111486 274713
rect 111452 274611 111486 274645
rect 112662 274679 112696 274713
rect 112662 274611 112696 274645
rect 112928 274649 112962 274683
rect 114138 274649 114172 274683
rect 114576 274648 114610 274682
rect 114576 274580 114610 274614
rect 114904 274648 114938 274682
rect 114904 274580 114938 274614
rect 115267 275724 115301 275758
rect 115267 275656 115301 275690
rect 115267 275588 115301 275622
rect 115267 275520 115301 275554
rect 115267 275452 115301 275486
rect 115595 275724 115629 275758
rect 115595 275656 115629 275690
rect 115595 275588 115629 275622
rect 115595 275520 115629 275554
rect 115595 275452 115629 275486
rect 116063 275747 116097 275781
rect 116063 275679 116097 275713
rect 117273 275747 117307 275781
rect 117273 275679 117307 275713
rect 117509 275759 117543 275793
rect 117509 275691 117543 275725
rect 118719 275759 118753 275793
rect 118719 275691 118753 275725
rect 116063 275323 116097 275357
rect 116063 275255 116097 275289
rect 117273 275323 117307 275357
rect 117509 275399 117543 275433
rect 117509 275331 117543 275365
rect 118719 275399 118753 275433
rect 118719 275331 118753 275365
rect 117273 275255 117307 275289
rect 115267 275056 115301 275090
rect 115267 274988 115301 275022
rect 115595 275056 115629 275090
rect 115595 274988 115629 275022
rect 117509 275039 117543 275073
rect 116033 274947 116067 274981
rect 117243 274947 117277 274981
rect 117509 274971 117543 275005
rect 118719 275039 118753 275073
rect 118719 274971 118753 275005
rect 115267 274648 115301 274682
rect 115267 274580 115301 274614
rect 115595 274648 115629 274682
rect 115595 274580 115629 274614
rect 116033 274649 116067 274683
rect 117243 274649 117277 274683
rect 117509 274679 117543 274713
rect 117509 274611 117543 274645
rect 118719 274679 118753 274713
rect 118719 274611 118753 274645
rect 111452 274093 111486 274127
rect 111452 274025 111486 274059
rect 112662 274093 112696 274127
rect 112662 274025 112696 274059
rect 112898 274081 112932 274115
rect 112898 274013 112932 274047
rect 114108 274081 114142 274115
rect 114108 274013 114142 274047
rect 111452 273733 111486 273767
rect 111452 273665 111486 273699
rect 112662 273733 112696 273767
rect 112662 273665 112696 273699
rect 112898 273657 112932 273691
rect 112898 273589 112932 273623
rect 114108 273657 114142 273691
rect 114108 273589 114142 273623
rect 114576 274058 114610 274092
rect 114576 273990 114610 274024
rect 114576 273922 114610 273956
rect 114576 273854 114610 273888
rect 114576 273786 114610 273820
rect 114904 274058 114938 274092
rect 114904 273990 114938 274024
rect 114904 273922 114938 273956
rect 114904 273854 114938 273888
rect 114904 273786 114938 273820
rect 111452 273373 111486 273407
rect 111452 273305 111486 273339
rect 112662 273373 112696 273407
rect 112662 273305 112696 273339
rect 112928 273281 112962 273315
rect 114138 273281 114172 273315
rect 114576 273390 114610 273424
rect 114576 273322 114610 273356
rect 114904 273390 114938 273424
rect 114904 273322 114938 273356
rect 111452 273013 111486 273047
rect 111452 272945 111486 272979
rect 112662 273013 112696 273047
rect 112662 272945 112696 272979
rect 112928 272983 112962 273017
rect 114138 272983 114172 273017
rect 114576 272982 114610 273016
rect 114576 272914 114610 272948
rect 114904 272982 114938 273016
rect 114904 272914 114938 272948
rect 115267 274058 115301 274092
rect 115267 273990 115301 274024
rect 115267 273922 115301 273956
rect 115267 273854 115301 273888
rect 115267 273786 115301 273820
rect 115595 274058 115629 274092
rect 115595 273990 115629 274024
rect 115595 273922 115629 273956
rect 115595 273854 115629 273888
rect 115595 273786 115629 273820
rect 116063 274081 116097 274115
rect 116063 274013 116097 274047
rect 117273 274081 117307 274115
rect 117273 274013 117307 274047
rect 117509 274093 117543 274127
rect 117509 274025 117543 274059
rect 118719 274093 118753 274127
rect 118719 274025 118753 274059
rect 116063 273657 116097 273691
rect 116063 273589 116097 273623
rect 117273 273657 117307 273691
rect 117509 273733 117543 273767
rect 117509 273665 117543 273699
rect 118719 273733 118753 273767
rect 118719 273665 118753 273699
rect 117273 273589 117307 273623
rect 115267 273390 115301 273424
rect 115267 273322 115301 273356
rect 115595 273390 115629 273424
rect 115595 273322 115629 273356
rect 117509 273373 117543 273407
rect 116033 273281 116067 273315
rect 117243 273281 117277 273315
rect 117509 273305 117543 273339
rect 118719 273373 118753 273407
rect 118719 273305 118753 273339
rect 115267 272982 115301 273016
rect 115267 272914 115301 272948
rect 115595 272982 115629 273016
rect 115595 272914 115629 272948
rect 116033 272983 116067 273017
rect 117243 272983 117277 273017
rect 117509 273013 117543 273047
rect 117509 272945 117543 272979
rect 118719 273013 118753 273047
rect 118719 272945 118753 272979
rect 115910 271962 115944 271996
rect 115978 271962 116012 271996
rect 116310 271962 116344 271996
rect 116378 271962 116412 271996
rect 116710 271962 116744 271996
rect 116778 271962 116812 271996
rect 117110 271962 117144 271996
rect 117178 271962 117212 271996
rect 117510 271962 117544 271996
rect 117578 271962 117612 271996
rect 117910 271962 117944 271996
rect 117978 271962 118012 271996
rect 118310 271962 118344 271996
rect 118378 271962 118412 271996
rect 118710 271962 118744 271996
rect 118778 271962 118812 271996
rect 112607 271353 112641 271387
rect 112675 271353 112709 271387
rect 113007 271353 113041 271387
rect 113075 271353 113109 271387
rect 113407 271353 113441 271387
rect 113475 271353 113509 271387
rect 113807 271353 113841 271387
rect 113875 271353 113909 271387
rect 112607 271025 112641 271059
rect 112675 271025 112709 271059
rect 113007 271025 113041 271059
rect 113075 271025 113109 271059
rect 113407 271025 113441 271059
rect 113475 271025 113509 271059
rect 113807 271025 113841 271059
rect 113875 271025 113909 271059
rect 114666 271324 114700 271358
rect 114734 271324 114768 271358
rect 115066 271324 115100 271358
rect 115134 271324 115168 271358
rect 114666 270996 114700 271030
rect 114734 270996 114768 271030
rect 115066 270996 115100 271030
rect 115134 270996 115168 271030
rect 115910 270752 115944 270786
rect 115978 270752 116012 270786
rect 116310 270752 116344 270786
rect 116378 270752 116412 270786
rect 116710 270752 116744 270786
rect 116778 270752 116812 270786
rect 117110 270752 117144 270786
rect 117178 270752 117212 270786
rect 117510 270752 117544 270786
rect 117578 270752 117612 270786
rect 117910 270752 117944 270786
rect 117978 270752 118012 270786
rect 118310 270752 118344 270786
rect 118378 270752 118412 270786
rect 118710 270752 118744 270786
rect 118778 270752 118812 270786
rect 112589 270262 112623 270296
rect 112657 270262 112691 270296
rect 112989 270262 113023 270296
rect 113057 270262 113091 270296
rect 113389 270262 113423 270296
rect 113457 270262 113491 270296
rect 113789 270262 113823 270296
rect 113857 270262 113891 270296
rect 114189 270262 114223 270296
rect 114257 270262 114291 270296
rect 114589 270262 114623 270296
rect 114657 270262 114691 270296
rect 114989 270262 115023 270296
rect 115057 270262 115091 270296
rect 115389 270262 115423 270296
rect 115457 270262 115491 270296
rect 115789 270262 115823 270296
rect 115857 270262 115891 270296
rect 116189 270262 116223 270296
rect 116257 270262 116291 270296
rect 116589 270262 116623 270296
rect 116657 270262 116691 270296
rect 116989 270262 117023 270296
rect 117057 270262 117091 270296
rect 117389 270262 117423 270296
rect 117457 270262 117491 270296
rect 117789 270262 117823 270296
rect 117857 270262 117891 270296
rect 118189 270262 118223 270296
rect 118257 270262 118291 270296
rect 118589 270262 118623 270296
rect 118657 270262 118691 270296
rect 112589 269052 112623 269086
rect 112657 269052 112691 269086
rect 112989 269052 113023 269086
rect 113057 269052 113091 269086
rect 113389 269052 113423 269086
rect 113457 269052 113491 269086
rect 113789 269052 113823 269086
rect 113857 269052 113891 269086
rect 114189 269052 114223 269086
rect 114257 269052 114291 269086
rect 114589 269052 114623 269086
rect 114657 269052 114691 269086
rect 114989 269052 115023 269086
rect 115057 269052 115091 269086
rect 115389 269052 115423 269086
rect 115457 269052 115491 269086
rect 115789 269052 115823 269086
rect 115857 269052 115891 269086
rect 116189 269052 116223 269086
rect 116257 269052 116291 269086
rect 116589 269052 116623 269086
rect 116657 269052 116691 269086
rect 116989 269052 117023 269086
rect 117057 269052 117091 269086
rect 117389 269052 117423 269086
rect 117457 269052 117491 269086
rect 117789 269052 117823 269086
rect 117857 269052 117891 269086
rect 118189 269052 118223 269086
rect 118257 269052 118291 269086
rect 118589 269052 118623 269086
rect 118657 269052 118691 269086
rect 120476 280684 120510 280718
rect 120544 280684 120578 280718
rect 120612 280684 120646 280718
rect 120680 280684 120714 280718
rect 120748 280684 120782 280718
rect 121176 280684 121210 280718
rect 121244 280684 121278 280718
rect 121312 280684 121346 280718
rect 121380 280684 121414 280718
rect 121448 280684 121482 280718
rect 120476 280456 120510 280490
rect 120544 280456 120578 280490
rect 120612 280456 120646 280490
rect 120680 280456 120714 280490
rect 120748 280456 120782 280490
rect 121176 280456 121210 280490
rect 121244 280456 121278 280490
rect 121312 280456 121346 280490
rect 121380 280456 121414 280490
rect 121448 280456 121482 280490
rect 120476 280300 120510 280334
rect 120544 280300 120578 280334
rect 120612 280300 120646 280334
rect 120680 280300 120714 280334
rect 120748 280300 120782 280334
rect 121176 280300 121210 280334
rect 121244 280300 121278 280334
rect 121312 280300 121346 280334
rect 121380 280300 121414 280334
rect 121448 280300 121482 280334
rect 120476 279672 120510 279706
rect 120544 279672 120578 279706
rect 120612 279672 120646 279706
rect 120680 279672 120714 279706
rect 120748 279672 120782 279706
rect 121176 279672 121210 279706
rect 121244 279672 121278 279706
rect 121312 279672 121346 279706
rect 121380 279672 121414 279706
rect 121448 279672 121482 279706
rect 120476 279516 120510 279550
rect 120544 279516 120578 279550
rect 120612 279516 120646 279550
rect 120680 279516 120714 279550
rect 120748 279516 120782 279550
rect 121176 279516 121210 279550
rect 121244 279516 121278 279550
rect 121312 279516 121346 279550
rect 121380 279516 121414 279550
rect 121448 279516 121482 279550
rect 120476 278888 120510 278922
rect 120544 278888 120578 278922
rect 120612 278888 120646 278922
rect 120680 278888 120714 278922
rect 120748 278888 120782 278922
rect 121176 278888 121210 278922
rect 121244 278888 121278 278922
rect 121312 278888 121346 278922
rect 121380 278888 121414 278922
rect 121448 278888 121482 278922
rect 122403 280470 122437 280504
rect 122471 280470 122505 280504
rect 122539 280470 122573 280504
rect 122607 280470 122641 280504
rect 122675 280470 122709 280504
rect 123103 280470 123137 280504
rect 123171 280470 123205 280504
rect 123239 280470 123273 280504
rect 123307 280470 123341 280504
rect 123375 280470 123409 280504
rect 122403 279842 122437 279876
rect 122471 279842 122505 279876
rect 122539 279842 122573 279876
rect 122607 279842 122641 279876
rect 122675 279842 122709 279876
rect 123103 279842 123137 279876
rect 123171 279842 123205 279876
rect 123239 279842 123273 279876
rect 123307 279842 123341 279876
rect 123375 279842 123409 279876
rect 122403 279686 122437 279720
rect 122471 279686 122505 279720
rect 122539 279686 122573 279720
rect 122607 279686 122641 279720
rect 122675 279686 122709 279720
rect 123103 279686 123137 279720
rect 123171 279686 123205 279720
rect 123239 279686 123273 279720
rect 123307 279686 123341 279720
rect 123375 279686 123409 279720
rect 122403 279058 122437 279092
rect 122471 279058 122505 279092
rect 122539 279058 122573 279092
rect 122607 279058 122641 279092
rect 122675 279058 122709 279092
rect 123103 279058 123137 279092
rect 123171 279058 123205 279092
rect 123239 279058 123273 279092
rect 123307 279058 123341 279092
rect 123375 279058 123409 279092
rect 120476 278732 120510 278766
rect 120544 278732 120578 278766
rect 120612 278732 120646 278766
rect 120680 278732 120714 278766
rect 120748 278732 120782 278766
rect 121176 278732 121210 278766
rect 121244 278732 121278 278766
rect 121312 278732 121346 278766
rect 121380 278732 121414 278766
rect 121448 278732 121482 278766
rect 120476 278104 120510 278138
rect 120544 278104 120578 278138
rect 120612 278104 120646 278138
rect 120680 278104 120714 278138
rect 120748 278104 120782 278138
rect 121176 278104 121210 278138
rect 121244 278104 121278 278138
rect 121312 278104 121346 278138
rect 121380 278104 121414 278138
rect 121448 278104 121482 278138
rect 120476 277948 120510 277982
rect 120544 277948 120578 277982
rect 120612 277948 120646 277982
rect 120680 277948 120714 277982
rect 120748 277948 120782 277982
rect 121176 277948 121210 277982
rect 121244 277948 121278 277982
rect 121312 277948 121346 277982
rect 121380 277948 121414 277982
rect 121448 277948 121482 277982
rect 120476 277320 120510 277354
rect 120544 277320 120578 277354
rect 120612 277320 120646 277354
rect 120680 277320 120714 277354
rect 120748 277320 120782 277354
rect 121176 277320 121210 277354
rect 121244 277320 121278 277354
rect 121312 277320 121346 277354
rect 121380 277320 121414 277354
rect 121448 277320 121482 277354
rect 120476 277164 120510 277198
rect 120544 277164 120578 277198
rect 120612 277164 120646 277198
rect 120680 277164 120714 277198
rect 120748 277164 120782 277198
rect 121176 277164 121210 277198
rect 121244 277164 121278 277198
rect 121312 277164 121346 277198
rect 121380 277164 121414 277198
rect 121448 277164 121482 277198
rect 120476 276536 120510 276570
rect 120544 276536 120578 276570
rect 120612 276536 120646 276570
rect 120680 276536 120714 276570
rect 120748 276536 120782 276570
rect 121176 276536 121210 276570
rect 121244 276536 121278 276570
rect 121312 276536 121346 276570
rect 121380 276536 121414 276570
rect 121448 276536 121482 276570
rect 120476 276380 120510 276414
rect 120544 276380 120578 276414
rect 120612 276380 120646 276414
rect 120680 276380 120714 276414
rect 120748 276380 120782 276414
rect 121176 276380 121210 276414
rect 121244 276380 121278 276414
rect 121312 276380 121346 276414
rect 121380 276380 121414 276414
rect 121448 276380 121482 276414
rect 120476 275752 120510 275786
rect 120544 275752 120578 275786
rect 120612 275752 120646 275786
rect 120680 275752 120714 275786
rect 120748 275752 120782 275786
rect 121176 275752 121210 275786
rect 121244 275752 121278 275786
rect 121312 275752 121346 275786
rect 121380 275752 121414 275786
rect 121448 275752 121482 275786
rect 120476 275596 120510 275630
rect 120544 275596 120578 275630
rect 120612 275596 120646 275630
rect 120680 275596 120714 275630
rect 120748 275596 120782 275630
rect 121176 275596 121210 275630
rect 121244 275596 121278 275630
rect 121312 275596 121346 275630
rect 121380 275596 121414 275630
rect 121448 275596 121482 275630
rect 122461 278313 122495 278347
rect 122529 278313 122563 278347
rect 122597 278313 122631 278347
rect 122665 278313 122699 278347
rect 122733 278313 122767 278347
rect 122801 278313 122835 278347
rect 122869 278313 122903 278347
rect 122937 278313 122971 278347
rect 123005 278313 123039 278347
rect 123073 278313 123107 278347
rect 123141 278313 123175 278347
rect 123209 278313 123243 278347
rect 123678 278127 123712 278161
rect 123746 278127 123780 278161
rect 123814 278127 123848 278161
rect 123882 278127 123916 278161
rect 123950 278127 123984 278161
rect 124018 278127 124052 278161
rect 124086 278127 124120 278161
rect 124154 278127 124188 278161
rect 122461 277711 122495 277745
rect 122529 277711 122563 277745
rect 122597 277711 122631 277745
rect 122665 277711 122699 277745
rect 122733 277711 122767 277745
rect 122801 277711 122835 277745
rect 122869 277711 122903 277745
rect 122937 277711 122971 277745
rect 123005 277711 123039 277745
rect 123073 277711 123107 277745
rect 123141 277711 123175 277745
rect 123209 277711 123243 277745
rect 122459 277547 122493 277581
rect 122527 277547 122561 277581
rect 122595 277547 122629 277581
rect 122663 277547 122697 277581
rect 122731 277547 122765 277581
rect 122799 277547 122833 277581
rect 122867 277547 122901 277581
rect 122935 277547 122969 277581
rect 123003 277547 123037 277581
rect 123071 277547 123105 277581
rect 123139 277547 123173 277581
rect 122459 277319 122493 277353
rect 122527 277319 122561 277353
rect 122595 277319 122629 277353
rect 122663 277319 122697 277353
rect 122731 277319 122765 277353
rect 122799 277319 122833 277353
rect 122867 277319 122901 277353
rect 122935 277319 122969 277353
rect 123003 277319 123037 277353
rect 123071 277319 123105 277353
rect 123139 277319 123173 277353
rect 123678 277313 123712 277347
rect 123746 277313 123780 277347
rect 123814 277313 123848 277347
rect 123882 277313 123916 277347
rect 123950 277313 123984 277347
rect 124018 277313 124052 277347
rect 124086 277313 124120 277347
rect 124154 277313 124188 277347
rect 122472 276715 122506 276749
rect 122540 276715 122574 276749
rect 122608 276715 122642 276749
rect 122676 276715 122710 276749
rect 122744 276715 122778 276749
rect 122812 276715 122846 276749
rect 122880 276715 122914 276749
rect 122948 276715 122982 276749
rect 123016 276715 123050 276749
rect 123084 276715 123118 276749
rect 123152 276715 123186 276749
rect 123220 276715 123254 276749
rect 123288 276715 123322 276749
rect 123356 276715 123390 276749
rect 123424 276715 123458 276749
rect 123492 276715 123526 276749
rect 123560 276715 123594 276749
rect 123628 276715 123662 276749
rect 123696 276715 123730 276749
rect 123764 276715 123798 276749
rect 122472 276411 122506 276445
rect 122540 276411 122574 276445
rect 122608 276411 122642 276445
rect 122676 276411 122710 276445
rect 122744 276411 122778 276445
rect 122812 276411 122846 276445
rect 122880 276411 122914 276445
rect 122948 276411 122982 276445
rect 123016 276411 123050 276445
rect 123084 276411 123118 276445
rect 123152 276411 123186 276445
rect 123220 276411 123254 276445
rect 123288 276411 123322 276445
rect 123356 276411 123390 276445
rect 123424 276411 123458 276445
rect 123492 276411 123526 276445
rect 123560 276411 123594 276445
rect 123628 276411 123662 276445
rect 123696 276411 123730 276445
rect 123764 276411 123798 276445
rect 122385 275744 122419 275778
rect 122913 275744 122947 275778
rect 123021 275744 123055 275778
rect 123549 275744 123583 275778
rect 123657 275744 123691 275778
rect 124185 275744 124219 275778
rect 124293 275744 124327 275778
rect 124821 275744 124855 275778
rect 120476 274968 120510 275002
rect 120544 274968 120578 275002
rect 120612 274968 120646 275002
rect 120680 274968 120714 275002
rect 120748 274968 120782 275002
rect 121176 274968 121210 275002
rect 121244 274968 121278 275002
rect 121312 274968 121346 275002
rect 121380 274968 121414 275002
rect 121448 274968 121482 275002
rect 120476 274812 120510 274846
rect 120544 274812 120578 274846
rect 120612 274812 120646 274846
rect 120680 274812 120714 274846
rect 120748 274812 120782 274846
rect 121176 274812 121210 274846
rect 121244 274812 121278 274846
rect 121312 274812 121346 274846
rect 121380 274812 121414 274846
rect 121448 274812 121482 274846
rect 122993 274900 123027 274934
rect 123061 274900 123095 274934
rect 123129 274900 123163 274934
rect 123197 274900 123231 274934
rect 123265 274900 123299 274934
rect 123333 274900 123367 274934
rect 123401 274900 123435 274934
rect 123469 274900 123503 274934
rect 123537 274900 123571 274934
rect 123605 274900 123639 274934
rect 123673 274900 123707 274934
rect 123741 274900 123775 274934
rect 123809 274900 123843 274934
rect 123877 274900 123911 274934
rect 122993 274590 123027 274624
rect 123061 274590 123095 274624
rect 123129 274590 123163 274624
rect 123197 274590 123231 274624
rect 123265 274590 123299 274624
rect 123333 274590 123367 274624
rect 123401 274590 123435 274624
rect 123469 274590 123503 274624
rect 123537 274590 123571 274624
rect 123605 274590 123639 274624
rect 123673 274590 123707 274624
rect 123741 274590 123775 274624
rect 123809 274590 123843 274624
rect 123877 274590 123911 274624
rect 120476 274184 120510 274218
rect 120544 274184 120578 274218
rect 120612 274184 120646 274218
rect 120680 274184 120714 274218
rect 120748 274184 120782 274218
rect 121176 274184 121210 274218
rect 121244 274184 121278 274218
rect 121312 274184 121346 274218
rect 121380 274184 121414 274218
rect 121448 274184 121482 274218
rect 120476 274028 120510 274062
rect 120544 274028 120578 274062
rect 120612 274028 120646 274062
rect 120680 274028 120714 274062
rect 120748 274028 120782 274062
rect 121176 274028 121210 274062
rect 121244 274028 121278 274062
rect 121312 274028 121346 274062
rect 121380 274028 121414 274062
rect 121448 274028 121482 274062
rect 122326 274316 122360 274350
rect 122394 274316 122428 274350
rect 122742 274316 122776 274350
rect 122810 274316 122844 274350
rect 123158 274316 123192 274350
rect 123226 274316 123260 274350
rect 123574 274316 123608 274350
rect 123642 274316 123676 274350
rect 123990 274316 124024 274350
rect 124058 274316 124092 274350
rect 124406 274316 124440 274350
rect 124474 274316 124508 274350
rect 122326 273706 122360 273740
rect 122394 273706 122428 273740
rect 122742 273706 122776 273740
rect 122810 273706 122844 273740
rect 123158 273706 123192 273740
rect 123226 273706 123260 273740
rect 123574 273706 123608 273740
rect 123642 273706 123676 273740
rect 123990 273706 124024 273740
rect 124058 273706 124092 273740
rect 124406 273706 124440 273740
rect 124474 273706 124508 273740
rect 120476 273400 120510 273434
rect 120544 273400 120578 273434
rect 120612 273400 120646 273434
rect 120680 273400 120714 273434
rect 120748 273400 120782 273434
rect 121176 273400 121210 273434
rect 121244 273400 121278 273434
rect 121312 273400 121346 273434
rect 121380 273400 121414 273434
rect 121448 273400 121482 273434
rect 120476 273244 120510 273278
rect 120544 273244 120578 273278
rect 120612 273244 120646 273278
rect 120680 273244 120714 273278
rect 120748 273244 120782 273278
rect 121176 273244 121210 273278
rect 121244 273244 121278 273278
rect 121312 273244 121346 273278
rect 121380 273244 121414 273278
rect 121448 273244 121482 273278
rect 120476 272616 120510 272650
rect 120544 272616 120578 272650
rect 120612 272616 120646 272650
rect 120680 272616 120714 272650
rect 120748 272616 120782 272650
rect 121176 272616 121210 272650
rect 121244 272616 121278 272650
rect 121312 272616 121346 272650
rect 121380 272616 121414 272650
rect 121448 272616 121482 272650
rect 120476 272460 120510 272494
rect 120544 272460 120578 272494
rect 120612 272460 120646 272494
rect 120680 272460 120714 272494
rect 120748 272460 120782 272494
rect 121176 272460 121210 272494
rect 121244 272460 121278 272494
rect 121312 272460 121346 272494
rect 121380 272460 121414 272494
rect 121448 272460 121482 272494
rect 120476 271832 120510 271866
rect 120544 271832 120578 271866
rect 120612 271832 120646 271866
rect 120680 271832 120714 271866
rect 120748 271832 120782 271866
rect 121176 271832 121210 271866
rect 121244 271832 121278 271866
rect 121312 271832 121346 271866
rect 121380 271832 121414 271866
rect 121448 271832 121482 271866
rect 120476 271676 120510 271710
rect 120544 271676 120578 271710
rect 120612 271676 120646 271710
rect 120680 271676 120714 271710
rect 120748 271676 120782 271710
rect 121176 271676 121210 271710
rect 121244 271676 121278 271710
rect 121312 271676 121346 271710
rect 121380 271676 121414 271710
rect 121448 271676 121482 271710
rect 120476 271048 120510 271082
rect 120544 271048 120578 271082
rect 120612 271048 120646 271082
rect 120680 271048 120714 271082
rect 120748 271048 120782 271082
rect 121176 271048 121210 271082
rect 121244 271048 121278 271082
rect 121312 271048 121346 271082
rect 121380 271048 121414 271082
rect 121448 271048 121482 271082
rect 120476 270892 120510 270926
rect 120544 270892 120578 270926
rect 120612 270892 120646 270926
rect 120680 270892 120714 270926
rect 120748 270892 120782 270926
rect 121176 270892 121210 270926
rect 121244 270892 121278 270926
rect 121312 270892 121346 270926
rect 121380 270892 121414 270926
rect 121448 270892 121482 270926
rect 120476 270264 120510 270298
rect 120544 270264 120578 270298
rect 120612 270264 120646 270298
rect 120680 270264 120714 270298
rect 120748 270264 120782 270298
rect 121176 270264 121210 270298
rect 121244 270264 121278 270298
rect 121312 270264 121346 270298
rect 121380 270264 121414 270298
rect 121448 270264 121482 270298
rect 120476 270108 120510 270142
rect 120544 270108 120578 270142
rect 120612 270108 120646 270142
rect 120680 270108 120714 270142
rect 120748 270108 120782 270142
rect 121176 270108 121210 270142
rect 121244 270108 121278 270142
rect 121312 270108 121346 270142
rect 121380 270108 121414 270142
rect 121448 270108 121482 270142
rect 120476 269480 120510 269514
rect 120544 269480 120578 269514
rect 120612 269480 120646 269514
rect 120680 269480 120714 269514
rect 120748 269480 120782 269514
rect 121176 269480 121210 269514
rect 121244 269480 121278 269514
rect 121312 269480 121346 269514
rect 121380 269480 121414 269514
rect 121448 269480 121482 269514
rect 120476 269324 120510 269358
rect 120544 269324 120578 269358
rect 120612 269324 120646 269358
rect 120680 269324 120714 269358
rect 120748 269324 120782 269358
rect 121176 269324 121210 269358
rect 121244 269324 121278 269358
rect 121312 269324 121346 269358
rect 121380 269324 121414 269358
rect 121448 269324 121482 269358
rect 120476 269096 120510 269130
rect 120544 269096 120578 269130
rect 120612 269096 120646 269130
rect 120680 269096 120714 269130
rect 120748 269096 120782 269130
rect 121176 269096 121210 269130
rect 121244 269096 121278 269130
rect 121312 269096 121346 269130
rect 121380 269096 121414 269130
rect 121448 269096 121482 269130
rect 122172 272860 122206 272894
rect 122240 272860 122274 272894
rect 122308 272860 122342 272894
rect 122376 272860 122410 272894
rect 122444 272860 122478 272894
rect 122872 272860 122906 272894
rect 122940 272860 122974 272894
rect 123008 272860 123042 272894
rect 123076 272860 123110 272894
rect 123144 272860 123178 272894
rect 122172 272632 122206 272666
rect 122240 272632 122274 272666
rect 122308 272632 122342 272666
rect 122376 272632 122410 272666
rect 122444 272632 122478 272666
rect 122872 272632 122906 272666
rect 122940 272632 122974 272666
rect 123008 272632 123042 272666
rect 123076 272632 123110 272666
rect 123144 272632 123178 272666
rect 122172 272476 122206 272510
rect 122240 272476 122274 272510
rect 122308 272476 122342 272510
rect 122376 272476 122410 272510
rect 122444 272476 122478 272510
rect 122872 272476 122906 272510
rect 122940 272476 122974 272510
rect 123008 272476 123042 272510
rect 123076 272476 123110 272510
rect 123144 272476 123178 272510
rect 122172 271848 122206 271882
rect 122240 271848 122274 271882
rect 122308 271848 122342 271882
rect 122376 271848 122410 271882
rect 122444 271848 122478 271882
rect 122872 271848 122906 271882
rect 122940 271848 122974 271882
rect 123008 271848 123042 271882
rect 123076 271848 123110 271882
rect 123144 271848 123178 271882
rect 122172 271692 122206 271726
rect 122240 271692 122274 271726
rect 122308 271692 122342 271726
rect 122376 271692 122410 271726
rect 122444 271692 122478 271726
rect 122872 271692 122906 271726
rect 122940 271692 122974 271726
rect 123008 271692 123042 271726
rect 123076 271692 123110 271726
rect 123144 271692 123178 271726
rect 122172 271064 122206 271098
rect 122240 271064 122274 271098
rect 122308 271064 122342 271098
rect 122376 271064 122410 271098
rect 122444 271064 122478 271098
rect 122872 271064 122906 271098
rect 122940 271064 122974 271098
rect 123008 271064 123042 271098
rect 123076 271064 123110 271098
rect 123144 271064 123178 271098
rect 122172 270908 122206 270942
rect 122240 270908 122274 270942
rect 122308 270908 122342 270942
rect 122376 270908 122410 270942
rect 122444 270908 122478 270942
rect 122872 270908 122906 270942
rect 122940 270908 122974 270942
rect 123008 270908 123042 270942
rect 123076 270908 123110 270942
rect 123144 270908 123178 270942
rect 122172 270280 122206 270314
rect 122240 270280 122274 270314
rect 122308 270280 122342 270314
rect 122376 270280 122410 270314
rect 122444 270280 122478 270314
rect 122872 270280 122906 270314
rect 122940 270280 122974 270314
rect 123008 270280 123042 270314
rect 123076 270280 123110 270314
rect 123144 270280 123178 270314
rect 122172 270124 122206 270158
rect 122240 270124 122274 270158
rect 122308 270124 122342 270158
rect 122376 270124 122410 270158
rect 122444 270124 122478 270158
rect 122872 270124 122906 270158
rect 122940 270124 122974 270158
rect 123008 270124 123042 270158
rect 123076 270124 123110 270158
rect 123144 270124 123178 270158
rect 122172 269496 122206 269530
rect 122240 269496 122274 269530
rect 122308 269496 122342 269530
rect 122376 269496 122410 269530
rect 122444 269496 122478 269530
rect 122872 269496 122906 269530
rect 122940 269496 122974 269530
rect 123008 269496 123042 269530
rect 123076 269496 123110 269530
rect 123144 269496 123178 269530
rect 122172 269340 122206 269374
rect 122240 269340 122274 269374
rect 122308 269340 122342 269374
rect 122376 269340 122410 269374
rect 122444 269340 122478 269374
rect 122872 269340 122906 269374
rect 122940 269340 122974 269374
rect 123008 269340 123042 269374
rect 123076 269340 123110 269374
rect 123144 269340 123178 269374
rect 122172 269112 122206 269146
rect 122240 269112 122274 269146
rect 122308 269112 122342 269146
rect 122376 269112 122410 269146
rect 122444 269112 122478 269146
rect 122872 269112 122906 269146
rect 122940 269112 122974 269146
rect 123008 269112 123042 269146
rect 123076 269112 123110 269146
rect 123144 269112 123178 269146
rect 124120 272437 124154 272471
rect 124120 272369 124154 272403
rect 124730 272437 124764 272471
rect 124730 272369 124764 272403
rect 124120 272021 124154 272055
rect 124120 271953 124154 271987
rect 124730 272021 124764 272055
rect 124730 271953 124764 271987
rect 124120 271605 124154 271639
rect 124120 271537 124154 271571
rect 124730 271605 124764 271639
rect 124730 271537 124764 271571
rect 124120 271189 124154 271223
rect 124120 271121 124154 271155
rect 124730 271189 124764 271223
rect 124730 271121 124764 271155
rect 124120 270773 124154 270807
rect 124120 270705 124154 270739
rect 124730 270773 124764 270807
rect 124730 270705 124764 270739
rect 124120 270357 124154 270391
rect 124120 270289 124154 270323
rect 124730 270357 124764 270391
rect 124730 270289 124764 270323
rect 124120 269941 124154 269975
rect 124120 269873 124154 269907
rect 124730 269941 124764 269975
rect 124730 269873 124764 269907
rect 124120 269525 124154 269559
rect 124120 269457 124154 269491
rect 124730 269525 124764 269559
rect 124730 269457 124764 269491
<< locali >>
rect 125105 281915 125658 281925
rect 105823 281315 125658 281915
rect 105976 281064 106456 281315
rect 105974 281045 106456 281064
rect 108743 281045 110315 281315
rect 111807 281179 118652 281315
rect 105974 281020 110315 281045
rect 105974 281017 106176 281020
rect 105974 280983 106000 281017
rect 106034 280986 106176 281017
rect 106210 280986 106244 281020
rect 106278 280986 106312 281020
rect 106346 280986 106380 281020
rect 106414 280986 106448 281020
rect 106482 280986 106516 281020
rect 106550 280986 106584 281020
rect 106618 280986 106652 281020
rect 106686 280986 106720 281020
rect 106754 280986 106788 281020
rect 106822 280986 106856 281020
rect 106890 280986 106924 281020
rect 106958 280986 106992 281020
rect 107026 280986 107060 281020
rect 107094 280986 107128 281020
rect 107162 280986 107196 281020
rect 107230 280986 107264 281020
rect 107298 280986 107332 281020
rect 107366 280986 107400 281020
rect 107434 280986 107468 281020
rect 107502 280986 107536 281020
rect 107570 280986 107604 281020
rect 107638 280986 107672 281020
rect 107706 280986 107740 281020
rect 107774 280986 107808 281020
rect 107842 280986 107876 281020
rect 107910 280986 107944 281020
rect 107978 280986 108012 281020
rect 108046 280986 108080 281020
rect 108114 280986 108148 281020
rect 108182 280986 108216 281020
rect 108250 280986 108284 281020
rect 108318 280986 108352 281020
rect 108386 280986 108420 281020
rect 108454 280986 108488 281020
rect 108522 280986 108556 281020
rect 108590 280986 108624 281020
rect 108658 280986 108692 281020
rect 108726 280986 108760 281020
rect 108794 280986 108828 281020
rect 108862 280986 108896 281020
rect 108930 280986 108964 281020
rect 108998 280986 109032 281020
rect 109066 280986 109100 281020
rect 109134 280986 109168 281020
rect 109202 280986 109236 281020
rect 109270 280986 109304 281020
rect 109338 280986 109372 281020
rect 109406 280986 109440 281020
rect 109474 280986 109508 281020
rect 109542 280986 109576 281020
rect 109610 280986 109644 281020
rect 109678 280986 109712 281020
rect 109746 280986 109780 281020
rect 109814 280986 109848 281020
rect 109882 280986 109916 281020
rect 109950 280986 109984 281020
rect 110018 280986 110052 281020
rect 110086 280986 110120 281020
rect 110154 280986 110188 281020
rect 110222 281005 110315 281020
rect 111046 281156 119159 281179
rect 122520 281165 125658 281315
rect 111046 281122 111264 281156
rect 111298 281122 111332 281156
rect 111366 281122 111400 281156
rect 111434 281122 111468 281156
rect 111502 281122 111536 281156
rect 111570 281122 111604 281156
rect 111638 281122 111672 281156
rect 111706 281122 111740 281156
rect 111774 281122 111808 281156
rect 111842 281122 111876 281156
rect 111910 281122 111944 281156
rect 111978 281122 112012 281156
rect 112046 281122 112080 281156
rect 112114 281122 112148 281156
rect 112182 281122 112216 281156
rect 112250 281122 112284 281156
rect 112318 281122 112352 281156
rect 112386 281122 112420 281156
rect 112454 281122 112488 281156
rect 112522 281122 112556 281156
rect 112590 281122 112624 281156
rect 112658 281122 112692 281156
rect 112726 281122 112760 281156
rect 112794 281122 112828 281156
rect 112862 281122 112896 281156
rect 112930 281122 112964 281156
rect 112998 281122 113032 281156
rect 113066 281122 113100 281156
rect 113134 281122 113168 281156
rect 113202 281122 113236 281156
rect 113270 281122 113304 281156
rect 113338 281122 113372 281156
rect 113406 281122 113440 281156
rect 113474 281122 113508 281156
rect 113542 281122 113576 281156
rect 113610 281122 113644 281156
rect 113678 281122 113712 281156
rect 113746 281122 113780 281156
rect 113814 281122 113848 281156
rect 113882 281122 113916 281156
rect 113950 281122 113984 281156
rect 114018 281122 114052 281156
rect 114086 281122 114120 281156
rect 114154 281122 114188 281156
rect 114222 281122 114256 281156
rect 114290 281122 114324 281156
rect 114358 281122 114392 281156
rect 114426 281122 114460 281156
rect 114494 281122 114528 281156
rect 114562 281122 114596 281156
rect 114630 281122 114664 281156
rect 114698 281122 114732 281156
rect 114766 281122 114800 281156
rect 114834 281122 114868 281156
rect 114902 281122 114936 281156
rect 114970 281122 115004 281156
rect 115038 281122 115072 281156
rect 115106 281122 115140 281156
rect 115174 281122 115208 281156
rect 115242 281122 115276 281156
rect 115310 281122 115344 281156
rect 115378 281122 115412 281156
rect 115446 281122 115480 281156
rect 115514 281122 115548 281156
rect 115582 281122 115616 281156
rect 115650 281122 115684 281156
rect 115718 281122 115752 281156
rect 115786 281122 115820 281156
rect 115854 281122 115888 281156
rect 115922 281122 115956 281156
rect 115990 281122 116024 281156
rect 116058 281122 116092 281156
rect 116126 281122 116160 281156
rect 116194 281122 116228 281156
rect 116262 281122 116296 281156
rect 116330 281122 116364 281156
rect 116398 281122 116432 281156
rect 116466 281122 116500 281156
rect 116534 281122 116568 281156
rect 116602 281122 116636 281156
rect 116670 281122 116704 281156
rect 116738 281122 116772 281156
rect 116806 281122 116840 281156
rect 116874 281122 116908 281156
rect 116942 281122 116976 281156
rect 117010 281122 117044 281156
rect 117078 281122 117112 281156
rect 117146 281122 117180 281156
rect 117214 281122 117248 281156
rect 117282 281122 117316 281156
rect 117350 281122 117384 281156
rect 117418 281122 117452 281156
rect 117486 281122 117520 281156
rect 117554 281122 117588 281156
rect 117622 281122 117656 281156
rect 117690 281122 117724 281156
rect 117758 281122 117792 281156
rect 117826 281122 117860 281156
rect 117894 281122 117928 281156
rect 117962 281122 117996 281156
rect 118030 281122 118064 281156
rect 118098 281122 118132 281156
rect 118166 281122 118200 281156
rect 118234 281122 118268 281156
rect 118302 281122 118336 281156
rect 118370 281122 118404 281156
rect 118438 281122 118472 281156
rect 118506 281122 118540 281156
rect 118574 281122 118608 281156
rect 118642 281122 118676 281156
rect 118710 281122 118744 281156
rect 118778 281122 118812 281156
rect 118846 281122 119159 281156
rect 111046 281102 119159 281122
rect 110222 280986 110313 281005
rect 106034 280983 110313 280986
rect 105974 280961 110313 280983
rect 105974 280949 106465 280961
rect 105974 280915 106000 280949
rect 106034 280915 106465 280949
rect 105974 280885 106465 280915
rect 105974 280881 106406 280885
rect 105974 280847 106000 280881
rect 106034 280859 106406 280881
rect 106034 280847 106149 280859
rect 105974 280825 106149 280847
rect 106183 280851 106406 280859
rect 106440 280851 106489 280885
rect 106183 280825 106345 280851
rect 105974 280813 106345 280825
rect 106666 280817 106711 280961
rect 106757 280851 106806 280885
rect 106840 280851 106889 280885
rect 107066 280817 107111 280961
rect 107157 280851 107206 280885
rect 107240 280851 107289 280885
rect 107466 280817 107511 280961
rect 107557 280851 107606 280885
rect 107640 280851 107689 280885
rect 107866 280817 107911 280961
rect 107957 280851 108006 280885
rect 108040 280851 108089 280885
rect 108357 280851 108406 280885
rect 108440 280851 108489 280885
rect 108535 280817 108580 280961
rect 108757 280851 108806 280885
rect 108840 280851 108889 280885
rect 108935 280817 108980 280961
rect 109157 280851 109206 280885
rect 109240 280851 109289 280885
rect 109335 280817 109380 280961
rect 109557 280851 109606 280885
rect 109640 280851 109689 280885
rect 109735 280817 109780 280961
rect 109980 280885 110313 280961
rect 109957 280851 110006 280885
rect 110040 280851 110313 280885
rect 110129 280841 110313 280851
rect 110129 280817 110255 280841
rect 105974 280779 106000 280813
rect 106034 280796 106345 280813
rect 106034 280791 106311 280796
rect 106034 280779 106149 280791
rect 105974 280757 106149 280779
rect 106183 280757 106311 280791
rect 105974 280754 106311 280757
rect 105974 280745 106345 280754
rect 105974 280711 106000 280745
rect 106034 280728 106345 280745
rect 106034 280723 106311 280728
rect 106034 280711 106149 280723
rect 105974 280689 106149 280711
rect 106183 280689 106311 280723
rect 105974 280682 106311 280689
rect 105974 280677 106345 280682
rect 105974 280643 106000 280677
rect 106034 280660 106345 280677
rect 106034 280655 106311 280660
rect 106034 280643 106149 280655
rect 105974 280621 106149 280643
rect 106183 280621 106311 280655
rect 105974 280610 106311 280621
rect 105974 280609 106345 280610
rect 105974 280575 106000 280609
rect 106034 280592 106345 280609
rect 106034 280587 106311 280592
rect 106034 280575 106149 280587
rect 105974 280553 106149 280575
rect 106183 280553 106311 280587
rect 105974 280541 106311 280553
rect 105974 280507 106000 280541
rect 106034 280538 106311 280541
rect 106034 280524 106345 280538
rect 106034 280519 106311 280524
rect 106034 280507 106149 280519
rect 105974 280485 106149 280507
rect 106183 280485 106311 280519
rect 105974 280473 106311 280485
rect 105974 280439 106000 280473
rect 106034 280466 106311 280473
rect 106034 280456 106345 280466
rect 106034 280451 106311 280456
rect 106034 280439 106149 280451
rect 105974 280417 106149 280439
rect 106183 280417 106311 280451
rect 105974 280405 106311 280417
rect 105974 280371 106000 280405
rect 106034 280394 106311 280405
rect 106034 280388 106345 280394
rect 106034 280383 106311 280388
rect 106034 280371 106149 280383
rect 105974 280349 106149 280371
rect 106183 280349 106311 280383
rect 105974 280337 106311 280349
rect 105974 280303 106000 280337
rect 106034 280322 106311 280337
rect 106034 280320 106345 280322
rect 106034 280315 106311 280320
rect 106034 280303 106149 280315
rect 105974 280281 106149 280303
rect 106183 280286 106311 280315
rect 106183 280284 106345 280286
rect 106183 280281 106311 280284
rect 105974 280269 106311 280281
rect 105974 280235 106000 280269
rect 106034 280247 106311 280269
rect 106034 280235 106149 280247
rect 105974 280213 106149 280235
rect 106183 280218 106311 280247
rect 106183 280213 106345 280218
rect 105974 280212 106345 280213
rect 105974 280201 106311 280212
rect 105974 280167 106000 280201
rect 106034 280179 106311 280201
rect 106034 280167 106149 280179
rect 105974 280145 106149 280167
rect 106183 280150 106311 280179
rect 106183 280145 106345 280150
rect 105974 280140 106345 280145
rect 105974 280133 106311 280140
rect 105974 280099 106000 280133
rect 106034 280111 106311 280133
rect 106034 280099 106149 280111
rect 105974 280077 106149 280099
rect 106183 280082 106311 280111
rect 106183 280077 106345 280082
rect 105974 280068 106345 280077
rect 105974 280065 106311 280068
rect 105974 280031 106000 280065
rect 106034 280043 106311 280065
rect 106034 280031 106149 280043
rect 105974 280009 106149 280031
rect 106183 280014 106311 280043
rect 106183 280009 106345 280014
rect 105974 279997 106345 280009
rect 105974 279963 106000 279997
rect 106034 279996 106345 279997
rect 106034 279975 106311 279996
rect 106034 279963 106149 279975
rect 105974 279941 106149 279963
rect 106183 279946 106311 279975
rect 106183 279941 106345 279946
rect 105974 279929 106345 279941
rect 105974 279895 106000 279929
rect 106034 279924 106345 279929
rect 106034 279907 106311 279924
rect 106034 279895 106149 279907
rect 105974 279873 106149 279895
rect 106183 279878 106311 279907
rect 106183 279873 106345 279878
rect 105974 279861 106345 279873
rect 105974 279827 106000 279861
rect 106034 279852 106345 279861
rect 106034 279839 106311 279852
rect 106034 279827 106149 279839
rect 105974 279805 106149 279827
rect 106183 279810 106311 279839
rect 106183 279805 106345 279810
rect 105974 279793 106345 279805
rect 105974 279759 106000 279793
rect 106034 279789 106345 279793
rect 106501 280796 106535 280817
rect 106501 280728 106535 280754
rect 106501 280660 106535 280682
rect 106501 280592 106535 280610
rect 106501 280524 106535 280538
rect 106501 280456 106535 280466
rect 106501 280388 106535 280394
rect 106501 280320 106535 280322
rect 106501 280284 106535 280286
rect 106501 280212 106535 280218
rect 106501 280140 106535 280150
rect 106501 280068 106535 280082
rect 106501 279996 106535 280014
rect 106501 279924 106535 279946
rect 106501 279852 106535 279878
rect 106501 279789 106535 279810
rect 106666 280796 106745 280817
rect 106666 280754 106711 280796
rect 106666 280728 106745 280754
rect 106666 280682 106711 280728
rect 106666 280660 106745 280682
rect 106666 280610 106711 280660
rect 106666 280592 106745 280610
rect 106666 280538 106711 280592
rect 106666 280524 106745 280538
rect 106666 280466 106711 280524
rect 106666 280456 106745 280466
rect 106666 280394 106711 280456
rect 106666 280388 106745 280394
rect 106666 280322 106711 280388
rect 106666 280320 106745 280322
rect 106666 280286 106711 280320
rect 106666 280284 106745 280286
rect 106666 280218 106711 280284
rect 106666 280212 106745 280218
rect 106666 280150 106711 280212
rect 106666 280140 106745 280150
rect 106666 280082 106711 280140
rect 106666 280068 106745 280082
rect 106666 280014 106711 280068
rect 106666 279996 106745 280014
rect 106666 279946 106711 279996
rect 106666 279924 106745 279946
rect 106666 279878 106711 279924
rect 106666 279852 106745 279878
rect 106666 279810 106711 279852
rect 106666 279789 106745 279810
rect 106901 280796 106935 280817
rect 106901 280728 106935 280754
rect 106901 280660 106935 280682
rect 106901 280592 106935 280610
rect 106901 280524 106935 280538
rect 106901 280456 106935 280466
rect 106901 280388 106935 280394
rect 106901 280320 106935 280322
rect 106901 280284 106935 280286
rect 106901 280212 106935 280218
rect 106901 280140 106935 280150
rect 106901 280068 106935 280082
rect 106901 279996 106935 280014
rect 106901 279924 106935 279946
rect 106901 279852 106935 279878
rect 106901 279789 106935 279810
rect 107066 280796 107145 280817
rect 107066 280754 107111 280796
rect 107066 280728 107145 280754
rect 107066 280682 107111 280728
rect 107066 280660 107145 280682
rect 107066 280610 107111 280660
rect 107066 280592 107145 280610
rect 107066 280538 107111 280592
rect 107066 280524 107145 280538
rect 107066 280466 107111 280524
rect 107066 280456 107145 280466
rect 107066 280394 107111 280456
rect 107066 280388 107145 280394
rect 107066 280322 107111 280388
rect 107066 280320 107145 280322
rect 107066 280286 107111 280320
rect 107066 280284 107145 280286
rect 107066 280218 107111 280284
rect 107066 280212 107145 280218
rect 107066 280150 107111 280212
rect 107066 280140 107145 280150
rect 107066 280082 107111 280140
rect 107066 280068 107145 280082
rect 107066 280014 107111 280068
rect 107066 279996 107145 280014
rect 107066 279946 107111 279996
rect 107066 279924 107145 279946
rect 107066 279878 107111 279924
rect 107066 279852 107145 279878
rect 107066 279810 107111 279852
rect 107066 279789 107145 279810
rect 107301 280796 107335 280817
rect 107301 280728 107335 280754
rect 107301 280660 107335 280682
rect 107301 280592 107335 280610
rect 107301 280524 107335 280538
rect 107301 280456 107335 280466
rect 107301 280388 107335 280394
rect 107301 280320 107335 280322
rect 107301 280284 107335 280286
rect 107301 280212 107335 280218
rect 107301 280140 107335 280150
rect 107301 280068 107335 280082
rect 107301 279996 107335 280014
rect 107301 279924 107335 279946
rect 107301 279852 107335 279878
rect 107301 279789 107335 279810
rect 107466 280796 107545 280817
rect 107466 280754 107511 280796
rect 107466 280728 107545 280754
rect 107466 280682 107511 280728
rect 107466 280660 107545 280682
rect 107466 280610 107511 280660
rect 107466 280592 107545 280610
rect 107466 280538 107511 280592
rect 107466 280524 107545 280538
rect 107466 280466 107511 280524
rect 107466 280456 107545 280466
rect 107466 280394 107511 280456
rect 107466 280388 107545 280394
rect 107466 280322 107511 280388
rect 107466 280320 107545 280322
rect 107466 280286 107511 280320
rect 107466 280284 107545 280286
rect 107466 280218 107511 280284
rect 107466 280212 107545 280218
rect 107466 280150 107511 280212
rect 107466 280140 107545 280150
rect 107466 280082 107511 280140
rect 107466 280068 107545 280082
rect 107466 280014 107511 280068
rect 107466 279996 107545 280014
rect 107466 279946 107511 279996
rect 107466 279924 107545 279946
rect 107466 279878 107511 279924
rect 107466 279852 107545 279878
rect 107466 279810 107511 279852
rect 107466 279789 107545 279810
rect 107701 280796 107735 280817
rect 107701 280728 107735 280754
rect 107701 280660 107735 280682
rect 107701 280592 107735 280610
rect 107701 280524 107735 280538
rect 107701 280456 107735 280466
rect 107701 280388 107735 280394
rect 107701 280320 107735 280322
rect 107701 280284 107735 280286
rect 107701 280212 107735 280218
rect 107701 280140 107735 280150
rect 107701 280068 107735 280082
rect 107701 279996 107735 280014
rect 107701 279924 107735 279946
rect 107701 279852 107735 279878
rect 107701 279789 107735 279810
rect 107866 280796 107945 280817
rect 107866 280754 107911 280796
rect 107866 280728 107945 280754
rect 107866 280682 107911 280728
rect 107866 280660 107945 280682
rect 107866 280610 107911 280660
rect 107866 280592 107945 280610
rect 107866 280538 107911 280592
rect 107866 280524 107945 280538
rect 107866 280466 107911 280524
rect 107866 280456 107945 280466
rect 107866 280394 107911 280456
rect 107866 280388 107945 280394
rect 107866 280322 107911 280388
rect 107866 280320 107945 280322
rect 107866 280286 107911 280320
rect 107866 280284 107945 280286
rect 107866 280218 107911 280284
rect 107866 280212 107945 280218
rect 107866 280150 107911 280212
rect 107866 280140 107945 280150
rect 107866 280082 107911 280140
rect 107866 280068 107945 280082
rect 107866 280014 107911 280068
rect 107866 279996 107945 280014
rect 107866 279946 107911 279996
rect 107866 279924 107945 279946
rect 107866 279878 107911 279924
rect 107866 279852 107945 279878
rect 107866 279810 107911 279852
rect 107866 279789 107945 279810
rect 108101 280796 108135 280817
rect 108101 280728 108135 280754
rect 108101 280660 108135 280682
rect 108101 280592 108135 280610
rect 108101 280524 108135 280538
rect 108101 280456 108135 280466
rect 108101 280388 108135 280394
rect 108101 280320 108135 280322
rect 108101 280284 108135 280286
rect 108101 280212 108135 280218
rect 108101 280140 108135 280150
rect 108101 280068 108135 280082
rect 108101 279996 108135 280014
rect 108101 279924 108135 279946
rect 108101 279852 108135 279878
rect 108101 279789 108135 279810
rect 108311 280796 108345 280817
rect 108311 280728 108345 280754
rect 108311 280660 108345 280682
rect 108311 280592 108345 280610
rect 108311 280524 108345 280538
rect 108311 280456 108345 280466
rect 108311 280388 108345 280394
rect 108311 280320 108345 280322
rect 108311 280284 108345 280286
rect 108311 280212 108345 280218
rect 108311 280140 108345 280150
rect 108311 280068 108345 280082
rect 108311 279996 108345 280014
rect 108311 279924 108345 279946
rect 108311 279852 108345 279878
rect 108311 279789 108345 279810
rect 108501 280796 108580 280817
rect 108535 280754 108580 280796
rect 108501 280728 108580 280754
rect 108535 280682 108580 280728
rect 108501 280660 108580 280682
rect 108535 280610 108580 280660
rect 108501 280592 108580 280610
rect 108535 280538 108580 280592
rect 108501 280524 108580 280538
rect 108535 280466 108580 280524
rect 108501 280456 108580 280466
rect 108535 280394 108580 280456
rect 108501 280388 108580 280394
rect 108535 280322 108580 280388
rect 108501 280320 108580 280322
rect 108535 280286 108580 280320
rect 108501 280284 108580 280286
rect 108535 280218 108580 280284
rect 108501 280212 108580 280218
rect 108535 280150 108580 280212
rect 108501 280140 108580 280150
rect 108535 280082 108580 280140
rect 108501 280068 108580 280082
rect 108535 280014 108580 280068
rect 108501 279996 108580 280014
rect 108535 279946 108580 279996
rect 108501 279924 108580 279946
rect 108535 279878 108580 279924
rect 108501 279852 108580 279878
rect 108535 279810 108580 279852
rect 108501 279789 108580 279810
rect 108711 280796 108745 280817
rect 108711 280728 108745 280754
rect 108711 280660 108745 280682
rect 108711 280592 108745 280610
rect 108711 280524 108745 280538
rect 108711 280456 108745 280466
rect 108711 280388 108745 280394
rect 108711 280320 108745 280322
rect 108711 280284 108745 280286
rect 108711 280212 108745 280218
rect 108711 280140 108745 280150
rect 108711 280068 108745 280082
rect 108711 279996 108745 280014
rect 108711 279924 108745 279946
rect 108711 279852 108745 279878
rect 108711 279789 108745 279810
rect 108901 280796 108980 280817
rect 108935 280754 108980 280796
rect 108901 280728 108980 280754
rect 108935 280682 108980 280728
rect 108901 280660 108980 280682
rect 108935 280610 108980 280660
rect 108901 280592 108980 280610
rect 108935 280538 108980 280592
rect 108901 280524 108980 280538
rect 108935 280466 108980 280524
rect 108901 280456 108980 280466
rect 108935 280394 108980 280456
rect 108901 280388 108980 280394
rect 108935 280322 108980 280388
rect 108901 280320 108980 280322
rect 108935 280286 108980 280320
rect 108901 280284 108980 280286
rect 108935 280218 108980 280284
rect 108901 280212 108980 280218
rect 108935 280150 108980 280212
rect 108901 280140 108980 280150
rect 108935 280082 108980 280140
rect 108901 280068 108980 280082
rect 108935 280014 108980 280068
rect 108901 279996 108980 280014
rect 108935 279946 108980 279996
rect 108901 279924 108980 279946
rect 108935 279878 108980 279924
rect 108901 279852 108980 279878
rect 108935 279810 108980 279852
rect 108901 279789 108980 279810
rect 109111 280796 109145 280817
rect 109111 280728 109145 280754
rect 109111 280660 109145 280682
rect 109111 280592 109145 280610
rect 109111 280524 109145 280538
rect 109111 280456 109145 280466
rect 109111 280388 109145 280394
rect 109111 280320 109145 280322
rect 109111 280284 109145 280286
rect 109111 280212 109145 280218
rect 109111 280140 109145 280150
rect 109111 280068 109145 280082
rect 109111 279996 109145 280014
rect 109111 279924 109145 279946
rect 109111 279852 109145 279878
rect 109111 279789 109145 279810
rect 109301 280796 109380 280817
rect 109335 280754 109380 280796
rect 109301 280728 109380 280754
rect 109335 280682 109380 280728
rect 109301 280660 109380 280682
rect 109335 280610 109380 280660
rect 109301 280592 109380 280610
rect 109335 280538 109380 280592
rect 109301 280524 109380 280538
rect 109335 280466 109380 280524
rect 109301 280456 109380 280466
rect 109335 280394 109380 280456
rect 109301 280388 109380 280394
rect 109335 280322 109380 280388
rect 109301 280320 109380 280322
rect 109335 280286 109380 280320
rect 109301 280284 109380 280286
rect 109335 280218 109380 280284
rect 109301 280212 109380 280218
rect 109335 280150 109380 280212
rect 109301 280140 109380 280150
rect 109335 280082 109380 280140
rect 109301 280068 109380 280082
rect 109335 280014 109380 280068
rect 109301 279996 109380 280014
rect 109335 279946 109380 279996
rect 109301 279924 109380 279946
rect 109335 279878 109380 279924
rect 109301 279852 109380 279878
rect 109335 279810 109380 279852
rect 109301 279789 109380 279810
rect 109511 280796 109545 280817
rect 109511 280728 109545 280754
rect 109511 280660 109545 280682
rect 109511 280592 109545 280610
rect 109511 280524 109545 280538
rect 109511 280456 109545 280466
rect 109511 280388 109545 280394
rect 109511 280320 109545 280322
rect 109511 280284 109545 280286
rect 109511 280212 109545 280218
rect 109511 280140 109545 280150
rect 109511 280068 109545 280082
rect 109511 279996 109545 280014
rect 109511 279924 109545 279946
rect 109511 279852 109545 279878
rect 109511 279789 109545 279810
rect 109701 280796 109780 280817
rect 109735 280754 109780 280796
rect 109701 280728 109780 280754
rect 109735 280682 109780 280728
rect 109701 280660 109780 280682
rect 109735 280610 109780 280660
rect 109701 280592 109780 280610
rect 109735 280538 109780 280592
rect 109701 280524 109780 280538
rect 109735 280466 109780 280524
rect 109701 280456 109780 280466
rect 109735 280394 109780 280456
rect 109701 280388 109780 280394
rect 109735 280322 109780 280388
rect 109701 280320 109780 280322
rect 109735 280286 109780 280320
rect 109701 280284 109780 280286
rect 109735 280218 109780 280284
rect 109701 280212 109780 280218
rect 109735 280150 109780 280212
rect 109701 280140 109780 280150
rect 109735 280082 109780 280140
rect 109701 280068 109780 280082
rect 109735 280014 109780 280068
rect 109701 279996 109780 280014
rect 109735 279946 109780 279996
rect 109701 279924 109780 279946
rect 109735 279878 109780 279924
rect 109701 279852 109780 279878
rect 109735 279810 109780 279852
rect 109701 279789 109780 279810
rect 109911 280796 109945 280817
rect 109911 280728 109945 280754
rect 109911 280660 109945 280682
rect 109911 280592 109945 280610
rect 109911 280524 109945 280538
rect 109911 280456 109945 280466
rect 109911 280388 109945 280394
rect 109911 280320 109945 280322
rect 109911 280284 109945 280286
rect 109911 280212 109945 280218
rect 109911 280140 109945 280150
rect 109911 280068 109945 280082
rect 109911 279996 109945 280014
rect 109911 279924 109945 279946
rect 109911 279852 109945 279878
rect 109911 279789 109945 279810
rect 110101 280807 110255 280817
rect 110289 280807 110313 280841
rect 110101 280796 110313 280807
rect 110135 280773 110313 280796
rect 110135 280754 110255 280773
rect 110101 280739 110255 280754
rect 110289 280739 110313 280773
rect 110101 280728 110313 280739
rect 110135 280705 110313 280728
rect 110135 280682 110255 280705
rect 110101 280671 110255 280682
rect 110289 280671 110313 280705
rect 110101 280660 110313 280671
rect 110135 280637 110313 280660
rect 110135 280610 110255 280637
rect 110101 280603 110255 280610
rect 110289 280603 110313 280637
rect 110101 280592 110313 280603
rect 110135 280569 110313 280592
rect 110135 280538 110255 280569
rect 110101 280535 110255 280538
rect 110289 280535 110313 280569
rect 110101 280524 110313 280535
rect 110135 280501 110313 280524
rect 110135 280467 110255 280501
rect 110289 280467 110313 280501
rect 110135 280466 110313 280467
rect 110101 280456 110313 280466
rect 110135 280433 110313 280456
rect 110135 280399 110255 280433
rect 110289 280399 110313 280433
rect 110135 280394 110313 280399
rect 110101 280388 110313 280394
rect 110135 280365 110313 280388
rect 110135 280331 110255 280365
rect 110289 280331 110313 280365
rect 110135 280322 110313 280331
rect 110101 280320 110313 280322
rect 110135 280297 110313 280320
rect 110135 280286 110255 280297
rect 110101 280284 110255 280286
rect 110135 280263 110255 280284
rect 110289 280263 110313 280297
rect 110135 280229 110313 280263
rect 110135 280218 110255 280229
rect 110101 280212 110255 280218
rect 110135 280195 110255 280212
rect 110289 280195 110313 280229
rect 110135 280161 110313 280195
rect 110135 280150 110255 280161
rect 110101 280140 110255 280150
rect 110135 280127 110255 280140
rect 110289 280127 110313 280161
rect 110135 280093 110313 280127
rect 110135 280082 110255 280093
rect 110101 280068 110255 280082
rect 110135 280059 110255 280068
rect 110289 280059 110313 280093
rect 110135 280025 110313 280059
rect 110135 280014 110255 280025
rect 110101 279996 110255 280014
rect 110135 279991 110255 279996
rect 110289 279991 110313 280025
rect 110135 279957 110313 279991
rect 110135 279946 110255 279957
rect 110101 279924 110255 279946
rect 110135 279923 110255 279924
rect 110289 279923 110313 279957
rect 110135 279889 110313 279923
rect 110135 279878 110255 279889
rect 110101 279855 110255 279878
rect 110289 279855 110313 279889
rect 110101 279852 110313 279855
rect 110135 279821 110313 279852
rect 110135 279810 110255 279821
rect 110101 279789 110255 279810
rect 106034 279771 106326 279789
rect 106034 279759 106149 279771
rect 105974 279737 106149 279759
rect 106183 279755 106326 279771
rect 106489 279755 106535 279789
rect 109911 279755 109957 279789
rect 110129 279787 110255 279789
rect 110289 279787 110313 279821
rect 106183 279737 106406 279755
rect 105974 279725 106406 279737
rect 105974 279691 106000 279725
rect 106034 279721 106406 279725
rect 106440 279721 106535 279755
rect 106757 279721 106806 279755
rect 106840 279721 106889 279755
rect 107157 279721 107206 279755
rect 107240 279721 107289 279755
rect 107557 279721 107606 279755
rect 107640 279721 107689 279755
rect 107957 279721 108006 279755
rect 108040 279721 108089 279755
rect 108357 279721 108406 279755
rect 108440 279721 108489 279755
rect 108757 279721 108806 279755
rect 108840 279721 108889 279755
rect 109157 279721 109206 279755
rect 109240 279721 109289 279755
rect 109557 279721 109606 279755
rect 109640 279721 109689 279755
rect 109911 279721 110006 279755
rect 110040 279747 110089 279755
rect 110129 279753 110313 279787
rect 110129 279747 110255 279753
rect 110040 279721 110255 279747
rect 106034 279691 106463 279721
rect 105974 279657 106463 279691
rect 106757 279687 109689 279721
rect 109982 279719 110255 279721
rect 110289 279719 110313 279753
rect 105974 279623 106000 279657
rect 106034 279625 106463 279657
rect 109982 279625 110313 279719
rect 106034 279623 110313 279625
rect 105974 279600 110313 279623
rect 105974 279589 106176 279600
rect 105974 279555 106000 279589
rect 106034 279566 106176 279589
rect 106210 279566 106244 279600
rect 106278 279566 106312 279600
rect 106346 279566 106380 279600
rect 106414 279566 106448 279600
rect 106482 279566 106516 279600
rect 106550 279566 106584 279600
rect 106618 279566 106652 279600
rect 106686 279566 106720 279600
rect 106754 279566 106788 279600
rect 106822 279566 106856 279600
rect 106890 279566 106924 279600
rect 106958 279566 106992 279600
rect 107026 279566 107060 279600
rect 107094 279566 107128 279600
rect 107162 279566 107196 279600
rect 107230 279566 107264 279600
rect 107298 279566 107332 279600
rect 107366 279566 107400 279600
rect 107434 279566 107468 279600
rect 107502 279566 107536 279600
rect 107570 279566 107604 279600
rect 107638 279566 107672 279600
rect 107706 279566 107740 279600
rect 107774 279566 107808 279600
rect 107842 279566 107876 279600
rect 107910 279566 107944 279600
rect 107978 279566 108012 279600
rect 108046 279566 108080 279600
rect 108114 279566 108148 279600
rect 108182 279566 108216 279600
rect 108250 279566 108284 279600
rect 108318 279566 108352 279600
rect 108386 279566 108420 279600
rect 108454 279566 108488 279600
rect 108522 279566 108556 279600
rect 108590 279566 108624 279600
rect 108658 279566 108692 279600
rect 108726 279566 108760 279600
rect 108794 279566 108828 279600
rect 108862 279566 108896 279600
rect 108930 279566 108964 279600
rect 108998 279566 109032 279600
rect 109066 279566 109100 279600
rect 109134 279566 109168 279600
rect 109202 279566 109236 279600
rect 109270 279566 109304 279600
rect 109338 279566 109372 279600
rect 109406 279566 109440 279600
rect 109474 279566 109508 279600
rect 109542 279566 109576 279600
rect 109610 279566 109644 279600
rect 109678 279566 109712 279600
rect 109746 279566 109780 279600
rect 109814 279566 109848 279600
rect 109882 279566 109916 279600
rect 109950 279566 109984 279600
rect 110018 279566 110052 279600
rect 110086 279566 110120 279600
rect 110154 279566 110188 279600
rect 110222 279566 110313 279600
rect 106034 279555 110313 279566
rect 105974 279549 110313 279555
rect 105974 279521 106060 279549
rect 106125 279541 110313 279549
rect 105974 279487 106000 279521
rect 106034 279487 106060 279521
rect 105974 279453 106060 279487
rect 105974 279419 106000 279453
rect 106034 279419 106060 279453
rect 105974 279385 106060 279419
rect 105974 279351 106000 279385
rect 106034 279351 106060 279385
rect 105974 279317 106060 279351
rect 105974 279283 106000 279317
rect 106034 279283 106060 279317
rect 105974 279249 106060 279283
rect 105974 279215 106000 279249
rect 106034 279215 106060 279249
rect 105974 279181 106060 279215
rect 105974 279147 106000 279181
rect 106034 279147 106060 279181
rect 105974 279113 106060 279147
rect 105974 279079 106000 279113
rect 106034 279079 106060 279113
rect 105974 279045 106060 279079
rect 105974 279011 106000 279045
rect 106034 279011 106060 279045
rect 105974 278977 106060 279011
rect 105974 278943 106000 278977
rect 106034 278943 106060 278977
rect 105974 278909 106060 278943
rect 105974 278875 106000 278909
rect 106034 278875 106060 278909
rect 105974 278841 106060 278875
rect 105974 278807 106000 278841
rect 106034 278807 106060 278841
rect 105974 278773 106060 278807
rect 105974 278739 106000 278773
rect 106034 278739 106060 278773
rect 105974 278705 106060 278739
rect 105974 278671 106000 278705
rect 106034 278671 106060 278705
rect 105974 278637 106060 278671
rect 105974 278603 106000 278637
rect 106034 278603 106060 278637
rect 105974 278569 106060 278603
rect 105974 278535 106000 278569
rect 106034 278535 106060 278569
rect 105974 278501 106060 278535
rect 105974 278467 106000 278501
rect 106034 278467 106060 278501
rect 105974 278433 106060 278467
rect 105974 278399 106000 278433
rect 106034 278399 106060 278433
rect 105974 278365 106060 278399
rect 105974 278331 106000 278365
rect 106034 278331 106060 278365
rect 105974 278297 106060 278331
rect 105974 278263 106000 278297
rect 106034 278263 106060 278297
rect 105974 278229 106060 278263
rect 105974 278195 106000 278229
rect 106034 278195 106060 278229
rect 105974 278161 106060 278195
rect 105974 278127 106000 278161
rect 106034 278127 106060 278161
rect 105974 278093 106060 278127
rect 105974 278059 106000 278093
rect 106034 278059 106060 278093
rect 105974 278025 106060 278059
rect 105974 277991 106000 278025
rect 106034 277991 106060 278025
rect 105974 277957 106060 277991
rect 105974 277923 106000 277957
rect 106034 277923 106060 277957
rect 106169 279188 106237 279222
rect 106271 279188 106305 279222
rect 106339 279188 106373 279222
rect 106407 279188 106441 279222
rect 106475 279188 106509 279222
rect 106543 279188 106577 279222
rect 106611 279188 106645 279222
rect 106679 279188 106713 279222
rect 106747 279188 106781 279222
rect 106815 279188 106849 279222
rect 106883 279188 106917 279222
rect 106951 279188 106985 279222
rect 107019 279188 107053 279222
rect 107087 279188 107121 279222
rect 107155 279188 107189 279222
rect 107223 279188 107257 279222
rect 107291 279188 107325 279222
rect 107359 279188 107393 279222
rect 107427 279188 107461 279222
rect 107495 279188 107529 279222
rect 107563 279188 107597 279222
rect 107631 279188 107665 279222
rect 107699 279188 107768 279222
rect 106169 279147 106203 279188
rect 106169 279079 106203 279113
rect 107734 279147 107768 279188
rect 109636 279185 110312 279541
rect 107734 279079 107768 279113
rect 106169 279011 106203 279045
rect 106364 279023 106380 279057
rect 106416 279023 106448 279057
rect 106488 279023 106516 279057
rect 106560 279023 106584 279057
rect 106632 279023 106652 279057
rect 106704 279023 106720 279057
rect 106776 279023 106788 279057
rect 106848 279023 106856 279057
rect 106920 279023 106924 279057
rect 107026 279023 107030 279057
rect 107094 279023 107102 279057
rect 107162 279023 107174 279057
rect 107230 279023 107246 279057
rect 107298 279023 107318 279057
rect 107366 279023 107390 279057
rect 107434 279023 107462 279057
rect 107502 279023 107534 279057
rect 107570 279023 107586 279057
rect 107734 279011 107768 279045
rect 106169 278943 106203 278977
rect 106169 278875 106203 278909
rect 106169 278807 106203 278841
rect 106169 278739 106203 278773
rect 106169 278671 106203 278705
rect 106169 278603 106203 278637
rect 106169 278535 106203 278569
rect 106169 278467 106203 278501
rect 106169 278399 106203 278433
rect 106169 278331 106203 278365
rect 106169 278263 106203 278297
rect 106169 278195 106203 278229
rect 106169 278127 106203 278161
rect 106275 278973 106321 279011
rect 106275 278935 106287 278973
rect 106275 278901 106321 278935
rect 106275 278867 106287 278901
rect 106275 278833 106321 278867
rect 106275 278795 106287 278833
rect 106275 278373 106321 278795
rect 107629 278973 107675 279011
rect 107663 278935 107675 278973
rect 107629 278901 107675 278935
rect 107663 278867 107675 278901
rect 107629 278833 107675 278867
rect 107663 278795 107675 278833
rect 106364 278711 106380 278745
rect 106416 278711 106448 278745
rect 106488 278711 106516 278745
rect 106560 278711 106584 278745
rect 106632 278711 106652 278745
rect 106704 278711 106720 278745
rect 106776 278711 106788 278745
rect 106848 278711 106856 278745
rect 106920 278711 106924 278745
rect 107026 278711 107030 278745
rect 107094 278711 107102 278745
rect 107162 278711 107174 278745
rect 107230 278711 107246 278745
rect 107298 278711 107318 278745
rect 107366 278711 107390 278745
rect 107434 278711 107462 278745
rect 107502 278711 107534 278745
rect 107570 278711 107586 278745
rect 106364 278423 106380 278457
rect 106416 278423 106448 278457
rect 106488 278423 106516 278457
rect 106560 278423 106584 278457
rect 106632 278423 106652 278457
rect 106704 278423 106720 278457
rect 106776 278423 106788 278457
rect 106848 278423 106856 278457
rect 106920 278423 106924 278457
rect 107026 278423 107030 278457
rect 107094 278423 107102 278457
rect 107162 278423 107174 278457
rect 107230 278423 107246 278457
rect 107298 278423 107318 278457
rect 107366 278423 107390 278457
rect 107434 278423 107462 278457
rect 107502 278423 107534 278457
rect 107570 278423 107586 278457
rect 106275 278335 106287 278373
rect 106275 278301 106321 278335
rect 106275 278267 106287 278301
rect 106275 278233 106321 278267
rect 106275 278195 106287 278233
rect 106275 278157 106321 278195
rect 107629 278373 107675 278795
rect 107663 278335 107675 278373
rect 107629 278301 107675 278335
rect 107663 278267 107675 278301
rect 107629 278233 107675 278267
rect 107663 278195 107675 278233
rect 107629 278157 107675 278195
rect 107734 278943 107768 278977
rect 107734 278875 107768 278909
rect 107734 278807 107768 278841
rect 107734 278739 107768 278773
rect 107734 278671 107768 278705
rect 107734 278603 107768 278637
rect 107734 278535 107768 278569
rect 107734 278467 107768 278501
rect 107734 278399 107768 278433
rect 107734 278331 107768 278365
rect 107734 278263 107768 278297
rect 107734 278195 107768 278229
rect 106364 278111 106380 278145
rect 106416 278111 106448 278145
rect 106488 278111 106516 278145
rect 106560 278111 106584 278145
rect 106632 278111 106652 278145
rect 106704 278111 106720 278145
rect 106776 278111 106788 278145
rect 106848 278111 106856 278145
rect 106920 278111 106924 278145
rect 107026 278111 107030 278145
rect 107094 278111 107102 278145
rect 107162 278111 107174 278145
rect 107230 278111 107246 278145
rect 107298 278111 107318 278145
rect 107366 278111 107390 278145
rect 107434 278111 107462 278145
rect 107502 278111 107534 278145
rect 107570 278111 107586 278145
rect 107734 278127 107768 278161
rect 106169 278059 106203 278093
rect 106169 277984 106203 278025
rect 106762 278053 107237 278111
rect 106762 277984 106966 278053
rect 107072 277984 107237 278053
rect 107734 278059 107768 278093
rect 107734 277984 107768 278025
rect 106169 277950 106237 277984
rect 106271 277950 106305 277984
rect 106339 277950 106373 277984
rect 106407 277950 106441 277984
rect 106475 277950 106509 277984
rect 106543 277950 106577 277984
rect 106611 277950 106645 277984
rect 106679 277950 106713 277984
rect 106747 277950 106781 277984
rect 106815 277950 106849 277984
rect 106883 277950 106917 277984
rect 106951 277950 106966 277984
rect 107087 277950 107121 277984
rect 107155 277950 107189 277984
rect 107223 277950 107257 277984
rect 107291 277950 107325 277984
rect 107359 277950 107393 277984
rect 107427 277950 107461 277984
rect 107495 277950 107529 277984
rect 107563 277950 107597 277984
rect 107631 277950 107665 277984
rect 107699 277950 107768 277984
rect 109617 279151 109733 279185
rect 109767 279151 109801 279185
rect 109835 279151 109869 279185
rect 109903 279151 109937 279185
rect 109971 279151 110005 279185
rect 110039 279151 110073 279185
rect 110107 279151 110312 279185
rect 109617 279071 109651 279151
rect 109777 279049 109795 279083
rect 109835 279049 109867 279083
rect 109903 279049 109937 279083
rect 109973 279049 110005 279083
rect 110045 279049 110063 279083
rect 110189 279071 110312 279151
rect 109617 279003 109651 279037
rect 110223 279037 110312 279071
rect 109617 278935 109651 278969
rect 109617 278867 109651 278901
rect 109617 278799 109651 278833
rect 109617 278731 109651 278765
rect 109617 278663 109651 278697
rect 109617 278595 109651 278629
rect 109617 278527 109651 278561
rect 109617 278459 109651 278493
rect 109617 278391 109651 278425
rect 109617 278323 109651 278357
rect 109617 278255 109651 278289
rect 109617 278187 109651 278221
rect 109617 278119 109651 278153
rect 109617 278051 109651 278085
rect 109617 277983 109651 278017
rect 105974 277889 106060 277923
rect 105974 277855 106000 277889
rect 106034 277855 106060 277889
rect 105974 277821 106060 277855
rect 105974 277787 106000 277821
rect 106034 277787 106060 277821
rect 105974 277753 106060 277787
rect 105974 277719 106000 277753
rect 106034 277719 106060 277753
rect 106902 277803 106966 277950
rect 107072 277803 107130 277950
rect 106902 277724 107130 277803
rect 109731 278985 109765 279015
rect 109731 278917 109765 278943
rect 109731 278849 109765 278871
rect 109731 278781 109765 278799
rect 109731 278713 109765 278727
rect 109731 278645 109765 278655
rect 109731 278577 109765 278583
rect 109731 278509 109765 278511
rect 109731 278473 109765 278475
rect 109731 278401 109765 278407
rect 109731 278329 109765 278339
rect 109731 278257 109765 278271
rect 109731 278185 109765 278203
rect 109731 278113 109765 278135
rect 109731 278041 109765 278067
rect 109731 277969 109765 277999
rect 110075 278985 110109 279015
rect 110075 278917 110109 278943
rect 110075 278849 110109 278871
rect 110075 278781 110109 278799
rect 110075 278713 110109 278727
rect 110075 278645 110109 278655
rect 110075 278577 110109 278583
rect 110075 278509 110109 278511
rect 110075 278473 110109 278475
rect 110075 278401 110109 278407
rect 110075 278329 110109 278339
rect 110075 278257 110109 278271
rect 110075 278185 110109 278203
rect 110075 278113 110109 278135
rect 110075 278041 110109 278067
rect 110075 277969 110109 277999
rect 110189 279003 110312 279037
rect 110223 278969 110312 279003
rect 110189 278935 110312 278969
rect 110223 278901 110312 278935
rect 110189 278867 110312 278901
rect 110223 278833 110312 278867
rect 110189 278799 110312 278833
rect 110223 278765 110312 278799
rect 110189 278731 110312 278765
rect 110223 278697 110312 278731
rect 110189 278663 110312 278697
rect 110223 278629 110312 278663
rect 110189 278595 110312 278629
rect 110223 278561 110312 278595
rect 110189 278527 110312 278561
rect 110223 278493 110312 278527
rect 110189 278459 110312 278493
rect 110223 278425 110312 278459
rect 110189 278391 110312 278425
rect 110223 278357 110312 278391
rect 110189 278323 110312 278357
rect 110223 278289 110312 278323
rect 110189 278255 110312 278289
rect 110223 278221 110312 278255
rect 110189 278187 110312 278221
rect 110223 278153 110312 278187
rect 110189 278119 110312 278153
rect 110223 278085 110312 278119
rect 110189 278051 110312 278085
rect 110223 278017 110312 278051
rect 110189 277983 110312 278017
rect 109617 277915 109651 277949
rect 110223 277949 110312 277983
rect 109777 277901 109795 277935
rect 109835 277901 109867 277935
rect 109903 277901 109937 277935
rect 109973 277901 110005 277935
rect 110045 277901 110063 277935
rect 110189 277915 110312 277949
rect 109617 277847 109651 277881
rect 110223 277881 110312 277915
rect 110189 277847 110312 277881
rect 109617 277779 109651 277813
rect 109777 277793 109795 277827
rect 109835 277793 109867 277827
rect 109903 277793 109937 277827
rect 109973 277793 110005 277827
rect 110045 277793 110063 277827
rect 110223 277813 110312 277847
rect 110189 277779 110312 277813
rect 105974 277685 106060 277719
rect 105974 277651 106000 277685
rect 106034 277651 106060 277685
rect 105974 277617 106060 277651
rect 105974 277583 106000 277617
rect 106034 277583 106060 277617
rect 105974 277549 106060 277583
rect 105974 277515 106000 277549
rect 106034 277515 106060 277549
rect 105974 277481 106060 277515
rect 105974 277447 106000 277481
rect 106034 277447 106060 277481
rect 105974 277413 106060 277447
rect 105974 277379 106000 277413
rect 106034 277379 106060 277413
rect 105974 277345 106060 277379
rect 105974 277311 106000 277345
rect 106034 277311 106060 277345
rect 109617 277711 109651 277745
rect 109617 277643 109651 277677
rect 109617 277575 109651 277609
rect 109617 277507 109651 277541
rect 109617 277439 109651 277473
rect 109617 277371 109651 277405
rect 105974 277277 106060 277311
rect 105974 277243 106000 277277
rect 106034 277243 106060 277277
rect 105974 277209 106060 277243
rect 105974 277175 106000 277209
rect 106034 277175 106060 277209
rect 105974 277141 106060 277175
rect 105974 277107 106000 277141
rect 106034 277107 106060 277141
rect 105974 277073 106060 277107
rect 105974 277039 106000 277073
rect 106034 277039 106060 277073
rect 105974 277005 106060 277039
rect 105974 276971 106000 277005
rect 106034 276971 106060 277005
rect 105974 276937 106060 276971
rect 105974 276903 106000 276937
rect 106034 276903 106060 276937
rect 106308 277290 106413 277324
rect 106447 277290 106481 277324
rect 106515 277290 106549 277324
rect 106583 277290 106617 277324
rect 106651 277290 106685 277324
rect 106719 277290 106753 277324
rect 106787 277290 106821 277324
rect 106855 277290 106889 277324
rect 106923 277290 106957 277324
rect 106991 277290 107025 277324
rect 107059 277290 107093 277324
rect 107127 277290 107161 277324
rect 107195 277290 107229 277324
rect 107263 277290 107297 277324
rect 107331 277290 107365 277324
rect 107399 277290 107433 277324
rect 107467 277290 107501 277324
rect 107535 277290 107569 277324
rect 107603 277290 107708 277324
rect 106308 277212 106342 277290
rect 107674 277212 107708 277290
rect 106308 277144 106342 277178
rect 106487 277176 106515 277210
rect 106557 277176 106583 277210
rect 106629 277176 106651 277210
rect 106701 277176 106719 277210
rect 106773 277176 106787 277210
rect 106845 277176 106855 277210
rect 106917 277176 106923 277210
rect 106989 277176 106991 277210
rect 107025 277176 107027 277210
rect 107093 277176 107099 277210
rect 107161 277176 107171 277210
rect 107229 277176 107243 277210
rect 107297 277176 107315 277210
rect 107365 277176 107387 277210
rect 107433 277176 107459 277210
rect 107501 277176 107529 277210
rect 106308 277076 106342 277110
rect 106410 277144 106444 277164
rect 106410 277090 106444 277110
rect 107572 277144 107606 277164
rect 107572 277090 107606 277110
rect 107674 277144 107708 277178
rect 106487 277044 106515 277078
rect 106557 277044 106583 277078
rect 106629 277044 106651 277078
rect 106701 277044 106719 277078
rect 106773 277044 106787 277078
rect 106845 277044 106855 277078
rect 106917 277044 106923 277078
rect 106989 277044 106991 277078
rect 107025 277044 107027 277078
rect 107093 277044 107099 277078
rect 107161 277044 107171 277078
rect 107229 277044 107243 277078
rect 107297 277044 107315 277078
rect 107365 277044 107387 277078
rect 107433 277044 107459 277078
rect 107501 277044 107529 277078
rect 107674 277076 107708 277110
rect 106308 276964 106342 277042
rect 106849 276964 107133 277044
rect 107674 276964 107708 277042
rect 106308 276930 106413 276964
rect 106447 276930 106481 276964
rect 106515 276930 106549 276964
rect 106583 276930 106617 276964
rect 106651 276930 106685 276964
rect 106719 276930 106753 276964
rect 106787 276930 106821 276964
rect 106855 276930 106889 276964
rect 106923 276930 106957 276964
rect 106991 276930 107025 276964
rect 107059 276930 107093 276964
rect 107127 276930 107161 276964
rect 107195 276930 107229 276964
rect 107263 276930 107297 276964
rect 107331 276930 107365 276964
rect 107399 276930 107433 276964
rect 107467 276930 107501 276964
rect 107535 276930 107569 276964
rect 107603 276930 107708 276964
rect 109617 277303 109651 277337
rect 109617 277235 109651 277269
rect 109617 277167 109651 277201
rect 109617 277099 109651 277133
rect 109617 277031 109651 277065
rect 109617 276963 109651 276997
rect 105974 276869 106060 276903
rect 105974 276835 106000 276869
rect 106034 276835 106060 276869
rect 105974 276801 106060 276835
rect 105974 276767 106000 276801
rect 106034 276767 106060 276801
rect 105974 276733 106060 276767
rect 105974 276699 106000 276733
rect 106034 276699 106060 276733
rect 105974 276665 106060 276699
rect 105974 276631 106000 276665
rect 106034 276631 106060 276665
rect 105974 276597 106060 276631
rect 105974 276563 106000 276597
rect 106034 276563 106060 276597
rect 105974 276529 106060 276563
rect 105974 276495 106000 276529
rect 106034 276495 106060 276529
rect 105974 276461 106060 276495
rect 105974 276427 106000 276461
rect 106034 276427 106060 276461
rect 105974 276393 106060 276427
rect 106719 276403 106985 276930
rect 109617 276895 109651 276929
rect 109617 276827 109651 276861
rect 109617 276759 109651 276793
rect 109617 276691 109651 276725
rect 109731 277729 109765 277759
rect 109731 277661 109765 277687
rect 109731 277593 109765 277615
rect 109731 277525 109765 277543
rect 109731 277457 109765 277471
rect 109731 277389 109765 277399
rect 109731 277321 109765 277327
rect 109731 277253 109765 277255
rect 109731 277217 109765 277219
rect 109731 277145 109765 277151
rect 109731 277073 109765 277083
rect 109731 277001 109765 277015
rect 109731 276929 109765 276947
rect 109731 276857 109765 276879
rect 109731 276785 109765 276811
rect 109731 276713 109765 276743
rect 110075 277729 110109 277759
rect 110075 277661 110109 277687
rect 110075 277593 110109 277615
rect 110075 277525 110109 277543
rect 110075 277457 110109 277471
rect 110075 277389 110109 277399
rect 110075 277321 110109 277327
rect 110075 277253 110109 277255
rect 110075 277217 110109 277219
rect 110075 277145 110109 277151
rect 110075 277073 110109 277083
rect 110075 277001 110109 277015
rect 110075 276929 110109 276947
rect 110075 276857 110109 276879
rect 110075 276785 110109 276811
rect 110075 276713 110109 276743
rect 110223 277745 110312 277779
rect 110189 277711 110312 277745
rect 110223 277677 110312 277711
rect 110189 277643 110312 277677
rect 110223 277609 110312 277643
rect 110189 277575 110312 277609
rect 110223 277541 110312 277575
rect 110189 277507 110312 277541
rect 110223 277473 110312 277507
rect 110189 277439 110312 277473
rect 110223 277405 110312 277439
rect 110189 277371 110312 277405
rect 110223 277337 110312 277371
rect 110189 277303 110312 277337
rect 110223 277269 110312 277303
rect 110189 277235 110312 277269
rect 110223 277201 110312 277235
rect 110189 277167 110312 277201
rect 110223 277133 110312 277167
rect 110189 277099 110312 277133
rect 110223 277065 110312 277099
rect 110189 277031 110312 277065
rect 110223 276997 110312 277031
rect 110189 276963 110312 276997
rect 110223 276929 110312 276963
rect 110189 276895 110312 276929
rect 110223 276861 110312 276895
rect 110189 276827 110312 276861
rect 110223 276793 110312 276827
rect 110189 276759 110312 276793
rect 110223 276725 110312 276759
rect 110189 276691 110312 276725
rect 109617 276577 109651 276657
rect 109777 276645 109795 276679
rect 109835 276645 109867 276679
rect 109903 276645 109937 276679
rect 109973 276645 110005 276679
rect 110045 276645 110063 276679
rect 110223 276657 110312 276691
rect 110189 276577 110312 276657
rect 109617 276543 109733 276577
rect 109767 276543 109801 276577
rect 109835 276543 109869 276577
rect 109903 276543 109937 276577
rect 109971 276543 110005 276577
rect 110039 276543 110073 276577
rect 110107 276553 110312 276577
rect 110107 276543 110224 276553
rect 105974 276359 106000 276393
rect 106034 276359 106060 276393
rect 105974 276325 106060 276359
rect 105974 276291 106000 276325
rect 106034 276291 106060 276325
rect 105974 276257 106060 276291
rect 105974 276223 106000 276257
rect 106034 276223 106060 276257
rect 105974 276189 106060 276223
rect 105974 276155 106000 276189
rect 106034 276155 106060 276189
rect 105974 276121 106060 276155
rect 105974 276087 106000 276121
rect 106034 276087 106060 276121
rect 105974 276053 106060 276087
rect 105974 276019 106000 276053
rect 106034 276019 106060 276053
rect 105974 275985 106060 276019
rect 105974 275951 106000 275985
rect 106034 275951 106060 275985
rect 105974 275917 106060 275951
rect 105974 275883 106000 275917
rect 106034 275883 106060 275917
rect 105974 275849 106060 275883
rect 105974 275815 106000 275849
rect 106034 275815 106060 275849
rect 105974 275781 106060 275815
rect 105974 275747 106000 275781
rect 106034 275747 106060 275781
rect 105974 275713 106060 275747
rect 105974 275679 106000 275713
rect 106034 275679 106060 275713
rect 105974 275645 106060 275679
rect 105974 275611 106000 275645
rect 106034 275611 106060 275645
rect 105974 275577 106060 275611
rect 105974 275543 106000 275577
rect 106034 275543 106060 275577
rect 105974 275509 106060 275543
rect 105974 275475 106000 275509
rect 106034 275475 106060 275509
rect 105974 275441 106060 275475
rect 105974 275407 106000 275441
rect 106034 275407 106060 275441
rect 105974 275373 106060 275407
rect 105974 275339 106000 275373
rect 106034 275339 106060 275373
rect 105974 275305 106060 275339
rect 105974 275271 106000 275305
rect 106034 275271 106060 275305
rect 105974 275237 106060 275271
rect 105974 275203 106000 275237
rect 106034 275203 106060 275237
rect 105974 275169 106060 275203
rect 105974 275135 106000 275169
rect 106034 275135 106060 275169
rect 105974 275101 106060 275135
rect 105974 275067 106000 275101
rect 106034 275067 106060 275101
rect 105974 275033 106060 275067
rect 105974 274999 106000 275033
rect 106034 274999 106060 275033
rect 105974 274965 106060 274999
rect 105974 274931 106000 274965
rect 106034 274931 106060 274965
rect 105974 274897 106060 274931
rect 105974 274863 106000 274897
rect 106034 274863 106060 274897
rect 105974 274829 106060 274863
rect 105974 274795 106000 274829
rect 106034 274795 106060 274829
rect 105974 274761 106060 274795
rect 105974 274727 106000 274761
rect 106034 274727 106060 274761
rect 106294 276272 106985 276403
rect 106294 274870 106409 276272
rect 106515 275934 106985 276272
rect 110145 276025 110224 276543
rect 110145 275991 110167 276025
rect 110201 275991 110224 276025
rect 110145 275957 110224 275991
rect 106515 275900 106797 275934
rect 106831 275900 106865 275934
rect 106899 275900 106933 275934
rect 106967 275900 107001 275934
rect 107035 275900 107069 275934
rect 107103 275900 107137 275934
rect 107171 275900 107205 275934
rect 107239 275900 107273 275934
rect 107307 275900 107341 275934
rect 107375 275900 107409 275934
rect 107443 275900 107477 275934
rect 107511 275900 107545 275934
rect 107579 275900 107613 275934
rect 107647 275900 107681 275934
rect 107715 275900 107749 275934
rect 107783 275900 107817 275934
rect 107851 275900 107885 275934
rect 107919 275900 107953 275934
rect 107987 275900 108021 275934
rect 108055 275900 108089 275934
rect 108123 275900 108157 275934
rect 108191 275900 108225 275934
rect 108259 275900 108293 275934
rect 108327 275900 108361 275934
rect 108395 275900 108429 275934
rect 108463 275900 108497 275934
rect 108531 275900 108565 275934
rect 108599 275900 108633 275934
rect 108667 275900 108701 275934
rect 108735 275900 108769 275934
rect 108803 275900 108837 275934
rect 108871 275900 108905 275934
rect 108939 275900 108973 275934
rect 109007 275900 109041 275934
rect 109075 275900 109109 275934
rect 109143 275900 109177 275934
rect 109211 275900 109245 275934
rect 109279 275900 109313 275934
rect 109347 275900 109381 275934
rect 109415 275900 109449 275934
rect 109483 275900 109517 275934
rect 109551 275900 109585 275934
rect 109619 275900 109653 275934
rect 109687 275900 109721 275934
rect 109755 275900 109847 275934
rect 106515 275850 106887 275900
rect 106515 275816 106706 275850
rect 106740 275816 106887 275850
rect 106515 275782 106887 275816
rect 106515 275748 106706 275782
rect 106740 275748 106887 275782
rect 106995 275759 107075 275900
rect 109498 275759 109578 275900
rect 109693 275850 109847 275900
rect 109693 275816 109813 275850
rect 109693 275782 109847 275816
rect 106515 275714 106887 275748
rect 106947 275725 106987 275759
rect 107023 275725 107057 275759
rect 107093 275725 107133 275759
rect 107447 275725 107487 275759
rect 107523 275725 107557 275759
rect 107593 275725 107633 275759
rect 107947 275725 107987 275759
rect 108023 275725 108057 275759
rect 108093 275725 108133 275759
rect 108447 275725 108487 275759
rect 108523 275725 108557 275759
rect 108593 275725 108633 275759
rect 108947 275725 108987 275759
rect 109023 275725 109057 275759
rect 109093 275725 109133 275759
rect 109447 275725 109487 275759
rect 109523 275725 109557 275759
rect 109593 275725 109633 275759
rect 109693 275748 109813 275782
rect 106515 275680 106706 275714
rect 106740 275713 106887 275714
rect 109693 275714 109847 275748
rect 109693 275713 109813 275714
rect 106740 275681 106904 275713
rect 106740 275680 106870 275681
rect 106515 275646 106870 275680
rect 106515 275612 106706 275646
rect 106740 275631 106870 275646
rect 106740 275613 106904 275631
rect 106740 275612 106870 275613
rect 106515 275578 106870 275612
rect 106515 275544 106706 275578
rect 106740 275559 106870 275578
rect 106740 275545 106904 275559
rect 106740 275544 106870 275545
rect 106515 275510 106870 275544
rect 106515 275476 106706 275510
rect 106740 275487 106870 275510
rect 106740 275477 106904 275487
rect 106740 275476 106870 275477
rect 106515 275442 106870 275476
rect 106515 275408 106706 275442
rect 106740 275415 106870 275442
rect 106740 275409 106904 275415
rect 106740 275408 106870 275409
rect 106515 275374 106870 275408
rect 106515 275340 106706 275374
rect 106740 275343 106870 275374
rect 106740 275341 106904 275343
rect 106740 275340 106870 275341
rect 106515 275307 106870 275340
rect 106515 275306 106904 275307
rect 106515 275272 106706 275306
rect 106740 275305 106904 275306
rect 106740 275272 106870 275305
rect 106515 275239 106870 275272
rect 106515 275238 106904 275239
rect 106515 275204 106706 275238
rect 106740 275233 106904 275238
rect 106740 275204 106870 275233
rect 106515 275171 106870 275204
rect 106515 275170 106904 275171
rect 106515 275136 106706 275170
rect 106740 275161 106904 275170
rect 106740 275136 106870 275161
rect 106515 275103 106870 275136
rect 106515 275102 106904 275103
rect 106515 275068 106706 275102
rect 106740 275089 106904 275102
rect 106740 275068 106870 275089
rect 106515 275035 106870 275068
rect 106515 275034 106904 275035
rect 106515 275000 106706 275034
rect 106740 275017 106904 275034
rect 106740 275000 106870 275017
rect 106515 274967 106870 275000
rect 106515 274966 106904 274967
rect 106515 274932 106706 274966
rect 106740 274935 106904 274966
rect 107176 275681 107210 275713
rect 107176 275613 107210 275631
rect 107176 275545 107210 275559
rect 107176 275477 107210 275487
rect 107176 275409 107210 275415
rect 107176 275341 107210 275343
rect 107176 275305 107210 275307
rect 107176 275233 107210 275239
rect 107176 275161 107210 275171
rect 107176 275089 107210 275103
rect 107176 275017 107210 275035
rect 107176 274935 107210 274967
rect 107370 275681 107404 275713
rect 107370 275613 107404 275631
rect 107370 275545 107404 275559
rect 107370 275477 107404 275487
rect 107370 275409 107404 275415
rect 107370 275341 107404 275343
rect 107370 275305 107404 275307
rect 107370 275233 107404 275239
rect 107370 275161 107404 275171
rect 107370 275089 107404 275103
rect 107370 275017 107404 275035
rect 107370 274935 107404 274967
rect 107676 275681 107710 275713
rect 107676 275613 107710 275631
rect 107676 275545 107710 275559
rect 107676 275477 107710 275487
rect 107676 275409 107710 275415
rect 107676 275341 107710 275343
rect 107676 275305 107710 275307
rect 107676 275233 107710 275239
rect 107676 275161 107710 275171
rect 107676 275089 107710 275103
rect 107676 275017 107710 275035
rect 107676 274935 107710 274967
rect 107870 275681 107904 275713
rect 107870 275613 107904 275631
rect 107870 275545 107904 275559
rect 107870 275477 107904 275487
rect 107870 275409 107904 275415
rect 107870 275341 107904 275343
rect 107870 275305 107904 275307
rect 107870 275233 107904 275239
rect 107870 275161 107904 275171
rect 107870 275089 107904 275103
rect 107870 275017 107904 275035
rect 107870 274935 107904 274967
rect 108176 275681 108210 275713
rect 108176 275613 108210 275631
rect 108176 275545 108210 275559
rect 108176 275477 108210 275487
rect 108176 275409 108210 275415
rect 108176 275341 108210 275343
rect 108176 275305 108210 275307
rect 108176 275233 108210 275239
rect 108176 275161 108210 275171
rect 108176 275089 108210 275103
rect 108176 275017 108210 275035
rect 108176 274935 108210 274967
rect 108370 275681 108404 275713
rect 108370 275613 108404 275631
rect 108370 275545 108404 275559
rect 108370 275477 108404 275487
rect 108370 275409 108404 275415
rect 108370 275341 108404 275343
rect 108370 275305 108404 275307
rect 108370 275233 108404 275239
rect 108370 275161 108404 275171
rect 108370 275089 108404 275103
rect 108370 275017 108404 275035
rect 108370 274935 108404 274967
rect 108676 275681 108710 275713
rect 108676 275613 108710 275631
rect 108676 275545 108710 275559
rect 108676 275477 108710 275487
rect 108676 275409 108710 275415
rect 108676 275341 108710 275343
rect 108676 275305 108710 275307
rect 108676 275233 108710 275239
rect 108676 275161 108710 275171
rect 108676 275089 108710 275103
rect 108676 275017 108710 275035
rect 108676 274935 108710 274967
rect 108870 275681 108904 275713
rect 108870 275613 108904 275631
rect 108870 275545 108904 275559
rect 108870 275477 108904 275487
rect 108870 275409 108904 275415
rect 108870 275341 108904 275343
rect 108870 275305 108904 275307
rect 108870 275233 108904 275239
rect 108870 275161 108904 275171
rect 108870 275089 108904 275103
rect 108870 275017 108904 275035
rect 108870 274935 108904 274967
rect 109176 275681 109210 275713
rect 109176 275613 109210 275631
rect 109176 275545 109210 275559
rect 109176 275477 109210 275487
rect 109176 275409 109210 275415
rect 109176 275341 109210 275343
rect 109176 275305 109210 275307
rect 109176 275233 109210 275239
rect 109176 275161 109210 275171
rect 109176 275089 109210 275103
rect 109176 275017 109210 275035
rect 109176 274935 109210 274967
rect 109370 275681 109404 275713
rect 109370 275613 109404 275631
rect 109370 275545 109404 275559
rect 109370 275477 109404 275487
rect 109370 275409 109404 275415
rect 109370 275341 109404 275343
rect 109370 275305 109404 275307
rect 109370 275233 109404 275239
rect 109370 275161 109404 275171
rect 109370 275089 109404 275103
rect 109370 275017 109404 275035
rect 109370 274935 109404 274967
rect 109676 275681 109813 275713
rect 109710 275680 109813 275681
rect 109710 275646 109847 275680
rect 109710 275631 109813 275646
rect 109676 275613 109813 275631
rect 109710 275612 109813 275613
rect 109710 275578 109847 275612
rect 109710 275559 109813 275578
rect 109676 275545 109813 275559
rect 109710 275544 109813 275545
rect 109710 275510 109847 275544
rect 109710 275487 109813 275510
rect 109676 275477 109813 275487
rect 109710 275476 109813 275477
rect 109710 275442 109847 275476
rect 109710 275415 109813 275442
rect 109676 275409 109813 275415
rect 109710 275408 109813 275409
rect 109710 275374 109847 275408
rect 109710 275343 109813 275374
rect 109676 275341 109813 275343
rect 109710 275340 109813 275341
rect 109710 275307 109847 275340
rect 109676 275306 109847 275307
rect 109676 275305 109813 275306
rect 109710 275272 109813 275305
rect 109710 275239 109847 275272
rect 109676 275238 109847 275239
rect 109676 275233 109813 275238
rect 109710 275204 109813 275233
rect 109710 275171 109847 275204
rect 109676 275170 109847 275171
rect 109676 275161 109813 275170
rect 109710 275136 109813 275161
rect 109710 275103 109847 275136
rect 109676 275102 109847 275103
rect 109676 275089 109813 275102
rect 109710 275068 109813 275089
rect 109710 275035 109847 275068
rect 109676 275034 109847 275035
rect 109676 275017 109813 275034
rect 109710 275000 109813 275017
rect 109710 274967 109847 275000
rect 109676 274966 109847 274967
rect 109676 274935 109813 274966
rect 106740 274932 106891 274935
rect 106515 274898 106891 274932
rect 109692 274932 109813 274935
rect 106515 274870 106706 274898
rect 106294 274864 106706 274870
rect 106740 274886 106891 274898
rect 106947 274889 106987 274923
rect 107023 274889 107057 274923
rect 107093 274889 107133 274923
rect 107447 274889 107487 274923
rect 107523 274889 107557 274923
rect 107593 274889 107633 274923
rect 107947 274889 107987 274923
rect 108023 274889 108057 274923
rect 108093 274889 108133 274923
rect 108447 274889 108487 274923
rect 108523 274889 108557 274923
rect 108593 274889 108633 274923
rect 108947 274889 108987 274923
rect 109023 274889 109057 274923
rect 109093 274889 109133 274923
rect 109447 274889 109487 274923
rect 109523 274889 109557 274923
rect 109593 274889 109633 274923
rect 106947 274886 109633 274889
rect 106740 274882 109633 274886
rect 109692 274898 109847 274932
rect 109692 274882 109813 274898
rect 106740 274864 109813 274882
rect 106294 274830 109847 274864
rect 106294 274796 106706 274830
rect 106740 274796 109813 274830
rect 106294 274747 109847 274796
rect 106294 274731 106797 274747
rect 105974 274693 106060 274727
rect 106706 274713 106797 274731
rect 106831 274713 106865 274747
rect 106899 274713 106933 274747
rect 106967 274713 107001 274747
rect 107035 274713 107069 274747
rect 107103 274713 107137 274747
rect 107171 274713 107205 274747
rect 107239 274713 107273 274747
rect 107307 274713 107341 274747
rect 107375 274713 107409 274747
rect 107443 274713 107477 274747
rect 107511 274713 107545 274747
rect 107579 274713 107613 274747
rect 107647 274713 107681 274747
rect 107715 274713 107749 274747
rect 107783 274713 107817 274747
rect 107851 274713 107885 274747
rect 107919 274713 107953 274747
rect 107987 274713 108021 274747
rect 108055 274713 108089 274747
rect 108123 274713 108157 274747
rect 108191 274713 108225 274747
rect 108259 274713 108293 274747
rect 108327 274713 108361 274747
rect 108395 274713 108429 274747
rect 108463 274713 108497 274747
rect 108531 274713 108565 274747
rect 108599 274713 108633 274747
rect 108667 274713 108701 274747
rect 108735 274713 108769 274747
rect 108803 274713 108837 274747
rect 108871 274713 108905 274747
rect 108939 274713 108973 274747
rect 109007 274713 109041 274747
rect 109075 274713 109109 274747
rect 109143 274713 109177 274747
rect 109211 274713 109245 274747
rect 109279 274713 109313 274747
rect 109347 274713 109381 274747
rect 109415 274713 109449 274747
rect 109483 274713 109517 274747
rect 109551 274713 109585 274747
rect 109619 274713 109653 274747
rect 109687 274713 109721 274747
rect 109755 274713 109847 274747
rect 110145 275923 110167 275957
rect 110201 275923 110224 275957
rect 110145 275889 110224 275923
rect 110145 275855 110167 275889
rect 110201 275855 110224 275889
rect 110145 275821 110224 275855
rect 110145 275787 110167 275821
rect 110201 275787 110224 275821
rect 110145 275753 110224 275787
rect 110145 275719 110167 275753
rect 110201 275719 110224 275753
rect 110145 275685 110224 275719
rect 110145 275651 110167 275685
rect 110201 275651 110224 275685
rect 110145 275617 110224 275651
rect 110145 275583 110167 275617
rect 110201 275583 110224 275617
rect 110145 275549 110224 275583
rect 110145 275515 110167 275549
rect 110201 275515 110224 275549
rect 110145 275481 110224 275515
rect 110145 275447 110167 275481
rect 110201 275447 110224 275481
rect 110145 275413 110224 275447
rect 110145 275379 110167 275413
rect 110201 275379 110224 275413
rect 110145 275345 110224 275379
rect 110145 275311 110167 275345
rect 110201 275311 110224 275345
rect 110145 275277 110224 275311
rect 110145 275243 110167 275277
rect 110201 275243 110224 275277
rect 110145 275209 110224 275243
rect 110145 275175 110167 275209
rect 110201 275175 110224 275209
rect 110145 275141 110224 275175
rect 110145 275107 110167 275141
rect 110201 275107 110224 275141
rect 110145 275073 110224 275107
rect 110145 275039 110167 275073
rect 110201 275039 110224 275073
rect 110145 275005 110224 275039
rect 110145 274971 110167 275005
rect 110201 274971 110224 275005
rect 110145 274937 110224 274971
rect 110145 274903 110167 274937
rect 110201 274903 110224 274937
rect 110145 274869 110224 274903
rect 110145 274835 110167 274869
rect 110201 274835 110224 274869
rect 110145 274801 110224 274835
rect 110145 274767 110167 274801
rect 110201 274767 110224 274801
rect 110145 274733 110224 274767
rect 105974 274659 106000 274693
rect 106034 274659 106060 274693
rect 105974 274619 106060 274659
rect 110145 274699 110167 274733
rect 110201 274699 110224 274733
rect 110145 274619 110224 274699
rect 105974 274590 110224 274619
rect 105974 274556 106117 274590
rect 106151 274556 106185 274590
rect 106219 274556 106253 274590
rect 106287 274556 106321 274590
rect 106355 274556 106389 274590
rect 106423 274556 106457 274590
rect 106491 274556 106525 274590
rect 106559 274556 106593 274590
rect 106627 274556 106661 274590
rect 106695 274556 106729 274590
rect 106763 274556 106797 274590
rect 106831 274556 106865 274590
rect 106899 274556 106933 274590
rect 106967 274556 107001 274590
rect 107035 274556 107069 274590
rect 107103 274556 107137 274590
rect 107171 274556 107205 274590
rect 107239 274556 107273 274590
rect 107307 274556 107341 274590
rect 107375 274556 107409 274590
rect 107443 274556 107477 274590
rect 107511 274556 107545 274590
rect 107579 274556 107613 274590
rect 107647 274556 107681 274590
rect 107715 274556 107749 274590
rect 107783 274556 107817 274590
rect 107851 274556 107885 274590
rect 107919 274556 107953 274590
rect 107987 274556 108021 274590
rect 108055 274556 108089 274590
rect 108123 274556 108157 274590
rect 108191 274556 108225 274590
rect 108259 274556 108293 274590
rect 108327 274556 108361 274590
rect 108395 274556 108429 274590
rect 108463 274556 108497 274590
rect 108531 274556 108565 274590
rect 108599 274556 108633 274590
rect 108667 274556 108701 274590
rect 108735 274556 108769 274590
rect 108803 274556 108837 274590
rect 108871 274556 108905 274590
rect 108939 274556 108973 274590
rect 109007 274556 109041 274590
rect 109075 274556 109109 274590
rect 109143 274556 109177 274590
rect 109211 274556 109245 274590
rect 109279 274556 109313 274590
rect 109347 274556 109381 274590
rect 109415 274556 109449 274590
rect 109483 274556 109517 274590
rect 109551 274556 109585 274590
rect 109619 274556 109653 274590
rect 109687 274556 109721 274590
rect 109755 274556 109789 274590
rect 109823 274556 109857 274590
rect 109891 274556 109925 274590
rect 109959 274556 109993 274590
rect 110027 274556 110061 274590
rect 110095 274556 110129 274590
rect 110163 274556 110224 274590
rect 105974 274527 110224 274556
rect 106281 272923 110259 272951
rect 106281 272898 106595 272923
rect 106281 270212 106285 272898
rect 106455 272821 106595 272898
rect 109961 272898 110259 272923
rect 109961 272821 110085 272898
rect 106455 272786 110085 272821
rect 106455 270334 106459 272786
rect 107343 272367 108250 272786
rect 109088 272568 109151 272602
rect 109185 272568 109219 272602
rect 109253 272568 109287 272602
rect 109321 272568 109355 272602
rect 109389 272568 109423 272602
rect 109457 272568 109491 272602
rect 109525 272568 109559 272602
rect 109593 272568 109627 272602
rect 109661 272568 109695 272602
rect 109729 272568 109763 272602
rect 109797 272568 109861 272602
rect 109088 272530 109122 272568
rect 109827 272530 109861 272568
rect 109088 272462 109122 272496
rect 109088 272394 109122 272428
rect 106715 272350 108803 272367
rect 106715 272321 106848 272350
rect 106715 272287 106735 272321
rect 106769 272316 106848 272321
rect 106882 272316 106977 272350
rect 107011 272316 107045 272350
rect 107079 272316 107113 272350
rect 107147 272316 107181 272350
rect 107215 272316 107249 272350
rect 107283 272316 107317 272350
rect 107351 272316 107385 272350
rect 107419 272316 107453 272350
rect 107487 272316 107521 272350
rect 107555 272316 107589 272350
rect 107623 272316 107657 272350
rect 107691 272316 107725 272350
rect 107759 272316 107793 272350
rect 107827 272316 107861 272350
rect 107895 272316 107929 272350
rect 107963 272316 107997 272350
rect 108031 272316 108065 272350
rect 108099 272316 108133 272350
rect 108167 272316 108201 272350
rect 108235 272316 108269 272350
rect 108303 272316 108337 272350
rect 108371 272316 108405 272350
rect 108439 272316 108473 272350
rect 108507 272316 108541 272350
rect 108575 272316 108609 272350
rect 108643 272321 108803 272350
rect 108643 272316 108749 272321
rect 106769 272299 108749 272316
rect 106769 272287 106789 272299
rect 106715 272253 106789 272287
rect 106715 272219 106735 272253
rect 106769 272219 106789 272253
rect 106715 272185 106789 272219
rect 106715 272151 106735 272185
rect 106769 272151 106789 272185
rect 108729 272287 108749 272299
rect 108783 272287 108803 272321
rect 108729 272253 108803 272287
rect 108729 272219 108749 272253
rect 108783 272219 108803 272253
rect 108729 272185 108803 272219
rect 108729 272151 108749 272185
rect 108783 272151 108803 272185
rect 106715 272117 106789 272151
rect 107459 272117 107480 272151
rect 107534 272117 107548 272151
rect 107606 272117 107616 272151
rect 107678 272117 107684 272151
rect 107750 272117 107752 272151
rect 107786 272117 107788 272151
rect 107854 272117 107860 272151
rect 107922 272117 107932 272151
rect 107990 272117 108004 272151
rect 108058 272117 108079 272151
rect 108729 272117 108803 272151
rect 106715 272083 106735 272117
rect 106769 272083 106789 272117
rect 108729 272083 108749 272117
rect 108783 272083 108803 272117
rect 106715 272049 106789 272083
rect 106715 272015 106735 272049
rect 106769 272015 106789 272049
rect 107413 272060 107447 272083
rect 106715 271981 106789 272015
rect 106981 272009 106997 272043
rect 107035 272009 107069 272043
rect 107103 272009 107137 272043
rect 107175 272009 107191 272043
rect 106715 271947 106735 271981
rect 106769 271975 106789 271981
rect 107413 271992 107447 271998
rect 106769 271947 106969 271975
rect 106715 271942 106969 271947
rect 106715 271913 106935 271942
rect 106715 271879 106735 271913
rect 106769 271906 106935 271913
rect 106769 271879 106969 271906
rect 106715 271872 106969 271879
rect 106715 271845 106935 271872
rect 106715 271811 106735 271845
rect 106769 271836 106935 271845
rect 106769 271811 106969 271836
rect 106715 271803 106969 271811
rect 107203 271942 107237 271975
rect 107203 271872 107237 271906
rect 107203 271803 107237 271836
rect 107413 271924 107447 271926
rect 107413 271888 107447 271890
rect 107413 271816 107447 271822
rect 106715 271777 106789 271803
rect 106715 271743 106735 271777
rect 106769 271743 106789 271777
rect 106715 271709 106789 271743
rect 106981 271735 106997 271769
rect 107035 271735 107069 271769
rect 107103 271735 107137 271769
rect 107175 271735 107191 271769
rect 107413 271731 107447 271754
rect 108091 272060 108125 272083
rect 108091 271992 108125 271998
rect 108091 271924 108125 271926
rect 108091 271888 108125 271890
rect 108091 271816 108125 271822
rect 108091 271731 108125 271754
rect 108729 272049 108803 272083
rect 108729 272015 108749 272049
rect 108783 272015 108803 272049
rect 108729 271981 108803 272015
rect 108729 271947 108749 271981
rect 108783 271947 108803 271981
rect 108729 271913 108803 271947
rect 108729 271879 108749 271913
rect 108783 271879 108803 271913
rect 108729 271845 108803 271879
rect 108729 271811 108749 271845
rect 108783 271811 108803 271845
rect 108729 271777 108803 271811
rect 108729 271743 108749 271777
rect 108783 271743 108803 271777
rect 106715 271675 106735 271709
rect 106769 271675 106789 271709
rect 108729 271709 108803 271743
rect 106715 271641 106789 271675
rect 107459 271663 107480 271697
rect 107534 271663 107548 271697
rect 107606 271663 107616 271697
rect 107678 271663 107684 271697
rect 107750 271663 107752 271697
rect 107786 271663 107788 271697
rect 107854 271663 107860 271697
rect 107922 271663 107932 271697
rect 107990 271663 108004 271697
rect 108058 271663 108079 271697
rect 108729 271675 108749 271709
rect 108783 271675 108803 271709
rect 106715 271607 106735 271641
rect 106769 271607 106789 271641
rect 106715 271573 106789 271607
rect 106715 271539 106735 271573
rect 106769 271539 106789 271573
rect 106715 271505 106789 271539
rect 108729 271641 108803 271675
rect 108729 271607 108749 271641
rect 108783 271607 108803 271641
rect 108729 271573 108803 271607
rect 108729 271539 108749 271573
rect 108783 271539 108803 271573
rect 106715 271471 106735 271505
rect 106769 271471 106789 271505
rect 107169 271501 107212 271535
rect 107250 271501 107280 271535
rect 107322 271501 107348 271535
rect 107394 271501 107416 271535
rect 107466 271501 107484 271535
rect 107538 271501 107552 271535
rect 107610 271501 107620 271535
rect 107682 271501 107688 271535
rect 107754 271501 107756 271535
rect 107790 271501 107792 271535
rect 107858 271501 107864 271535
rect 107926 271501 107936 271535
rect 107994 271501 108008 271535
rect 108062 271501 108080 271535
rect 108130 271501 108152 271535
rect 108198 271501 108224 271535
rect 108266 271501 108296 271535
rect 108334 271501 108377 271535
rect 108729 271505 108803 271539
rect 106715 271437 106789 271471
rect 106715 271403 106735 271437
rect 106769 271403 106789 271437
rect 106715 271369 106789 271403
rect 106715 271335 106735 271369
rect 106769 271335 106789 271369
rect 106715 271301 106789 271335
rect 107101 271453 107135 271489
rect 107101 271383 107135 271417
rect 107101 271311 107135 271347
rect 108411 271453 108445 271489
rect 108411 271383 108445 271417
rect 108411 271311 108445 271347
rect 108729 271471 108749 271505
rect 108783 271471 108803 271505
rect 108729 271437 108803 271471
rect 108729 271403 108749 271437
rect 108783 271403 108803 271437
rect 108729 271369 108803 271403
rect 108729 271335 108749 271369
rect 108783 271335 108803 271369
rect 106715 271267 106735 271301
rect 106769 271267 106789 271301
rect 108729 271301 108803 271335
rect 106715 271233 106789 271267
rect 107169 271265 107212 271299
rect 107250 271265 107280 271299
rect 107322 271265 107348 271299
rect 107394 271265 107416 271299
rect 107466 271265 107484 271299
rect 107538 271265 107552 271299
rect 107610 271265 107620 271299
rect 107682 271265 107688 271299
rect 107754 271265 107756 271299
rect 107790 271265 107792 271299
rect 107858 271265 107864 271299
rect 107926 271265 107936 271299
rect 107994 271265 108008 271299
rect 108062 271265 108080 271299
rect 108130 271265 108152 271299
rect 108198 271265 108224 271299
rect 108266 271265 108296 271299
rect 108334 271265 108377 271299
rect 108729 271267 108749 271301
rect 108783 271267 108803 271301
rect 106715 271199 106735 271233
rect 106769 271199 106789 271233
rect 106715 271165 106789 271199
rect 108729 271233 108803 271267
rect 108729 271199 108749 271233
rect 108783 271199 108803 271233
rect 108729 271165 108803 271199
rect 106715 271131 106735 271165
rect 106769 271131 106789 271165
rect 107169 271131 107212 271165
rect 107250 271131 107280 271165
rect 107322 271131 107348 271165
rect 107394 271131 107416 271165
rect 107466 271131 107484 271165
rect 107538 271131 107552 271165
rect 107610 271131 107620 271165
rect 107682 271131 107688 271165
rect 107754 271131 107756 271165
rect 107790 271131 107792 271165
rect 107858 271131 107864 271165
rect 107926 271131 107936 271165
rect 107994 271131 108008 271165
rect 108062 271131 108080 271165
rect 108130 271131 108152 271165
rect 108198 271131 108224 271165
rect 108266 271131 108296 271165
rect 108334 271131 108377 271165
rect 108729 271131 108749 271165
rect 108783 271131 108803 271165
rect 106715 271097 106789 271131
rect 106715 271063 106735 271097
rect 106769 271063 106789 271097
rect 106715 271029 106789 271063
rect 106715 270995 106735 271029
rect 106769 270995 106789 271029
rect 106715 270961 106789 270995
rect 106715 270927 106735 270961
rect 106769 270927 106789 270961
rect 107101 271083 107135 271119
rect 107101 271013 107135 271047
rect 107101 270941 107135 270977
rect 108411 271083 108445 271119
rect 108411 271013 108445 271047
rect 108411 270941 108445 270977
rect 108729 271097 108803 271131
rect 108729 271063 108749 271097
rect 108783 271063 108803 271097
rect 108729 271029 108803 271063
rect 109088 272326 109122 272360
rect 109088 272258 109122 272292
rect 109088 272190 109122 272224
rect 109088 272122 109122 272156
rect 109088 272054 109122 272088
rect 109088 271986 109122 272020
rect 109088 271918 109122 271952
rect 109088 271850 109122 271884
rect 109088 271782 109122 271816
rect 109088 271714 109122 271748
rect 109088 271646 109122 271680
rect 109088 271578 109122 271612
rect 109088 271510 109122 271544
rect 109088 271442 109122 271476
rect 109088 271374 109122 271408
rect 109088 271306 109122 271340
rect 109088 271238 109122 271272
rect 109088 271170 109122 271204
rect 109088 271102 109122 271136
rect 109088 271034 109122 271068
rect 108729 270995 108749 271029
rect 108783 270995 108803 271029
rect 108729 270961 108803 270995
rect 106715 270893 106789 270927
rect 107169 270895 107212 270929
rect 107250 270895 107280 270929
rect 107322 270895 107348 270929
rect 107394 270895 107416 270929
rect 107466 270895 107484 270929
rect 107538 270895 107552 270929
rect 107610 270895 107620 270929
rect 107682 270895 107688 270929
rect 107754 270895 107756 270929
rect 107790 270895 107792 270929
rect 107858 270895 107864 270929
rect 107926 270895 107936 270929
rect 107994 270895 108008 270929
rect 108062 270895 108080 270929
rect 108130 270895 108152 270929
rect 108198 270895 108224 270929
rect 108266 270895 108296 270929
rect 108334 270895 108377 270929
rect 108729 270927 108749 270961
rect 108783 270927 108803 270961
rect 106715 270859 106735 270893
rect 106769 270859 106789 270893
rect 106715 270825 106789 270859
rect 106715 270791 106735 270825
rect 106769 270801 106789 270825
rect 108729 270893 108803 270927
rect 108729 270859 108749 270893
rect 108783 270859 108803 270893
rect 108729 270825 108803 270859
rect 108729 270801 108749 270825
rect 106769 270791 108749 270801
rect 108783 270791 108803 270825
rect 108947 271000 109088 271029
rect 108947 270974 109122 271000
rect 108947 270940 109009 270974
rect 109043 270966 109122 270974
rect 109043 270940 109088 270966
rect 108947 270932 109088 270940
rect 108947 270902 109122 270932
rect 108947 270868 109009 270902
rect 109043 270898 109122 270902
rect 109043 270868 109088 270898
rect 108947 270864 109088 270868
rect 108947 270830 109122 270864
rect 108947 270811 109088 270830
rect 106715 270784 108803 270791
rect 106715 270750 106875 270784
rect 106909 270750 106943 270784
rect 106977 270750 107011 270784
rect 107045 270750 107079 270784
rect 107113 270750 107147 270784
rect 107181 270750 107215 270784
rect 107249 270750 107283 270784
rect 107317 270750 107351 270784
rect 107385 270750 107419 270784
rect 107453 270750 107487 270784
rect 107521 270750 107555 270784
rect 107589 270750 107623 270784
rect 107657 270750 107691 270784
rect 107725 270750 107759 270784
rect 107793 270750 107827 270784
rect 107861 270750 107895 270784
rect 107929 270750 107963 270784
rect 107997 270750 108031 270784
rect 108065 270750 108099 270784
rect 108133 270750 108167 270784
rect 108201 270750 108235 270784
rect 108269 270750 108303 270784
rect 108337 270750 108371 270784
rect 108405 270750 108439 270784
rect 108473 270750 108507 270784
rect 108541 270750 108575 270784
rect 108609 270750 108643 270784
rect 108677 270750 108803 270784
rect 106715 270733 108803 270750
rect 109088 270762 109122 270796
rect 107329 270334 108364 270733
rect 109088 270694 109122 270728
rect 109088 270626 109122 270660
rect 109394 272473 109458 272507
rect 109492 272473 109556 272507
rect 109394 272411 109428 272473
rect 109394 272339 109428 272365
rect 109394 272267 109428 272297
rect 109394 272195 109428 272229
rect 109394 272127 109428 272161
rect 109394 272059 109428 272089
rect 109394 271991 109428 272017
rect 109394 271923 109428 271945
rect 109394 271855 109428 271873
rect 109394 271787 109428 271801
rect 109394 271719 109428 271729
rect 109394 271651 109428 271657
rect 109394 271583 109428 271585
rect 109394 271547 109428 271549
rect 109394 271475 109428 271481
rect 109394 271403 109428 271413
rect 109394 271331 109428 271345
rect 109394 271259 109428 271277
rect 109394 271187 109428 271209
rect 109394 271115 109428 271141
rect 109394 271043 109428 271073
rect 109394 270971 109428 271005
rect 109394 270903 109428 270937
rect 109394 270835 109428 270865
rect 109394 270767 109428 270793
rect 109394 270659 109428 270721
rect 109522 272411 109556 272473
rect 109522 272339 109556 272365
rect 109522 272267 109556 272297
rect 109522 272195 109556 272229
rect 109522 272127 109556 272161
rect 109522 272059 109556 272089
rect 109522 271991 109556 272017
rect 109522 271923 109556 271945
rect 109522 271855 109556 271873
rect 109522 271787 109556 271801
rect 109522 271719 109556 271729
rect 109522 271651 109556 271657
rect 109522 271583 109556 271585
rect 109522 271547 109556 271549
rect 109522 271475 109556 271481
rect 109522 271403 109556 271413
rect 109522 271331 109556 271345
rect 109522 271259 109556 271277
rect 109522 271187 109556 271209
rect 109522 271115 109556 271141
rect 109522 271043 109556 271073
rect 109522 270971 109556 271005
rect 109522 270903 109556 270937
rect 109522 270835 109556 270865
rect 109522 270767 109556 270793
rect 109522 270659 109556 270721
rect 109394 270625 109458 270659
rect 109492 270625 109556 270659
rect 109827 272462 109861 272496
rect 109827 272394 109861 272428
rect 109827 272326 109861 272360
rect 109827 272258 109861 272292
rect 109827 272190 109861 272224
rect 109827 272122 109861 272156
rect 109827 272054 109861 272088
rect 109827 271986 109861 272020
rect 109827 271918 109861 271952
rect 109827 271850 109861 271884
rect 109827 271782 109861 271816
rect 109827 271714 109861 271748
rect 109827 271646 109861 271680
rect 109827 271578 109861 271612
rect 109827 271510 109861 271544
rect 109827 271442 109861 271476
rect 109827 271374 109861 271408
rect 109827 271306 109861 271340
rect 109827 271238 109861 271272
rect 109827 271170 109861 271204
rect 109827 271102 109861 271136
rect 109827 271034 109861 271068
rect 109827 270966 109861 271000
rect 109827 270898 109861 270932
rect 109827 270830 109861 270864
rect 109827 270762 109861 270796
rect 109827 270694 109861 270728
rect 109827 270626 109861 270660
rect 109088 270555 109122 270592
rect 109827 270555 109861 270592
rect 109088 270521 109151 270555
rect 109185 270521 109219 270555
rect 109253 270521 109287 270555
rect 109321 270521 109355 270555
rect 109389 270521 109423 270555
rect 109457 270521 109491 270555
rect 109525 270521 109559 270555
rect 109593 270521 109627 270555
rect 109661 270521 109695 270555
rect 109729 270521 109763 270555
rect 109797 270521 109861 270555
rect 110081 270334 110085 272786
rect 106455 270306 110085 270334
rect 106455 270212 106585 270306
rect 106281 270204 106585 270212
rect 109951 270212 110085 270306
rect 110255 270212 110259 272898
rect 111046 272704 111072 281102
rect 111174 281099 119031 281102
rect 111174 272704 111200 281099
rect 113036 280904 114022 281099
rect 114455 280929 114537 280963
rect 114571 280929 114605 280963
rect 114639 280929 114673 280963
rect 114707 280929 114741 280963
rect 114775 280929 114809 280963
rect 114843 280929 114877 280963
rect 114911 280929 114945 280963
rect 114979 280929 115226 280963
rect 115260 280929 115294 280963
rect 115328 280929 115362 280963
rect 115396 280929 115430 280963
rect 115464 280929 115498 280963
rect 115532 280929 115566 280963
rect 115600 280929 115634 280963
rect 115668 280929 115750 280963
rect 111520 280866 112814 280902
rect 113036 280900 114246 280904
rect 113036 280899 114353 280900
rect 111520 280832 111547 280866
rect 111587 280832 111615 280866
rect 111659 280832 111683 280866
rect 111731 280832 111751 280866
rect 111803 280832 111819 280866
rect 111875 280832 111887 280866
rect 111947 280832 111955 280866
rect 112019 280832 112023 280866
rect 112125 280832 112129 280866
rect 112193 280832 112201 280866
rect 112261 280832 112273 280866
rect 112329 280832 112345 280866
rect 112397 280832 112417 280866
rect 112465 280832 112489 280866
rect 112533 280832 112561 280866
rect 112601 280832 112628 280866
rect 111452 280793 111486 280820
rect 111452 280723 111486 280757
rect 111452 280660 111486 280687
rect 112662 280793 112696 280820
rect 112662 280723 112696 280757
rect 112662 280660 112696 280687
rect 111520 280614 111547 280648
rect 111587 280614 111615 280648
rect 111659 280614 111683 280648
rect 111731 280614 111751 280648
rect 111803 280614 111819 280648
rect 111875 280614 111887 280648
rect 111947 280614 111955 280648
rect 112019 280614 112023 280648
rect 112125 280614 112129 280648
rect 112193 280614 112201 280648
rect 112261 280614 112273 280648
rect 112329 280614 112345 280648
rect 112397 280614 112417 280648
rect 112465 280614 112489 280648
rect 112533 280614 112561 280648
rect 112601 280614 112628 280648
rect 111334 280578 112628 280614
rect 112772 280582 112814 280866
rect 112966 280876 114353 280899
rect 112966 280874 114243 280876
rect 112966 280840 112993 280874
rect 113033 280840 113061 280874
rect 113105 280840 113129 280874
rect 113177 280840 113197 280874
rect 113249 280840 113265 280874
rect 113321 280840 113333 280874
rect 113393 280840 113401 280874
rect 113465 280840 113469 280874
rect 113571 280840 113575 280874
rect 113639 280840 113647 280874
rect 113707 280840 113719 280874
rect 113775 280840 113791 280874
rect 113843 280840 113863 280874
rect 113911 280840 113935 280874
rect 113979 280840 114007 280874
rect 114047 280870 114243 280874
rect 114047 280840 114074 280870
rect 112898 280781 112932 280828
rect 112898 280711 112932 280745
rect 112898 280628 112932 280675
rect 114108 280781 114142 280828
rect 114108 280711 114142 280745
rect 114108 280628 114142 280675
rect 114210 280774 114243 280870
rect 114345 280774 114353 280876
rect 114210 280750 114353 280774
rect 114455 280897 114489 280929
rect 114455 280829 114489 280863
rect 114652 280849 114862 280929
rect 114652 280815 114672 280849
rect 114738 280815 114740 280849
rect 114774 280815 114776 280849
rect 114842 280815 114862 280849
rect 114652 280814 114862 280815
rect 115027 280897 115178 280929
rect 115061 280863 115144 280897
rect 115027 280829 115178 280863
rect 114455 280761 114489 280795
rect 112966 280582 112993 280616
rect 113033 280582 113061 280616
rect 113105 280582 113129 280616
rect 113177 280582 113197 280616
rect 113249 280582 113265 280616
rect 113321 280582 113333 280616
rect 113393 280582 113401 280616
rect 113465 280582 113469 280616
rect 113571 280582 113575 280616
rect 113639 280582 113647 280616
rect 113707 280582 113719 280616
rect 113775 280582 113791 280616
rect 113843 280582 113863 280616
rect 113911 280582 113935 280616
rect 113979 280582 114007 280616
rect 114047 280582 114074 280616
rect 111334 280254 111376 280578
rect 112772 280548 114074 280582
rect 112772 280542 112832 280548
rect 111520 280506 112832 280542
rect 111520 280472 111547 280506
rect 111587 280472 111615 280506
rect 111659 280472 111683 280506
rect 111731 280472 111751 280506
rect 111803 280472 111819 280506
rect 111875 280472 111887 280506
rect 111947 280472 111955 280506
rect 112019 280472 112023 280506
rect 112125 280472 112129 280506
rect 112193 280472 112201 280506
rect 112261 280472 112273 280506
rect 112329 280472 112345 280506
rect 112397 280472 112417 280506
rect 112465 280472 112489 280506
rect 112533 280472 112561 280506
rect 112601 280472 112628 280506
rect 111452 280433 111486 280460
rect 111452 280363 111486 280397
rect 111452 280300 111486 280327
rect 112662 280433 112696 280460
rect 112662 280363 112696 280397
rect 112662 280300 112696 280327
rect 111520 280254 111547 280288
rect 111587 280254 111615 280288
rect 111659 280254 111683 280288
rect 111731 280254 111751 280288
rect 111803 280254 111819 280288
rect 111875 280254 111887 280288
rect 111947 280254 111955 280288
rect 112019 280254 112023 280288
rect 112125 280254 112129 280288
rect 112193 280254 112201 280288
rect 112261 280254 112273 280288
rect 112329 280254 112345 280288
rect 112397 280254 112417 280288
rect 112465 280254 112489 280288
rect 112533 280254 112561 280288
rect 112601 280254 112628 280288
rect 111334 280218 112628 280254
rect 111334 279894 111376 280218
rect 112772 280182 112832 280506
rect 114210 280484 114246 280750
rect 112966 280450 114246 280484
rect 114455 280693 114489 280727
rect 114455 280625 114489 280659
rect 114455 280557 114489 280591
rect 114455 280489 114489 280523
rect 112966 280416 112993 280450
rect 113033 280416 113061 280450
rect 113105 280416 113129 280450
rect 113177 280416 113197 280450
rect 113249 280416 113265 280450
rect 113321 280416 113333 280450
rect 113393 280416 113401 280450
rect 113465 280416 113469 280450
rect 113571 280416 113575 280450
rect 113639 280416 113647 280450
rect 113707 280416 113719 280450
rect 113775 280416 113791 280450
rect 113843 280416 113863 280450
rect 113911 280416 113935 280450
rect 113979 280416 114007 280450
rect 114047 280416 114074 280450
rect 114455 280421 114489 280455
rect 112898 280357 112932 280404
rect 112898 280287 112932 280321
rect 112898 280204 112932 280251
rect 114108 280357 114142 280404
rect 114108 280287 114142 280321
rect 114108 280204 114142 280251
rect 114455 280353 114489 280387
rect 114455 280285 114489 280319
rect 114455 280217 114489 280251
rect 111520 280160 112832 280182
rect 112966 280160 112993 280192
rect 111520 280158 112993 280160
rect 113033 280158 113061 280192
rect 113105 280158 113129 280192
rect 113177 280158 113197 280192
rect 113249 280158 113265 280192
rect 113321 280158 113333 280192
rect 113393 280158 113401 280192
rect 113465 280158 113469 280192
rect 113571 280158 113575 280192
rect 113639 280158 113647 280192
rect 113707 280158 113719 280192
rect 113775 280158 113791 280192
rect 113843 280158 113863 280192
rect 113911 280158 113935 280192
rect 113979 280158 114007 280192
rect 114047 280158 114074 280192
rect 111520 280146 114074 280158
rect 111520 280112 111547 280146
rect 111587 280112 111615 280146
rect 111659 280112 111683 280146
rect 111731 280112 111751 280146
rect 111803 280112 111819 280146
rect 111875 280112 111887 280146
rect 111947 280112 111955 280146
rect 112019 280112 112023 280146
rect 112125 280112 112129 280146
rect 112193 280112 112201 280146
rect 112261 280112 112273 280146
rect 112329 280112 112345 280146
rect 112397 280112 112417 280146
rect 112465 280112 112489 280146
rect 112533 280112 112561 280146
rect 112601 280112 112628 280146
rect 112744 280143 114074 280146
rect 114455 280149 114489 280183
rect 112744 280126 114396 280143
rect 111452 280073 111486 280100
rect 111452 280003 111486 280037
rect 111452 279940 111486 279967
rect 112662 280073 112696 280100
rect 112662 280003 112696 280037
rect 112662 279940 112696 279967
rect 111520 279894 111547 279928
rect 111587 279894 111615 279928
rect 111659 279894 111683 279928
rect 111731 279894 111751 279928
rect 111803 279894 111819 279928
rect 111875 279894 111887 279928
rect 111947 279894 111955 279928
rect 112019 279894 112023 279928
rect 112125 279894 112129 279928
rect 112193 279894 112201 279928
rect 112261 279894 112273 279928
rect 112329 279894 112345 279928
rect 112397 279894 112417 279928
rect 112465 279894 112489 279928
rect 112533 279894 112561 279928
rect 112601 279894 112628 279928
rect 111334 279858 112628 279894
rect 111334 279534 111376 279858
rect 112744 279822 112780 280126
rect 113892 280107 114396 280126
rect 111520 279786 112780 279822
rect 112832 280048 113264 280082
rect 112832 280040 113023 280048
rect 112832 279786 112872 280040
rect 112996 280014 113023 280040
rect 113063 280014 113091 280048
rect 113135 280014 113159 280048
rect 113207 280014 113227 280048
rect 113279 280014 113295 280048
rect 113351 280014 113363 280048
rect 113423 280014 113431 280048
rect 113495 280014 113499 280048
rect 113601 280014 113605 280048
rect 113669 280014 113677 280048
rect 113737 280014 113749 280048
rect 113805 280014 113821 280048
rect 113873 280014 113893 280048
rect 113941 280014 113965 280048
rect 114009 280014 114037 280048
rect 114077 280014 114104 280048
rect 112928 279979 112962 280002
rect 112928 279922 112962 279945
rect 114138 279979 114172 280002
rect 114138 279922 114172 279945
rect 114324 279951 114396 280107
rect 114324 279917 114342 279951
rect 114376 279917 114396 279951
rect 112996 279882 113023 279910
rect 112994 279876 113023 279882
rect 113063 279876 113091 279910
rect 113135 279876 113159 279910
rect 113207 279876 113227 279910
rect 113279 279876 113295 279910
rect 113351 279876 113363 279910
rect 113423 279876 113431 279910
rect 113495 279876 113499 279910
rect 113601 279876 113605 279910
rect 113669 279876 113677 279910
rect 113737 279876 113749 279910
rect 113805 279876 113821 279910
rect 113873 279876 113893 279910
rect 113941 279876 113965 279910
rect 114009 279876 114037 279910
rect 114077 279882 114104 279910
rect 114077 279876 114274 279882
rect 112994 279836 114274 279876
rect 114324 279869 114396 279917
rect 114455 280081 114489 280115
rect 114455 280013 114489 280047
rect 114455 279945 114489 279979
rect 114576 280764 114610 280803
rect 114576 280692 114610 280722
rect 114576 280620 114610 280654
rect 114576 280552 114610 280586
rect 114576 280484 114610 280514
rect 114576 280275 114610 280442
rect 114904 280764 114938 280803
rect 114904 280692 114938 280722
rect 114904 280620 114938 280654
rect 114904 280552 114938 280586
rect 114904 280484 114938 280514
rect 114653 280357 114672 280391
rect 114738 280357 114740 280391
rect 114774 280357 114776 280391
rect 114842 280357 114861 280391
rect 114904 280311 114938 280442
rect 115061 280795 115144 280829
rect 115343 280849 115553 280929
rect 115343 280815 115363 280849
rect 115429 280815 115431 280849
rect 115465 280815 115467 280849
rect 115533 280815 115553 280849
rect 115343 280814 115553 280815
rect 115716 280897 115750 280929
rect 116183 280904 117169 281099
rect 115959 280900 117169 280904
rect 115716 280829 115750 280863
rect 115027 280761 115178 280795
rect 115061 280727 115144 280761
rect 115027 280693 115178 280727
rect 115061 280659 115144 280693
rect 115027 280625 115178 280659
rect 115061 280591 115144 280625
rect 115027 280557 115178 280591
rect 115061 280523 115144 280557
rect 115027 280489 115178 280523
rect 115061 280455 115144 280489
rect 115027 280421 115178 280455
rect 115061 280387 115144 280421
rect 115027 280353 115178 280387
rect 115061 280319 115144 280353
rect 114865 280277 114970 280311
rect 114865 280275 114899 280277
rect 114576 280243 114899 280275
rect 114933 280243 114970 280277
rect 114576 280227 114970 280243
rect 114576 280090 114610 280227
rect 114865 280204 114970 280227
rect 115027 280285 115178 280319
rect 115267 280764 115301 280803
rect 115267 280692 115301 280722
rect 115267 280620 115301 280654
rect 115267 280552 115301 280586
rect 115267 280484 115301 280514
rect 115267 280311 115301 280442
rect 115595 280764 115629 280803
rect 115595 280692 115629 280722
rect 115595 280620 115629 280654
rect 115595 280552 115629 280586
rect 115595 280484 115629 280514
rect 115344 280357 115363 280391
rect 115429 280357 115431 280391
rect 115465 280357 115467 280391
rect 115533 280357 115552 280391
rect 115061 280251 115144 280285
rect 115027 280217 115178 280251
rect 114653 280129 114672 280163
rect 114738 280129 114740 280163
rect 114774 280129 114776 280163
rect 114842 280129 114861 280163
rect 114576 280020 114610 280054
rect 114576 279957 114610 279984
rect 114904 280090 114938 280204
rect 114904 280020 114938 280054
rect 114904 279957 114938 279984
rect 115061 280183 115144 280217
rect 115235 280277 115340 280311
rect 115235 280243 115271 280277
rect 115305 280275 115340 280277
rect 115595 280275 115629 280442
rect 115305 280243 115629 280275
rect 115235 280227 115629 280243
rect 115235 280204 115340 280227
rect 115027 280149 115178 280183
rect 115061 280115 115144 280149
rect 115027 280081 115178 280115
rect 115061 280047 115144 280081
rect 115027 280013 115178 280047
rect 115061 279979 115144 280013
rect 115027 279945 115178 279979
rect 115267 280090 115301 280204
rect 115344 280129 115363 280163
rect 115429 280129 115431 280163
rect 115465 280129 115467 280163
rect 115533 280129 115552 280163
rect 115267 280020 115301 280054
rect 115267 279957 115301 279984
rect 115595 280090 115629 280227
rect 115595 280020 115629 280054
rect 115595 279957 115629 279984
rect 115716 280761 115750 280795
rect 115852 280899 117169 280900
rect 115852 280876 117239 280899
rect 115852 280774 115860 280876
rect 115962 280874 117239 280876
rect 115962 280870 116158 280874
rect 115962 280774 115995 280870
rect 116131 280840 116158 280870
rect 116198 280840 116226 280874
rect 116270 280840 116294 280874
rect 116342 280840 116362 280874
rect 116414 280840 116430 280874
rect 116486 280840 116498 280874
rect 116558 280840 116566 280874
rect 116630 280840 116634 280874
rect 116736 280840 116740 280874
rect 116804 280840 116812 280874
rect 116872 280840 116884 280874
rect 116940 280840 116956 280874
rect 117008 280840 117028 280874
rect 117076 280840 117100 280874
rect 117144 280840 117172 280874
rect 117212 280840 117239 280874
rect 117391 280866 118685 280902
rect 115852 280750 115995 280774
rect 115716 280693 115750 280727
rect 115716 280625 115750 280659
rect 115716 280557 115750 280591
rect 115716 280489 115750 280523
rect 115716 280421 115750 280455
rect 115959 280484 115995 280750
rect 116063 280781 116097 280828
rect 116063 280711 116097 280745
rect 116063 280628 116097 280675
rect 117273 280781 117307 280828
rect 117273 280711 117307 280745
rect 117273 280628 117307 280675
rect 116131 280582 116158 280616
rect 116198 280582 116226 280616
rect 116270 280582 116294 280616
rect 116342 280582 116362 280616
rect 116414 280582 116430 280616
rect 116486 280582 116498 280616
rect 116558 280582 116566 280616
rect 116630 280582 116634 280616
rect 116736 280582 116740 280616
rect 116804 280582 116812 280616
rect 116872 280582 116884 280616
rect 116940 280582 116956 280616
rect 117008 280582 117028 280616
rect 117076 280582 117100 280616
rect 117144 280582 117172 280616
rect 117212 280582 117239 280616
rect 117391 280582 117433 280866
rect 117577 280832 117604 280866
rect 117644 280832 117672 280866
rect 117716 280832 117740 280866
rect 117788 280832 117808 280866
rect 117860 280832 117876 280866
rect 117932 280832 117944 280866
rect 118004 280832 118012 280866
rect 118076 280832 118080 280866
rect 118182 280832 118186 280866
rect 118250 280832 118258 280866
rect 118318 280832 118330 280866
rect 118386 280832 118402 280866
rect 118454 280832 118474 280866
rect 118522 280832 118546 280866
rect 118590 280832 118618 280866
rect 118658 280832 118685 280866
rect 117509 280793 117543 280820
rect 117509 280723 117543 280757
rect 117509 280660 117543 280687
rect 118719 280793 118753 280820
rect 118719 280723 118753 280757
rect 118719 280660 118753 280687
rect 116131 280548 117433 280582
rect 117577 280614 117604 280648
rect 117644 280614 117672 280648
rect 117716 280614 117740 280648
rect 117788 280614 117808 280648
rect 117860 280614 117876 280648
rect 117932 280614 117944 280648
rect 118004 280614 118012 280648
rect 118076 280614 118080 280648
rect 118182 280614 118186 280648
rect 118250 280614 118258 280648
rect 118318 280614 118330 280648
rect 118386 280614 118402 280648
rect 118454 280614 118474 280648
rect 118522 280614 118546 280648
rect 118590 280614 118618 280648
rect 118658 280614 118685 280648
rect 117577 280578 118871 280614
rect 117373 280542 117433 280548
rect 117373 280506 118685 280542
rect 115959 280450 117239 280484
rect 116131 280416 116158 280450
rect 116198 280416 116226 280450
rect 116270 280416 116294 280450
rect 116342 280416 116362 280450
rect 116414 280416 116430 280450
rect 116486 280416 116498 280450
rect 116558 280416 116566 280450
rect 116630 280416 116634 280450
rect 116736 280416 116740 280450
rect 116804 280416 116812 280450
rect 116872 280416 116884 280450
rect 116940 280416 116956 280450
rect 117008 280416 117028 280450
rect 117076 280416 117100 280450
rect 117144 280416 117172 280450
rect 117212 280416 117239 280450
rect 115716 280353 115750 280387
rect 115716 280285 115750 280319
rect 115716 280217 115750 280251
rect 116063 280357 116097 280404
rect 116063 280287 116097 280321
rect 116063 280204 116097 280251
rect 117273 280357 117307 280404
rect 117273 280287 117307 280321
rect 117273 280204 117307 280251
rect 115716 280149 115750 280183
rect 116131 280158 116158 280192
rect 116198 280158 116226 280192
rect 116270 280158 116294 280192
rect 116342 280158 116362 280192
rect 116414 280158 116430 280192
rect 116486 280158 116498 280192
rect 116558 280158 116566 280192
rect 116630 280158 116634 280192
rect 116736 280158 116740 280192
rect 116804 280158 116812 280192
rect 116872 280158 116884 280192
rect 116940 280158 116956 280192
rect 117008 280158 117028 280192
rect 117076 280158 117100 280192
rect 117144 280158 117172 280192
rect 117212 280160 117239 280192
rect 117373 280182 117433 280506
rect 117577 280472 117604 280506
rect 117644 280472 117672 280506
rect 117716 280472 117740 280506
rect 117788 280472 117808 280506
rect 117860 280472 117876 280506
rect 117932 280472 117944 280506
rect 118004 280472 118012 280506
rect 118076 280472 118080 280506
rect 118182 280472 118186 280506
rect 118250 280472 118258 280506
rect 118318 280472 118330 280506
rect 118386 280472 118402 280506
rect 118454 280472 118474 280506
rect 118522 280472 118546 280506
rect 118590 280472 118618 280506
rect 118658 280472 118685 280506
rect 117509 280433 117543 280460
rect 117509 280363 117543 280397
rect 117509 280300 117543 280327
rect 118719 280433 118753 280460
rect 118719 280363 118753 280397
rect 118719 280300 118753 280327
rect 117577 280254 117604 280288
rect 117644 280254 117672 280288
rect 117716 280254 117740 280288
rect 117788 280254 117808 280288
rect 117860 280254 117876 280288
rect 117932 280254 117944 280288
rect 118004 280254 118012 280288
rect 118076 280254 118080 280288
rect 118182 280254 118186 280288
rect 118250 280254 118258 280288
rect 118318 280254 118330 280288
rect 118386 280254 118402 280288
rect 118454 280254 118474 280288
rect 118522 280254 118546 280288
rect 118590 280254 118618 280288
rect 118658 280254 118685 280288
rect 118829 280254 118871 280578
rect 117577 280218 118871 280254
rect 117373 280160 118685 280182
rect 117212 280158 118685 280160
rect 116131 280146 118685 280158
rect 116131 280143 117461 280146
rect 115716 280081 115750 280115
rect 115716 280013 115750 280047
rect 115716 279945 115750 279979
rect 114455 279877 114489 279911
rect 111520 279752 111547 279786
rect 111587 279752 111615 279786
rect 111659 279752 111683 279786
rect 111731 279752 111751 279786
rect 111803 279752 111819 279786
rect 111875 279752 111887 279786
rect 111947 279752 111955 279786
rect 112019 279752 112023 279786
rect 112125 279752 112129 279786
rect 112193 279752 112201 279786
rect 112261 279752 112273 279786
rect 112329 279752 112345 279786
rect 112397 279752 112417 279786
rect 112465 279752 112489 279786
rect 112533 279752 112561 279786
rect 112601 279752 112628 279786
rect 112832 279750 113216 279786
rect 112832 279746 113023 279750
rect 111452 279713 111486 279740
rect 111452 279643 111486 279677
rect 111452 279580 111486 279607
rect 112662 279713 112696 279740
rect 112832 279718 112872 279746
rect 112996 279716 113023 279746
rect 113063 279716 113091 279750
rect 113135 279716 113159 279750
rect 113207 279716 113227 279750
rect 113279 279716 113295 279750
rect 113351 279716 113363 279750
rect 113423 279716 113431 279750
rect 113495 279716 113499 279750
rect 113601 279716 113605 279750
rect 113669 279716 113677 279750
rect 113737 279716 113749 279750
rect 113805 279716 113821 279750
rect 113873 279716 113893 279750
rect 113941 279716 113965 279750
rect 114009 279716 114037 279750
rect 114077 279716 114104 279750
rect 112662 279643 112696 279677
rect 112928 279681 112962 279704
rect 112928 279624 112962 279647
rect 114138 279681 114172 279704
rect 114138 279624 114172 279647
rect 112662 279580 112696 279607
rect 112996 279578 113023 279612
rect 113063 279578 113091 279612
rect 113135 279578 113159 279612
rect 113207 279578 113227 279612
rect 113279 279578 113295 279612
rect 113351 279578 113363 279612
rect 113423 279578 113431 279612
rect 113495 279578 113499 279612
rect 113601 279578 113605 279612
rect 113669 279578 113677 279612
rect 113737 279578 113749 279612
rect 113805 279578 113821 279612
rect 113873 279578 113893 279612
rect 113941 279578 113965 279612
rect 114009 279578 114037 279612
rect 114077 279578 114104 279612
rect 114234 279578 114274 279836
rect 114653 279911 114672 279945
rect 114738 279911 114740 279945
rect 114774 279911 114776 279945
rect 114842 279911 114861 279945
rect 114653 279874 114709 279911
rect 114805 279876 114861 279911
rect 115061 279911 115144 279945
rect 115027 279877 115178 279911
rect 114455 279809 114489 279843
rect 114455 279741 114489 279775
rect 114455 279673 114489 279707
rect 114455 279605 114489 279639
rect 112994 279571 114455 279578
rect 111520 279534 111547 279568
rect 111587 279534 111615 279568
rect 111659 279534 111683 279568
rect 111731 279534 111751 279568
rect 111803 279534 111819 279568
rect 111875 279534 111887 279568
rect 111947 279534 111955 279568
rect 112019 279534 112023 279568
rect 112125 279534 112129 279568
rect 112193 279534 112201 279568
rect 112261 279534 112273 279568
rect 112329 279534 112345 279568
rect 112397 279534 112417 279568
rect 112465 279534 112489 279568
rect 112533 279534 112561 279568
rect 112601 279534 112628 279568
rect 111334 279498 112628 279534
rect 112994 279537 114489 279571
rect 114538 279835 114709 279874
rect 114804 279854 114991 279876
rect 114538 279709 114576 279835
rect 114804 279820 114899 279854
rect 114933 279820 114991 279854
rect 114804 279791 114991 279820
rect 115061 279843 115144 279877
rect 115344 279911 115363 279945
rect 115429 279911 115431 279945
rect 115465 279911 115467 279945
rect 115533 279911 115552 279945
rect 115344 279876 115400 279911
rect 115027 279809 115178 279843
rect 114653 279721 114672 279755
rect 114738 279721 114740 279755
rect 114774 279721 114776 279755
rect 114842 279721 114861 279755
rect 114938 279709 114975 279791
rect 114538 279682 114610 279709
rect 114538 279646 114576 279682
rect 114538 279612 114610 279646
rect 114538 279576 114576 279612
rect 114538 279549 114610 279576
rect 114904 279682 114975 279709
rect 114938 279646 114975 279682
rect 114904 279612 114975 279646
rect 114938 279576 114975 279612
rect 114904 279549 114975 279576
rect 115061 279775 115144 279809
rect 115214 279854 115401 279876
rect 115214 279820 115271 279854
rect 115305 279820 115401 279854
rect 115496 279874 115552 279911
rect 115716 279877 115750 279911
rect 115496 279835 115667 279874
rect 115214 279791 115401 279820
rect 115027 279741 115178 279775
rect 115061 279707 115144 279741
rect 115027 279673 115178 279707
rect 115061 279639 115144 279673
rect 115027 279605 115178 279639
rect 115061 279571 115144 279605
rect 115027 279537 115178 279571
rect 115230 279709 115267 279791
rect 115344 279721 115363 279755
rect 115429 279721 115431 279755
rect 115465 279721 115467 279755
rect 115533 279721 115552 279755
rect 115629 279709 115667 279835
rect 115230 279682 115301 279709
rect 115230 279646 115267 279682
rect 115230 279612 115301 279646
rect 115230 279576 115267 279612
rect 115230 279549 115301 279576
rect 115595 279682 115667 279709
rect 115629 279646 115667 279682
rect 115595 279612 115667 279646
rect 115629 279576 115667 279612
rect 115595 279549 115667 279576
rect 115809 280126 117461 280143
rect 115809 280107 116313 280126
rect 115809 279951 115881 280107
rect 116941 280048 117373 280082
rect 116101 280014 116128 280048
rect 116168 280014 116196 280048
rect 116240 280014 116264 280048
rect 116312 280014 116332 280048
rect 116384 280014 116400 280048
rect 116456 280014 116468 280048
rect 116528 280014 116536 280048
rect 116600 280014 116604 280048
rect 116706 280014 116710 280048
rect 116774 280014 116782 280048
rect 116842 280014 116854 280048
rect 116910 280014 116926 280048
rect 116978 280014 116998 280048
rect 117046 280014 117070 280048
rect 117114 280014 117142 280048
rect 117182 280040 117373 280048
rect 117182 280014 117209 280040
rect 115809 279917 115828 279951
rect 115862 279917 115881 279951
rect 116033 279979 116067 280002
rect 116033 279922 116067 279945
rect 117243 279979 117277 280002
rect 117243 279922 117277 279945
rect 115809 279869 115881 279917
rect 116101 279882 116128 279910
rect 115931 279876 116128 279882
rect 116168 279876 116196 279910
rect 116240 279876 116264 279910
rect 116312 279876 116332 279910
rect 116384 279876 116400 279910
rect 116456 279876 116468 279910
rect 116528 279876 116536 279910
rect 116600 279876 116604 279910
rect 116706 279876 116710 279910
rect 116774 279876 116782 279910
rect 116842 279876 116854 279910
rect 116910 279876 116926 279910
rect 116978 279876 116998 279910
rect 117046 279876 117070 279910
rect 117114 279876 117142 279910
rect 117182 279882 117209 279910
rect 117182 279876 117211 279882
rect 115716 279809 115750 279843
rect 115716 279741 115750 279775
rect 115716 279673 115750 279707
rect 115716 279605 115750 279639
rect 115931 279836 117211 279876
rect 115931 279578 115971 279836
rect 117333 279786 117373 280040
rect 117425 279822 117461 280126
rect 117577 280112 117604 280146
rect 117644 280112 117672 280146
rect 117716 280112 117740 280146
rect 117788 280112 117808 280146
rect 117860 280112 117876 280146
rect 117932 280112 117944 280146
rect 118004 280112 118012 280146
rect 118076 280112 118080 280146
rect 118182 280112 118186 280146
rect 118250 280112 118258 280146
rect 118318 280112 118330 280146
rect 118386 280112 118402 280146
rect 118454 280112 118474 280146
rect 118522 280112 118546 280146
rect 118590 280112 118618 280146
rect 118658 280112 118685 280146
rect 117509 280073 117543 280100
rect 117509 280003 117543 280037
rect 117509 279940 117543 279967
rect 118719 280073 118753 280100
rect 118719 280003 118753 280037
rect 118719 279940 118753 279967
rect 117577 279894 117604 279928
rect 117644 279894 117672 279928
rect 117716 279894 117740 279928
rect 117788 279894 117808 279928
rect 117860 279894 117876 279928
rect 117932 279894 117944 279928
rect 118004 279894 118012 279928
rect 118076 279894 118080 279928
rect 118182 279894 118186 279928
rect 118250 279894 118258 279928
rect 118318 279894 118330 279928
rect 118386 279894 118402 279928
rect 118454 279894 118474 279928
rect 118522 279894 118546 279928
rect 118590 279894 118618 279928
rect 118658 279894 118685 279928
rect 118829 279894 118871 280218
rect 117577 279858 118871 279894
rect 117425 279786 118685 279822
rect 116989 279750 117373 279786
rect 117577 279752 117604 279786
rect 117644 279752 117672 279786
rect 117716 279752 117740 279786
rect 117788 279752 117808 279786
rect 117860 279752 117876 279786
rect 117932 279752 117944 279786
rect 118004 279752 118012 279786
rect 118076 279752 118080 279786
rect 118182 279752 118186 279786
rect 118250 279752 118258 279786
rect 118318 279752 118330 279786
rect 118386 279752 118402 279786
rect 118454 279752 118474 279786
rect 118522 279752 118546 279786
rect 118590 279752 118618 279786
rect 118658 279752 118685 279786
rect 116101 279716 116128 279750
rect 116168 279716 116196 279750
rect 116240 279716 116264 279750
rect 116312 279716 116332 279750
rect 116384 279716 116400 279750
rect 116456 279716 116468 279750
rect 116528 279716 116536 279750
rect 116600 279716 116604 279750
rect 116706 279716 116710 279750
rect 116774 279716 116782 279750
rect 116842 279716 116854 279750
rect 116910 279716 116926 279750
rect 116978 279716 116998 279750
rect 117046 279716 117070 279750
rect 117114 279716 117142 279750
rect 117182 279746 117373 279750
rect 117182 279716 117209 279746
rect 117333 279718 117373 279746
rect 117509 279713 117543 279740
rect 116033 279681 116067 279704
rect 116033 279624 116067 279647
rect 117243 279681 117277 279704
rect 117243 279624 117277 279647
rect 117509 279643 117543 279677
rect 116101 279578 116128 279612
rect 116168 279578 116196 279612
rect 116240 279578 116264 279612
rect 116312 279578 116332 279612
rect 116384 279578 116400 279612
rect 116456 279578 116468 279612
rect 116528 279578 116536 279612
rect 116600 279578 116604 279612
rect 116706 279578 116710 279612
rect 116774 279578 116782 279612
rect 116842 279578 116854 279612
rect 116910 279578 116926 279612
rect 116978 279578 116998 279612
rect 117046 279578 117070 279612
rect 117114 279578 117142 279612
rect 117182 279578 117209 279612
rect 117509 279580 117543 279607
rect 118719 279713 118753 279740
rect 118719 279643 118753 279677
rect 118719 279580 118753 279607
rect 115750 279571 117211 279578
rect 115716 279537 117211 279571
rect 112994 279532 114455 279537
rect 114653 279503 114672 279537
rect 114738 279503 114740 279537
rect 114774 279503 114776 279537
rect 114842 279503 114861 279537
rect 115061 279503 115144 279537
rect 115344 279503 115363 279537
rect 115429 279503 115431 279537
rect 115465 279503 115467 279537
rect 115533 279503 115552 279537
rect 115750 279532 117211 279537
rect 117577 279534 117604 279568
rect 117644 279534 117672 279568
rect 117716 279534 117740 279568
rect 117788 279534 117808 279568
rect 117860 279534 117876 279568
rect 117932 279534 117944 279568
rect 118004 279534 118012 279568
rect 118076 279534 118080 279568
rect 118182 279534 118186 279568
rect 118250 279534 118258 279568
rect 118318 279534 118330 279568
rect 118386 279534 118402 279568
rect 118454 279534 118474 279568
rect 118522 279534 118546 279568
rect 118590 279534 118618 279568
rect 118658 279534 118685 279568
rect 118829 279534 118871 279858
rect 114455 279469 114489 279503
rect 115027 279487 115178 279503
rect 113982 279425 114266 279430
rect 111312 279399 114266 279425
rect 111312 279397 114034 279399
rect 114068 279397 114106 279399
rect 114140 279397 114178 279399
rect 114212 279397 114266 279399
rect 111312 279363 111340 279397
rect 111374 279363 111408 279397
rect 111442 279363 111476 279397
rect 111510 279363 111544 279397
rect 111578 279363 111612 279397
rect 111646 279363 111680 279397
rect 111714 279363 111748 279397
rect 111782 279363 111816 279397
rect 111850 279363 111884 279397
rect 111918 279363 111952 279397
rect 111986 279363 112020 279397
rect 112054 279363 112088 279397
rect 112122 279363 112156 279397
rect 112190 279363 112224 279397
rect 112258 279363 112292 279397
rect 112326 279363 112360 279397
rect 112394 279363 112428 279397
rect 112462 279363 112496 279397
rect 112530 279363 112564 279397
rect 112598 279363 112632 279397
rect 112666 279363 112700 279397
rect 112734 279363 112768 279397
rect 112802 279363 112836 279397
rect 112870 279363 112904 279397
rect 112938 279363 112972 279397
rect 113006 279363 113040 279397
rect 113074 279363 113108 279397
rect 113142 279363 113176 279397
rect 113210 279363 113244 279397
rect 113278 279363 113312 279397
rect 113346 279363 113380 279397
rect 113414 279363 113448 279397
rect 113482 279363 113516 279397
rect 113550 279363 113584 279397
rect 113618 279363 113652 279397
rect 113686 279363 113720 279397
rect 113754 279363 113788 279397
rect 113822 279363 113856 279397
rect 113890 279363 113924 279397
rect 113958 279363 113992 279397
rect 114026 279365 114034 279397
rect 114094 279365 114106 279397
rect 114162 279365 114178 279397
rect 114026 279363 114060 279365
rect 114094 279363 114128 279365
rect 114162 279363 114196 279365
rect 114230 279363 114266 279397
rect 114455 279403 114489 279435
rect 114930 279469 115275 279487
rect 114930 279435 115027 279469
rect 115061 279435 115144 279469
rect 115178 279435 115275 279469
rect 114930 279403 115275 279435
rect 115716 279469 115750 279503
rect 117577 279498 118871 279534
rect 115716 279403 115750 279435
rect 114455 279369 114537 279403
rect 114571 279369 114605 279403
rect 114639 279369 114673 279403
rect 114707 279369 114741 279403
rect 114775 279369 114809 279403
rect 114843 279369 114877 279403
rect 114911 279369 114945 279403
rect 114979 279369 115226 279403
rect 115260 279369 115294 279403
rect 115328 279369 115362 279403
rect 115396 279369 115430 279403
rect 115464 279369 115498 279403
rect 115532 279369 115566 279403
rect 115600 279369 115634 279403
rect 115668 279369 115750 279403
rect 115939 279425 116223 279430
rect 115939 279399 118893 279425
rect 115939 279397 115992 279399
rect 116026 279397 116064 279399
rect 116098 279397 116136 279399
rect 116170 279397 118893 279399
rect 111312 279335 114266 279363
rect 113036 279330 114266 279335
rect 113036 279238 114022 279330
rect 115061 279297 115144 279369
rect 115939 279363 115975 279397
rect 116026 279365 116043 279397
rect 116098 279365 116111 279397
rect 116170 279365 116179 279397
rect 116009 279363 116043 279365
rect 116077 279363 116111 279365
rect 116145 279363 116179 279365
rect 116213 279363 116247 279397
rect 116281 279363 116315 279397
rect 116349 279363 116383 279397
rect 116417 279363 116451 279397
rect 116485 279363 116519 279397
rect 116553 279363 116587 279397
rect 116621 279363 116655 279397
rect 116689 279363 116723 279397
rect 116757 279363 116791 279397
rect 116825 279363 116859 279397
rect 116893 279363 116927 279397
rect 116961 279363 116995 279397
rect 117029 279363 117063 279397
rect 117097 279363 117131 279397
rect 117165 279363 117199 279397
rect 117233 279363 117267 279397
rect 117301 279363 117335 279397
rect 117369 279363 117403 279397
rect 117437 279363 117471 279397
rect 117505 279363 117539 279397
rect 117573 279363 117607 279397
rect 117641 279363 117675 279397
rect 117709 279363 117743 279397
rect 117777 279363 117811 279397
rect 117845 279363 117879 279397
rect 117913 279363 117947 279397
rect 117981 279363 118015 279397
rect 118049 279363 118083 279397
rect 118117 279363 118151 279397
rect 118185 279363 118219 279397
rect 118253 279363 118287 279397
rect 118321 279363 118355 279397
rect 118389 279363 118423 279397
rect 118457 279363 118491 279397
rect 118525 279363 118559 279397
rect 118593 279363 118627 279397
rect 118661 279363 118695 279397
rect 118729 279363 118763 279397
rect 118797 279363 118831 279397
rect 118865 279363 118893 279397
rect 115939 279335 118893 279363
rect 115939 279330 117169 279335
rect 114455 279263 114537 279297
rect 114571 279263 114605 279297
rect 114639 279263 114673 279297
rect 114707 279263 114741 279297
rect 114775 279263 114809 279297
rect 114843 279263 114877 279297
rect 114911 279263 114945 279297
rect 114979 279263 115226 279297
rect 115260 279263 115294 279297
rect 115328 279263 115362 279297
rect 115396 279263 115430 279297
rect 115464 279263 115498 279297
rect 115532 279263 115566 279297
rect 115600 279263 115634 279297
rect 115668 279263 115750 279297
rect 111520 279200 112814 279236
rect 113036 279234 114246 279238
rect 113036 279233 114353 279234
rect 111520 279166 111547 279200
rect 111587 279166 111615 279200
rect 111659 279166 111683 279200
rect 111731 279166 111751 279200
rect 111803 279166 111819 279200
rect 111875 279166 111887 279200
rect 111947 279166 111955 279200
rect 112019 279166 112023 279200
rect 112125 279166 112129 279200
rect 112193 279166 112201 279200
rect 112261 279166 112273 279200
rect 112329 279166 112345 279200
rect 112397 279166 112417 279200
rect 112465 279166 112489 279200
rect 112533 279166 112561 279200
rect 112601 279166 112628 279200
rect 111452 279127 111486 279154
rect 111452 279057 111486 279091
rect 111452 278994 111486 279021
rect 112662 279127 112696 279154
rect 112662 279057 112696 279091
rect 112662 278994 112696 279021
rect 111520 278948 111547 278982
rect 111587 278948 111615 278982
rect 111659 278948 111683 278982
rect 111731 278948 111751 278982
rect 111803 278948 111819 278982
rect 111875 278948 111887 278982
rect 111947 278948 111955 278982
rect 112019 278948 112023 278982
rect 112125 278948 112129 278982
rect 112193 278948 112201 278982
rect 112261 278948 112273 278982
rect 112329 278948 112345 278982
rect 112397 278948 112417 278982
rect 112465 278948 112489 278982
rect 112533 278948 112561 278982
rect 112601 278948 112628 278982
rect 111334 278912 112628 278948
rect 112772 278916 112814 279200
rect 112966 279210 114353 279233
rect 112966 279208 114243 279210
rect 112966 279174 112993 279208
rect 113033 279174 113061 279208
rect 113105 279174 113129 279208
rect 113177 279174 113197 279208
rect 113249 279174 113265 279208
rect 113321 279174 113333 279208
rect 113393 279174 113401 279208
rect 113465 279174 113469 279208
rect 113571 279174 113575 279208
rect 113639 279174 113647 279208
rect 113707 279174 113719 279208
rect 113775 279174 113791 279208
rect 113843 279174 113863 279208
rect 113911 279174 113935 279208
rect 113979 279174 114007 279208
rect 114047 279204 114243 279208
rect 114047 279174 114074 279204
rect 112898 279115 112932 279162
rect 112898 279045 112932 279079
rect 112898 278962 112932 279009
rect 114108 279115 114142 279162
rect 114108 279045 114142 279079
rect 114108 278962 114142 279009
rect 114210 279108 114243 279204
rect 114345 279108 114353 279210
rect 114210 279084 114353 279108
rect 114455 279231 114489 279263
rect 114455 279163 114489 279197
rect 114652 279183 114862 279263
rect 114652 279149 114672 279183
rect 114738 279149 114740 279183
rect 114774 279149 114776 279183
rect 114842 279149 114862 279183
rect 114652 279148 114862 279149
rect 115027 279231 115178 279263
rect 115061 279197 115144 279231
rect 115027 279163 115178 279197
rect 114455 279095 114489 279129
rect 112966 278916 112993 278950
rect 113033 278916 113061 278950
rect 113105 278916 113129 278950
rect 113177 278916 113197 278950
rect 113249 278916 113265 278950
rect 113321 278916 113333 278950
rect 113393 278916 113401 278950
rect 113465 278916 113469 278950
rect 113571 278916 113575 278950
rect 113639 278916 113647 278950
rect 113707 278916 113719 278950
rect 113775 278916 113791 278950
rect 113843 278916 113863 278950
rect 113911 278916 113935 278950
rect 113979 278916 114007 278950
rect 114047 278916 114074 278950
rect 111334 278588 111376 278912
rect 112772 278882 114074 278916
rect 112772 278876 112832 278882
rect 111520 278840 112832 278876
rect 111520 278806 111547 278840
rect 111587 278806 111615 278840
rect 111659 278806 111683 278840
rect 111731 278806 111751 278840
rect 111803 278806 111819 278840
rect 111875 278806 111887 278840
rect 111947 278806 111955 278840
rect 112019 278806 112023 278840
rect 112125 278806 112129 278840
rect 112193 278806 112201 278840
rect 112261 278806 112273 278840
rect 112329 278806 112345 278840
rect 112397 278806 112417 278840
rect 112465 278806 112489 278840
rect 112533 278806 112561 278840
rect 112601 278806 112628 278840
rect 111452 278767 111486 278794
rect 111452 278697 111486 278731
rect 111452 278634 111486 278661
rect 112662 278767 112696 278794
rect 112662 278697 112696 278731
rect 112662 278634 112696 278661
rect 111520 278588 111547 278622
rect 111587 278588 111615 278622
rect 111659 278588 111683 278622
rect 111731 278588 111751 278622
rect 111803 278588 111819 278622
rect 111875 278588 111887 278622
rect 111947 278588 111955 278622
rect 112019 278588 112023 278622
rect 112125 278588 112129 278622
rect 112193 278588 112201 278622
rect 112261 278588 112273 278622
rect 112329 278588 112345 278622
rect 112397 278588 112417 278622
rect 112465 278588 112489 278622
rect 112533 278588 112561 278622
rect 112601 278588 112628 278622
rect 111334 278552 112628 278588
rect 111334 278228 111376 278552
rect 112772 278516 112832 278840
rect 114210 278818 114246 279084
rect 112966 278784 114246 278818
rect 114455 279027 114489 279061
rect 114455 278959 114489 278993
rect 114455 278891 114489 278925
rect 114455 278823 114489 278857
rect 112966 278750 112993 278784
rect 113033 278750 113061 278784
rect 113105 278750 113129 278784
rect 113177 278750 113197 278784
rect 113249 278750 113265 278784
rect 113321 278750 113333 278784
rect 113393 278750 113401 278784
rect 113465 278750 113469 278784
rect 113571 278750 113575 278784
rect 113639 278750 113647 278784
rect 113707 278750 113719 278784
rect 113775 278750 113791 278784
rect 113843 278750 113863 278784
rect 113911 278750 113935 278784
rect 113979 278750 114007 278784
rect 114047 278750 114074 278784
rect 114455 278755 114489 278789
rect 112898 278691 112932 278738
rect 112898 278621 112932 278655
rect 112898 278538 112932 278585
rect 114108 278691 114142 278738
rect 114108 278621 114142 278655
rect 114108 278538 114142 278585
rect 114455 278687 114489 278721
rect 114455 278619 114489 278653
rect 114455 278551 114489 278585
rect 111520 278494 112832 278516
rect 112966 278494 112993 278526
rect 111520 278492 112993 278494
rect 113033 278492 113061 278526
rect 113105 278492 113129 278526
rect 113177 278492 113197 278526
rect 113249 278492 113265 278526
rect 113321 278492 113333 278526
rect 113393 278492 113401 278526
rect 113465 278492 113469 278526
rect 113571 278492 113575 278526
rect 113639 278492 113647 278526
rect 113707 278492 113719 278526
rect 113775 278492 113791 278526
rect 113843 278492 113863 278526
rect 113911 278492 113935 278526
rect 113979 278492 114007 278526
rect 114047 278492 114074 278526
rect 111520 278480 114074 278492
rect 111520 278446 111547 278480
rect 111587 278446 111615 278480
rect 111659 278446 111683 278480
rect 111731 278446 111751 278480
rect 111803 278446 111819 278480
rect 111875 278446 111887 278480
rect 111947 278446 111955 278480
rect 112019 278446 112023 278480
rect 112125 278446 112129 278480
rect 112193 278446 112201 278480
rect 112261 278446 112273 278480
rect 112329 278446 112345 278480
rect 112397 278446 112417 278480
rect 112465 278446 112489 278480
rect 112533 278446 112561 278480
rect 112601 278446 112628 278480
rect 112744 278477 114074 278480
rect 114455 278483 114489 278517
rect 112744 278460 114396 278477
rect 111452 278407 111486 278434
rect 111452 278337 111486 278371
rect 111452 278274 111486 278301
rect 112662 278407 112696 278434
rect 112662 278337 112696 278371
rect 112662 278274 112696 278301
rect 111520 278228 111547 278262
rect 111587 278228 111615 278262
rect 111659 278228 111683 278262
rect 111731 278228 111751 278262
rect 111803 278228 111819 278262
rect 111875 278228 111887 278262
rect 111947 278228 111955 278262
rect 112019 278228 112023 278262
rect 112125 278228 112129 278262
rect 112193 278228 112201 278262
rect 112261 278228 112273 278262
rect 112329 278228 112345 278262
rect 112397 278228 112417 278262
rect 112465 278228 112489 278262
rect 112533 278228 112561 278262
rect 112601 278228 112628 278262
rect 111334 278192 112628 278228
rect 111334 277868 111376 278192
rect 112744 278156 112780 278460
rect 113892 278441 114396 278460
rect 111520 278120 112780 278156
rect 112832 278382 113264 278416
rect 112832 278374 113023 278382
rect 112832 278120 112872 278374
rect 112996 278348 113023 278374
rect 113063 278348 113091 278382
rect 113135 278348 113159 278382
rect 113207 278348 113227 278382
rect 113279 278348 113295 278382
rect 113351 278348 113363 278382
rect 113423 278348 113431 278382
rect 113495 278348 113499 278382
rect 113601 278348 113605 278382
rect 113669 278348 113677 278382
rect 113737 278348 113749 278382
rect 113805 278348 113821 278382
rect 113873 278348 113893 278382
rect 113941 278348 113965 278382
rect 114009 278348 114037 278382
rect 114077 278348 114104 278382
rect 112928 278313 112962 278336
rect 112928 278256 112962 278279
rect 114138 278313 114172 278336
rect 114138 278256 114172 278279
rect 114324 278285 114396 278441
rect 114324 278251 114342 278285
rect 114376 278251 114396 278285
rect 112996 278216 113023 278244
rect 112994 278210 113023 278216
rect 113063 278210 113091 278244
rect 113135 278210 113159 278244
rect 113207 278210 113227 278244
rect 113279 278210 113295 278244
rect 113351 278210 113363 278244
rect 113423 278210 113431 278244
rect 113495 278210 113499 278244
rect 113601 278210 113605 278244
rect 113669 278210 113677 278244
rect 113737 278210 113749 278244
rect 113805 278210 113821 278244
rect 113873 278210 113893 278244
rect 113941 278210 113965 278244
rect 114009 278210 114037 278244
rect 114077 278216 114104 278244
rect 114077 278210 114274 278216
rect 112994 278170 114274 278210
rect 114324 278203 114396 278251
rect 114455 278415 114489 278449
rect 114455 278347 114489 278381
rect 114455 278279 114489 278313
rect 114576 279098 114610 279137
rect 114576 279026 114610 279056
rect 114576 278954 114610 278988
rect 114576 278886 114610 278920
rect 114576 278818 114610 278848
rect 114576 278609 114610 278776
rect 114904 279098 114938 279137
rect 114904 279026 114938 279056
rect 114904 278954 114938 278988
rect 114904 278886 114938 278920
rect 114904 278818 114938 278848
rect 114653 278691 114672 278725
rect 114738 278691 114740 278725
rect 114774 278691 114776 278725
rect 114842 278691 114861 278725
rect 114904 278645 114938 278776
rect 115061 279129 115144 279163
rect 115343 279183 115553 279263
rect 115343 279149 115363 279183
rect 115429 279149 115431 279183
rect 115465 279149 115467 279183
rect 115533 279149 115553 279183
rect 115343 279148 115553 279149
rect 115716 279231 115750 279263
rect 116183 279238 117169 279330
rect 115959 279234 117169 279238
rect 115716 279163 115750 279197
rect 115027 279095 115178 279129
rect 115061 279061 115144 279095
rect 115027 279027 115178 279061
rect 115061 278993 115144 279027
rect 115027 278959 115178 278993
rect 115061 278925 115144 278959
rect 115027 278891 115178 278925
rect 115061 278857 115144 278891
rect 115027 278823 115178 278857
rect 115061 278789 115144 278823
rect 115027 278755 115178 278789
rect 115061 278721 115144 278755
rect 115027 278687 115178 278721
rect 115061 278653 115144 278687
rect 114865 278611 114970 278645
rect 114865 278609 114899 278611
rect 114576 278577 114899 278609
rect 114933 278577 114970 278611
rect 114576 278561 114970 278577
rect 114576 278424 114610 278561
rect 114865 278538 114970 278561
rect 115027 278619 115178 278653
rect 115267 279098 115301 279137
rect 115267 279026 115301 279056
rect 115267 278954 115301 278988
rect 115267 278886 115301 278920
rect 115267 278818 115301 278848
rect 115267 278645 115301 278776
rect 115595 279098 115629 279137
rect 115595 279026 115629 279056
rect 115595 278954 115629 278988
rect 115595 278886 115629 278920
rect 115595 278818 115629 278848
rect 115344 278691 115363 278725
rect 115429 278691 115431 278725
rect 115465 278691 115467 278725
rect 115533 278691 115552 278725
rect 115061 278585 115144 278619
rect 115027 278551 115178 278585
rect 114653 278463 114672 278497
rect 114738 278463 114740 278497
rect 114774 278463 114776 278497
rect 114842 278463 114861 278497
rect 114576 278354 114610 278388
rect 114576 278291 114610 278318
rect 114904 278424 114938 278538
rect 114904 278354 114938 278388
rect 114904 278291 114938 278318
rect 115061 278517 115144 278551
rect 115235 278611 115340 278645
rect 115235 278577 115271 278611
rect 115305 278609 115340 278611
rect 115595 278609 115629 278776
rect 115305 278577 115629 278609
rect 115235 278561 115629 278577
rect 115235 278538 115340 278561
rect 115027 278483 115178 278517
rect 115061 278449 115144 278483
rect 115027 278415 115178 278449
rect 115061 278381 115144 278415
rect 115027 278347 115178 278381
rect 115061 278313 115144 278347
rect 115027 278279 115178 278313
rect 115267 278424 115301 278538
rect 115344 278463 115363 278497
rect 115429 278463 115431 278497
rect 115465 278463 115467 278497
rect 115533 278463 115552 278497
rect 115267 278354 115301 278388
rect 115267 278291 115301 278318
rect 115595 278424 115629 278561
rect 115595 278354 115629 278388
rect 115595 278291 115629 278318
rect 115716 279095 115750 279129
rect 115852 279233 117169 279234
rect 115852 279210 117239 279233
rect 115852 279108 115860 279210
rect 115962 279208 117239 279210
rect 115962 279204 116158 279208
rect 115962 279108 115995 279204
rect 116131 279174 116158 279204
rect 116198 279174 116226 279208
rect 116270 279174 116294 279208
rect 116342 279174 116362 279208
rect 116414 279174 116430 279208
rect 116486 279174 116498 279208
rect 116558 279174 116566 279208
rect 116630 279174 116634 279208
rect 116736 279174 116740 279208
rect 116804 279174 116812 279208
rect 116872 279174 116884 279208
rect 116940 279174 116956 279208
rect 117008 279174 117028 279208
rect 117076 279174 117100 279208
rect 117144 279174 117172 279208
rect 117212 279174 117239 279208
rect 117391 279200 118685 279236
rect 115852 279084 115995 279108
rect 115716 279027 115750 279061
rect 115716 278959 115750 278993
rect 115716 278891 115750 278925
rect 115716 278823 115750 278857
rect 115716 278755 115750 278789
rect 115959 278818 115995 279084
rect 116063 279115 116097 279162
rect 116063 279045 116097 279079
rect 116063 278962 116097 279009
rect 117273 279115 117307 279162
rect 117273 279045 117307 279079
rect 117273 278962 117307 279009
rect 116131 278916 116158 278950
rect 116198 278916 116226 278950
rect 116270 278916 116294 278950
rect 116342 278916 116362 278950
rect 116414 278916 116430 278950
rect 116486 278916 116498 278950
rect 116558 278916 116566 278950
rect 116630 278916 116634 278950
rect 116736 278916 116740 278950
rect 116804 278916 116812 278950
rect 116872 278916 116884 278950
rect 116940 278916 116956 278950
rect 117008 278916 117028 278950
rect 117076 278916 117100 278950
rect 117144 278916 117172 278950
rect 117212 278916 117239 278950
rect 117391 278916 117433 279200
rect 117577 279166 117604 279200
rect 117644 279166 117672 279200
rect 117716 279166 117740 279200
rect 117788 279166 117808 279200
rect 117860 279166 117876 279200
rect 117932 279166 117944 279200
rect 118004 279166 118012 279200
rect 118076 279166 118080 279200
rect 118182 279166 118186 279200
rect 118250 279166 118258 279200
rect 118318 279166 118330 279200
rect 118386 279166 118402 279200
rect 118454 279166 118474 279200
rect 118522 279166 118546 279200
rect 118590 279166 118618 279200
rect 118658 279166 118685 279200
rect 117509 279127 117543 279154
rect 117509 279057 117543 279091
rect 117509 278994 117543 279021
rect 118719 279127 118753 279154
rect 118719 279057 118753 279091
rect 118719 278994 118753 279021
rect 116131 278882 117433 278916
rect 117577 278948 117604 278982
rect 117644 278948 117672 278982
rect 117716 278948 117740 278982
rect 117788 278948 117808 278982
rect 117860 278948 117876 278982
rect 117932 278948 117944 278982
rect 118004 278948 118012 278982
rect 118076 278948 118080 278982
rect 118182 278948 118186 278982
rect 118250 278948 118258 278982
rect 118318 278948 118330 278982
rect 118386 278948 118402 278982
rect 118454 278948 118474 278982
rect 118522 278948 118546 278982
rect 118590 278948 118618 278982
rect 118658 278948 118685 278982
rect 117577 278912 118871 278948
rect 117373 278876 117433 278882
rect 117373 278840 118685 278876
rect 115959 278784 117239 278818
rect 116131 278750 116158 278784
rect 116198 278750 116226 278784
rect 116270 278750 116294 278784
rect 116342 278750 116362 278784
rect 116414 278750 116430 278784
rect 116486 278750 116498 278784
rect 116558 278750 116566 278784
rect 116630 278750 116634 278784
rect 116736 278750 116740 278784
rect 116804 278750 116812 278784
rect 116872 278750 116884 278784
rect 116940 278750 116956 278784
rect 117008 278750 117028 278784
rect 117076 278750 117100 278784
rect 117144 278750 117172 278784
rect 117212 278750 117239 278784
rect 115716 278687 115750 278721
rect 115716 278619 115750 278653
rect 115716 278551 115750 278585
rect 116063 278691 116097 278738
rect 116063 278621 116097 278655
rect 116063 278538 116097 278585
rect 117273 278691 117307 278738
rect 117273 278621 117307 278655
rect 117273 278538 117307 278585
rect 115716 278483 115750 278517
rect 116131 278492 116158 278526
rect 116198 278492 116226 278526
rect 116270 278492 116294 278526
rect 116342 278492 116362 278526
rect 116414 278492 116430 278526
rect 116486 278492 116498 278526
rect 116558 278492 116566 278526
rect 116630 278492 116634 278526
rect 116736 278492 116740 278526
rect 116804 278492 116812 278526
rect 116872 278492 116884 278526
rect 116940 278492 116956 278526
rect 117008 278492 117028 278526
rect 117076 278492 117100 278526
rect 117144 278492 117172 278526
rect 117212 278494 117239 278526
rect 117373 278516 117433 278840
rect 117577 278806 117604 278840
rect 117644 278806 117672 278840
rect 117716 278806 117740 278840
rect 117788 278806 117808 278840
rect 117860 278806 117876 278840
rect 117932 278806 117944 278840
rect 118004 278806 118012 278840
rect 118076 278806 118080 278840
rect 118182 278806 118186 278840
rect 118250 278806 118258 278840
rect 118318 278806 118330 278840
rect 118386 278806 118402 278840
rect 118454 278806 118474 278840
rect 118522 278806 118546 278840
rect 118590 278806 118618 278840
rect 118658 278806 118685 278840
rect 117509 278767 117543 278794
rect 117509 278697 117543 278731
rect 117509 278634 117543 278661
rect 118719 278767 118753 278794
rect 118719 278697 118753 278731
rect 118719 278634 118753 278661
rect 117577 278588 117604 278622
rect 117644 278588 117672 278622
rect 117716 278588 117740 278622
rect 117788 278588 117808 278622
rect 117860 278588 117876 278622
rect 117932 278588 117944 278622
rect 118004 278588 118012 278622
rect 118076 278588 118080 278622
rect 118182 278588 118186 278622
rect 118250 278588 118258 278622
rect 118318 278588 118330 278622
rect 118386 278588 118402 278622
rect 118454 278588 118474 278622
rect 118522 278588 118546 278622
rect 118590 278588 118618 278622
rect 118658 278588 118685 278622
rect 118829 278588 118871 278912
rect 117577 278552 118871 278588
rect 117373 278494 118685 278516
rect 117212 278492 118685 278494
rect 116131 278480 118685 278492
rect 116131 278477 117461 278480
rect 115716 278415 115750 278449
rect 115716 278347 115750 278381
rect 115716 278279 115750 278313
rect 114455 278211 114489 278245
rect 111520 278086 111547 278120
rect 111587 278086 111615 278120
rect 111659 278086 111683 278120
rect 111731 278086 111751 278120
rect 111803 278086 111819 278120
rect 111875 278086 111887 278120
rect 111947 278086 111955 278120
rect 112019 278086 112023 278120
rect 112125 278086 112129 278120
rect 112193 278086 112201 278120
rect 112261 278086 112273 278120
rect 112329 278086 112345 278120
rect 112397 278086 112417 278120
rect 112465 278086 112489 278120
rect 112533 278086 112561 278120
rect 112601 278086 112628 278120
rect 112832 278084 113216 278120
rect 112832 278080 113023 278084
rect 111452 278047 111486 278074
rect 111452 277977 111486 278011
rect 111452 277914 111486 277941
rect 112662 278047 112696 278074
rect 112832 278052 112872 278080
rect 112996 278050 113023 278080
rect 113063 278050 113091 278084
rect 113135 278050 113159 278084
rect 113207 278050 113227 278084
rect 113279 278050 113295 278084
rect 113351 278050 113363 278084
rect 113423 278050 113431 278084
rect 113495 278050 113499 278084
rect 113601 278050 113605 278084
rect 113669 278050 113677 278084
rect 113737 278050 113749 278084
rect 113805 278050 113821 278084
rect 113873 278050 113893 278084
rect 113941 278050 113965 278084
rect 114009 278050 114037 278084
rect 114077 278050 114104 278084
rect 112662 277977 112696 278011
rect 112928 278015 112962 278038
rect 112928 277958 112962 277981
rect 114138 278015 114172 278038
rect 114138 277958 114172 277981
rect 112662 277914 112696 277941
rect 112996 277912 113023 277946
rect 113063 277912 113091 277946
rect 113135 277912 113159 277946
rect 113207 277912 113227 277946
rect 113279 277912 113295 277946
rect 113351 277912 113363 277946
rect 113423 277912 113431 277946
rect 113495 277912 113499 277946
rect 113601 277912 113605 277946
rect 113669 277912 113677 277946
rect 113737 277912 113749 277946
rect 113805 277912 113821 277946
rect 113873 277912 113893 277946
rect 113941 277912 113965 277946
rect 114009 277912 114037 277946
rect 114077 277912 114104 277946
rect 114234 277912 114274 278170
rect 114653 278245 114672 278279
rect 114738 278245 114740 278279
rect 114774 278245 114776 278279
rect 114842 278245 114861 278279
rect 114653 278208 114709 278245
rect 114805 278210 114861 278245
rect 115061 278245 115144 278279
rect 115027 278211 115178 278245
rect 114455 278143 114489 278177
rect 114455 278075 114489 278109
rect 114455 278007 114489 278041
rect 114455 277939 114489 277973
rect 112994 277905 114455 277912
rect 111520 277868 111547 277902
rect 111587 277868 111615 277902
rect 111659 277868 111683 277902
rect 111731 277868 111751 277902
rect 111803 277868 111819 277902
rect 111875 277868 111887 277902
rect 111947 277868 111955 277902
rect 112019 277868 112023 277902
rect 112125 277868 112129 277902
rect 112193 277868 112201 277902
rect 112261 277868 112273 277902
rect 112329 277868 112345 277902
rect 112397 277868 112417 277902
rect 112465 277868 112489 277902
rect 112533 277868 112561 277902
rect 112601 277868 112628 277902
rect 111334 277832 112628 277868
rect 112994 277871 114489 277905
rect 114538 278169 114709 278208
rect 114804 278188 114991 278210
rect 114538 278043 114576 278169
rect 114804 278154 114899 278188
rect 114933 278154 114991 278188
rect 114804 278125 114991 278154
rect 115061 278177 115144 278211
rect 115344 278245 115363 278279
rect 115429 278245 115431 278279
rect 115465 278245 115467 278279
rect 115533 278245 115552 278279
rect 115344 278210 115400 278245
rect 115027 278143 115178 278177
rect 114653 278055 114672 278089
rect 114738 278055 114740 278089
rect 114774 278055 114776 278089
rect 114842 278055 114861 278089
rect 114938 278043 114975 278125
rect 114538 278016 114610 278043
rect 114538 277980 114576 278016
rect 114538 277946 114610 277980
rect 114538 277910 114576 277946
rect 114538 277883 114610 277910
rect 114904 278016 114975 278043
rect 114938 277980 114975 278016
rect 114904 277946 114975 277980
rect 114938 277910 114975 277946
rect 114904 277883 114975 277910
rect 115061 278109 115144 278143
rect 115214 278188 115401 278210
rect 115214 278154 115271 278188
rect 115305 278154 115401 278188
rect 115496 278208 115552 278245
rect 115716 278211 115750 278245
rect 115496 278169 115667 278208
rect 115214 278125 115401 278154
rect 115027 278075 115178 278109
rect 115061 278041 115144 278075
rect 115027 278007 115178 278041
rect 115061 277973 115144 278007
rect 115027 277939 115178 277973
rect 115061 277905 115144 277939
rect 115027 277871 115178 277905
rect 115230 278043 115267 278125
rect 115344 278055 115363 278089
rect 115429 278055 115431 278089
rect 115465 278055 115467 278089
rect 115533 278055 115552 278089
rect 115629 278043 115667 278169
rect 115230 278016 115301 278043
rect 115230 277980 115267 278016
rect 115230 277946 115301 277980
rect 115230 277910 115267 277946
rect 115230 277883 115301 277910
rect 115595 278016 115667 278043
rect 115629 277980 115667 278016
rect 115595 277946 115667 277980
rect 115629 277910 115667 277946
rect 115595 277883 115667 277910
rect 115809 278460 117461 278477
rect 115809 278441 116313 278460
rect 115809 278285 115881 278441
rect 116941 278382 117373 278416
rect 116101 278348 116128 278382
rect 116168 278348 116196 278382
rect 116240 278348 116264 278382
rect 116312 278348 116332 278382
rect 116384 278348 116400 278382
rect 116456 278348 116468 278382
rect 116528 278348 116536 278382
rect 116600 278348 116604 278382
rect 116706 278348 116710 278382
rect 116774 278348 116782 278382
rect 116842 278348 116854 278382
rect 116910 278348 116926 278382
rect 116978 278348 116998 278382
rect 117046 278348 117070 278382
rect 117114 278348 117142 278382
rect 117182 278374 117373 278382
rect 117182 278348 117209 278374
rect 115809 278251 115828 278285
rect 115862 278251 115881 278285
rect 116033 278313 116067 278336
rect 116033 278256 116067 278279
rect 117243 278313 117277 278336
rect 117243 278256 117277 278279
rect 115809 278203 115881 278251
rect 116101 278216 116128 278244
rect 115931 278210 116128 278216
rect 116168 278210 116196 278244
rect 116240 278210 116264 278244
rect 116312 278210 116332 278244
rect 116384 278210 116400 278244
rect 116456 278210 116468 278244
rect 116528 278210 116536 278244
rect 116600 278210 116604 278244
rect 116706 278210 116710 278244
rect 116774 278210 116782 278244
rect 116842 278210 116854 278244
rect 116910 278210 116926 278244
rect 116978 278210 116998 278244
rect 117046 278210 117070 278244
rect 117114 278210 117142 278244
rect 117182 278216 117209 278244
rect 117182 278210 117211 278216
rect 115716 278143 115750 278177
rect 115716 278075 115750 278109
rect 115716 278007 115750 278041
rect 115716 277939 115750 277973
rect 115931 278170 117211 278210
rect 115931 277912 115971 278170
rect 117333 278120 117373 278374
rect 117425 278156 117461 278460
rect 117577 278446 117604 278480
rect 117644 278446 117672 278480
rect 117716 278446 117740 278480
rect 117788 278446 117808 278480
rect 117860 278446 117876 278480
rect 117932 278446 117944 278480
rect 118004 278446 118012 278480
rect 118076 278446 118080 278480
rect 118182 278446 118186 278480
rect 118250 278446 118258 278480
rect 118318 278446 118330 278480
rect 118386 278446 118402 278480
rect 118454 278446 118474 278480
rect 118522 278446 118546 278480
rect 118590 278446 118618 278480
rect 118658 278446 118685 278480
rect 117509 278407 117543 278434
rect 117509 278337 117543 278371
rect 117509 278274 117543 278301
rect 118719 278407 118753 278434
rect 118719 278337 118753 278371
rect 118719 278274 118753 278301
rect 117577 278228 117604 278262
rect 117644 278228 117672 278262
rect 117716 278228 117740 278262
rect 117788 278228 117808 278262
rect 117860 278228 117876 278262
rect 117932 278228 117944 278262
rect 118004 278228 118012 278262
rect 118076 278228 118080 278262
rect 118182 278228 118186 278262
rect 118250 278228 118258 278262
rect 118318 278228 118330 278262
rect 118386 278228 118402 278262
rect 118454 278228 118474 278262
rect 118522 278228 118546 278262
rect 118590 278228 118618 278262
rect 118658 278228 118685 278262
rect 118829 278228 118871 278552
rect 117577 278192 118871 278228
rect 117425 278120 118685 278156
rect 116989 278084 117373 278120
rect 117577 278086 117604 278120
rect 117644 278086 117672 278120
rect 117716 278086 117740 278120
rect 117788 278086 117808 278120
rect 117860 278086 117876 278120
rect 117932 278086 117944 278120
rect 118004 278086 118012 278120
rect 118076 278086 118080 278120
rect 118182 278086 118186 278120
rect 118250 278086 118258 278120
rect 118318 278086 118330 278120
rect 118386 278086 118402 278120
rect 118454 278086 118474 278120
rect 118522 278086 118546 278120
rect 118590 278086 118618 278120
rect 118658 278086 118685 278120
rect 116101 278050 116128 278084
rect 116168 278050 116196 278084
rect 116240 278050 116264 278084
rect 116312 278050 116332 278084
rect 116384 278050 116400 278084
rect 116456 278050 116468 278084
rect 116528 278050 116536 278084
rect 116600 278050 116604 278084
rect 116706 278050 116710 278084
rect 116774 278050 116782 278084
rect 116842 278050 116854 278084
rect 116910 278050 116926 278084
rect 116978 278050 116998 278084
rect 117046 278050 117070 278084
rect 117114 278050 117142 278084
rect 117182 278080 117373 278084
rect 117182 278050 117209 278080
rect 117333 278052 117373 278080
rect 117509 278047 117543 278074
rect 116033 278015 116067 278038
rect 116033 277958 116067 277981
rect 117243 278015 117277 278038
rect 117243 277958 117277 277981
rect 117509 277977 117543 278011
rect 116101 277912 116128 277946
rect 116168 277912 116196 277946
rect 116240 277912 116264 277946
rect 116312 277912 116332 277946
rect 116384 277912 116400 277946
rect 116456 277912 116468 277946
rect 116528 277912 116536 277946
rect 116600 277912 116604 277946
rect 116706 277912 116710 277946
rect 116774 277912 116782 277946
rect 116842 277912 116854 277946
rect 116910 277912 116926 277946
rect 116978 277912 116998 277946
rect 117046 277912 117070 277946
rect 117114 277912 117142 277946
rect 117182 277912 117209 277946
rect 117509 277914 117543 277941
rect 118719 278047 118753 278074
rect 118719 277977 118753 278011
rect 118719 277914 118753 277941
rect 115750 277905 117211 277912
rect 115716 277871 117211 277905
rect 112994 277866 114455 277871
rect 114653 277837 114672 277871
rect 114738 277837 114740 277871
rect 114774 277837 114776 277871
rect 114842 277837 114861 277871
rect 115061 277837 115144 277871
rect 115344 277837 115363 277871
rect 115429 277837 115431 277871
rect 115465 277837 115467 277871
rect 115533 277837 115552 277871
rect 115750 277866 117211 277871
rect 117577 277868 117604 277902
rect 117644 277868 117672 277902
rect 117716 277868 117740 277902
rect 117788 277868 117808 277902
rect 117860 277868 117876 277902
rect 117932 277868 117944 277902
rect 118004 277868 118012 277902
rect 118076 277868 118080 277902
rect 118182 277868 118186 277902
rect 118250 277868 118258 277902
rect 118318 277868 118330 277902
rect 118386 277868 118402 277902
rect 118454 277868 118474 277902
rect 118522 277868 118546 277902
rect 118590 277868 118618 277902
rect 118658 277868 118685 277902
rect 118829 277868 118871 278192
rect 114455 277803 114489 277837
rect 115027 277821 115178 277837
rect 113982 277759 114266 277764
rect 111312 277733 114266 277759
rect 111312 277731 114034 277733
rect 114068 277731 114106 277733
rect 114140 277731 114178 277733
rect 114212 277731 114266 277733
rect 111312 277697 111340 277731
rect 111374 277697 111408 277731
rect 111442 277697 111476 277731
rect 111510 277697 111544 277731
rect 111578 277697 111612 277731
rect 111646 277697 111680 277731
rect 111714 277697 111748 277731
rect 111782 277697 111816 277731
rect 111850 277697 111884 277731
rect 111918 277697 111952 277731
rect 111986 277697 112020 277731
rect 112054 277697 112088 277731
rect 112122 277697 112156 277731
rect 112190 277697 112224 277731
rect 112258 277697 112292 277731
rect 112326 277697 112360 277731
rect 112394 277697 112428 277731
rect 112462 277697 112496 277731
rect 112530 277697 112564 277731
rect 112598 277697 112632 277731
rect 112666 277697 112700 277731
rect 112734 277697 112768 277731
rect 112802 277697 112836 277731
rect 112870 277697 112904 277731
rect 112938 277697 112972 277731
rect 113006 277697 113040 277731
rect 113074 277697 113108 277731
rect 113142 277697 113176 277731
rect 113210 277697 113244 277731
rect 113278 277697 113312 277731
rect 113346 277697 113380 277731
rect 113414 277697 113448 277731
rect 113482 277697 113516 277731
rect 113550 277697 113584 277731
rect 113618 277697 113652 277731
rect 113686 277697 113720 277731
rect 113754 277697 113788 277731
rect 113822 277697 113856 277731
rect 113890 277697 113924 277731
rect 113958 277697 113992 277731
rect 114026 277699 114034 277731
rect 114094 277699 114106 277731
rect 114162 277699 114178 277731
rect 114026 277697 114060 277699
rect 114094 277697 114128 277699
rect 114162 277697 114196 277699
rect 114230 277697 114266 277731
rect 114455 277737 114489 277769
rect 114930 277803 115275 277821
rect 114930 277769 115027 277803
rect 115061 277769 115144 277803
rect 115178 277769 115275 277803
rect 114930 277737 115275 277769
rect 115716 277803 115750 277837
rect 117577 277832 118871 277868
rect 115716 277737 115750 277769
rect 114455 277703 114537 277737
rect 114571 277703 114605 277737
rect 114639 277703 114673 277737
rect 114707 277703 114741 277737
rect 114775 277703 114809 277737
rect 114843 277703 114877 277737
rect 114911 277703 114945 277737
rect 114979 277703 115226 277737
rect 115260 277703 115294 277737
rect 115328 277703 115362 277737
rect 115396 277703 115430 277737
rect 115464 277703 115498 277737
rect 115532 277703 115566 277737
rect 115600 277703 115634 277737
rect 115668 277703 115750 277737
rect 115939 277759 116223 277764
rect 115939 277733 118893 277759
rect 115939 277731 115992 277733
rect 116026 277731 116064 277733
rect 116098 277731 116136 277733
rect 116170 277731 118893 277733
rect 111312 277669 114266 277697
rect 113036 277664 114266 277669
rect 113036 277572 114022 277664
rect 115061 277631 115144 277703
rect 115939 277697 115975 277731
rect 116026 277699 116043 277731
rect 116098 277699 116111 277731
rect 116170 277699 116179 277731
rect 116009 277697 116043 277699
rect 116077 277697 116111 277699
rect 116145 277697 116179 277699
rect 116213 277697 116247 277731
rect 116281 277697 116315 277731
rect 116349 277697 116383 277731
rect 116417 277697 116451 277731
rect 116485 277697 116519 277731
rect 116553 277697 116587 277731
rect 116621 277697 116655 277731
rect 116689 277697 116723 277731
rect 116757 277697 116791 277731
rect 116825 277697 116859 277731
rect 116893 277697 116927 277731
rect 116961 277697 116995 277731
rect 117029 277697 117063 277731
rect 117097 277697 117131 277731
rect 117165 277697 117199 277731
rect 117233 277697 117267 277731
rect 117301 277697 117335 277731
rect 117369 277697 117403 277731
rect 117437 277697 117471 277731
rect 117505 277697 117539 277731
rect 117573 277697 117607 277731
rect 117641 277697 117675 277731
rect 117709 277697 117743 277731
rect 117777 277697 117811 277731
rect 117845 277697 117879 277731
rect 117913 277697 117947 277731
rect 117981 277697 118015 277731
rect 118049 277697 118083 277731
rect 118117 277697 118151 277731
rect 118185 277697 118219 277731
rect 118253 277697 118287 277731
rect 118321 277697 118355 277731
rect 118389 277697 118423 277731
rect 118457 277697 118491 277731
rect 118525 277697 118559 277731
rect 118593 277697 118627 277731
rect 118661 277697 118695 277731
rect 118729 277697 118763 277731
rect 118797 277697 118831 277731
rect 118865 277697 118893 277731
rect 115939 277669 118893 277697
rect 115939 277664 117169 277669
rect 114455 277597 114537 277631
rect 114571 277597 114605 277631
rect 114639 277597 114673 277631
rect 114707 277597 114741 277631
rect 114775 277597 114809 277631
rect 114843 277597 114877 277631
rect 114911 277597 114945 277631
rect 114979 277597 115226 277631
rect 115260 277597 115294 277631
rect 115328 277597 115362 277631
rect 115396 277597 115430 277631
rect 115464 277597 115498 277631
rect 115532 277597 115566 277631
rect 115600 277597 115634 277631
rect 115668 277597 115750 277631
rect 111520 277534 112814 277570
rect 113036 277568 114246 277572
rect 113036 277567 114353 277568
rect 111520 277500 111547 277534
rect 111587 277500 111615 277534
rect 111659 277500 111683 277534
rect 111731 277500 111751 277534
rect 111803 277500 111819 277534
rect 111875 277500 111887 277534
rect 111947 277500 111955 277534
rect 112019 277500 112023 277534
rect 112125 277500 112129 277534
rect 112193 277500 112201 277534
rect 112261 277500 112273 277534
rect 112329 277500 112345 277534
rect 112397 277500 112417 277534
rect 112465 277500 112489 277534
rect 112533 277500 112561 277534
rect 112601 277500 112628 277534
rect 111452 277461 111486 277488
rect 111452 277391 111486 277425
rect 111452 277328 111486 277355
rect 112662 277461 112696 277488
rect 112662 277391 112696 277425
rect 112662 277328 112696 277355
rect 111520 277282 111547 277316
rect 111587 277282 111615 277316
rect 111659 277282 111683 277316
rect 111731 277282 111751 277316
rect 111803 277282 111819 277316
rect 111875 277282 111887 277316
rect 111947 277282 111955 277316
rect 112019 277282 112023 277316
rect 112125 277282 112129 277316
rect 112193 277282 112201 277316
rect 112261 277282 112273 277316
rect 112329 277282 112345 277316
rect 112397 277282 112417 277316
rect 112465 277282 112489 277316
rect 112533 277282 112561 277316
rect 112601 277282 112628 277316
rect 111334 277246 112628 277282
rect 112772 277250 112814 277534
rect 112966 277544 114353 277567
rect 112966 277542 114243 277544
rect 112966 277508 112993 277542
rect 113033 277508 113061 277542
rect 113105 277508 113129 277542
rect 113177 277508 113197 277542
rect 113249 277508 113265 277542
rect 113321 277508 113333 277542
rect 113393 277508 113401 277542
rect 113465 277508 113469 277542
rect 113571 277508 113575 277542
rect 113639 277508 113647 277542
rect 113707 277508 113719 277542
rect 113775 277508 113791 277542
rect 113843 277508 113863 277542
rect 113911 277508 113935 277542
rect 113979 277508 114007 277542
rect 114047 277538 114243 277542
rect 114047 277508 114074 277538
rect 112898 277449 112932 277496
rect 112898 277379 112932 277413
rect 112898 277296 112932 277343
rect 114108 277449 114142 277496
rect 114108 277379 114142 277413
rect 114108 277296 114142 277343
rect 114210 277442 114243 277538
rect 114345 277442 114353 277544
rect 114210 277418 114353 277442
rect 114455 277565 114489 277597
rect 114455 277497 114489 277531
rect 114652 277517 114862 277597
rect 114652 277483 114672 277517
rect 114738 277483 114740 277517
rect 114774 277483 114776 277517
rect 114842 277483 114862 277517
rect 114652 277482 114862 277483
rect 115027 277565 115178 277597
rect 115061 277531 115144 277565
rect 115027 277497 115178 277531
rect 114455 277429 114489 277463
rect 112966 277250 112993 277284
rect 113033 277250 113061 277284
rect 113105 277250 113129 277284
rect 113177 277250 113197 277284
rect 113249 277250 113265 277284
rect 113321 277250 113333 277284
rect 113393 277250 113401 277284
rect 113465 277250 113469 277284
rect 113571 277250 113575 277284
rect 113639 277250 113647 277284
rect 113707 277250 113719 277284
rect 113775 277250 113791 277284
rect 113843 277250 113863 277284
rect 113911 277250 113935 277284
rect 113979 277250 114007 277284
rect 114047 277250 114074 277284
rect 111334 276922 111376 277246
rect 112772 277216 114074 277250
rect 112772 277210 112832 277216
rect 111520 277174 112832 277210
rect 111520 277140 111547 277174
rect 111587 277140 111615 277174
rect 111659 277140 111683 277174
rect 111731 277140 111751 277174
rect 111803 277140 111819 277174
rect 111875 277140 111887 277174
rect 111947 277140 111955 277174
rect 112019 277140 112023 277174
rect 112125 277140 112129 277174
rect 112193 277140 112201 277174
rect 112261 277140 112273 277174
rect 112329 277140 112345 277174
rect 112397 277140 112417 277174
rect 112465 277140 112489 277174
rect 112533 277140 112561 277174
rect 112601 277140 112628 277174
rect 111452 277101 111486 277128
rect 111452 277031 111486 277065
rect 111452 276968 111486 276995
rect 112662 277101 112696 277128
rect 112662 277031 112696 277065
rect 112662 276968 112696 276995
rect 111520 276922 111547 276956
rect 111587 276922 111615 276956
rect 111659 276922 111683 276956
rect 111731 276922 111751 276956
rect 111803 276922 111819 276956
rect 111875 276922 111887 276956
rect 111947 276922 111955 276956
rect 112019 276922 112023 276956
rect 112125 276922 112129 276956
rect 112193 276922 112201 276956
rect 112261 276922 112273 276956
rect 112329 276922 112345 276956
rect 112397 276922 112417 276956
rect 112465 276922 112489 276956
rect 112533 276922 112561 276956
rect 112601 276922 112628 276956
rect 111334 276886 112628 276922
rect 111334 276562 111376 276886
rect 112772 276850 112832 277174
rect 114210 277152 114246 277418
rect 112966 277118 114246 277152
rect 114455 277361 114489 277395
rect 114455 277293 114489 277327
rect 114455 277225 114489 277259
rect 114455 277157 114489 277191
rect 112966 277084 112993 277118
rect 113033 277084 113061 277118
rect 113105 277084 113129 277118
rect 113177 277084 113197 277118
rect 113249 277084 113265 277118
rect 113321 277084 113333 277118
rect 113393 277084 113401 277118
rect 113465 277084 113469 277118
rect 113571 277084 113575 277118
rect 113639 277084 113647 277118
rect 113707 277084 113719 277118
rect 113775 277084 113791 277118
rect 113843 277084 113863 277118
rect 113911 277084 113935 277118
rect 113979 277084 114007 277118
rect 114047 277084 114074 277118
rect 114455 277089 114489 277123
rect 112898 277025 112932 277072
rect 112898 276955 112932 276989
rect 112898 276872 112932 276919
rect 114108 277025 114142 277072
rect 114108 276955 114142 276989
rect 114108 276872 114142 276919
rect 114455 277021 114489 277055
rect 114455 276953 114489 276987
rect 114455 276885 114489 276919
rect 111520 276828 112832 276850
rect 112966 276828 112993 276860
rect 111520 276826 112993 276828
rect 113033 276826 113061 276860
rect 113105 276826 113129 276860
rect 113177 276826 113197 276860
rect 113249 276826 113265 276860
rect 113321 276826 113333 276860
rect 113393 276826 113401 276860
rect 113465 276826 113469 276860
rect 113571 276826 113575 276860
rect 113639 276826 113647 276860
rect 113707 276826 113719 276860
rect 113775 276826 113791 276860
rect 113843 276826 113863 276860
rect 113911 276826 113935 276860
rect 113979 276826 114007 276860
rect 114047 276826 114074 276860
rect 111520 276814 114074 276826
rect 111520 276780 111547 276814
rect 111587 276780 111615 276814
rect 111659 276780 111683 276814
rect 111731 276780 111751 276814
rect 111803 276780 111819 276814
rect 111875 276780 111887 276814
rect 111947 276780 111955 276814
rect 112019 276780 112023 276814
rect 112125 276780 112129 276814
rect 112193 276780 112201 276814
rect 112261 276780 112273 276814
rect 112329 276780 112345 276814
rect 112397 276780 112417 276814
rect 112465 276780 112489 276814
rect 112533 276780 112561 276814
rect 112601 276780 112628 276814
rect 112744 276811 114074 276814
rect 114455 276817 114489 276851
rect 112744 276794 114396 276811
rect 111452 276741 111486 276768
rect 111452 276671 111486 276705
rect 111452 276608 111486 276635
rect 112662 276741 112696 276768
rect 112662 276671 112696 276705
rect 112662 276608 112696 276635
rect 111520 276562 111547 276596
rect 111587 276562 111615 276596
rect 111659 276562 111683 276596
rect 111731 276562 111751 276596
rect 111803 276562 111819 276596
rect 111875 276562 111887 276596
rect 111947 276562 111955 276596
rect 112019 276562 112023 276596
rect 112125 276562 112129 276596
rect 112193 276562 112201 276596
rect 112261 276562 112273 276596
rect 112329 276562 112345 276596
rect 112397 276562 112417 276596
rect 112465 276562 112489 276596
rect 112533 276562 112561 276596
rect 112601 276562 112628 276596
rect 111334 276526 112628 276562
rect 111334 276202 111376 276526
rect 112744 276490 112780 276794
rect 113892 276775 114396 276794
rect 111520 276454 112780 276490
rect 112832 276716 113264 276750
rect 112832 276708 113023 276716
rect 112832 276454 112872 276708
rect 112996 276682 113023 276708
rect 113063 276682 113091 276716
rect 113135 276682 113159 276716
rect 113207 276682 113227 276716
rect 113279 276682 113295 276716
rect 113351 276682 113363 276716
rect 113423 276682 113431 276716
rect 113495 276682 113499 276716
rect 113601 276682 113605 276716
rect 113669 276682 113677 276716
rect 113737 276682 113749 276716
rect 113805 276682 113821 276716
rect 113873 276682 113893 276716
rect 113941 276682 113965 276716
rect 114009 276682 114037 276716
rect 114077 276682 114104 276716
rect 112928 276647 112962 276670
rect 112928 276590 112962 276613
rect 114138 276647 114172 276670
rect 114138 276590 114172 276613
rect 114324 276619 114396 276775
rect 114324 276585 114342 276619
rect 114376 276585 114396 276619
rect 112996 276550 113023 276578
rect 112994 276544 113023 276550
rect 113063 276544 113091 276578
rect 113135 276544 113159 276578
rect 113207 276544 113227 276578
rect 113279 276544 113295 276578
rect 113351 276544 113363 276578
rect 113423 276544 113431 276578
rect 113495 276544 113499 276578
rect 113601 276544 113605 276578
rect 113669 276544 113677 276578
rect 113737 276544 113749 276578
rect 113805 276544 113821 276578
rect 113873 276544 113893 276578
rect 113941 276544 113965 276578
rect 114009 276544 114037 276578
rect 114077 276550 114104 276578
rect 114077 276544 114274 276550
rect 112994 276504 114274 276544
rect 114324 276537 114396 276585
rect 114455 276749 114489 276783
rect 114455 276681 114489 276715
rect 114455 276613 114489 276647
rect 114576 277432 114610 277471
rect 114576 277360 114610 277390
rect 114576 277288 114610 277322
rect 114576 277220 114610 277254
rect 114576 277152 114610 277182
rect 114576 276943 114610 277110
rect 114904 277432 114938 277471
rect 114904 277360 114938 277390
rect 114904 277288 114938 277322
rect 114904 277220 114938 277254
rect 114904 277152 114938 277182
rect 114653 277025 114672 277059
rect 114738 277025 114740 277059
rect 114774 277025 114776 277059
rect 114842 277025 114861 277059
rect 114904 276979 114938 277110
rect 115061 277463 115144 277497
rect 115343 277517 115553 277597
rect 115343 277483 115363 277517
rect 115429 277483 115431 277517
rect 115465 277483 115467 277517
rect 115533 277483 115553 277517
rect 115343 277482 115553 277483
rect 115716 277565 115750 277597
rect 116183 277572 117169 277664
rect 115959 277568 117169 277572
rect 115716 277497 115750 277531
rect 115027 277429 115178 277463
rect 115061 277395 115144 277429
rect 115027 277361 115178 277395
rect 115061 277327 115144 277361
rect 115027 277293 115178 277327
rect 115061 277259 115144 277293
rect 115027 277225 115178 277259
rect 115061 277191 115144 277225
rect 115027 277157 115178 277191
rect 115061 277123 115144 277157
rect 115027 277089 115178 277123
rect 115061 277055 115144 277089
rect 115027 277021 115178 277055
rect 115061 276987 115144 277021
rect 114865 276945 114970 276979
rect 114865 276943 114899 276945
rect 114576 276911 114899 276943
rect 114933 276911 114970 276945
rect 114576 276895 114970 276911
rect 114576 276758 114610 276895
rect 114865 276872 114970 276895
rect 115027 276953 115178 276987
rect 115267 277432 115301 277471
rect 115267 277360 115301 277390
rect 115267 277288 115301 277322
rect 115267 277220 115301 277254
rect 115267 277152 115301 277182
rect 115267 276979 115301 277110
rect 115595 277432 115629 277471
rect 115595 277360 115629 277390
rect 115595 277288 115629 277322
rect 115595 277220 115629 277254
rect 115595 277152 115629 277182
rect 115344 277025 115363 277059
rect 115429 277025 115431 277059
rect 115465 277025 115467 277059
rect 115533 277025 115552 277059
rect 115061 276919 115144 276953
rect 115027 276885 115178 276919
rect 114653 276797 114672 276831
rect 114738 276797 114740 276831
rect 114774 276797 114776 276831
rect 114842 276797 114861 276831
rect 114576 276688 114610 276722
rect 114576 276625 114610 276652
rect 114904 276758 114938 276872
rect 114904 276688 114938 276722
rect 114904 276625 114938 276652
rect 115061 276851 115144 276885
rect 115235 276945 115340 276979
rect 115235 276911 115271 276945
rect 115305 276943 115340 276945
rect 115595 276943 115629 277110
rect 115305 276911 115629 276943
rect 115235 276895 115629 276911
rect 115235 276872 115340 276895
rect 115027 276817 115178 276851
rect 115061 276783 115144 276817
rect 115027 276749 115178 276783
rect 115061 276715 115144 276749
rect 115027 276681 115178 276715
rect 115061 276647 115144 276681
rect 115027 276613 115178 276647
rect 115267 276758 115301 276872
rect 115344 276797 115363 276831
rect 115429 276797 115431 276831
rect 115465 276797 115467 276831
rect 115533 276797 115552 276831
rect 115267 276688 115301 276722
rect 115267 276625 115301 276652
rect 115595 276758 115629 276895
rect 115595 276688 115629 276722
rect 115595 276625 115629 276652
rect 115716 277429 115750 277463
rect 115852 277567 117169 277568
rect 115852 277544 117239 277567
rect 115852 277442 115860 277544
rect 115962 277542 117239 277544
rect 115962 277538 116158 277542
rect 115962 277442 115995 277538
rect 116131 277508 116158 277538
rect 116198 277508 116226 277542
rect 116270 277508 116294 277542
rect 116342 277508 116362 277542
rect 116414 277508 116430 277542
rect 116486 277508 116498 277542
rect 116558 277508 116566 277542
rect 116630 277508 116634 277542
rect 116736 277508 116740 277542
rect 116804 277508 116812 277542
rect 116872 277508 116884 277542
rect 116940 277508 116956 277542
rect 117008 277508 117028 277542
rect 117076 277508 117100 277542
rect 117144 277508 117172 277542
rect 117212 277508 117239 277542
rect 117391 277534 118685 277570
rect 115852 277418 115995 277442
rect 115716 277361 115750 277395
rect 115716 277293 115750 277327
rect 115716 277225 115750 277259
rect 115716 277157 115750 277191
rect 115716 277089 115750 277123
rect 115959 277152 115995 277418
rect 116063 277449 116097 277496
rect 116063 277379 116097 277413
rect 116063 277296 116097 277343
rect 117273 277449 117307 277496
rect 117273 277379 117307 277413
rect 117273 277296 117307 277343
rect 116131 277250 116158 277284
rect 116198 277250 116226 277284
rect 116270 277250 116294 277284
rect 116342 277250 116362 277284
rect 116414 277250 116430 277284
rect 116486 277250 116498 277284
rect 116558 277250 116566 277284
rect 116630 277250 116634 277284
rect 116736 277250 116740 277284
rect 116804 277250 116812 277284
rect 116872 277250 116884 277284
rect 116940 277250 116956 277284
rect 117008 277250 117028 277284
rect 117076 277250 117100 277284
rect 117144 277250 117172 277284
rect 117212 277250 117239 277284
rect 117391 277250 117433 277534
rect 117577 277500 117604 277534
rect 117644 277500 117672 277534
rect 117716 277500 117740 277534
rect 117788 277500 117808 277534
rect 117860 277500 117876 277534
rect 117932 277500 117944 277534
rect 118004 277500 118012 277534
rect 118076 277500 118080 277534
rect 118182 277500 118186 277534
rect 118250 277500 118258 277534
rect 118318 277500 118330 277534
rect 118386 277500 118402 277534
rect 118454 277500 118474 277534
rect 118522 277500 118546 277534
rect 118590 277500 118618 277534
rect 118658 277500 118685 277534
rect 117509 277461 117543 277488
rect 117509 277391 117543 277425
rect 117509 277328 117543 277355
rect 118719 277461 118753 277488
rect 118719 277391 118753 277425
rect 118719 277328 118753 277355
rect 116131 277216 117433 277250
rect 117577 277282 117604 277316
rect 117644 277282 117672 277316
rect 117716 277282 117740 277316
rect 117788 277282 117808 277316
rect 117860 277282 117876 277316
rect 117932 277282 117944 277316
rect 118004 277282 118012 277316
rect 118076 277282 118080 277316
rect 118182 277282 118186 277316
rect 118250 277282 118258 277316
rect 118318 277282 118330 277316
rect 118386 277282 118402 277316
rect 118454 277282 118474 277316
rect 118522 277282 118546 277316
rect 118590 277282 118618 277316
rect 118658 277282 118685 277316
rect 117577 277246 118871 277282
rect 117373 277210 117433 277216
rect 117373 277174 118685 277210
rect 115959 277118 117239 277152
rect 116131 277084 116158 277118
rect 116198 277084 116226 277118
rect 116270 277084 116294 277118
rect 116342 277084 116362 277118
rect 116414 277084 116430 277118
rect 116486 277084 116498 277118
rect 116558 277084 116566 277118
rect 116630 277084 116634 277118
rect 116736 277084 116740 277118
rect 116804 277084 116812 277118
rect 116872 277084 116884 277118
rect 116940 277084 116956 277118
rect 117008 277084 117028 277118
rect 117076 277084 117100 277118
rect 117144 277084 117172 277118
rect 117212 277084 117239 277118
rect 115716 277021 115750 277055
rect 115716 276953 115750 276987
rect 115716 276885 115750 276919
rect 116063 277025 116097 277072
rect 116063 276955 116097 276989
rect 116063 276872 116097 276919
rect 117273 277025 117307 277072
rect 117273 276955 117307 276989
rect 117273 276872 117307 276919
rect 115716 276817 115750 276851
rect 116131 276826 116158 276860
rect 116198 276826 116226 276860
rect 116270 276826 116294 276860
rect 116342 276826 116362 276860
rect 116414 276826 116430 276860
rect 116486 276826 116498 276860
rect 116558 276826 116566 276860
rect 116630 276826 116634 276860
rect 116736 276826 116740 276860
rect 116804 276826 116812 276860
rect 116872 276826 116884 276860
rect 116940 276826 116956 276860
rect 117008 276826 117028 276860
rect 117076 276826 117100 276860
rect 117144 276826 117172 276860
rect 117212 276828 117239 276860
rect 117373 276850 117433 277174
rect 117577 277140 117604 277174
rect 117644 277140 117672 277174
rect 117716 277140 117740 277174
rect 117788 277140 117808 277174
rect 117860 277140 117876 277174
rect 117932 277140 117944 277174
rect 118004 277140 118012 277174
rect 118076 277140 118080 277174
rect 118182 277140 118186 277174
rect 118250 277140 118258 277174
rect 118318 277140 118330 277174
rect 118386 277140 118402 277174
rect 118454 277140 118474 277174
rect 118522 277140 118546 277174
rect 118590 277140 118618 277174
rect 118658 277140 118685 277174
rect 117509 277101 117543 277128
rect 117509 277031 117543 277065
rect 117509 276968 117543 276995
rect 118719 277101 118753 277128
rect 118719 277031 118753 277065
rect 118719 276968 118753 276995
rect 117577 276922 117604 276956
rect 117644 276922 117672 276956
rect 117716 276922 117740 276956
rect 117788 276922 117808 276956
rect 117860 276922 117876 276956
rect 117932 276922 117944 276956
rect 118004 276922 118012 276956
rect 118076 276922 118080 276956
rect 118182 276922 118186 276956
rect 118250 276922 118258 276956
rect 118318 276922 118330 276956
rect 118386 276922 118402 276956
rect 118454 276922 118474 276956
rect 118522 276922 118546 276956
rect 118590 276922 118618 276956
rect 118658 276922 118685 276956
rect 118829 276922 118871 277246
rect 117577 276886 118871 276922
rect 117373 276828 118685 276850
rect 117212 276826 118685 276828
rect 116131 276814 118685 276826
rect 116131 276811 117461 276814
rect 115716 276749 115750 276783
rect 115716 276681 115750 276715
rect 115716 276613 115750 276647
rect 114455 276545 114489 276579
rect 111520 276420 111547 276454
rect 111587 276420 111615 276454
rect 111659 276420 111683 276454
rect 111731 276420 111751 276454
rect 111803 276420 111819 276454
rect 111875 276420 111887 276454
rect 111947 276420 111955 276454
rect 112019 276420 112023 276454
rect 112125 276420 112129 276454
rect 112193 276420 112201 276454
rect 112261 276420 112273 276454
rect 112329 276420 112345 276454
rect 112397 276420 112417 276454
rect 112465 276420 112489 276454
rect 112533 276420 112561 276454
rect 112601 276420 112628 276454
rect 112832 276418 113216 276454
rect 112832 276414 113023 276418
rect 111452 276381 111486 276408
rect 111452 276311 111486 276345
rect 111452 276248 111486 276275
rect 112662 276381 112696 276408
rect 112832 276386 112872 276414
rect 112996 276384 113023 276414
rect 113063 276384 113091 276418
rect 113135 276384 113159 276418
rect 113207 276384 113227 276418
rect 113279 276384 113295 276418
rect 113351 276384 113363 276418
rect 113423 276384 113431 276418
rect 113495 276384 113499 276418
rect 113601 276384 113605 276418
rect 113669 276384 113677 276418
rect 113737 276384 113749 276418
rect 113805 276384 113821 276418
rect 113873 276384 113893 276418
rect 113941 276384 113965 276418
rect 114009 276384 114037 276418
rect 114077 276384 114104 276418
rect 112662 276311 112696 276345
rect 112928 276349 112962 276372
rect 112928 276292 112962 276315
rect 114138 276349 114172 276372
rect 114138 276292 114172 276315
rect 112662 276248 112696 276275
rect 112996 276246 113023 276280
rect 113063 276246 113091 276280
rect 113135 276246 113159 276280
rect 113207 276246 113227 276280
rect 113279 276246 113295 276280
rect 113351 276246 113363 276280
rect 113423 276246 113431 276280
rect 113495 276246 113499 276280
rect 113601 276246 113605 276280
rect 113669 276246 113677 276280
rect 113737 276246 113749 276280
rect 113805 276246 113821 276280
rect 113873 276246 113893 276280
rect 113941 276246 113965 276280
rect 114009 276246 114037 276280
rect 114077 276246 114104 276280
rect 114234 276246 114274 276504
rect 114653 276579 114672 276613
rect 114738 276579 114740 276613
rect 114774 276579 114776 276613
rect 114842 276579 114861 276613
rect 114653 276542 114709 276579
rect 114805 276544 114861 276579
rect 115061 276579 115144 276613
rect 115027 276545 115178 276579
rect 114455 276477 114489 276511
rect 114455 276409 114489 276443
rect 114455 276341 114489 276375
rect 114455 276273 114489 276307
rect 112994 276239 114455 276246
rect 111520 276202 111547 276236
rect 111587 276202 111615 276236
rect 111659 276202 111683 276236
rect 111731 276202 111751 276236
rect 111803 276202 111819 276236
rect 111875 276202 111887 276236
rect 111947 276202 111955 276236
rect 112019 276202 112023 276236
rect 112125 276202 112129 276236
rect 112193 276202 112201 276236
rect 112261 276202 112273 276236
rect 112329 276202 112345 276236
rect 112397 276202 112417 276236
rect 112465 276202 112489 276236
rect 112533 276202 112561 276236
rect 112601 276202 112628 276236
rect 111334 276166 112628 276202
rect 112994 276205 114489 276239
rect 114538 276503 114709 276542
rect 114804 276522 114991 276544
rect 114538 276377 114576 276503
rect 114804 276488 114899 276522
rect 114933 276488 114991 276522
rect 114804 276459 114991 276488
rect 115061 276511 115144 276545
rect 115344 276579 115363 276613
rect 115429 276579 115431 276613
rect 115465 276579 115467 276613
rect 115533 276579 115552 276613
rect 115344 276544 115400 276579
rect 115027 276477 115178 276511
rect 114653 276389 114672 276423
rect 114738 276389 114740 276423
rect 114774 276389 114776 276423
rect 114842 276389 114861 276423
rect 114938 276377 114975 276459
rect 114538 276350 114610 276377
rect 114538 276314 114576 276350
rect 114538 276280 114610 276314
rect 114538 276244 114576 276280
rect 114538 276217 114610 276244
rect 114904 276350 114975 276377
rect 114938 276314 114975 276350
rect 114904 276280 114975 276314
rect 114938 276244 114975 276280
rect 114904 276217 114975 276244
rect 115061 276443 115144 276477
rect 115214 276522 115401 276544
rect 115214 276488 115271 276522
rect 115305 276488 115401 276522
rect 115496 276542 115552 276579
rect 115716 276545 115750 276579
rect 115496 276503 115667 276542
rect 115214 276459 115401 276488
rect 115027 276409 115178 276443
rect 115061 276375 115144 276409
rect 115027 276341 115178 276375
rect 115061 276307 115144 276341
rect 115027 276273 115178 276307
rect 115061 276239 115144 276273
rect 115027 276205 115178 276239
rect 115230 276377 115267 276459
rect 115344 276389 115363 276423
rect 115429 276389 115431 276423
rect 115465 276389 115467 276423
rect 115533 276389 115552 276423
rect 115629 276377 115667 276503
rect 115230 276350 115301 276377
rect 115230 276314 115267 276350
rect 115230 276280 115301 276314
rect 115230 276244 115267 276280
rect 115230 276217 115301 276244
rect 115595 276350 115667 276377
rect 115629 276314 115667 276350
rect 115595 276280 115667 276314
rect 115629 276244 115667 276280
rect 115595 276217 115667 276244
rect 115809 276794 117461 276811
rect 115809 276775 116313 276794
rect 115809 276619 115881 276775
rect 116941 276716 117373 276750
rect 116101 276682 116128 276716
rect 116168 276682 116196 276716
rect 116240 276682 116264 276716
rect 116312 276682 116332 276716
rect 116384 276682 116400 276716
rect 116456 276682 116468 276716
rect 116528 276682 116536 276716
rect 116600 276682 116604 276716
rect 116706 276682 116710 276716
rect 116774 276682 116782 276716
rect 116842 276682 116854 276716
rect 116910 276682 116926 276716
rect 116978 276682 116998 276716
rect 117046 276682 117070 276716
rect 117114 276682 117142 276716
rect 117182 276708 117373 276716
rect 117182 276682 117209 276708
rect 115809 276585 115828 276619
rect 115862 276585 115881 276619
rect 116033 276647 116067 276670
rect 116033 276590 116067 276613
rect 117243 276647 117277 276670
rect 117243 276590 117277 276613
rect 115809 276537 115881 276585
rect 116101 276550 116128 276578
rect 115931 276544 116128 276550
rect 116168 276544 116196 276578
rect 116240 276544 116264 276578
rect 116312 276544 116332 276578
rect 116384 276544 116400 276578
rect 116456 276544 116468 276578
rect 116528 276544 116536 276578
rect 116600 276544 116604 276578
rect 116706 276544 116710 276578
rect 116774 276544 116782 276578
rect 116842 276544 116854 276578
rect 116910 276544 116926 276578
rect 116978 276544 116998 276578
rect 117046 276544 117070 276578
rect 117114 276544 117142 276578
rect 117182 276550 117209 276578
rect 117182 276544 117211 276550
rect 115716 276477 115750 276511
rect 115716 276409 115750 276443
rect 115716 276341 115750 276375
rect 115716 276273 115750 276307
rect 115931 276504 117211 276544
rect 115931 276246 115971 276504
rect 117333 276454 117373 276708
rect 117425 276490 117461 276794
rect 117577 276780 117604 276814
rect 117644 276780 117672 276814
rect 117716 276780 117740 276814
rect 117788 276780 117808 276814
rect 117860 276780 117876 276814
rect 117932 276780 117944 276814
rect 118004 276780 118012 276814
rect 118076 276780 118080 276814
rect 118182 276780 118186 276814
rect 118250 276780 118258 276814
rect 118318 276780 118330 276814
rect 118386 276780 118402 276814
rect 118454 276780 118474 276814
rect 118522 276780 118546 276814
rect 118590 276780 118618 276814
rect 118658 276780 118685 276814
rect 117509 276741 117543 276768
rect 117509 276671 117543 276705
rect 117509 276608 117543 276635
rect 118719 276741 118753 276768
rect 118719 276671 118753 276705
rect 118719 276608 118753 276635
rect 117577 276562 117604 276596
rect 117644 276562 117672 276596
rect 117716 276562 117740 276596
rect 117788 276562 117808 276596
rect 117860 276562 117876 276596
rect 117932 276562 117944 276596
rect 118004 276562 118012 276596
rect 118076 276562 118080 276596
rect 118182 276562 118186 276596
rect 118250 276562 118258 276596
rect 118318 276562 118330 276596
rect 118386 276562 118402 276596
rect 118454 276562 118474 276596
rect 118522 276562 118546 276596
rect 118590 276562 118618 276596
rect 118658 276562 118685 276596
rect 118829 276562 118871 276886
rect 117577 276526 118871 276562
rect 117425 276454 118685 276490
rect 116989 276418 117373 276454
rect 117577 276420 117604 276454
rect 117644 276420 117672 276454
rect 117716 276420 117740 276454
rect 117788 276420 117808 276454
rect 117860 276420 117876 276454
rect 117932 276420 117944 276454
rect 118004 276420 118012 276454
rect 118076 276420 118080 276454
rect 118182 276420 118186 276454
rect 118250 276420 118258 276454
rect 118318 276420 118330 276454
rect 118386 276420 118402 276454
rect 118454 276420 118474 276454
rect 118522 276420 118546 276454
rect 118590 276420 118618 276454
rect 118658 276420 118685 276454
rect 116101 276384 116128 276418
rect 116168 276384 116196 276418
rect 116240 276384 116264 276418
rect 116312 276384 116332 276418
rect 116384 276384 116400 276418
rect 116456 276384 116468 276418
rect 116528 276384 116536 276418
rect 116600 276384 116604 276418
rect 116706 276384 116710 276418
rect 116774 276384 116782 276418
rect 116842 276384 116854 276418
rect 116910 276384 116926 276418
rect 116978 276384 116998 276418
rect 117046 276384 117070 276418
rect 117114 276384 117142 276418
rect 117182 276414 117373 276418
rect 117182 276384 117209 276414
rect 117333 276386 117373 276414
rect 117509 276381 117543 276408
rect 116033 276349 116067 276372
rect 116033 276292 116067 276315
rect 117243 276349 117277 276372
rect 117243 276292 117277 276315
rect 117509 276311 117543 276345
rect 116101 276246 116128 276280
rect 116168 276246 116196 276280
rect 116240 276246 116264 276280
rect 116312 276246 116332 276280
rect 116384 276246 116400 276280
rect 116456 276246 116468 276280
rect 116528 276246 116536 276280
rect 116600 276246 116604 276280
rect 116706 276246 116710 276280
rect 116774 276246 116782 276280
rect 116842 276246 116854 276280
rect 116910 276246 116926 276280
rect 116978 276246 116998 276280
rect 117046 276246 117070 276280
rect 117114 276246 117142 276280
rect 117182 276246 117209 276280
rect 117509 276248 117543 276275
rect 118719 276381 118753 276408
rect 118719 276311 118753 276345
rect 118719 276248 118753 276275
rect 115750 276239 117211 276246
rect 115716 276205 117211 276239
rect 112994 276200 114455 276205
rect 114653 276171 114672 276205
rect 114738 276171 114740 276205
rect 114774 276171 114776 276205
rect 114842 276171 114861 276205
rect 115061 276171 115144 276205
rect 115344 276171 115363 276205
rect 115429 276171 115431 276205
rect 115465 276171 115467 276205
rect 115533 276171 115552 276205
rect 115750 276200 117211 276205
rect 117577 276202 117604 276236
rect 117644 276202 117672 276236
rect 117716 276202 117740 276236
rect 117788 276202 117808 276236
rect 117860 276202 117876 276236
rect 117932 276202 117944 276236
rect 118004 276202 118012 276236
rect 118076 276202 118080 276236
rect 118182 276202 118186 276236
rect 118250 276202 118258 276236
rect 118318 276202 118330 276236
rect 118386 276202 118402 276236
rect 118454 276202 118474 276236
rect 118522 276202 118546 276236
rect 118590 276202 118618 276236
rect 118658 276202 118685 276236
rect 118829 276202 118871 276526
rect 114455 276137 114489 276171
rect 115027 276155 115178 276171
rect 113982 276093 114266 276098
rect 111312 276067 114266 276093
rect 111312 276065 114034 276067
rect 114068 276065 114106 276067
rect 114140 276065 114178 276067
rect 114212 276065 114266 276067
rect 111312 276031 111340 276065
rect 111374 276031 111408 276065
rect 111442 276031 111476 276065
rect 111510 276031 111544 276065
rect 111578 276031 111612 276065
rect 111646 276031 111680 276065
rect 111714 276031 111748 276065
rect 111782 276031 111816 276065
rect 111850 276031 111884 276065
rect 111918 276031 111952 276065
rect 111986 276031 112020 276065
rect 112054 276031 112088 276065
rect 112122 276031 112156 276065
rect 112190 276031 112224 276065
rect 112258 276031 112292 276065
rect 112326 276031 112360 276065
rect 112394 276031 112428 276065
rect 112462 276031 112496 276065
rect 112530 276031 112564 276065
rect 112598 276031 112632 276065
rect 112666 276031 112700 276065
rect 112734 276031 112768 276065
rect 112802 276031 112836 276065
rect 112870 276031 112904 276065
rect 112938 276031 112972 276065
rect 113006 276031 113040 276065
rect 113074 276031 113108 276065
rect 113142 276031 113176 276065
rect 113210 276031 113244 276065
rect 113278 276031 113312 276065
rect 113346 276031 113380 276065
rect 113414 276031 113448 276065
rect 113482 276031 113516 276065
rect 113550 276031 113584 276065
rect 113618 276031 113652 276065
rect 113686 276031 113720 276065
rect 113754 276031 113788 276065
rect 113822 276031 113856 276065
rect 113890 276031 113924 276065
rect 113958 276031 113992 276065
rect 114026 276033 114034 276065
rect 114094 276033 114106 276065
rect 114162 276033 114178 276065
rect 114026 276031 114060 276033
rect 114094 276031 114128 276033
rect 114162 276031 114196 276033
rect 114230 276031 114266 276065
rect 114455 276071 114489 276103
rect 114930 276137 115275 276155
rect 114930 276103 115027 276137
rect 115061 276103 115144 276137
rect 115178 276103 115275 276137
rect 114930 276071 115275 276103
rect 115716 276137 115750 276171
rect 117577 276166 118871 276202
rect 115716 276071 115750 276103
rect 114455 276037 114537 276071
rect 114571 276037 114605 276071
rect 114639 276037 114673 276071
rect 114707 276037 114741 276071
rect 114775 276037 114809 276071
rect 114843 276037 114877 276071
rect 114911 276037 114945 276071
rect 114979 276037 115226 276071
rect 115260 276037 115294 276071
rect 115328 276037 115362 276071
rect 115396 276037 115430 276071
rect 115464 276037 115498 276071
rect 115532 276037 115566 276071
rect 115600 276037 115634 276071
rect 115668 276037 115750 276071
rect 115939 276093 116223 276098
rect 115939 276067 118893 276093
rect 115939 276065 115992 276067
rect 116026 276065 116064 276067
rect 116098 276065 116136 276067
rect 116170 276065 118893 276067
rect 111312 276003 114266 276031
rect 113036 275998 114266 276003
rect 113036 275906 114022 275998
rect 115061 275965 115144 276037
rect 115939 276031 115975 276065
rect 116026 276033 116043 276065
rect 116098 276033 116111 276065
rect 116170 276033 116179 276065
rect 116009 276031 116043 276033
rect 116077 276031 116111 276033
rect 116145 276031 116179 276033
rect 116213 276031 116247 276065
rect 116281 276031 116315 276065
rect 116349 276031 116383 276065
rect 116417 276031 116451 276065
rect 116485 276031 116519 276065
rect 116553 276031 116587 276065
rect 116621 276031 116655 276065
rect 116689 276031 116723 276065
rect 116757 276031 116791 276065
rect 116825 276031 116859 276065
rect 116893 276031 116927 276065
rect 116961 276031 116995 276065
rect 117029 276031 117063 276065
rect 117097 276031 117131 276065
rect 117165 276031 117199 276065
rect 117233 276031 117267 276065
rect 117301 276031 117335 276065
rect 117369 276031 117403 276065
rect 117437 276031 117471 276065
rect 117505 276031 117539 276065
rect 117573 276031 117607 276065
rect 117641 276031 117675 276065
rect 117709 276031 117743 276065
rect 117777 276031 117811 276065
rect 117845 276031 117879 276065
rect 117913 276031 117947 276065
rect 117981 276031 118015 276065
rect 118049 276031 118083 276065
rect 118117 276031 118151 276065
rect 118185 276031 118219 276065
rect 118253 276031 118287 276065
rect 118321 276031 118355 276065
rect 118389 276031 118423 276065
rect 118457 276031 118491 276065
rect 118525 276031 118559 276065
rect 118593 276031 118627 276065
rect 118661 276031 118695 276065
rect 118729 276031 118763 276065
rect 118797 276031 118831 276065
rect 118865 276031 118893 276065
rect 115939 276003 118893 276031
rect 115939 275998 117169 276003
rect 114455 275931 114537 275965
rect 114571 275931 114605 275965
rect 114639 275931 114673 275965
rect 114707 275931 114741 275965
rect 114775 275931 114809 275965
rect 114843 275931 114877 275965
rect 114911 275931 114945 275965
rect 114979 275931 115226 275965
rect 115260 275931 115294 275965
rect 115328 275931 115362 275965
rect 115396 275931 115430 275965
rect 115464 275931 115498 275965
rect 115532 275931 115566 275965
rect 115600 275931 115634 275965
rect 115668 275931 115750 275965
rect 111520 275868 112814 275904
rect 113036 275902 114246 275906
rect 113036 275901 114353 275902
rect 111520 275834 111547 275868
rect 111587 275834 111615 275868
rect 111659 275834 111683 275868
rect 111731 275834 111751 275868
rect 111803 275834 111819 275868
rect 111875 275834 111887 275868
rect 111947 275834 111955 275868
rect 112019 275834 112023 275868
rect 112125 275834 112129 275868
rect 112193 275834 112201 275868
rect 112261 275834 112273 275868
rect 112329 275834 112345 275868
rect 112397 275834 112417 275868
rect 112465 275834 112489 275868
rect 112533 275834 112561 275868
rect 112601 275834 112628 275868
rect 111452 275795 111486 275822
rect 111452 275725 111486 275759
rect 111452 275662 111486 275689
rect 112662 275795 112696 275822
rect 112662 275725 112696 275759
rect 112662 275662 112696 275689
rect 111520 275616 111547 275650
rect 111587 275616 111615 275650
rect 111659 275616 111683 275650
rect 111731 275616 111751 275650
rect 111803 275616 111819 275650
rect 111875 275616 111887 275650
rect 111947 275616 111955 275650
rect 112019 275616 112023 275650
rect 112125 275616 112129 275650
rect 112193 275616 112201 275650
rect 112261 275616 112273 275650
rect 112329 275616 112345 275650
rect 112397 275616 112417 275650
rect 112465 275616 112489 275650
rect 112533 275616 112561 275650
rect 112601 275616 112628 275650
rect 111334 275580 112628 275616
rect 112772 275584 112814 275868
rect 112966 275878 114353 275901
rect 112966 275876 114243 275878
rect 112966 275842 112993 275876
rect 113033 275842 113061 275876
rect 113105 275842 113129 275876
rect 113177 275842 113197 275876
rect 113249 275842 113265 275876
rect 113321 275842 113333 275876
rect 113393 275842 113401 275876
rect 113465 275842 113469 275876
rect 113571 275842 113575 275876
rect 113639 275842 113647 275876
rect 113707 275842 113719 275876
rect 113775 275842 113791 275876
rect 113843 275842 113863 275876
rect 113911 275842 113935 275876
rect 113979 275842 114007 275876
rect 114047 275872 114243 275876
rect 114047 275842 114074 275872
rect 112898 275783 112932 275830
rect 112898 275713 112932 275747
rect 112898 275630 112932 275677
rect 114108 275783 114142 275830
rect 114108 275713 114142 275747
rect 114108 275630 114142 275677
rect 114210 275776 114243 275872
rect 114345 275776 114353 275878
rect 114210 275752 114353 275776
rect 114455 275899 114489 275931
rect 114455 275831 114489 275865
rect 114652 275851 114862 275931
rect 114652 275817 114672 275851
rect 114738 275817 114740 275851
rect 114774 275817 114776 275851
rect 114842 275817 114862 275851
rect 114652 275816 114862 275817
rect 115027 275899 115178 275931
rect 115061 275865 115144 275899
rect 115027 275831 115178 275865
rect 114455 275763 114489 275797
rect 112966 275584 112993 275618
rect 113033 275584 113061 275618
rect 113105 275584 113129 275618
rect 113177 275584 113197 275618
rect 113249 275584 113265 275618
rect 113321 275584 113333 275618
rect 113393 275584 113401 275618
rect 113465 275584 113469 275618
rect 113571 275584 113575 275618
rect 113639 275584 113647 275618
rect 113707 275584 113719 275618
rect 113775 275584 113791 275618
rect 113843 275584 113863 275618
rect 113911 275584 113935 275618
rect 113979 275584 114007 275618
rect 114047 275584 114074 275618
rect 111334 275256 111376 275580
rect 112772 275550 114074 275584
rect 112772 275544 112832 275550
rect 111520 275508 112832 275544
rect 111520 275474 111547 275508
rect 111587 275474 111615 275508
rect 111659 275474 111683 275508
rect 111731 275474 111751 275508
rect 111803 275474 111819 275508
rect 111875 275474 111887 275508
rect 111947 275474 111955 275508
rect 112019 275474 112023 275508
rect 112125 275474 112129 275508
rect 112193 275474 112201 275508
rect 112261 275474 112273 275508
rect 112329 275474 112345 275508
rect 112397 275474 112417 275508
rect 112465 275474 112489 275508
rect 112533 275474 112561 275508
rect 112601 275474 112628 275508
rect 111452 275435 111486 275462
rect 111452 275365 111486 275399
rect 111452 275302 111486 275329
rect 112662 275435 112696 275462
rect 112662 275365 112696 275399
rect 112662 275302 112696 275329
rect 111520 275256 111547 275290
rect 111587 275256 111615 275290
rect 111659 275256 111683 275290
rect 111731 275256 111751 275290
rect 111803 275256 111819 275290
rect 111875 275256 111887 275290
rect 111947 275256 111955 275290
rect 112019 275256 112023 275290
rect 112125 275256 112129 275290
rect 112193 275256 112201 275290
rect 112261 275256 112273 275290
rect 112329 275256 112345 275290
rect 112397 275256 112417 275290
rect 112465 275256 112489 275290
rect 112533 275256 112561 275290
rect 112601 275256 112628 275290
rect 111334 275220 112628 275256
rect 111334 274896 111376 275220
rect 112772 275184 112832 275508
rect 114210 275486 114246 275752
rect 112966 275452 114246 275486
rect 114455 275695 114489 275729
rect 114455 275627 114489 275661
rect 114455 275559 114489 275593
rect 114455 275491 114489 275525
rect 112966 275418 112993 275452
rect 113033 275418 113061 275452
rect 113105 275418 113129 275452
rect 113177 275418 113197 275452
rect 113249 275418 113265 275452
rect 113321 275418 113333 275452
rect 113393 275418 113401 275452
rect 113465 275418 113469 275452
rect 113571 275418 113575 275452
rect 113639 275418 113647 275452
rect 113707 275418 113719 275452
rect 113775 275418 113791 275452
rect 113843 275418 113863 275452
rect 113911 275418 113935 275452
rect 113979 275418 114007 275452
rect 114047 275418 114074 275452
rect 114455 275423 114489 275457
rect 112898 275359 112932 275406
rect 112898 275289 112932 275323
rect 112898 275206 112932 275253
rect 114108 275359 114142 275406
rect 114108 275289 114142 275323
rect 114108 275206 114142 275253
rect 114455 275355 114489 275389
rect 114455 275287 114489 275321
rect 114455 275219 114489 275253
rect 111520 275162 112832 275184
rect 112966 275162 112993 275194
rect 111520 275160 112993 275162
rect 113033 275160 113061 275194
rect 113105 275160 113129 275194
rect 113177 275160 113197 275194
rect 113249 275160 113265 275194
rect 113321 275160 113333 275194
rect 113393 275160 113401 275194
rect 113465 275160 113469 275194
rect 113571 275160 113575 275194
rect 113639 275160 113647 275194
rect 113707 275160 113719 275194
rect 113775 275160 113791 275194
rect 113843 275160 113863 275194
rect 113911 275160 113935 275194
rect 113979 275160 114007 275194
rect 114047 275160 114074 275194
rect 111520 275148 114074 275160
rect 111520 275114 111547 275148
rect 111587 275114 111615 275148
rect 111659 275114 111683 275148
rect 111731 275114 111751 275148
rect 111803 275114 111819 275148
rect 111875 275114 111887 275148
rect 111947 275114 111955 275148
rect 112019 275114 112023 275148
rect 112125 275114 112129 275148
rect 112193 275114 112201 275148
rect 112261 275114 112273 275148
rect 112329 275114 112345 275148
rect 112397 275114 112417 275148
rect 112465 275114 112489 275148
rect 112533 275114 112561 275148
rect 112601 275114 112628 275148
rect 112744 275145 114074 275148
rect 114455 275151 114489 275185
rect 112744 275128 114396 275145
rect 111452 275075 111486 275102
rect 111452 275005 111486 275039
rect 111452 274942 111486 274969
rect 112662 275075 112696 275102
rect 112662 275005 112696 275039
rect 112662 274942 112696 274969
rect 111520 274896 111547 274930
rect 111587 274896 111615 274930
rect 111659 274896 111683 274930
rect 111731 274896 111751 274930
rect 111803 274896 111819 274930
rect 111875 274896 111887 274930
rect 111947 274896 111955 274930
rect 112019 274896 112023 274930
rect 112125 274896 112129 274930
rect 112193 274896 112201 274930
rect 112261 274896 112273 274930
rect 112329 274896 112345 274930
rect 112397 274896 112417 274930
rect 112465 274896 112489 274930
rect 112533 274896 112561 274930
rect 112601 274896 112628 274930
rect 111334 274860 112628 274896
rect 111334 274536 111376 274860
rect 112744 274824 112780 275128
rect 113892 275109 114396 275128
rect 111520 274788 112780 274824
rect 112832 275050 113264 275084
rect 112832 275042 113023 275050
rect 112832 274788 112872 275042
rect 112996 275016 113023 275042
rect 113063 275016 113091 275050
rect 113135 275016 113159 275050
rect 113207 275016 113227 275050
rect 113279 275016 113295 275050
rect 113351 275016 113363 275050
rect 113423 275016 113431 275050
rect 113495 275016 113499 275050
rect 113601 275016 113605 275050
rect 113669 275016 113677 275050
rect 113737 275016 113749 275050
rect 113805 275016 113821 275050
rect 113873 275016 113893 275050
rect 113941 275016 113965 275050
rect 114009 275016 114037 275050
rect 114077 275016 114104 275050
rect 112928 274981 112962 275004
rect 112928 274924 112962 274947
rect 114138 274981 114172 275004
rect 114138 274924 114172 274947
rect 114324 274953 114396 275109
rect 114324 274919 114342 274953
rect 114376 274919 114396 274953
rect 112996 274884 113023 274912
rect 112994 274878 113023 274884
rect 113063 274878 113091 274912
rect 113135 274878 113159 274912
rect 113207 274878 113227 274912
rect 113279 274878 113295 274912
rect 113351 274878 113363 274912
rect 113423 274878 113431 274912
rect 113495 274878 113499 274912
rect 113601 274878 113605 274912
rect 113669 274878 113677 274912
rect 113737 274878 113749 274912
rect 113805 274878 113821 274912
rect 113873 274878 113893 274912
rect 113941 274878 113965 274912
rect 114009 274878 114037 274912
rect 114077 274884 114104 274912
rect 114077 274878 114274 274884
rect 112994 274838 114274 274878
rect 114324 274871 114396 274919
rect 114455 275083 114489 275117
rect 114455 275015 114489 275049
rect 114455 274947 114489 274981
rect 114576 275766 114610 275805
rect 114576 275694 114610 275724
rect 114576 275622 114610 275656
rect 114576 275554 114610 275588
rect 114576 275486 114610 275516
rect 114576 275277 114610 275444
rect 114904 275766 114938 275805
rect 114904 275694 114938 275724
rect 114904 275622 114938 275656
rect 114904 275554 114938 275588
rect 114904 275486 114938 275516
rect 114653 275359 114672 275393
rect 114738 275359 114740 275393
rect 114774 275359 114776 275393
rect 114842 275359 114861 275393
rect 114904 275313 114938 275444
rect 115061 275797 115144 275831
rect 115343 275851 115553 275931
rect 115343 275817 115363 275851
rect 115429 275817 115431 275851
rect 115465 275817 115467 275851
rect 115533 275817 115553 275851
rect 115343 275816 115553 275817
rect 115716 275899 115750 275931
rect 116183 275906 117169 275998
rect 115959 275902 117169 275906
rect 115716 275831 115750 275865
rect 115027 275763 115178 275797
rect 115061 275729 115144 275763
rect 115027 275695 115178 275729
rect 115061 275661 115144 275695
rect 115027 275627 115178 275661
rect 115061 275593 115144 275627
rect 115027 275559 115178 275593
rect 115061 275525 115144 275559
rect 115027 275491 115178 275525
rect 115061 275457 115144 275491
rect 115027 275423 115178 275457
rect 115061 275389 115144 275423
rect 115027 275355 115178 275389
rect 115061 275321 115144 275355
rect 114865 275279 114970 275313
rect 114865 275277 114899 275279
rect 114576 275245 114899 275277
rect 114933 275245 114970 275279
rect 114576 275229 114970 275245
rect 114576 275092 114610 275229
rect 114865 275206 114970 275229
rect 115027 275287 115178 275321
rect 115267 275766 115301 275805
rect 115267 275694 115301 275724
rect 115267 275622 115301 275656
rect 115267 275554 115301 275588
rect 115267 275486 115301 275516
rect 115267 275313 115301 275444
rect 115595 275766 115629 275805
rect 115595 275694 115629 275724
rect 115595 275622 115629 275656
rect 115595 275554 115629 275588
rect 115595 275486 115629 275516
rect 115344 275359 115363 275393
rect 115429 275359 115431 275393
rect 115465 275359 115467 275393
rect 115533 275359 115552 275393
rect 115061 275253 115144 275287
rect 115027 275219 115178 275253
rect 114653 275131 114672 275165
rect 114738 275131 114740 275165
rect 114774 275131 114776 275165
rect 114842 275131 114861 275165
rect 114576 275022 114610 275056
rect 114576 274959 114610 274986
rect 114904 275092 114938 275206
rect 114904 275022 114938 275056
rect 114904 274959 114938 274986
rect 115061 275185 115144 275219
rect 115235 275279 115340 275313
rect 115235 275245 115271 275279
rect 115305 275277 115340 275279
rect 115595 275277 115629 275444
rect 115305 275245 115629 275277
rect 115235 275229 115629 275245
rect 115235 275206 115340 275229
rect 115027 275151 115178 275185
rect 115061 275117 115144 275151
rect 115027 275083 115178 275117
rect 115061 275049 115144 275083
rect 115027 275015 115178 275049
rect 115061 274981 115144 275015
rect 115027 274947 115178 274981
rect 115267 275092 115301 275206
rect 115344 275131 115363 275165
rect 115429 275131 115431 275165
rect 115465 275131 115467 275165
rect 115533 275131 115552 275165
rect 115267 275022 115301 275056
rect 115267 274959 115301 274986
rect 115595 275092 115629 275229
rect 115595 275022 115629 275056
rect 115595 274959 115629 274986
rect 115716 275763 115750 275797
rect 115852 275901 117169 275902
rect 115852 275878 117239 275901
rect 115852 275776 115860 275878
rect 115962 275876 117239 275878
rect 115962 275872 116158 275876
rect 115962 275776 115995 275872
rect 116131 275842 116158 275872
rect 116198 275842 116226 275876
rect 116270 275842 116294 275876
rect 116342 275842 116362 275876
rect 116414 275842 116430 275876
rect 116486 275842 116498 275876
rect 116558 275842 116566 275876
rect 116630 275842 116634 275876
rect 116736 275842 116740 275876
rect 116804 275842 116812 275876
rect 116872 275842 116884 275876
rect 116940 275842 116956 275876
rect 117008 275842 117028 275876
rect 117076 275842 117100 275876
rect 117144 275842 117172 275876
rect 117212 275842 117239 275876
rect 117391 275868 118685 275904
rect 115852 275752 115995 275776
rect 115716 275695 115750 275729
rect 115716 275627 115750 275661
rect 115716 275559 115750 275593
rect 115716 275491 115750 275525
rect 115716 275423 115750 275457
rect 115959 275486 115995 275752
rect 116063 275783 116097 275830
rect 116063 275713 116097 275747
rect 116063 275630 116097 275677
rect 117273 275783 117307 275830
rect 117273 275713 117307 275747
rect 117273 275630 117307 275677
rect 116131 275584 116158 275618
rect 116198 275584 116226 275618
rect 116270 275584 116294 275618
rect 116342 275584 116362 275618
rect 116414 275584 116430 275618
rect 116486 275584 116498 275618
rect 116558 275584 116566 275618
rect 116630 275584 116634 275618
rect 116736 275584 116740 275618
rect 116804 275584 116812 275618
rect 116872 275584 116884 275618
rect 116940 275584 116956 275618
rect 117008 275584 117028 275618
rect 117076 275584 117100 275618
rect 117144 275584 117172 275618
rect 117212 275584 117239 275618
rect 117391 275584 117433 275868
rect 117577 275834 117604 275868
rect 117644 275834 117672 275868
rect 117716 275834 117740 275868
rect 117788 275834 117808 275868
rect 117860 275834 117876 275868
rect 117932 275834 117944 275868
rect 118004 275834 118012 275868
rect 118076 275834 118080 275868
rect 118182 275834 118186 275868
rect 118250 275834 118258 275868
rect 118318 275834 118330 275868
rect 118386 275834 118402 275868
rect 118454 275834 118474 275868
rect 118522 275834 118546 275868
rect 118590 275834 118618 275868
rect 118658 275834 118685 275868
rect 117509 275795 117543 275822
rect 117509 275725 117543 275759
rect 117509 275662 117543 275689
rect 118719 275795 118753 275822
rect 118719 275725 118753 275759
rect 118719 275662 118753 275689
rect 116131 275550 117433 275584
rect 117577 275616 117604 275650
rect 117644 275616 117672 275650
rect 117716 275616 117740 275650
rect 117788 275616 117808 275650
rect 117860 275616 117876 275650
rect 117932 275616 117944 275650
rect 118004 275616 118012 275650
rect 118076 275616 118080 275650
rect 118182 275616 118186 275650
rect 118250 275616 118258 275650
rect 118318 275616 118330 275650
rect 118386 275616 118402 275650
rect 118454 275616 118474 275650
rect 118522 275616 118546 275650
rect 118590 275616 118618 275650
rect 118658 275616 118685 275650
rect 117577 275580 118871 275616
rect 117373 275544 117433 275550
rect 117373 275508 118685 275544
rect 115959 275452 117239 275486
rect 116131 275418 116158 275452
rect 116198 275418 116226 275452
rect 116270 275418 116294 275452
rect 116342 275418 116362 275452
rect 116414 275418 116430 275452
rect 116486 275418 116498 275452
rect 116558 275418 116566 275452
rect 116630 275418 116634 275452
rect 116736 275418 116740 275452
rect 116804 275418 116812 275452
rect 116872 275418 116884 275452
rect 116940 275418 116956 275452
rect 117008 275418 117028 275452
rect 117076 275418 117100 275452
rect 117144 275418 117172 275452
rect 117212 275418 117239 275452
rect 115716 275355 115750 275389
rect 115716 275287 115750 275321
rect 115716 275219 115750 275253
rect 116063 275359 116097 275406
rect 116063 275289 116097 275323
rect 116063 275206 116097 275253
rect 117273 275359 117307 275406
rect 117273 275289 117307 275323
rect 117273 275206 117307 275253
rect 115716 275151 115750 275185
rect 116131 275160 116158 275194
rect 116198 275160 116226 275194
rect 116270 275160 116294 275194
rect 116342 275160 116362 275194
rect 116414 275160 116430 275194
rect 116486 275160 116498 275194
rect 116558 275160 116566 275194
rect 116630 275160 116634 275194
rect 116736 275160 116740 275194
rect 116804 275160 116812 275194
rect 116872 275160 116884 275194
rect 116940 275160 116956 275194
rect 117008 275160 117028 275194
rect 117076 275160 117100 275194
rect 117144 275160 117172 275194
rect 117212 275162 117239 275194
rect 117373 275184 117433 275508
rect 117577 275474 117604 275508
rect 117644 275474 117672 275508
rect 117716 275474 117740 275508
rect 117788 275474 117808 275508
rect 117860 275474 117876 275508
rect 117932 275474 117944 275508
rect 118004 275474 118012 275508
rect 118076 275474 118080 275508
rect 118182 275474 118186 275508
rect 118250 275474 118258 275508
rect 118318 275474 118330 275508
rect 118386 275474 118402 275508
rect 118454 275474 118474 275508
rect 118522 275474 118546 275508
rect 118590 275474 118618 275508
rect 118658 275474 118685 275508
rect 117509 275435 117543 275462
rect 117509 275365 117543 275399
rect 117509 275302 117543 275329
rect 118719 275435 118753 275462
rect 118719 275365 118753 275399
rect 118719 275302 118753 275329
rect 117577 275256 117604 275290
rect 117644 275256 117672 275290
rect 117716 275256 117740 275290
rect 117788 275256 117808 275290
rect 117860 275256 117876 275290
rect 117932 275256 117944 275290
rect 118004 275256 118012 275290
rect 118076 275256 118080 275290
rect 118182 275256 118186 275290
rect 118250 275256 118258 275290
rect 118318 275256 118330 275290
rect 118386 275256 118402 275290
rect 118454 275256 118474 275290
rect 118522 275256 118546 275290
rect 118590 275256 118618 275290
rect 118658 275256 118685 275290
rect 118829 275256 118871 275580
rect 117577 275220 118871 275256
rect 117373 275162 118685 275184
rect 117212 275160 118685 275162
rect 116131 275148 118685 275160
rect 116131 275145 117461 275148
rect 115716 275083 115750 275117
rect 115716 275015 115750 275049
rect 115716 274947 115750 274981
rect 114455 274879 114489 274913
rect 111520 274754 111547 274788
rect 111587 274754 111615 274788
rect 111659 274754 111683 274788
rect 111731 274754 111751 274788
rect 111803 274754 111819 274788
rect 111875 274754 111887 274788
rect 111947 274754 111955 274788
rect 112019 274754 112023 274788
rect 112125 274754 112129 274788
rect 112193 274754 112201 274788
rect 112261 274754 112273 274788
rect 112329 274754 112345 274788
rect 112397 274754 112417 274788
rect 112465 274754 112489 274788
rect 112533 274754 112561 274788
rect 112601 274754 112628 274788
rect 112832 274752 113216 274788
rect 112832 274748 113023 274752
rect 111452 274715 111486 274742
rect 111452 274645 111486 274679
rect 111452 274582 111486 274609
rect 112662 274715 112696 274742
rect 112832 274720 112872 274748
rect 112996 274718 113023 274748
rect 113063 274718 113091 274752
rect 113135 274718 113159 274752
rect 113207 274718 113227 274752
rect 113279 274718 113295 274752
rect 113351 274718 113363 274752
rect 113423 274718 113431 274752
rect 113495 274718 113499 274752
rect 113601 274718 113605 274752
rect 113669 274718 113677 274752
rect 113737 274718 113749 274752
rect 113805 274718 113821 274752
rect 113873 274718 113893 274752
rect 113941 274718 113965 274752
rect 114009 274718 114037 274752
rect 114077 274718 114104 274752
rect 112662 274645 112696 274679
rect 112928 274683 112962 274706
rect 112928 274626 112962 274649
rect 114138 274683 114172 274706
rect 114138 274626 114172 274649
rect 112662 274582 112696 274609
rect 112996 274580 113023 274614
rect 113063 274580 113091 274614
rect 113135 274580 113159 274614
rect 113207 274580 113227 274614
rect 113279 274580 113295 274614
rect 113351 274580 113363 274614
rect 113423 274580 113431 274614
rect 113495 274580 113499 274614
rect 113601 274580 113605 274614
rect 113669 274580 113677 274614
rect 113737 274580 113749 274614
rect 113805 274580 113821 274614
rect 113873 274580 113893 274614
rect 113941 274580 113965 274614
rect 114009 274580 114037 274614
rect 114077 274580 114104 274614
rect 114234 274580 114274 274838
rect 114653 274913 114672 274947
rect 114738 274913 114740 274947
rect 114774 274913 114776 274947
rect 114842 274913 114861 274947
rect 114653 274876 114709 274913
rect 114805 274878 114861 274913
rect 115061 274913 115144 274947
rect 115027 274879 115178 274913
rect 114455 274811 114489 274845
rect 114455 274743 114489 274777
rect 114455 274675 114489 274709
rect 114455 274607 114489 274641
rect 112994 274573 114455 274580
rect 111520 274536 111547 274570
rect 111587 274536 111615 274570
rect 111659 274536 111683 274570
rect 111731 274536 111751 274570
rect 111803 274536 111819 274570
rect 111875 274536 111887 274570
rect 111947 274536 111955 274570
rect 112019 274536 112023 274570
rect 112125 274536 112129 274570
rect 112193 274536 112201 274570
rect 112261 274536 112273 274570
rect 112329 274536 112345 274570
rect 112397 274536 112417 274570
rect 112465 274536 112489 274570
rect 112533 274536 112561 274570
rect 112601 274536 112628 274570
rect 111334 274500 112628 274536
rect 112994 274539 114489 274573
rect 114538 274837 114709 274876
rect 114804 274856 114991 274878
rect 114538 274711 114576 274837
rect 114804 274822 114899 274856
rect 114933 274822 114991 274856
rect 114804 274793 114991 274822
rect 115061 274845 115144 274879
rect 115344 274913 115363 274947
rect 115429 274913 115431 274947
rect 115465 274913 115467 274947
rect 115533 274913 115552 274947
rect 115344 274878 115400 274913
rect 115027 274811 115178 274845
rect 114653 274723 114672 274757
rect 114738 274723 114740 274757
rect 114774 274723 114776 274757
rect 114842 274723 114861 274757
rect 114938 274711 114975 274793
rect 114538 274684 114610 274711
rect 114538 274648 114576 274684
rect 114538 274614 114610 274648
rect 114538 274578 114576 274614
rect 114538 274551 114610 274578
rect 114904 274684 114975 274711
rect 114938 274648 114975 274684
rect 114904 274614 114975 274648
rect 114938 274578 114975 274614
rect 114904 274551 114975 274578
rect 115061 274777 115144 274811
rect 115214 274856 115401 274878
rect 115214 274822 115271 274856
rect 115305 274822 115401 274856
rect 115496 274876 115552 274913
rect 115716 274879 115750 274913
rect 115496 274837 115667 274876
rect 115214 274793 115401 274822
rect 115027 274743 115178 274777
rect 115061 274709 115144 274743
rect 115027 274675 115178 274709
rect 115061 274641 115144 274675
rect 115027 274607 115178 274641
rect 115061 274573 115144 274607
rect 115027 274539 115178 274573
rect 115230 274711 115267 274793
rect 115344 274723 115363 274757
rect 115429 274723 115431 274757
rect 115465 274723 115467 274757
rect 115533 274723 115552 274757
rect 115629 274711 115667 274837
rect 115230 274684 115301 274711
rect 115230 274648 115267 274684
rect 115230 274614 115301 274648
rect 115230 274578 115267 274614
rect 115230 274551 115301 274578
rect 115595 274684 115667 274711
rect 115629 274648 115667 274684
rect 115595 274614 115667 274648
rect 115629 274578 115667 274614
rect 115595 274551 115667 274578
rect 115809 275128 117461 275145
rect 115809 275109 116313 275128
rect 115809 274953 115881 275109
rect 116941 275050 117373 275084
rect 116101 275016 116128 275050
rect 116168 275016 116196 275050
rect 116240 275016 116264 275050
rect 116312 275016 116332 275050
rect 116384 275016 116400 275050
rect 116456 275016 116468 275050
rect 116528 275016 116536 275050
rect 116600 275016 116604 275050
rect 116706 275016 116710 275050
rect 116774 275016 116782 275050
rect 116842 275016 116854 275050
rect 116910 275016 116926 275050
rect 116978 275016 116998 275050
rect 117046 275016 117070 275050
rect 117114 275016 117142 275050
rect 117182 275042 117373 275050
rect 117182 275016 117209 275042
rect 115809 274919 115828 274953
rect 115862 274919 115881 274953
rect 116033 274981 116067 275004
rect 116033 274924 116067 274947
rect 117243 274981 117277 275004
rect 117243 274924 117277 274947
rect 115809 274871 115881 274919
rect 116101 274884 116128 274912
rect 115931 274878 116128 274884
rect 116168 274878 116196 274912
rect 116240 274878 116264 274912
rect 116312 274878 116332 274912
rect 116384 274878 116400 274912
rect 116456 274878 116468 274912
rect 116528 274878 116536 274912
rect 116600 274878 116604 274912
rect 116706 274878 116710 274912
rect 116774 274878 116782 274912
rect 116842 274878 116854 274912
rect 116910 274878 116926 274912
rect 116978 274878 116998 274912
rect 117046 274878 117070 274912
rect 117114 274878 117142 274912
rect 117182 274884 117209 274912
rect 117182 274878 117211 274884
rect 115716 274811 115750 274845
rect 115716 274743 115750 274777
rect 115716 274675 115750 274709
rect 115716 274607 115750 274641
rect 115931 274838 117211 274878
rect 115931 274580 115971 274838
rect 117333 274788 117373 275042
rect 117425 274824 117461 275128
rect 117577 275114 117604 275148
rect 117644 275114 117672 275148
rect 117716 275114 117740 275148
rect 117788 275114 117808 275148
rect 117860 275114 117876 275148
rect 117932 275114 117944 275148
rect 118004 275114 118012 275148
rect 118076 275114 118080 275148
rect 118182 275114 118186 275148
rect 118250 275114 118258 275148
rect 118318 275114 118330 275148
rect 118386 275114 118402 275148
rect 118454 275114 118474 275148
rect 118522 275114 118546 275148
rect 118590 275114 118618 275148
rect 118658 275114 118685 275148
rect 117509 275075 117543 275102
rect 117509 275005 117543 275039
rect 117509 274942 117543 274969
rect 118719 275075 118753 275102
rect 118719 275005 118753 275039
rect 118719 274942 118753 274969
rect 117577 274896 117604 274930
rect 117644 274896 117672 274930
rect 117716 274896 117740 274930
rect 117788 274896 117808 274930
rect 117860 274896 117876 274930
rect 117932 274896 117944 274930
rect 118004 274896 118012 274930
rect 118076 274896 118080 274930
rect 118182 274896 118186 274930
rect 118250 274896 118258 274930
rect 118318 274896 118330 274930
rect 118386 274896 118402 274930
rect 118454 274896 118474 274930
rect 118522 274896 118546 274930
rect 118590 274896 118618 274930
rect 118658 274896 118685 274930
rect 118829 274896 118871 275220
rect 117577 274860 118871 274896
rect 117425 274788 118685 274824
rect 116989 274752 117373 274788
rect 117577 274754 117604 274788
rect 117644 274754 117672 274788
rect 117716 274754 117740 274788
rect 117788 274754 117808 274788
rect 117860 274754 117876 274788
rect 117932 274754 117944 274788
rect 118004 274754 118012 274788
rect 118076 274754 118080 274788
rect 118182 274754 118186 274788
rect 118250 274754 118258 274788
rect 118318 274754 118330 274788
rect 118386 274754 118402 274788
rect 118454 274754 118474 274788
rect 118522 274754 118546 274788
rect 118590 274754 118618 274788
rect 118658 274754 118685 274788
rect 116101 274718 116128 274752
rect 116168 274718 116196 274752
rect 116240 274718 116264 274752
rect 116312 274718 116332 274752
rect 116384 274718 116400 274752
rect 116456 274718 116468 274752
rect 116528 274718 116536 274752
rect 116600 274718 116604 274752
rect 116706 274718 116710 274752
rect 116774 274718 116782 274752
rect 116842 274718 116854 274752
rect 116910 274718 116926 274752
rect 116978 274718 116998 274752
rect 117046 274718 117070 274752
rect 117114 274718 117142 274752
rect 117182 274748 117373 274752
rect 117182 274718 117209 274748
rect 117333 274720 117373 274748
rect 117509 274715 117543 274742
rect 116033 274683 116067 274706
rect 116033 274626 116067 274649
rect 117243 274683 117277 274706
rect 117243 274626 117277 274649
rect 117509 274645 117543 274679
rect 116101 274580 116128 274614
rect 116168 274580 116196 274614
rect 116240 274580 116264 274614
rect 116312 274580 116332 274614
rect 116384 274580 116400 274614
rect 116456 274580 116468 274614
rect 116528 274580 116536 274614
rect 116600 274580 116604 274614
rect 116706 274580 116710 274614
rect 116774 274580 116782 274614
rect 116842 274580 116854 274614
rect 116910 274580 116926 274614
rect 116978 274580 116998 274614
rect 117046 274580 117070 274614
rect 117114 274580 117142 274614
rect 117182 274580 117209 274614
rect 117509 274582 117543 274609
rect 118719 274715 118753 274742
rect 118719 274645 118753 274679
rect 118719 274582 118753 274609
rect 115750 274573 117211 274580
rect 115716 274539 117211 274573
rect 112994 274534 114455 274539
rect 114653 274505 114672 274539
rect 114738 274505 114740 274539
rect 114774 274505 114776 274539
rect 114842 274505 114861 274539
rect 115061 274505 115144 274539
rect 115344 274505 115363 274539
rect 115429 274505 115431 274539
rect 115465 274505 115467 274539
rect 115533 274505 115552 274539
rect 115750 274534 117211 274539
rect 117577 274536 117604 274570
rect 117644 274536 117672 274570
rect 117716 274536 117740 274570
rect 117788 274536 117808 274570
rect 117860 274536 117876 274570
rect 117932 274536 117944 274570
rect 118004 274536 118012 274570
rect 118076 274536 118080 274570
rect 118182 274536 118186 274570
rect 118250 274536 118258 274570
rect 118318 274536 118330 274570
rect 118386 274536 118402 274570
rect 118454 274536 118474 274570
rect 118522 274536 118546 274570
rect 118590 274536 118618 274570
rect 118658 274536 118685 274570
rect 118829 274536 118871 274860
rect 114455 274471 114489 274505
rect 115027 274489 115178 274505
rect 113982 274427 114266 274432
rect 111312 274401 114266 274427
rect 111312 274399 114034 274401
rect 114068 274399 114106 274401
rect 114140 274399 114178 274401
rect 114212 274399 114266 274401
rect 111312 274365 111340 274399
rect 111374 274365 111408 274399
rect 111442 274365 111476 274399
rect 111510 274365 111544 274399
rect 111578 274365 111612 274399
rect 111646 274365 111680 274399
rect 111714 274365 111748 274399
rect 111782 274365 111816 274399
rect 111850 274365 111884 274399
rect 111918 274365 111952 274399
rect 111986 274365 112020 274399
rect 112054 274365 112088 274399
rect 112122 274365 112156 274399
rect 112190 274365 112224 274399
rect 112258 274365 112292 274399
rect 112326 274365 112360 274399
rect 112394 274365 112428 274399
rect 112462 274365 112496 274399
rect 112530 274365 112564 274399
rect 112598 274365 112632 274399
rect 112666 274365 112700 274399
rect 112734 274365 112768 274399
rect 112802 274365 112836 274399
rect 112870 274365 112904 274399
rect 112938 274365 112972 274399
rect 113006 274365 113040 274399
rect 113074 274365 113108 274399
rect 113142 274365 113176 274399
rect 113210 274365 113244 274399
rect 113278 274365 113312 274399
rect 113346 274365 113380 274399
rect 113414 274365 113448 274399
rect 113482 274365 113516 274399
rect 113550 274365 113584 274399
rect 113618 274365 113652 274399
rect 113686 274365 113720 274399
rect 113754 274365 113788 274399
rect 113822 274365 113856 274399
rect 113890 274365 113924 274399
rect 113958 274365 113992 274399
rect 114026 274367 114034 274399
rect 114094 274367 114106 274399
rect 114162 274367 114178 274399
rect 114026 274365 114060 274367
rect 114094 274365 114128 274367
rect 114162 274365 114196 274367
rect 114230 274365 114266 274399
rect 114455 274405 114489 274437
rect 114930 274471 115275 274489
rect 114930 274437 115027 274471
rect 115061 274437 115144 274471
rect 115178 274437 115275 274471
rect 114930 274405 115275 274437
rect 115716 274471 115750 274505
rect 117577 274500 118871 274536
rect 115716 274405 115750 274437
rect 114455 274371 114537 274405
rect 114571 274371 114605 274405
rect 114639 274371 114673 274405
rect 114707 274371 114741 274405
rect 114775 274371 114809 274405
rect 114843 274371 114877 274405
rect 114911 274371 114945 274405
rect 114979 274371 115226 274405
rect 115260 274371 115294 274405
rect 115328 274371 115362 274405
rect 115396 274371 115430 274405
rect 115464 274371 115498 274405
rect 115532 274371 115566 274405
rect 115600 274371 115634 274405
rect 115668 274371 115750 274405
rect 115939 274427 116223 274432
rect 115939 274401 118893 274427
rect 115939 274399 115992 274401
rect 116026 274399 116064 274401
rect 116098 274399 116136 274401
rect 116170 274399 118893 274401
rect 111312 274337 114266 274365
rect 113036 274332 114266 274337
rect 113036 274240 114022 274332
rect 115061 274299 115144 274371
rect 115939 274365 115975 274399
rect 116026 274367 116043 274399
rect 116098 274367 116111 274399
rect 116170 274367 116179 274399
rect 116009 274365 116043 274367
rect 116077 274365 116111 274367
rect 116145 274365 116179 274367
rect 116213 274365 116247 274399
rect 116281 274365 116315 274399
rect 116349 274365 116383 274399
rect 116417 274365 116451 274399
rect 116485 274365 116519 274399
rect 116553 274365 116587 274399
rect 116621 274365 116655 274399
rect 116689 274365 116723 274399
rect 116757 274365 116791 274399
rect 116825 274365 116859 274399
rect 116893 274365 116927 274399
rect 116961 274365 116995 274399
rect 117029 274365 117063 274399
rect 117097 274365 117131 274399
rect 117165 274365 117199 274399
rect 117233 274365 117267 274399
rect 117301 274365 117335 274399
rect 117369 274365 117403 274399
rect 117437 274365 117471 274399
rect 117505 274365 117539 274399
rect 117573 274365 117607 274399
rect 117641 274365 117675 274399
rect 117709 274365 117743 274399
rect 117777 274365 117811 274399
rect 117845 274365 117879 274399
rect 117913 274365 117947 274399
rect 117981 274365 118015 274399
rect 118049 274365 118083 274399
rect 118117 274365 118151 274399
rect 118185 274365 118219 274399
rect 118253 274365 118287 274399
rect 118321 274365 118355 274399
rect 118389 274365 118423 274399
rect 118457 274365 118491 274399
rect 118525 274365 118559 274399
rect 118593 274365 118627 274399
rect 118661 274365 118695 274399
rect 118729 274365 118763 274399
rect 118797 274365 118831 274399
rect 118865 274365 118893 274399
rect 115939 274337 118893 274365
rect 115939 274332 117169 274337
rect 114455 274265 114537 274299
rect 114571 274265 114605 274299
rect 114639 274265 114673 274299
rect 114707 274265 114741 274299
rect 114775 274265 114809 274299
rect 114843 274265 114877 274299
rect 114911 274265 114945 274299
rect 114979 274265 115226 274299
rect 115260 274265 115294 274299
rect 115328 274265 115362 274299
rect 115396 274265 115430 274299
rect 115464 274265 115498 274299
rect 115532 274265 115566 274299
rect 115600 274265 115634 274299
rect 115668 274265 115750 274299
rect 111520 274202 112814 274238
rect 113036 274236 114246 274240
rect 113036 274235 114353 274236
rect 111520 274168 111547 274202
rect 111587 274168 111615 274202
rect 111659 274168 111683 274202
rect 111731 274168 111751 274202
rect 111803 274168 111819 274202
rect 111875 274168 111887 274202
rect 111947 274168 111955 274202
rect 112019 274168 112023 274202
rect 112125 274168 112129 274202
rect 112193 274168 112201 274202
rect 112261 274168 112273 274202
rect 112329 274168 112345 274202
rect 112397 274168 112417 274202
rect 112465 274168 112489 274202
rect 112533 274168 112561 274202
rect 112601 274168 112628 274202
rect 111452 274129 111486 274156
rect 111452 274059 111486 274093
rect 111452 273996 111486 274023
rect 112662 274129 112696 274156
rect 112662 274059 112696 274093
rect 112662 273996 112696 274023
rect 111520 273950 111547 273984
rect 111587 273950 111615 273984
rect 111659 273950 111683 273984
rect 111731 273950 111751 273984
rect 111803 273950 111819 273984
rect 111875 273950 111887 273984
rect 111947 273950 111955 273984
rect 112019 273950 112023 273984
rect 112125 273950 112129 273984
rect 112193 273950 112201 273984
rect 112261 273950 112273 273984
rect 112329 273950 112345 273984
rect 112397 273950 112417 273984
rect 112465 273950 112489 273984
rect 112533 273950 112561 273984
rect 112601 273950 112628 273984
rect 111334 273914 112628 273950
rect 112772 273918 112814 274202
rect 112966 274212 114353 274235
rect 112966 274210 114243 274212
rect 112966 274176 112993 274210
rect 113033 274176 113061 274210
rect 113105 274176 113129 274210
rect 113177 274176 113197 274210
rect 113249 274176 113265 274210
rect 113321 274176 113333 274210
rect 113393 274176 113401 274210
rect 113465 274176 113469 274210
rect 113571 274176 113575 274210
rect 113639 274176 113647 274210
rect 113707 274176 113719 274210
rect 113775 274176 113791 274210
rect 113843 274176 113863 274210
rect 113911 274176 113935 274210
rect 113979 274176 114007 274210
rect 114047 274206 114243 274210
rect 114047 274176 114074 274206
rect 112898 274117 112932 274164
rect 112898 274047 112932 274081
rect 112898 273964 112932 274011
rect 114108 274117 114142 274164
rect 114108 274047 114142 274081
rect 114108 273964 114142 274011
rect 114210 274110 114243 274206
rect 114345 274110 114353 274212
rect 114210 274086 114353 274110
rect 114455 274233 114489 274265
rect 114455 274165 114489 274199
rect 114652 274185 114862 274265
rect 114652 274151 114672 274185
rect 114738 274151 114740 274185
rect 114774 274151 114776 274185
rect 114842 274151 114862 274185
rect 114652 274150 114862 274151
rect 115027 274233 115178 274265
rect 115061 274199 115144 274233
rect 115027 274165 115178 274199
rect 114455 274097 114489 274131
rect 112966 273918 112993 273952
rect 113033 273918 113061 273952
rect 113105 273918 113129 273952
rect 113177 273918 113197 273952
rect 113249 273918 113265 273952
rect 113321 273918 113333 273952
rect 113393 273918 113401 273952
rect 113465 273918 113469 273952
rect 113571 273918 113575 273952
rect 113639 273918 113647 273952
rect 113707 273918 113719 273952
rect 113775 273918 113791 273952
rect 113843 273918 113863 273952
rect 113911 273918 113935 273952
rect 113979 273918 114007 273952
rect 114047 273918 114074 273952
rect 111334 273590 111376 273914
rect 112772 273884 114074 273918
rect 112772 273878 112832 273884
rect 111520 273842 112832 273878
rect 111520 273808 111547 273842
rect 111587 273808 111615 273842
rect 111659 273808 111683 273842
rect 111731 273808 111751 273842
rect 111803 273808 111819 273842
rect 111875 273808 111887 273842
rect 111947 273808 111955 273842
rect 112019 273808 112023 273842
rect 112125 273808 112129 273842
rect 112193 273808 112201 273842
rect 112261 273808 112273 273842
rect 112329 273808 112345 273842
rect 112397 273808 112417 273842
rect 112465 273808 112489 273842
rect 112533 273808 112561 273842
rect 112601 273808 112628 273842
rect 111452 273769 111486 273796
rect 111452 273699 111486 273733
rect 111452 273636 111486 273663
rect 112662 273769 112696 273796
rect 112662 273699 112696 273733
rect 112662 273636 112696 273663
rect 111520 273590 111547 273624
rect 111587 273590 111615 273624
rect 111659 273590 111683 273624
rect 111731 273590 111751 273624
rect 111803 273590 111819 273624
rect 111875 273590 111887 273624
rect 111947 273590 111955 273624
rect 112019 273590 112023 273624
rect 112125 273590 112129 273624
rect 112193 273590 112201 273624
rect 112261 273590 112273 273624
rect 112329 273590 112345 273624
rect 112397 273590 112417 273624
rect 112465 273590 112489 273624
rect 112533 273590 112561 273624
rect 112601 273590 112628 273624
rect 111334 273554 112628 273590
rect 111334 273230 111376 273554
rect 112772 273518 112832 273842
rect 114210 273820 114246 274086
rect 112966 273786 114246 273820
rect 114455 274029 114489 274063
rect 114455 273961 114489 273995
rect 114455 273893 114489 273927
rect 114455 273825 114489 273859
rect 112966 273752 112993 273786
rect 113033 273752 113061 273786
rect 113105 273752 113129 273786
rect 113177 273752 113197 273786
rect 113249 273752 113265 273786
rect 113321 273752 113333 273786
rect 113393 273752 113401 273786
rect 113465 273752 113469 273786
rect 113571 273752 113575 273786
rect 113639 273752 113647 273786
rect 113707 273752 113719 273786
rect 113775 273752 113791 273786
rect 113843 273752 113863 273786
rect 113911 273752 113935 273786
rect 113979 273752 114007 273786
rect 114047 273752 114074 273786
rect 114455 273757 114489 273791
rect 112898 273693 112932 273740
rect 112898 273623 112932 273657
rect 112898 273540 112932 273587
rect 114108 273693 114142 273740
rect 114108 273623 114142 273657
rect 114108 273540 114142 273587
rect 114455 273689 114489 273723
rect 114455 273621 114489 273655
rect 114455 273553 114489 273587
rect 111520 273496 112832 273518
rect 112966 273496 112993 273528
rect 111520 273494 112993 273496
rect 113033 273494 113061 273528
rect 113105 273494 113129 273528
rect 113177 273494 113197 273528
rect 113249 273494 113265 273528
rect 113321 273494 113333 273528
rect 113393 273494 113401 273528
rect 113465 273494 113469 273528
rect 113571 273494 113575 273528
rect 113639 273494 113647 273528
rect 113707 273494 113719 273528
rect 113775 273494 113791 273528
rect 113843 273494 113863 273528
rect 113911 273494 113935 273528
rect 113979 273494 114007 273528
rect 114047 273494 114074 273528
rect 111520 273482 114074 273494
rect 111520 273448 111547 273482
rect 111587 273448 111615 273482
rect 111659 273448 111683 273482
rect 111731 273448 111751 273482
rect 111803 273448 111819 273482
rect 111875 273448 111887 273482
rect 111947 273448 111955 273482
rect 112019 273448 112023 273482
rect 112125 273448 112129 273482
rect 112193 273448 112201 273482
rect 112261 273448 112273 273482
rect 112329 273448 112345 273482
rect 112397 273448 112417 273482
rect 112465 273448 112489 273482
rect 112533 273448 112561 273482
rect 112601 273448 112628 273482
rect 112744 273479 114074 273482
rect 114455 273485 114489 273519
rect 112744 273462 114396 273479
rect 111452 273409 111486 273436
rect 111452 273339 111486 273373
rect 111452 273276 111486 273303
rect 112662 273409 112696 273436
rect 112662 273339 112696 273373
rect 112662 273276 112696 273303
rect 111520 273230 111547 273264
rect 111587 273230 111615 273264
rect 111659 273230 111683 273264
rect 111731 273230 111751 273264
rect 111803 273230 111819 273264
rect 111875 273230 111887 273264
rect 111947 273230 111955 273264
rect 112019 273230 112023 273264
rect 112125 273230 112129 273264
rect 112193 273230 112201 273264
rect 112261 273230 112273 273264
rect 112329 273230 112345 273264
rect 112397 273230 112417 273264
rect 112465 273230 112489 273264
rect 112533 273230 112561 273264
rect 112601 273230 112628 273264
rect 111334 273194 112628 273230
rect 111334 272870 111376 273194
rect 112744 273158 112780 273462
rect 113892 273443 114396 273462
rect 111520 273122 112780 273158
rect 112832 273384 113264 273418
rect 112832 273376 113023 273384
rect 112832 273122 112872 273376
rect 112996 273350 113023 273376
rect 113063 273350 113091 273384
rect 113135 273350 113159 273384
rect 113207 273350 113227 273384
rect 113279 273350 113295 273384
rect 113351 273350 113363 273384
rect 113423 273350 113431 273384
rect 113495 273350 113499 273384
rect 113601 273350 113605 273384
rect 113669 273350 113677 273384
rect 113737 273350 113749 273384
rect 113805 273350 113821 273384
rect 113873 273350 113893 273384
rect 113941 273350 113965 273384
rect 114009 273350 114037 273384
rect 114077 273350 114104 273384
rect 112928 273315 112962 273338
rect 112928 273258 112962 273281
rect 114138 273315 114172 273338
rect 114138 273258 114172 273281
rect 114324 273287 114396 273443
rect 114324 273253 114342 273287
rect 114376 273253 114396 273287
rect 112996 273218 113023 273246
rect 112994 273212 113023 273218
rect 113063 273212 113091 273246
rect 113135 273212 113159 273246
rect 113207 273212 113227 273246
rect 113279 273212 113295 273246
rect 113351 273212 113363 273246
rect 113423 273212 113431 273246
rect 113495 273212 113499 273246
rect 113601 273212 113605 273246
rect 113669 273212 113677 273246
rect 113737 273212 113749 273246
rect 113805 273212 113821 273246
rect 113873 273212 113893 273246
rect 113941 273212 113965 273246
rect 114009 273212 114037 273246
rect 114077 273218 114104 273246
rect 114077 273212 114274 273218
rect 112994 273172 114274 273212
rect 114324 273205 114396 273253
rect 114455 273417 114489 273451
rect 114455 273349 114489 273383
rect 114455 273281 114489 273315
rect 114576 274100 114610 274139
rect 114576 274028 114610 274058
rect 114576 273956 114610 273990
rect 114576 273888 114610 273922
rect 114576 273820 114610 273850
rect 114576 273611 114610 273778
rect 114904 274100 114938 274139
rect 114904 274028 114938 274058
rect 114904 273956 114938 273990
rect 114904 273888 114938 273922
rect 114904 273820 114938 273850
rect 114653 273693 114672 273727
rect 114738 273693 114740 273727
rect 114774 273693 114776 273727
rect 114842 273693 114861 273727
rect 114904 273647 114938 273778
rect 115061 274131 115144 274165
rect 115343 274185 115553 274265
rect 115343 274151 115363 274185
rect 115429 274151 115431 274185
rect 115465 274151 115467 274185
rect 115533 274151 115553 274185
rect 115343 274150 115553 274151
rect 115716 274233 115750 274265
rect 116183 274240 117169 274332
rect 115959 274236 117169 274240
rect 115716 274165 115750 274199
rect 115027 274097 115178 274131
rect 115061 274063 115144 274097
rect 115027 274029 115178 274063
rect 115061 273995 115144 274029
rect 115027 273961 115178 273995
rect 115061 273927 115144 273961
rect 115027 273893 115178 273927
rect 115061 273859 115144 273893
rect 115027 273825 115178 273859
rect 115061 273791 115144 273825
rect 115027 273757 115178 273791
rect 115061 273723 115144 273757
rect 115027 273689 115178 273723
rect 115061 273655 115144 273689
rect 114865 273613 114970 273647
rect 114865 273611 114899 273613
rect 114576 273579 114899 273611
rect 114933 273579 114970 273613
rect 114576 273563 114970 273579
rect 114576 273426 114610 273563
rect 114865 273540 114970 273563
rect 115027 273621 115178 273655
rect 115267 274100 115301 274139
rect 115267 274028 115301 274058
rect 115267 273956 115301 273990
rect 115267 273888 115301 273922
rect 115267 273820 115301 273850
rect 115267 273647 115301 273778
rect 115595 274100 115629 274139
rect 115595 274028 115629 274058
rect 115595 273956 115629 273990
rect 115595 273888 115629 273922
rect 115595 273820 115629 273850
rect 115344 273693 115363 273727
rect 115429 273693 115431 273727
rect 115465 273693 115467 273727
rect 115533 273693 115552 273727
rect 115061 273587 115144 273621
rect 115027 273553 115178 273587
rect 114653 273465 114672 273499
rect 114738 273465 114740 273499
rect 114774 273465 114776 273499
rect 114842 273465 114861 273499
rect 114576 273356 114610 273390
rect 114576 273293 114610 273320
rect 114904 273426 114938 273540
rect 114904 273356 114938 273390
rect 114904 273293 114938 273320
rect 115061 273519 115144 273553
rect 115235 273613 115340 273647
rect 115235 273579 115271 273613
rect 115305 273611 115340 273613
rect 115595 273611 115629 273778
rect 115305 273579 115629 273611
rect 115235 273563 115629 273579
rect 115235 273540 115340 273563
rect 115027 273485 115178 273519
rect 115061 273451 115144 273485
rect 115027 273417 115178 273451
rect 115061 273383 115144 273417
rect 115027 273349 115178 273383
rect 115061 273315 115144 273349
rect 115027 273281 115178 273315
rect 115267 273426 115301 273540
rect 115344 273465 115363 273499
rect 115429 273465 115431 273499
rect 115465 273465 115467 273499
rect 115533 273465 115552 273499
rect 115267 273356 115301 273390
rect 115267 273293 115301 273320
rect 115595 273426 115629 273563
rect 115595 273356 115629 273390
rect 115595 273293 115629 273320
rect 115716 274097 115750 274131
rect 115852 274235 117169 274236
rect 115852 274212 117239 274235
rect 115852 274110 115860 274212
rect 115962 274210 117239 274212
rect 115962 274206 116158 274210
rect 115962 274110 115995 274206
rect 116131 274176 116158 274206
rect 116198 274176 116226 274210
rect 116270 274176 116294 274210
rect 116342 274176 116362 274210
rect 116414 274176 116430 274210
rect 116486 274176 116498 274210
rect 116558 274176 116566 274210
rect 116630 274176 116634 274210
rect 116736 274176 116740 274210
rect 116804 274176 116812 274210
rect 116872 274176 116884 274210
rect 116940 274176 116956 274210
rect 117008 274176 117028 274210
rect 117076 274176 117100 274210
rect 117144 274176 117172 274210
rect 117212 274176 117239 274210
rect 117391 274202 118685 274238
rect 115852 274086 115995 274110
rect 115716 274029 115750 274063
rect 115716 273961 115750 273995
rect 115716 273893 115750 273927
rect 115716 273825 115750 273859
rect 115716 273757 115750 273791
rect 115959 273820 115995 274086
rect 116063 274117 116097 274164
rect 116063 274047 116097 274081
rect 116063 273964 116097 274011
rect 117273 274117 117307 274164
rect 117273 274047 117307 274081
rect 117273 273964 117307 274011
rect 116131 273918 116158 273952
rect 116198 273918 116226 273952
rect 116270 273918 116294 273952
rect 116342 273918 116362 273952
rect 116414 273918 116430 273952
rect 116486 273918 116498 273952
rect 116558 273918 116566 273952
rect 116630 273918 116634 273952
rect 116736 273918 116740 273952
rect 116804 273918 116812 273952
rect 116872 273918 116884 273952
rect 116940 273918 116956 273952
rect 117008 273918 117028 273952
rect 117076 273918 117100 273952
rect 117144 273918 117172 273952
rect 117212 273918 117239 273952
rect 117391 273918 117433 274202
rect 117577 274168 117604 274202
rect 117644 274168 117672 274202
rect 117716 274168 117740 274202
rect 117788 274168 117808 274202
rect 117860 274168 117876 274202
rect 117932 274168 117944 274202
rect 118004 274168 118012 274202
rect 118076 274168 118080 274202
rect 118182 274168 118186 274202
rect 118250 274168 118258 274202
rect 118318 274168 118330 274202
rect 118386 274168 118402 274202
rect 118454 274168 118474 274202
rect 118522 274168 118546 274202
rect 118590 274168 118618 274202
rect 118658 274168 118685 274202
rect 117509 274129 117543 274156
rect 117509 274059 117543 274093
rect 117509 273996 117543 274023
rect 118719 274129 118753 274156
rect 118719 274059 118753 274093
rect 118719 273996 118753 274023
rect 116131 273884 117433 273918
rect 117577 273950 117604 273984
rect 117644 273950 117672 273984
rect 117716 273950 117740 273984
rect 117788 273950 117808 273984
rect 117860 273950 117876 273984
rect 117932 273950 117944 273984
rect 118004 273950 118012 273984
rect 118076 273950 118080 273984
rect 118182 273950 118186 273984
rect 118250 273950 118258 273984
rect 118318 273950 118330 273984
rect 118386 273950 118402 273984
rect 118454 273950 118474 273984
rect 118522 273950 118546 273984
rect 118590 273950 118618 273984
rect 118658 273950 118685 273984
rect 117577 273914 118871 273950
rect 117373 273878 117433 273884
rect 117373 273842 118685 273878
rect 115959 273786 117239 273820
rect 116131 273752 116158 273786
rect 116198 273752 116226 273786
rect 116270 273752 116294 273786
rect 116342 273752 116362 273786
rect 116414 273752 116430 273786
rect 116486 273752 116498 273786
rect 116558 273752 116566 273786
rect 116630 273752 116634 273786
rect 116736 273752 116740 273786
rect 116804 273752 116812 273786
rect 116872 273752 116884 273786
rect 116940 273752 116956 273786
rect 117008 273752 117028 273786
rect 117076 273752 117100 273786
rect 117144 273752 117172 273786
rect 117212 273752 117239 273786
rect 115716 273689 115750 273723
rect 115716 273621 115750 273655
rect 115716 273553 115750 273587
rect 116063 273693 116097 273740
rect 116063 273623 116097 273657
rect 116063 273540 116097 273587
rect 117273 273693 117307 273740
rect 117273 273623 117307 273657
rect 117273 273540 117307 273587
rect 115716 273485 115750 273519
rect 116131 273494 116158 273528
rect 116198 273494 116226 273528
rect 116270 273494 116294 273528
rect 116342 273494 116362 273528
rect 116414 273494 116430 273528
rect 116486 273494 116498 273528
rect 116558 273494 116566 273528
rect 116630 273494 116634 273528
rect 116736 273494 116740 273528
rect 116804 273494 116812 273528
rect 116872 273494 116884 273528
rect 116940 273494 116956 273528
rect 117008 273494 117028 273528
rect 117076 273494 117100 273528
rect 117144 273494 117172 273528
rect 117212 273496 117239 273528
rect 117373 273518 117433 273842
rect 117577 273808 117604 273842
rect 117644 273808 117672 273842
rect 117716 273808 117740 273842
rect 117788 273808 117808 273842
rect 117860 273808 117876 273842
rect 117932 273808 117944 273842
rect 118004 273808 118012 273842
rect 118076 273808 118080 273842
rect 118182 273808 118186 273842
rect 118250 273808 118258 273842
rect 118318 273808 118330 273842
rect 118386 273808 118402 273842
rect 118454 273808 118474 273842
rect 118522 273808 118546 273842
rect 118590 273808 118618 273842
rect 118658 273808 118685 273842
rect 117509 273769 117543 273796
rect 117509 273699 117543 273733
rect 117509 273636 117543 273663
rect 118719 273769 118753 273796
rect 118719 273699 118753 273733
rect 118719 273636 118753 273663
rect 117577 273590 117604 273624
rect 117644 273590 117672 273624
rect 117716 273590 117740 273624
rect 117788 273590 117808 273624
rect 117860 273590 117876 273624
rect 117932 273590 117944 273624
rect 118004 273590 118012 273624
rect 118076 273590 118080 273624
rect 118182 273590 118186 273624
rect 118250 273590 118258 273624
rect 118318 273590 118330 273624
rect 118386 273590 118402 273624
rect 118454 273590 118474 273624
rect 118522 273590 118546 273624
rect 118590 273590 118618 273624
rect 118658 273590 118685 273624
rect 118829 273590 118871 273914
rect 117577 273554 118871 273590
rect 117373 273496 118685 273518
rect 117212 273494 118685 273496
rect 116131 273482 118685 273494
rect 116131 273479 117461 273482
rect 115716 273417 115750 273451
rect 115716 273349 115750 273383
rect 115716 273281 115750 273315
rect 114455 273213 114489 273247
rect 111520 273088 111547 273122
rect 111587 273088 111615 273122
rect 111659 273088 111683 273122
rect 111731 273088 111751 273122
rect 111803 273088 111819 273122
rect 111875 273088 111887 273122
rect 111947 273088 111955 273122
rect 112019 273088 112023 273122
rect 112125 273088 112129 273122
rect 112193 273088 112201 273122
rect 112261 273088 112273 273122
rect 112329 273088 112345 273122
rect 112397 273088 112417 273122
rect 112465 273088 112489 273122
rect 112533 273088 112561 273122
rect 112601 273088 112628 273122
rect 112832 273086 113216 273122
rect 112832 273082 113023 273086
rect 111452 273049 111486 273076
rect 111452 272979 111486 273013
rect 111452 272916 111486 272943
rect 112662 273049 112696 273076
rect 112832 273054 112872 273082
rect 112996 273052 113023 273082
rect 113063 273052 113091 273086
rect 113135 273052 113159 273086
rect 113207 273052 113227 273086
rect 113279 273052 113295 273086
rect 113351 273052 113363 273086
rect 113423 273052 113431 273086
rect 113495 273052 113499 273086
rect 113601 273052 113605 273086
rect 113669 273052 113677 273086
rect 113737 273052 113749 273086
rect 113805 273052 113821 273086
rect 113873 273052 113893 273086
rect 113941 273052 113965 273086
rect 114009 273052 114037 273086
rect 114077 273052 114104 273086
rect 112662 272979 112696 273013
rect 112928 273017 112962 273040
rect 112928 272960 112962 272983
rect 114138 273017 114172 273040
rect 114138 272960 114172 272983
rect 112662 272916 112696 272943
rect 112996 272914 113023 272948
rect 113063 272914 113091 272948
rect 113135 272914 113159 272948
rect 113207 272914 113227 272948
rect 113279 272914 113295 272948
rect 113351 272914 113363 272948
rect 113423 272914 113431 272948
rect 113495 272914 113499 272948
rect 113601 272914 113605 272948
rect 113669 272914 113677 272948
rect 113737 272914 113749 272948
rect 113805 272914 113821 272948
rect 113873 272914 113893 272948
rect 113941 272914 113965 272948
rect 114009 272914 114037 272948
rect 114077 272914 114104 272948
rect 114234 272914 114274 273172
rect 114653 273247 114672 273281
rect 114738 273247 114740 273281
rect 114774 273247 114776 273281
rect 114842 273247 114861 273281
rect 114653 273210 114709 273247
rect 114805 273212 114861 273247
rect 115061 273247 115144 273281
rect 115027 273213 115178 273247
rect 114455 273145 114489 273179
rect 114455 273077 114489 273111
rect 114455 273009 114489 273043
rect 114455 272941 114489 272975
rect 112994 272907 114455 272914
rect 111520 272870 111547 272904
rect 111587 272870 111615 272904
rect 111659 272870 111683 272904
rect 111731 272870 111751 272904
rect 111803 272870 111819 272904
rect 111875 272870 111887 272904
rect 111947 272870 111955 272904
rect 112019 272870 112023 272904
rect 112125 272870 112129 272904
rect 112193 272870 112201 272904
rect 112261 272870 112273 272904
rect 112329 272870 112345 272904
rect 112397 272870 112417 272904
rect 112465 272870 112489 272904
rect 112533 272870 112561 272904
rect 112601 272870 112628 272904
rect 111334 272834 112628 272870
rect 112994 272873 114489 272907
rect 114538 273171 114709 273210
rect 114804 273190 114991 273212
rect 114538 273045 114576 273171
rect 114804 273156 114899 273190
rect 114933 273156 114991 273190
rect 114804 273127 114991 273156
rect 115061 273179 115144 273213
rect 115344 273247 115363 273281
rect 115429 273247 115431 273281
rect 115465 273247 115467 273281
rect 115533 273247 115552 273281
rect 115344 273212 115400 273247
rect 115027 273145 115178 273179
rect 114653 273057 114672 273091
rect 114738 273057 114740 273091
rect 114774 273057 114776 273091
rect 114842 273057 114861 273091
rect 114938 273045 114975 273127
rect 114538 273018 114610 273045
rect 114538 272982 114576 273018
rect 114538 272948 114610 272982
rect 114538 272912 114576 272948
rect 114538 272885 114610 272912
rect 114904 273018 114975 273045
rect 114938 272982 114975 273018
rect 114904 272948 114975 272982
rect 114938 272912 114975 272948
rect 114904 272885 114975 272912
rect 115061 273111 115144 273145
rect 115214 273190 115401 273212
rect 115214 273156 115271 273190
rect 115305 273156 115401 273190
rect 115496 273210 115552 273247
rect 115716 273213 115750 273247
rect 115496 273171 115667 273210
rect 115214 273127 115401 273156
rect 115027 273077 115178 273111
rect 115061 273043 115144 273077
rect 115027 273009 115178 273043
rect 115061 272975 115144 273009
rect 115027 272941 115178 272975
rect 115061 272907 115144 272941
rect 115027 272873 115178 272907
rect 115230 273045 115267 273127
rect 115344 273057 115363 273091
rect 115429 273057 115431 273091
rect 115465 273057 115467 273091
rect 115533 273057 115552 273091
rect 115629 273045 115667 273171
rect 115230 273018 115301 273045
rect 115230 272982 115267 273018
rect 115230 272948 115301 272982
rect 115230 272912 115267 272948
rect 115230 272885 115301 272912
rect 115595 273018 115667 273045
rect 115629 272982 115667 273018
rect 115595 272948 115667 272982
rect 115629 272912 115667 272948
rect 115595 272885 115667 272912
rect 115809 273462 117461 273479
rect 115809 273443 116313 273462
rect 115809 273287 115881 273443
rect 116941 273384 117373 273418
rect 116101 273350 116128 273384
rect 116168 273350 116196 273384
rect 116240 273350 116264 273384
rect 116312 273350 116332 273384
rect 116384 273350 116400 273384
rect 116456 273350 116468 273384
rect 116528 273350 116536 273384
rect 116600 273350 116604 273384
rect 116706 273350 116710 273384
rect 116774 273350 116782 273384
rect 116842 273350 116854 273384
rect 116910 273350 116926 273384
rect 116978 273350 116998 273384
rect 117046 273350 117070 273384
rect 117114 273350 117142 273384
rect 117182 273376 117373 273384
rect 117182 273350 117209 273376
rect 115809 273253 115828 273287
rect 115862 273253 115881 273287
rect 116033 273315 116067 273338
rect 116033 273258 116067 273281
rect 117243 273315 117277 273338
rect 117243 273258 117277 273281
rect 115809 273205 115881 273253
rect 116101 273218 116128 273246
rect 115931 273212 116128 273218
rect 116168 273212 116196 273246
rect 116240 273212 116264 273246
rect 116312 273212 116332 273246
rect 116384 273212 116400 273246
rect 116456 273212 116468 273246
rect 116528 273212 116536 273246
rect 116600 273212 116604 273246
rect 116706 273212 116710 273246
rect 116774 273212 116782 273246
rect 116842 273212 116854 273246
rect 116910 273212 116926 273246
rect 116978 273212 116998 273246
rect 117046 273212 117070 273246
rect 117114 273212 117142 273246
rect 117182 273218 117209 273246
rect 117182 273212 117211 273218
rect 115716 273145 115750 273179
rect 115716 273077 115750 273111
rect 115716 273009 115750 273043
rect 115716 272941 115750 272975
rect 115931 273172 117211 273212
rect 115931 272914 115971 273172
rect 117333 273122 117373 273376
rect 117425 273158 117461 273462
rect 117577 273448 117604 273482
rect 117644 273448 117672 273482
rect 117716 273448 117740 273482
rect 117788 273448 117808 273482
rect 117860 273448 117876 273482
rect 117932 273448 117944 273482
rect 118004 273448 118012 273482
rect 118076 273448 118080 273482
rect 118182 273448 118186 273482
rect 118250 273448 118258 273482
rect 118318 273448 118330 273482
rect 118386 273448 118402 273482
rect 118454 273448 118474 273482
rect 118522 273448 118546 273482
rect 118590 273448 118618 273482
rect 118658 273448 118685 273482
rect 117509 273409 117543 273436
rect 117509 273339 117543 273373
rect 117509 273276 117543 273303
rect 118719 273409 118753 273436
rect 118719 273339 118753 273373
rect 118719 273276 118753 273303
rect 117577 273230 117604 273264
rect 117644 273230 117672 273264
rect 117716 273230 117740 273264
rect 117788 273230 117808 273264
rect 117860 273230 117876 273264
rect 117932 273230 117944 273264
rect 118004 273230 118012 273264
rect 118076 273230 118080 273264
rect 118182 273230 118186 273264
rect 118250 273230 118258 273264
rect 118318 273230 118330 273264
rect 118386 273230 118402 273264
rect 118454 273230 118474 273264
rect 118522 273230 118546 273264
rect 118590 273230 118618 273264
rect 118658 273230 118685 273264
rect 118829 273230 118871 273554
rect 117577 273194 118871 273230
rect 117425 273122 118685 273158
rect 116989 273086 117373 273122
rect 117577 273088 117604 273122
rect 117644 273088 117672 273122
rect 117716 273088 117740 273122
rect 117788 273088 117808 273122
rect 117860 273088 117876 273122
rect 117932 273088 117944 273122
rect 118004 273088 118012 273122
rect 118076 273088 118080 273122
rect 118182 273088 118186 273122
rect 118250 273088 118258 273122
rect 118318 273088 118330 273122
rect 118386 273088 118402 273122
rect 118454 273088 118474 273122
rect 118522 273088 118546 273122
rect 118590 273088 118618 273122
rect 118658 273088 118685 273122
rect 116101 273052 116128 273086
rect 116168 273052 116196 273086
rect 116240 273052 116264 273086
rect 116312 273052 116332 273086
rect 116384 273052 116400 273086
rect 116456 273052 116468 273086
rect 116528 273052 116536 273086
rect 116600 273052 116604 273086
rect 116706 273052 116710 273086
rect 116774 273052 116782 273086
rect 116842 273052 116854 273086
rect 116910 273052 116926 273086
rect 116978 273052 116998 273086
rect 117046 273052 117070 273086
rect 117114 273052 117142 273086
rect 117182 273082 117373 273086
rect 117182 273052 117209 273082
rect 117333 273054 117373 273082
rect 117509 273049 117543 273076
rect 116033 273017 116067 273040
rect 116033 272960 116067 272983
rect 117243 273017 117277 273040
rect 117243 272960 117277 272983
rect 117509 272979 117543 273013
rect 116101 272914 116128 272948
rect 116168 272914 116196 272948
rect 116240 272914 116264 272948
rect 116312 272914 116332 272948
rect 116384 272914 116400 272948
rect 116456 272914 116468 272948
rect 116528 272914 116536 272948
rect 116600 272914 116604 272948
rect 116706 272914 116710 272948
rect 116774 272914 116782 272948
rect 116842 272914 116854 272948
rect 116910 272914 116926 272948
rect 116978 272914 116998 272948
rect 117046 272914 117070 272948
rect 117114 272914 117142 272948
rect 117182 272914 117209 272948
rect 117509 272916 117543 272943
rect 118719 273049 118753 273076
rect 118719 272979 118753 273013
rect 118719 272916 118753 272943
rect 115750 272907 117211 272914
rect 115716 272873 117211 272907
rect 112994 272868 114455 272873
rect 114653 272839 114672 272873
rect 114738 272839 114740 272873
rect 114774 272839 114776 272873
rect 114842 272839 114861 272873
rect 115061 272839 115144 272873
rect 115344 272839 115363 272873
rect 115429 272839 115431 272873
rect 115465 272839 115467 272873
rect 115533 272839 115552 272873
rect 115750 272868 117211 272873
rect 117577 272870 117604 272904
rect 117644 272870 117672 272904
rect 117716 272870 117740 272904
rect 117788 272870 117808 272904
rect 117860 272870 117876 272904
rect 117932 272870 117944 272904
rect 118004 272870 118012 272904
rect 118076 272870 118080 272904
rect 118182 272870 118186 272904
rect 118250 272870 118258 272904
rect 118318 272870 118330 272904
rect 118386 272870 118402 272904
rect 118454 272870 118474 272904
rect 118522 272870 118546 272904
rect 118590 272870 118618 272904
rect 118658 272870 118685 272904
rect 118829 272870 118871 273194
rect 114455 272805 114489 272839
rect 115027 272825 115178 272839
rect 113982 272761 114266 272766
rect 111046 272683 111200 272704
rect 111312 272735 114266 272761
rect 111312 272733 114034 272735
rect 114068 272733 114106 272735
rect 114140 272733 114178 272735
rect 114212 272733 114266 272735
rect 111312 272699 111340 272733
rect 111374 272699 111408 272733
rect 111442 272699 111476 272733
rect 111510 272699 111544 272733
rect 111578 272699 111612 272733
rect 111646 272699 111680 272733
rect 111714 272699 111748 272733
rect 111782 272699 111816 272733
rect 111850 272699 111884 272733
rect 111918 272699 111952 272733
rect 111986 272699 112020 272733
rect 112054 272699 112088 272733
rect 112122 272699 112156 272733
rect 112190 272699 112224 272733
rect 112258 272699 112292 272733
rect 112326 272699 112360 272733
rect 112394 272699 112428 272733
rect 112462 272699 112496 272733
rect 112530 272699 112564 272733
rect 112598 272699 112632 272733
rect 112666 272699 112700 272733
rect 112734 272699 112768 272733
rect 112802 272699 112836 272733
rect 112870 272699 112904 272733
rect 112938 272699 112972 272733
rect 113006 272699 113040 272733
rect 113074 272699 113108 272733
rect 113142 272699 113176 272733
rect 113210 272699 113244 272733
rect 113278 272699 113312 272733
rect 113346 272699 113380 272733
rect 113414 272699 113448 272733
rect 113482 272699 113516 272733
rect 113550 272699 113584 272733
rect 113618 272699 113652 272733
rect 113686 272699 113720 272733
rect 113754 272699 113788 272733
rect 113822 272699 113856 272733
rect 113890 272699 113924 272733
rect 113958 272699 113992 272733
rect 114026 272701 114034 272733
rect 114094 272701 114106 272733
rect 114162 272701 114178 272733
rect 114026 272699 114060 272701
rect 114094 272699 114128 272701
rect 114162 272699 114196 272701
rect 114230 272699 114266 272733
rect 114455 272739 114489 272771
rect 114928 272805 115275 272825
rect 114928 272771 115027 272805
rect 115061 272771 115144 272805
rect 115178 272771 115275 272805
rect 114928 272766 115275 272771
rect 114928 272739 115016 272766
rect 114455 272705 114537 272739
rect 114571 272705 114605 272739
rect 114639 272705 114673 272739
rect 114707 272705 114741 272739
rect 114775 272705 114809 272739
rect 114843 272705 114877 272739
rect 114911 272705 114945 272739
rect 114979 272705 115016 272739
rect 111312 272671 114266 272699
rect 109951 270204 110259 270212
rect 106281 270169 110259 270204
rect 111939 272249 112069 272265
rect 112673 272249 113101 272671
rect 113982 272666 114266 272671
rect 114928 272444 115016 272705
rect 115194 272739 115275 272766
rect 115716 272805 115750 272839
rect 117577 272834 118871 272870
rect 115716 272739 115750 272771
rect 115194 272705 115226 272739
rect 115260 272705 115294 272739
rect 115328 272705 115362 272739
rect 115396 272705 115430 272739
rect 115464 272705 115498 272739
rect 115532 272705 115566 272739
rect 115600 272705 115634 272739
rect 115668 272705 115750 272739
rect 115939 272761 116223 272766
rect 119005 272762 119031 281099
rect 118762 272761 119031 272762
rect 115939 272735 119031 272761
rect 115939 272733 115992 272735
rect 116026 272733 116064 272735
rect 116098 272733 116136 272735
rect 116170 272733 119031 272735
rect 115194 272444 115275 272705
rect 115939 272699 115975 272733
rect 116026 272701 116043 272733
rect 116098 272701 116111 272733
rect 116170 272701 116179 272733
rect 116009 272699 116043 272701
rect 116077 272699 116111 272701
rect 116145 272699 116179 272701
rect 116213 272699 116247 272733
rect 116281 272699 116315 272733
rect 116349 272699 116383 272733
rect 116417 272699 116451 272733
rect 116485 272699 116519 272733
rect 116553 272699 116587 272733
rect 116621 272699 116655 272733
rect 116689 272699 116723 272733
rect 116757 272699 116791 272733
rect 116825 272699 116859 272733
rect 116893 272699 116927 272733
rect 116961 272699 116995 272733
rect 117029 272699 117063 272733
rect 117097 272699 117131 272733
rect 117165 272699 117199 272733
rect 117233 272699 117267 272733
rect 117301 272699 117335 272733
rect 117369 272699 117403 272733
rect 117437 272699 117471 272733
rect 117505 272699 117539 272733
rect 117573 272699 117607 272733
rect 117641 272699 117675 272733
rect 117709 272699 117743 272733
rect 117777 272699 117811 272733
rect 117845 272699 117879 272733
rect 117913 272699 117947 272733
rect 117981 272699 118015 272733
rect 118049 272699 118083 272733
rect 118117 272699 118151 272733
rect 118185 272699 118219 272733
rect 118253 272699 118287 272733
rect 118321 272699 118355 272733
rect 118389 272699 118423 272733
rect 118457 272699 118491 272733
rect 118525 272699 118559 272733
rect 118593 272699 118627 272733
rect 118661 272699 118695 272733
rect 118729 272699 118763 272733
rect 118797 272699 118831 272733
rect 118865 272704 119031 272733
rect 119133 272704 119159 281102
rect 118865 272699 119159 272704
rect 115939 272683 119159 272699
rect 119938 281139 125658 281165
rect 119938 281059 120256 281139
rect 115939 272671 119158 272683
rect 115939 272666 116223 272671
rect 114928 272372 115275 272444
rect 116523 272249 119158 272671
rect 111939 272247 119158 272249
rect 107329 268607 108364 270169
rect 111939 268677 111953 272247
rect 112055 272238 119035 272247
rect 112055 272136 112178 272238
rect 118944 272136 119035 272238
rect 112055 272125 119035 272136
rect 112055 268826 112069 272125
rect 116590 272098 118192 272125
rect 113800 271981 114102 272051
rect 113800 271731 113863 271981
rect 114041 271731 114102 271981
rect 114984 272036 115601 272048
rect 114984 271996 118841 272036
rect 114984 271984 115908 271996
rect 114984 271950 115019 271984
rect 115053 271950 115091 271984
rect 115125 271950 115163 271984
rect 115197 271950 115235 271984
rect 115269 271950 115307 271984
rect 115341 271950 115379 271984
rect 115413 271950 115451 271984
rect 115485 271950 115523 271984
rect 115557 271981 115908 271984
rect 115557 271950 115601 271981
rect 114984 271886 115601 271950
rect 113800 271668 114102 271731
rect 112307 271634 112391 271668
rect 112425 271634 112459 271668
rect 112493 271634 112527 271668
rect 112561 271634 112595 271668
rect 112629 271634 112663 271668
rect 112697 271634 112731 271668
rect 112765 271634 112799 271668
rect 112833 271634 112867 271668
rect 112901 271634 112935 271668
rect 112969 271634 113003 271668
rect 113037 271634 113071 271668
rect 113105 271634 113139 271668
rect 113173 271634 113207 271668
rect 113241 271634 113275 271668
rect 113309 271634 113343 271668
rect 113377 271634 113411 271668
rect 113445 271634 113479 271668
rect 113513 271634 113547 271668
rect 113581 271634 113615 271668
rect 113649 271634 113683 271668
rect 113717 271634 113751 271668
rect 113785 271634 113819 271668
rect 113853 271634 113887 271668
rect 113921 271634 113955 271668
rect 113989 271634 114023 271668
rect 114057 271634 114091 271668
rect 114125 271634 114210 271668
rect 112307 271582 112341 271634
rect 112307 271514 112341 271548
rect 113068 271601 113461 271634
rect 113068 271567 113100 271601
rect 113134 271567 113172 271601
rect 113206 271567 113244 271601
rect 113278 271567 113316 271601
rect 113350 271567 113388 271601
rect 113422 271567 113461 271601
rect 113068 271524 113461 271567
rect 114176 271582 114210 271634
rect 114329 271567 114389 271588
rect 114210 271554 114389 271567
rect 114423 271554 114457 271588
rect 114491 271554 114525 271588
rect 114559 271554 114593 271588
rect 114627 271554 114661 271588
rect 114695 271554 114729 271588
rect 114763 271554 114797 271588
rect 114831 271554 114865 271588
rect 114899 271554 114933 271588
rect 114967 271554 115001 271588
rect 115035 271554 115069 271588
rect 115103 271554 115137 271588
rect 115171 271554 115205 271588
rect 115239 271554 115273 271588
rect 115307 271554 115341 271588
rect 115375 271554 115409 271588
rect 115443 271554 115503 271588
rect 114210 271548 114363 271554
rect 112307 271446 112341 271480
rect 112307 271378 112341 271412
rect 114176 271514 114363 271548
rect 114210 271503 114363 271514
rect 114210 271480 114329 271503
rect 114176 271469 114329 271480
rect 114176 271446 114363 271469
rect 114210 271435 114363 271446
rect 114210 271412 114329 271435
rect 114176 271401 114329 271412
rect 112578 271353 112605 271387
rect 112641 271353 112675 271387
rect 112711 271353 113005 271387
rect 113041 271353 113075 271387
rect 113111 271353 113405 271387
rect 113441 271353 113475 271387
rect 113511 271353 113805 271387
rect 113841 271353 113875 271387
rect 113911 271353 113938 271387
rect 114176 271378 114363 271401
rect 112307 271310 112341 271344
rect 112307 271242 112341 271276
rect 112307 271174 112341 271208
rect 112307 271106 112341 271140
rect 112532 271291 112566 271310
rect 112532 271223 112566 271225
rect 112532 271187 112566 271189
rect 112532 271102 112566 271121
rect 112750 271291 112784 271310
rect 112750 271223 112784 271225
rect 112750 271187 112784 271189
rect 112750 271102 112784 271121
rect 112307 271038 112341 271072
rect 112838 271059 112886 271353
rect 112932 271291 112966 271310
rect 112932 271223 112966 271225
rect 112932 271187 112966 271189
rect 112932 271102 112966 271121
rect 113150 271291 113184 271310
rect 113150 271223 113184 271225
rect 113150 271187 113184 271189
rect 113150 271102 113184 271121
rect 113332 271291 113366 271310
rect 113332 271223 113366 271225
rect 113332 271187 113366 271189
rect 113332 271102 113366 271121
rect 113550 271291 113584 271310
rect 113550 271223 113584 271225
rect 113550 271187 113584 271189
rect 113550 271102 113584 271121
rect 113634 271059 113682 271353
rect 114210 271367 114363 271378
rect 114210 271344 114329 271367
rect 114176 271333 114329 271344
rect 114176 271310 114363 271333
rect 114637 271324 114664 271358
rect 114700 271324 114734 271358
rect 114770 271324 114797 271358
rect 113732 271291 113766 271310
rect 113732 271223 113766 271225
rect 113732 271187 113766 271189
rect 113732 271102 113766 271121
rect 113950 271291 113984 271310
rect 113950 271223 113984 271225
rect 113950 271187 113984 271189
rect 113950 271102 113984 271121
rect 114210 271299 114363 271310
rect 114210 271276 114329 271299
rect 114176 271265 114329 271276
rect 114176 271242 114363 271265
rect 114210 271231 114363 271242
rect 114210 271208 114329 271231
rect 114176 271197 114329 271208
rect 114176 271174 114363 271197
rect 114210 271163 114363 271174
rect 114210 271140 114329 271163
rect 114176 271129 114329 271140
rect 114176 271106 114363 271129
rect 114210 271095 114363 271106
rect 114210 271072 114329 271095
rect 114176 271061 114329 271072
rect 114591 271262 114625 271281
rect 114591 271194 114625 271196
rect 114591 271158 114625 271160
rect 114591 271073 114625 271092
rect 114809 271279 114843 271281
rect 114890 271279 114942 271554
rect 115469 271503 115503 271554
rect 115469 271435 115503 271469
rect 115337 271373 115382 271375
rect 115060 271358 115382 271373
rect 115037 271324 115064 271358
rect 115100 271324 115134 271358
rect 115170 271331 115382 271358
rect 115170 271324 115197 271331
rect 114991 271279 115025 271281
rect 114809 271262 115025 271279
rect 114843 271229 114991 271262
rect 114809 271194 114843 271196
rect 114809 271158 114843 271160
rect 114809 271073 114843 271092
rect 114991 271194 115025 271196
rect 114991 271158 115025 271160
rect 114991 271073 115025 271092
rect 115209 271262 115243 271281
rect 115209 271194 115243 271196
rect 115209 271158 115243 271160
rect 115209 271073 115243 271092
rect 112578 271025 112605 271059
rect 112641 271025 112675 271059
rect 112711 271025 113005 271059
rect 113041 271025 113075 271059
rect 113111 271025 113405 271059
rect 113441 271025 113475 271059
rect 113511 271025 113805 271059
rect 113841 271025 113875 271059
rect 113911 271025 113938 271059
rect 114176 271038 114363 271061
rect 112307 270970 112341 271004
rect 112307 270902 112341 270936
rect 112307 270817 112341 270868
rect 114210 271027 114363 271038
rect 114210 271004 114329 271027
rect 114176 270993 114329 271004
rect 114637 270996 114664 271030
rect 114700 270996 114734 271030
rect 114770 270996 115064 271030
rect 115100 270996 115134 271030
rect 115170 271014 115197 271030
rect 115337 271014 115382 271331
rect 115170 270996 115382 271014
rect 114176 270970 114363 270993
rect 115074 270973 115382 270996
rect 115469 271367 115503 271401
rect 115469 271299 115503 271333
rect 115469 271231 115503 271265
rect 115469 271163 115503 271197
rect 115469 271095 115503 271129
rect 115469 271027 115503 271061
rect 115074 270972 115369 270973
rect 114210 270959 114363 270970
rect 114210 270936 114329 270959
rect 114176 270925 114329 270936
rect 114176 270902 114363 270925
rect 114210 270891 114363 270902
rect 114210 270868 114329 270891
rect 114176 270857 114329 270868
rect 114176 270817 114363 270857
rect 112307 270783 112391 270817
rect 112425 270783 112459 270817
rect 112493 270783 112527 270817
rect 112561 270783 112595 270817
rect 112629 270783 112663 270817
rect 112697 270783 112731 270817
rect 112765 270783 112799 270817
rect 112833 270783 112867 270817
rect 112901 270783 112935 270817
rect 112969 270783 113003 270817
rect 113037 270783 113071 270817
rect 113105 270783 113139 270817
rect 113173 270783 113207 270817
rect 113241 270783 113275 270817
rect 113309 270783 113343 270817
rect 113377 270783 113411 270817
rect 113445 270783 113479 270817
rect 113513 270783 113547 270817
rect 113581 270783 113615 270817
rect 113649 270783 113683 270817
rect 113717 270783 113751 270817
rect 113785 270783 113819 270817
rect 113853 270783 113887 270817
rect 113921 270783 113955 270817
rect 113989 270783 114023 270817
rect 114057 270783 114091 270817
rect 114125 270806 114363 270817
rect 115469 270959 115503 270993
rect 115469 270891 115503 270925
rect 115469 270806 115503 270857
rect 114125 270789 114389 270806
rect 114125 270783 114210 270789
rect 114329 270772 114389 270789
rect 114423 270772 114457 270806
rect 114491 270772 114525 270806
rect 114559 270772 114593 270806
rect 114627 270772 114661 270806
rect 114695 270772 114729 270806
rect 114763 270772 114797 270806
rect 114831 270772 114865 270806
rect 114899 270772 114933 270806
rect 114967 270772 115001 270806
rect 115035 270772 115069 270806
rect 115103 270772 115137 270806
rect 115171 270772 115205 270806
rect 115239 270772 115273 270806
rect 115307 270772 115341 270806
rect 115375 270772 115409 270806
rect 115443 270772 115503 270806
rect 115648 270763 115700 271981
rect 115881 271962 115908 271981
rect 115944 271962 115978 271996
rect 116014 271962 116308 271996
rect 116344 271962 116378 271996
rect 116414 271962 116708 271996
rect 116744 271962 116778 271996
rect 116814 271962 117108 271996
rect 117144 271962 117178 271996
rect 117214 271962 117508 271996
rect 117544 271962 117578 271996
rect 117614 271962 117908 271996
rect 117944 271962 117978 271996
rect 118014 271962 118308 271996
rect 118344 271962 118378 271996
rect 118414 271962 118708 271996
rect 118744 271962 118778 271996
rect 118814 271962 118841 271996
rect 115835 271901 115869 271928
rect 115835 271833 115869 271861
rect 115835 271765 115869 271789
rect 115835 271697 115869 271717
rect 115835 271629 115869 271645
rect 115835 271561 115869 271573
rect 115835 271493 115869 271501
rect 115835 271425 115869 271429
rect 115835 271319 115869 271323
rect 115835 271247 115869 271255
rect 115835 271175 115869 271187
rect 115835 271103 115869 271119
rect 115835 271031 115869 271051
rect 115835 270959 115869 270983
rect 115835 270887 115869 270915
rect 115835 270820 115869 270847
rect 116053 271901 116087 271928
rect 116053 271833 116087 271861
rect 116053 271765 116087 271789
rect 116053 271697 116087 271717
rect 116053 271629 116087 271645
rect 116053 271561 116087 271573
rect 116053 271493 116087 271501
rect 116053 271425 116087 271429
rect 116053 271319 116087 271323
rect 116053 271247 116087 271255
rect 116053 271175 116087 271187
rect 116053 271103 116087 271119
rect 116053 271031 116087 271051
rect 116053 270959 116087 270983
rect 116053 270887 116087 270915
rect 116053 270820 116087 270847
rect 116235 271901 116269 271928
rect 116235 271833 116269 271861
rect 116235 271765 116269 271789
rect 116235 271697 116269 271717
rect 116235 271629 116269 271645
rect 116235 271561 116269 271573
rect 116235 271493 116269 271501
rect 116235 271425 116269 271429
rect 116235 271319 116269 271323
rect 116235 271247 116269 271255
rect 116235 271175 116269 271187
rect 116235 271103 116269 271119
rect 116235 271031 116269 271051
rect 116235 270959 116269 270983
rect 116235 270887 116269 270915
rect 116235 270820 116269 270847
rect 116453 271901 116487 271928
rect 116453 271833 116487 271861
rect 116453 271765 116487 271789
rect 116453 271697 116487 271717
rect 116453 271629 116487 271645
rect 116453 271561 116487 271573
rect 116453 271493 116487 271501
rect 116453 271425 116487 271429
rect 116453 271319 116487 271323
rect 116453 271247 116487 271255
rect 116453 271175 116487 271187
rect 116453 271103 116487 271119
rect 116453 271031 116487 271051
rect 116453 270959 116487 270983
rect 116453 270887 116487 270915
rect 116453 270820 116487 270847
rect 116635 271901 116669 271928
rect 116635 271833 116669 271861
rect 116635 271765 116669 271789
rect 116635 271697 116669 271717
rect 116635 271629 116669 271645
rect 116635 271561 116669 271573
rect 116635 271493 116669 271501
rect 116635 271425 116669 271429
rect 116635 271319 116669 271323
rect 116635 271247 116669 271255
rect 116635 271175 116669 271187
rect 116635 271103 116669 271119
rect 116635 271031 116669 271051
rect 116635 270959 116669 270983
rect 116635 270887 116669 270915
rect 116635 270820 116669 270847
rect 116853 271901 116887 271928
rect 116853 271833 116887 271861
rect 116853 271765 116887 271789
rect 116853 271697 116887 271717
rect 116853 271629 116887 271645
rect 116853 271561 116887 271573
rect 116853 271493 116887 271501
rect 116853 271425 116887 271429
rect 116853 271319 116887 271323
rect 116853 271247 116887 271255
rect 116853 271175 116887 271187
rect 116853 271103 116887 271119
rect 116853 271031 116887 271051
rect 116853 270959 116887 270983
rect 116853 270887 116887 270915
rect 116853 270820 116887 270847
rect 117035 271901 117069 271928
rect 117035 271833 117069 271861
rect 117035 271765 117069 271789
rect 117035 271697 117069 271717
rect 117035 271629 117069 271645
rect 117035 271561 117069 271573
rect 117035 271493 117069 271501
rect 117035 271425 117069 271429
rect 117035 271319 117069 271323
rect 117035 271247 117069 271255
rect 117035 271175 117069 271187
rect 117035 271103 117069 271119
rect 117035 271031 117069 271051
rect 117035 270959 117069 270983
rect 117035 270887 117069 270915
rect 117035 270820 117069 270847
rect 117253 271901 117287 271928
rect 117253 271833 117287 271861
rect 117253 271765 117287 271789
rect 117253 271697 117287 271717
rect 117253 271629 117287 271645
rect 117253 271561 117287 271573
rect 117253 271493 117287 271501
rect 117253 271425 117287 271429
rect 117253 271319 117287 271323
rect 117253 271247 117287 271255
rect 117253 271175 117287 271187
rect 117253 271103 117287 271119
rect 117253 271031 117287 271051
rect 117253 270959 117287 270983
rect 117253 270887 117287 270915
rect 117253 270820 117287 270847
rect 117435 271901 117469 271928
rect 117435 271833 117469 271861
rect 117435 271765 117469 271789
rect 117435 271697 117469 271717
rect 117435 271629 117469 271645
rect 117435 271561 117469 271573
rect 117435 271493 117469 271501
rect 117435 271425 117469 271429
rect 117435 271319 117469 271323
rect 117435 271247 117469 271255
rect 117435 271175 117469 271187
rect 117435 271103 117469 271119
rect 117435 271031 117469 271051
rect 117435 270959 117469 270983
rect 117435 270887 117469 270915
rect 117435 270820 117469 270847
rect 117653 271901 117687 271928
rect 117653 271833 117687 271861
rect 117653 271765 117687 271789
rect 117653 271697 117687 271717
rect 117653 271629 117687 271645
rect 117653 271561 117687 271573
rect 117653 271493 117687 271501
rect 117653 271425 117687 271429
rect 117653 271319 117687 271323
rect 117653 271247 117687 271255
rect 117653 271175 117687 271187
rect 117653 271103 117687 271119
rect 117653 271031 117687 271051
rect 117653 270959 117687 270983
rect 117653 270887 117687 270915
rect 117653 270820 117687 270847
rect 117835 271901 117869 271928
rect 117835 271833 117869 271861
rect 117835 271765 117869 271789
rect 117835 271697 117869 271717
rect 117835 271629 117869 271645
rect 117835 271561 117869 271573
rect 117835 271493 117869 271501
rect 117835 271425 117869 271429
rect 117835 271319 117869 271323
rect 117835 271247 117869 271255
rect 117835 271175 117869 271187
rect 117835 271103 117869 271119
rect 117835 271031 117869 271051
rect 117835 270959 117869 270983
rect 117835 270887 117869 270915
rect 117835 270820 117869 270847
rect 118053 271901 118087 271928
rect 118053 271833 118087 271861
rect 118053 271765 118087 271789
rect 118053 271697 118087 271717
rect 118053 271629 118087 271645
rect 118053 271561 118087 271573
rect 118053 271493 118087 271501
rect 118053 271425 118087 271429
rect 118053 271319 118087 271323
rect 118053 271247 118087 271255
rect 118053 271175 118087 271187
rect 118053 271103 118087 271119
rect 118053 271031 118087 271051
rect 118053 270959 118087 270983
rect 118053 270887 118087 270915
rect 118053 270820 118087 270847
rect 118235 271901 118269 271928
rect 118235 271833 118269 271861
rect 118235 271765 118269 271789
rect 118235 271697 118269 271717
rect 118235 271629 118269 271645
rect 118235 271561 118269 271573
rect 118235 271493 118269 271501
rect 118235 271425 118269 271429
rect 118235 271319 118269 271323
rect 118235 271247 118269 271255
rect 118235 271175 118269 271187
rect 118235 271103 118269 271119
rect 118235 271031 118269 271051
rect 118235 270959 118269 270983
rect 118235 270887 118269 270915
rect 118235 270820 118269 270847
rect 118453 271901 118487 271928
rect 118453 271833 118487 271861
rect 118453 271765 118487 271789
rect 118453 271697 118487 271717
rect 118453 271629 118487 271645
rect 118453 271561 118487 271573
rect 118453 271493 118487 271501
rect 118453 271425 118487 271429
rect 118453 271319 118487 271323
rect 118453 271247 118487 271255
rect 118453 271175 118487 271187
rect 118453 271103 118487 271119
rect 118453 271031 118487 271051
rect 118453 270959 118487 270983
rect 118453 270887 118487 270915
rect 118453 270820 118487 270847
rect 118635 271901 118669 271928
rect 118635 271833 118669 271861
rect 118635 271765 118669 271789
rect 118635 271697 118669 271717
rect 118635 271629 118669 271645
rect 118635 271561 118669 271573
rect 118635 271493 118669 271501
rect 118635 271425 118669 271429
rect 118635 271319 118669 271323
rect 118635 271247 118669 271255
rect 118635 271175 118669 271187
rect 118635 271103 118669 271119
rect 118635 271031 118669 271051
rect 118635 270959 118669 270983
rect 118635 270887 118669 270915
rect 118635 270820 118669 270847
rect 118853 271901 118887 271928
rect 118853 271833 118887 271861
rect 118853 271765 118887 271789
rect 118853 271697 118887 271717
rect 118853 271629 118887 271645
rect 118853 271561 118887 271573
rect 118853 271493 118887 271501
rect 118853 271425 118887 271429
rect 118853 271319 118887 271323
rect 118853 271247 118887 271255
rect 118853 271175 118887 271187
rect 118853 271103 118887 271119
rect 118853 271031 118887 271051
rect 118853 270959 118887 270983
rect 118853 270887 118887 270915
rect 118853 270820 118887 270847
rect 115881 270763 115908 270786
rect 115648 270752 115908 270763
rect 115944 270752 115978 270786
rect 116014 270752 116308 270786
rect 116344 270752 116378 270786
rect 116414 270752 116708 270786
rect 116744 270752 116778 270786
rect 116814 270752 117108 270786
rect 117144 270752 117178 270786
rect 117214 270752 117508 270786
rect 117544 270752 117578 270786
rect 117614 270752 117908 270786
rect 117944 270752 117978 270786
rect 118014 270752 118308 270786
rect 118344 270752 118378 270786
rect 118414 270752 118708 270786
rect 118744 270752 118778 270786
rect 118814 270752 118841 270786
rect 115648 270715 118841 270752
rect 115648 270714 115700 270715
rect 114050 270641 114542 270693
rect 114050 270607 114096 270641
rect 114130 270607 114168 270641
rect 114202 270607 114240 270641
rect 114274 270607 114312 270641
rect 114346 270607 114384 270641
rect 114418 270607 114456 270641
rect 114490 270607 114542 270641
rect 114050 270545 114542 270607
rect 114364 270296 114537 270545
rect 118418 270296 118934 270326
rect 112560 270262 112587 270296
rect 112623 270262 112657 270296
rect 112693 270262 112987 270296
rect 113023 270262 113057 270296
rect 113093 270262 113387 270296
rect 113423 270262 113457 270296
rect 113493 270262 113787 270296
rect 113823 270262 113857 270296
rect 113893 270262 114187 270296
rect 114223 270262 114257 270296
rect 114293 270262 114587 270296
rect 114623 270262 114657 270296
rect 114693 270262 114987 270296
rect 115023 270262 115057 270296
rect 115093 270262 115387 270296
rect 115423 270262 115457 270296
rect 115493 270262 115787 270296
rect 115823 270262 115857 270296
rect 115893 270262 116187 270296
rect 116223 270262 116257 270296
rect 116293 270262 116587 270296
rect 116623 270262 116657 270296
rect 116693 270262 116987 270296
rect 117023 270262 117057 270296
rect 117093 270262 117387 270296
rect 117423 270262 117457 270296
rect 117493 270262 117787 270296
rect 117823 270262 117857 270296
rect 117893 270262 118187 270296
rect 118223 270262 118257 270296
rect 118293 270262 118587 270296
rect 118623 270262 118657 270296
rect 118693 270288 118934 270296
rect 118693 270262 118720 270288
rect 112514 270201 112548 270228
rect 112514 270133 112548 270161
rect 112514 270065 112548 270089
rect 112514 269997 112548 270017
rect 112514 269929 112548 269945
rect 112514 269861 112548 269873
rect 112514 269793 112548 269801
rect 112514 269725 112548 269729
rect 112514 269619 112548 269623
rect 112514 269547 112548 269555
rect 112514 269475 112548 269487
rect 112514 269403 112548 269419
rect 112514 269331 112548 269351
rect 112514 269259 112548 269283
rect 112514 269187 112548 269215
rect 112514 269120 112548 269147
rect 112732 270201 112766 270228
rect 112732 270133 112766 270161
rect 112732 270065 112766 270089
rect 112732 269997 112766 270017
rect 112732 269929 112766 269945
rect 112732 269861 112766 269873
rect 112732 269793 112766 269801
rect 112732 269725 112766 269729
rect 112732 269619 112766 269623
rect 112732 269547 112766 269555
rect 112732 269475 112766 269487
rect 112732 269403 112766 269419
rect 112732 269331 112766 269351
rect 112732 269259 112766 269283
rect 112732 269187 112766 269215
rect 112732 269120 112766 269147
rect 112914 270201 112948 270228
rect 112914 270133 112948 270161
rect 112914 270065 112948 270089
rect 112914 269997 112948 270017
rect 112914 269929 112948 269945
rect 112914 269861 112948 269873
rect 112914 269793 112948 269801
rect 112914 269725 112948 269729
rect 112914 269619 112948 269623
rect 112914 269547 112948 269555
rect 112914 269475 112948 269487
rect 112914 269403 112948 269419
rect 112914 269331 112948 269351
rect 112914 269259 112948 269283
rect 112914 269187 112948 269215
rect 112914 269120 112948 269147
rect 113132 270201 113166 270228
rect 113132 270133 113166 270161
rect 113132 270065 113166 270089
rect 113132 269997 113166 270017
rect 113132 269929 113166 269945
rect 113132 269861 113166 269873
rect 113132 269793 113166 269801
rect 113132 269725 113166 269729
rect 113132 269619 113166 269623
rect 113132 269547 113166 269555
rect 113132 269475 113166 269487
rect 113132 269403 113166 269419
rect 113132 269331 113166 269351
rect 113132 269259 113166 269283
rect 113132 269187 113166 269215
rect 113132 269120 113166 269147
rect 113314 270201 113348 270228
rect 113314 270133 113348 270161
rect 113314 270065 113348 270089
rect 113314 269997 113348 270017
rect 113314 269929 113348 269945
rect 113314 269861 113348 269873
rect 113314 269793 113348 269801
rect 113314 269725 113348 269729
rect 113314 269619 113348 269623
rect 113314 269547 113348 269555
rect 113314 269475 113348 269487
rect 113314 269403 113348 269419
rect 113314 269331 113348 269351
rect 113314 269259 113348 269283
rect 113314 269187 113348 269215
rect 113314 269120 113348 269147
rect 113532 270201 113566 270228
rect 113532 270133 113566 270161
rect 113532 270065 113566 270089
rect 113532 269997 113566 270017
rect 113532 269929 113566 269945
rect 113532 269861 113566 269873
rect 113532 269793 113566 269801
rect 113532 269725 113566 269729
rect 113532 269619 113566 269623
rect 113532 269547 113566 269555
rect 113532 269475 113566 269487
rect 113532 269403 113566 269419
rect 113532 269331 113566 269351
rect 113532 269259 113566 269283
rect 113532 269187 113566 269215
rect 113532 269120 113566 269147
rect 113714 270201 113748 270228
rect 113714 270133 113748 270161
rect 113714 270065 113748 270089
rect 113714 269997 113748 270017
rect 113714 269929 113748 269945
rect 113714 269861 113748 269873
rect 113714 269793 113748 269801
rect 113714 269725 113748 269729
rect 113714 269619 113748 269623
rect 113714 269547 113748 269555
rect 113714 269475 113748 269487
rect 113714 269403 113748 269419
rect 113714 269331 113748 269351
rect 113714 269259 113748 269283
rect 113714 269187 113748 269215
rect 113714 269120 113748 269147
rect 113932 270201 113966 270228
rect 113932 270133 113966 270161
rect 113932 270065 113966 270089
rect 113932 269997 113966 270017
rect 113932 269929 113966 269945
rect 113932 269861 113966 269873
rect 113932 269793 113966 269801
rect 113932 269725 113966 269729
rect 113932 269619 113966 269623
rect 113932 269547 113966 269555
rect 113932 269475 113966 269487
rect 113932 269403 113966 269419
rect 113932 269331 113966 269351
rect 113932 269259 113966 269283
rect 113932 269187 113966 269215
rect 113932 269120 113966 269147
rect 114114 270201 114148 270228
rect 114114 270133 114148 270161
rect 114114 270065 114148 270089
rect 114114 269997 114148 270017
rect 114114 269929 114148 269945
rect 114114 269861 114148 269873
rect 114114 269793 114148 269801
rect 114114 269725 114148 269729
rect 114114 269619 114148 269623
rect 114114 269547 114148 269555
rect 114114 269475 114148 269487
rect 114114 269403 114148 269419
rect 114114 269331 114148 269351
rect 114114 269259 114148 269283
rect 114114 269187 114148 269215
rect 114114 269120 114148 269147
rect 114332 270201 114366 270228
rect 114332 270133 114366 270161
rect 114332 270065 114366 270089
rect 114332 269997 114366 270017
rect 114332 269929 114366 269945
rect 114332 269861 114366 269873
rect 114332 269793 114366 269801
rect 114332 269725 114366 269729
rect 114332 269619 114366 269623
rect 114332 269547 114366 269555
rect 114332 269475 114366 269487
rect 114332 269403 114366 269419
rect 114332 269331 114366 269351
rect 114332 269259 114366 269283
rect 114332 269187 114366 269215
rect 114332 269120 114366 269147
rect 114514 270201 114548 270228
rect 114514 270133 114548 270161
rect 114514 270065 114548 270089
rect 114514 269997 114548 270017
rect 114514 269929 114548 269945
rect 114514 269861 114548 269873
rect 114514 269793 114548 269801
rect 114514 269725 114548 269729
rect 114514 269619 114548 269623
rect 114514 269547 114548 269555
rect 114514 269475 114548 269487
rect 114514 269403 114548 269419
rect 114514 269331 114548 269351
rect 114514 269259 114548 269283
rect 114514 269187 114548 269215
rect 114514 269120 114548 269147
rect 114732 270201 114766 270228
rect 114732 270133 114766 270161
rect 114732 270065 114766 270089
rect 114732 269997 114766 270017
rect 114732 269929 114766 269945
rect 114732 269861 114766 269873
rect 114732 269793 114766 269801
rect 114732 269725 114766 269729
rect 114732 269619 114766 269623
rect 114732 269547 114766 269555
rect 114732 269475 114766 269487
rect 114732 269403 114766 269419
rect 114732 269331 114766 269351
rect 114732 269259 114766 269283
rect 114732 269187 114766 269215
rect 114732 269120 114766 269147
rect 114914 270201 114948 270228
rect 114914 270133 114948 270161
rect 114914 270065 114948 270089
rect 114914 269997 114948 270017
rect 114914 269929 114948 269945
rect 114914 269861 114948 269873
rect 114914 269793 114948 269801
rect 114914 269725 114948 269729
rect 114914 269619 114948 269623
rect 114914 269547 114948 269555
rect 114914 269475 114948 269487
rect 114914 269403 114948 269419
rect 114914 269331 114948 269351
rect 114914 269259 114948 269283
rect 114914 269187 114948 269215
rect 114914 269120 114948 269147
rect 115132 270201 115166 270228
rect 115132 270133 115166 270161
rect 115132 270065 115166 270089
rect 115132 269997 115166 270017
rect 115132 269929 115166 269945
rect 115132 269861 115166 269873
rect 115132 269793 115166 269801
rect 115132 269725 115166 269729
rect 115132 269619 115166 269623
rect 115132 269547 115166 269555
rect 115132 269475 115166 269487
rect 115132 269403 115166 269419
rect 115132 269331 115166 269351
rect 115132 269259 115166 269283
rect 115132 269187 115166 269215
rect 115132 269120 115166 269147
rect 115314 270201 115348 270228
rect 115314 270133 115348 270161
rect 115314 270065 115348 270089
rect 115314 269997 115348 270017
rect 115314 269929 115348 269945
rect 115314 269861 115348 269873
rect 115314 269793 115348 269801
rect 115314 269725 115348 269729
rect 115314 269619 115348 269623
rect 115314 269547 115348 269555
rect 115314 269475 115348 269487
rect 115314 269403 115348 269419
rect 115314 269331 115348 269351
rect 115314 269259 115348 269283
rect 115314 269187 115348 269215
rect 115314 269120 115348 269147
rect 115532 270201 115566 270228
rect 115532 270133 115566 270161
rect 115532 270065 115566 270089
rect 115532 269997 115566 270017
rect 115532 269929 115566 269945
rect 115532 269861 115566 269873
rect 115532 269793 115566 269801
rect 115532 269725 115566 269729
rect 115532 269619 115566 269623
rect 115532 269547 115566 269555
rect 115532 269475 115566 269487
rect 115532 269403 115566 269419
rect 115532 269331 115566 269351
rect 115532 269259 115566 269283
rect 115532 269187 115566 269215
rect 115532 269120 115566 269147
rect 115714 270201 115748 270228
rect 115714 270133 115748 270161
rect 115714 270065 115748 270089
rect 115714 269997 115748 270017
rect 115714 269929 115748 269945
rect 115714 269861 115748 269873
rect 115714 269793 115748 269801
rect 115714 269725 115748 269729
rect 115714 269619 115748 269623
rect 115714 269547 115748 269555
rect 115714 269475 115748 269487
rect 115714 269403 115748 269419
rect 115714 269331 115748 269351
rect 115714 269259 115748 269283
rect 115714 269187 115748 269215
rect 115714 269120 115748 269147
rect 115932 270201 115966 270228
rect 115932 270133 115966 270161
rect 115932 270065 115966 270089
rect 115932 269997 115966 270017
rect 115932 269929 115966 269945
rect 115932 269861 115966 269873
rect 115932 269793 115966 269801
rect 115932 269725 115966 269729
rect 115932 269619 115966 269623
rect 115932 269547 115966 269555
rect 115932 269475 115966 269487
rect 115932 269403 115966 269419
rect 115932 269331 115966 269351
rect 115932 269259 115966 269283
rect 115932 269187 115966 269215
rect 115932 269120 115966 269147
rect 116114 270201 116148 270228
rect 116114 270133 116148 270161
rect 116114 270065 116148 270089
rect 116114 269997 116148 270017
rect 116114 269929 116148 269945
rect 116114 269861 116148 269873
rect 116114 269793 116148 269801
rect 116114 269725 116148 269729
rect 116114 269619 116148 269623
rect 116114 269547 116148 269555
rect 116114 269475 116148 269487
rect 116114 269403 116148 269419
rect 116114 269331 116148 269351
rect 116114 269259 116148 269283
rect 116114 269187 116148 269215
rect 116114 269120 116148 269147
rect 116332 270201 116366 270228
rect 116332 270133 116366 270161
rect 116332 270065 116366 270089
rect 116332 269997 116366 270017
rect 116332 269929 116366 269945
rect 116332 269861 116366 269873
rect 116332 269793 116366 269801
rect 116332 269725 116366 269729
rect 116332 269619 116366 269623
rect 116332 269547 116366 269555
rect 116332 269475 116366 269487
rect 116332 269403 116366 269419
rect 116332 269331 116366 269351
rect 116332 269259 116366 269283
rect 116332 269187 116366 269215
rect 116332 269120 116366 269147
rect 116514 270201 116548 270228
rect 116514 270133 116548 270161
rect 116514 270065 116548 270089
rect 116514 269997 116548 270017
rect 116514 269929 116548 269945
rect 116514 269861 116548 269873
rect 116514 269793 116548 269801
rect 116514 269725 116548 269729
rect 116514 269619 116548 269623
rect 116514 269547 116548 269555
rect 116514 269475 116548 269487
rect 116514 269403 116548 269419
rect 116514 269331 116548 269351
rect 116514 269259 116548 269283
rect 116514 269187 116548 269215
rect 116514 269120 116548 269147
rect 116732 270201 116766 270228
rect 116732 270133 116766 270161
rect 116732 270065 116766 270089
rect 116732 269997 116766 270017
rect 116732 269929 116766 269945
rect 116732 269861 116766 269873
rect 116732 269793 116766 269801
rect 116732 269725 116766 269729
rect 116732 269619 116766 269623
rect 116732 269547 116766 269555
rect 116732 269475 116766 269487
rect 116732 269403 116766 269419
rect 116732 269331 116766 269351
rect 116732 269259 116766 269283
rect 116732 269187 116766 269215
rect 116732 269120 116766 269147
rect 116914 270201 116948 270228
rect 116914 270133 116948 270161
rect 116914 270065 116948 270089
rect 116914 269997 116948 270017
rect 116914 269929 116948 269945
rect 116914 269861 116948 269873
rect 116914 269793 116948 269801
rect 116914 269725 116948 269729
rect 116914 269619 116948 269623
rect 116914 269547 116948 269555
rect 116914 269475 116948 269487
rect 116914 269403 116948 269419
rect 116914 269331 116948 269351
rect 116914 269259 116948 269283
rect 116914 269187 116948 269215
rect 116914 269120 116948 269147
rect 117132 270201 117166 270228
rect 117132 270133 117166 270161
rect 117132 270065 117166 270089
rect 117132 269997 117166 270017
rect 117132 269929 117166 269945
rect 117132 269861 117166 269873
rect 117132 269793 117166 269801
rect 117132 269725 117166 269729
rect 117132 269619 117166 269623
rect 117132 269547 117166 269555
rect 117132 269475 117166 269487
rect 117132 269403 117166 269419
rect 117132 269331 117166 269351
rect 117132 269259 117166 269283
rect 117132 269187 117166 269215
rect 117132 269120 117166 269147
rect 117314 270201 117348 270228
rect 117314 270133 117348 270161
rect 117314 270065 117348 270089
rect 117314 269997 117348 270017
rect 117314 269929 117348 269945
rect 117314 269861 117348 269873
rect 117314 269793 117348 269801
rect 117314 269725 117348 269729
rect 117314 269619 117348 269623
rect 117314 269547 117348 269555
rect 117314 269475 117348 269487
rect 117314 269403 117348 269419
rect 117314 269331 117348 269351
rect 117314 269259 117348 269283
rect 117314 269187 117348 269215
rect 117314 269120 117348 269147
rect 117532 270201 117566 270228
rect 117532 270133 117566 270161
rect 117532 270065 117566 270089
rect 117532 269997 117566 270017
rect 117532 269929 117566 269945
rect 117532 269861 117566 269873
rect 117532 269793 117566 269801
rect 117532 269725 117566 269729
rect 117532 269619 117566 269623
rect 117532 269547 117566 269555
rect 117532 269475 117566 269487
rect 117532 269403 117566 269419
rect 117532 269331 117566 269351
rect 117532 269259 117566 269283
rect 117532 269187 117566 269215
rect 117532 269120 117566 269147
rect 117714 270201 117748 270228
rect 117714 270133 117748 270161
rect 117714 270065 117748 270089
rect 117714 269997 117748 270017
rect 117714 269929 117748 269945
rect 117714 269861 117748 269873
rect 117714 269793 117748 269801
rect 117714 269725 117748 269729
rect 117714 269619 117748 269623
rect 117714 269547 117748 269555
rect 117714 269475 117748 269487
rect 117714 269403 117748 269419
rect 117714 269331 117748 269351
rect 117714 269259 117748 269283
rect 117714 269187 117748 269215
rect 117714 269120 117748 269147
rect 117932 270201 117966 270228
rect 117932 270133 117966 270161
rect 117932 270065 117966 270089
rect 117932 269997 117966 270017
rect 117932 269929 117966 269945
rect 117932 269861 117966 269873
rect 117932 269793 117966 269801
rect 117932 269725 117966 269729
rect 117932 269619 117966 269623
rect 117932 269547 117966 269555
rect 117932 269475 117966 269487
rect 117932 269403 117966 269419
rect 117932 269331 117966 269351
rect 117932 269259 117966 269283
rect 117932 269187 117966 269215
rect 117932 269120 117966 269147
rect 118114 270201 118148 270228
rect 118114 270133 118148 270161
rect 118114 270065 118148 270089
rect 118114 269997 118148 270017
rect 118114 269929 118148 269945
rect 118114 269861 118148 269873
rect 118114 269793 118148 269801
rect 118114 269725 118148 269729
rect 118114 269619 118148 269623
rect 118114 269547 118148 269555
rect 118114 269475 118148 269487
rect 118114 269403 118148 269419
rect 118114 269331 118148 269351
rect 118114 269259 118148 269283
rect 118114 269187 118148 269215
rect 118114 269120 118148 269147
rect 118332 270201 118366 270228
rect 118332 270133 118366 270161
rect 118332 270065 118366 270089
rect 118332 269997 118366 270017
rect 118332 269929 118366 269945
rect 118332 269861 118366 269873
rect 118332 269793 118366 269801
rect 118332 269725 118366 269729
rect 118332 269619 118366 269623
rect 118332 269547 118366 269555
rect 118332 269475 118366 269487
rect 118332 269403 118366 269419
rect 118332 269331 118366 269351
rect 118332 269259 118366 269283
rect 118332 269187 118366 269215
rect 118332 269120 118366 269147
rect 118514 270201 118548 270228
rect 118514 270133 118548 270161
rect 118514 270065 118548 270089
rect 118514 269997 118548 270017
rect 118514 269929 118548 269945
rect 118514 269861 118548 269873
rect 118514 269793 118548 269801
rect 118514 269725 118548 269729
rect 118514 269619 118548 269623
rect 118514 269547 118548 269555
rect 118514 269475 118548 269487
rect 118514 269403 118548 269419
rect 118514 269331 118548 269351
rect 118514 269259 118548 269283
rect 118514 269187 118548 269215
rect 118514 269120 118548 269147
rect 118732 270201 118766 270228
rect 118732 270133 118766 270161
rect 118732 270065 118766 270089
rect 118732 269997 118766 270017
rect 118732 269929 118766 269945
rect 118732 269861 118766 269873
rect 118732 269793 118766 269801
rect 118732 269725 118766 269729
rect 118732 269619 118766 269623
rect 118732 269547 118766 269555
rect 118732 269475 118766 269487
rect 118732 269403 118766 269419
rect 118732 269331 118766 269351
rect 118732 269259 118766 269283
rect 118732 269187 118766 269215
rect 118732 269120 118766 269147
rect 112560 269052 112587 269086
rect 112623 269052 112657 269086
rect 112693 269052 112987 269086
rect 113023 269052 113057 269086
rect 113093 269052 113387 269086
rect 113423 269052 113457 269086
rect 113493 269052 113787 269086
rect 113823 269052 113857 269086
rect 113893 269052 114187 269086
rect 114223 269052 114257 269086
rect 114293 269052 114587 269086
rect 114623 269052 114657 269086
rect 114693 269052 114987 269086
rect 115023 269052 115057 269086
rect 115093 269052 115387 269086
rect 115423 269052 115457 269086
rect 115493 269052 115787 269086
rect 115823 269052 115857 269086
rect 115893 269052 116187 269086
rect 116223 269052 116257 269086
rect 116293 269052 116587 269086
rect 116623 269052 116657 269086
rect 116693 269052 116987 269086
rect 117023 269052 117057 269086
rect 117093 269052 117387 269086
rect 117423 269052 117457 269086
rect 117493 269052 117787 269086
rect 117823 269052 117857 269086
rect 117893 269052 118187 269086
rect 118223 269052 118257 269086
rect 118293 269052 118587 269086
rect 118623 269052 118657 269086
rect 118693 269055 118720 269086
rect 118882 269055 118934 270288
rect 118693 269052 118934 269055
rect 118416 269017 118934 269052
rect 114230 268868 117626 268907
rect 114230 268826 114345 268868
rect 112055 268815 114345 268826
rect 117475 268826 117626 268868
rect 119021 268826 119035 272125
rect 117475 268815 119035 268826
rect 112055 268713 112171 268815
rect 118937 268713 119035 268815
rect 112055 268677 119035 268713
rect 119137 272179 119158 272247
rect 119137 268677 119151 272179
rect 119938 268785 119970 281059
rect 120072 281037 120256 281059
rect 125118 281037 125658 281139
rect 120072 281012 125658 281037
rect 120072 268861 120104 281012
rect 125047 280856 125658 281012
rect 120237 280779 120319 280813
rect 120353 280779 120387 280813
rect 120421 280779 120455 280813
rect 120489 280779 120523 280813
rect 120557 280779 120591 280813
rect 120625 280779 120659 280813
rect 120693 280779 120727 280813
rect 120761 280779 120795 280813
rect 120829 280779 120863 280813
rect 120897 280779 120931 280813
rect 120965 280779 120999 280813
rect 121033 280779 121067 280813
rect 121101 280779 121135 280813
rect 121169 280779 121203 280813
rect 121237 280779 121271 280813
rect 121305 280779 121339 280813
rect 121373 280779 121407 280813
rect 121441 280779 121475 280813
rect 121509 280779 121543 280813
rect 121577 280779 121611 280813
rect 121645 280800 121728 280813
rect 121645 280779 121960 280800
rect 120237 280726 121960 280779
rect 120271 280718 121694 280726
rect 120271 280692 120468 280718
rect 120237 280684 120468 280692
rect 120510 280684 120540 280718
rect 120578 280684 120612 280718
rect 120646 280684 120680 280718
rect 120718 280684 120748 280718
rect 120790 280713 121168 280718
rect 120790 280684 120875 280713
rect 120237 280658 120429 280684
rect 120271 280641 120429 280658
rect 120829 280641 120875 280684
rect 120271 280624 120417 280641
rect 120237 280604 120417 280624
rect 120237 280590 120383 280604
rect 120271 280570 120383 280590
rect 120271 280556 120417 280570
rect 120237 280533 120417 280556
rect 120841 280604 120875 280641
rect 120841 280533 120875 280570
rect 121083 280684 121168 280713
rect 121210 280684 121240 280718
rect 121278 280684 121312 280718
rect 121346 280684 121380 280718
rect 121418 280684 121448 280718
rect 121490 280692 121694 280718
rect 121728 280692 121960 280726
rect 121490 280684 121960 280692
rect 121083 280641 121129 280684
rect 121529 280658 121960 280684
rect 121529 280641 121694 280658
rect 121083 280604 121117 280641
rect 121083 280533 121117 280570
rect 121541 280624 121694 280641
rect 121728 280624 121960 280658
rect 121541 280604 121960 280624
rect 121575 280590 121960 280604
rect 121575 280570 121694 280590
rect 121541 280556 121694 280570
rect 121728 280556 121960 280590
rect 121541 280545 121960 280556
rect 121541 280533 121575 280545
rect 120237 280522 120395 280533
rect 120271 280488 120395 280522
rect 121694 280522 121960 280545
rect 120237 280454 120395 280488
rect 120429 280456 120468 280490
rect 120510 280456 120540 280490
rect 120578 280456 120612 280490
rect 120646 280456 120680 280490
rect 120718 280456 120748 280490
rect 120790 280456 120829 280490
rect 121129 280456 121168 280490
rect 121210 280456 121240 280490
rect 121278 280456 121312 280490
rect 121346 280456 121380 280490
rect 121418 280456 121448 280490
rect 121490 280456 121529 280490
rect 121728 280488 121960 280522
rect 120271 280420 120395 280454
rect 120237 280386 120395 280420
rect 120271 280352 120395 280386
rect 120237 280318 120395 280352
rect 121694 280454 121960 280488
rect 121728 280420 121960 280454
rect 121694 280386 121960 280420
rect 121728 280352 121960 280386
rect 120271 280284 120395 280318
rect 120429 280300 120468 280334
rect 120510 280300 120540 280334
rect 120578 280300 120612 280334
rect 120646 280300 120680 280334
rect 120718 280300 120748 280334
rect 120790 280300 120829 280334
rect 121129 280300 121168 280334
rect 121210 280300 121240 280334
rect 121278 280300 121312 280334
rect 121346 280300 121380 280334
rect 121418 280300 121448 280334
rect 121490 280300 121529 280334
rect 121694 280318 121960 280352
rect 120237 280257 120395 280284
rect 121728 280284 121960 280318
rect 120237 280250 120417 280257
rect 120271 280236 120417 280250
rect 120271 280216 120383 280236
rect 120237 280190 120383 280216
rect 120237 280182 120417 280190
rect 120271 280164 120417 280182
rect 120271 280148 120383 280164
rect 120237 280122 120383 280148
rect 120237 280114 120417 280122
rect 120271 280092 120417 280114
rect 120271 280080 120383 280092
rect 120237 280054 120383 280080
rect 120237 280046 120417 280054
rect 120271 280020 120417 280046
rect 120271 280012 120383 280020
rect 120237 279986 120383 280012
rect 120237 279978 120417 279986
rect 120271 279952 120417 279978
rect 120271 279944 120383 279952
rect 120237 279914 120383 279944
rect 120237 279910 120417 279914
rect 120271 279884 120417 279910
rect 120271 279876 120383 279884
rect 120237 279842 120383 279876
rect 120271 279816 120417 279842
rect 120271 279808 120383 279816
rect 120237 279774 120383 279808
rect 120271 279770 120383 279774
rect 120271 279749 120417 279770
rect 120841 280236 120875 280257
rect 120841 280164 120875 280190
rect 120841 280092 120875 280122
rect 120841 280020 120875 280054
rect 120841 279952 120875 279986
rect 120841 279884 120875 279914
rect 120841 279816 120875 279842
rect 120841 279749 120875 279770
rect 121083 280236 121117 280257
rect 121083 280164 121117 280190
rect 121083 280092 121117 280122
rect 121083 280020 121117 280054
rect 121083 279952 121117 279986
rect 121083 279884 121117 279914
rect 121083 279816 121117 279842
rect 121083 279749 121117 279770
rect 121541 280236 121575 280257
rect 121541 280164 121575 280190
rect 121541 280092 121575 280122
rect 121541 280020 121575 280054
rect 121541 279952 121575 279986
rect 121541 279884 121575 279914
rect 121541 279816 121575 279842
rect 121541 279749 121575 279770
rect 121694 280250 121960 280284
rect 121728 280216 121960 280250
rect 121694 280182 121960 280216
rect 121728 280148 121960 280182
rect 121694 280114 121960 280148
rect 121728 280080 121960 280114
rect 121694 280046 121960 280080
rect 121728 280012 121960 280046
rect 121694 279988 121960 280012
rect 122178 280574 122245 280608
rect 122279 280574 122313 280608
rect 122347 280574 122381 280608
rect 122415 280574 122449 280608
rect 122483 280574 122517 280608
rect 122551 280574 122585 280608
rect 122619 280574 122653 280608
rect 122687 280574 122721 280608
rect 122755 280574 122789 280608
rect 122823 280574 122857 280608
rect 122891 280574 122925 280608
rect 122959 280574 122993 280608
rect 123027 280574 123061 280608
rect 123095 280574 123129 280608
rect 123163 280574 123197 280608
rect 123231 280574 123265 280608
rect 123299 280574 123333 280608
rect 123367 280574 123401 280608
rect 123435 280574 123469 280608
rect 123503 280574 123537 280608
rect 123571 280574 123638 280608
rect 122178 280518 122212 280574
rect 123604 280518 123638 280574
rect 122178 280450 122212 280484
rect 122356 280470 122395 280504
rect 122437 280470 122467 280504
rect 122505 280470 122539 280504
rect 122573 280470 122607 280504
rect 122645 280470 122675 280504
rect 122717 280470 122756 280504
rect 123056 280470 123095 280504
rect 123137 280470 123167 280504
rect 123205 280470 123239 280504
rect 123273 280470 123307 280504
rect 123345 280470 123375 280504
rect 123417 280470 123456 280504
rect 123604 280450 123638 280484
rect 122212 280416 122344 280427
rect 122178 280406 122344 280416
rect 122178 280382 122310 280406
rect 122212 280360 122310 280382
rect 122212 280348 122344 280360
rect 122178 280334 122344 280348
rect 122178 280314 122310 280334
rect 122212 280292 122310 280314
rect 122212 280280 122344 280292
rect 122178 280262 122344 280280
rect 122178 280246 122310 280262
rect 122212 280224 122310 280246
rect 122212 280212 122344 280224
rect 122178 280190 122344 280212
rect 122178 280178 122310 280190
rect 122212 280156 122310 280178
rect 122212 280144 122344 280156
rect 122178 280122 122344 280144
rect 122178 280110 122310 280122
rect 122212 280084 122310 280110
rect 122212 280076 122344 280084
rect 122178 280054 122344 280076
rect 122178 280042 122310 280054
rect 122212 280012 122310 280042
rect 122212 280008 122344 280012
rect 122178 279988 122344 280008
rect 121694 279986 122344 279988
rect 121694 279978 122310 279986
rect 121728 279974 122310 279978
rect 121728 279944 122178 279974
rect 121694 279940 122178 279944
rect 122212 279940 122310 279974
rect 121694 279919 122344 279940
rect 122768 280406 122802 280427
rect 122768 280334 122802 280360
rect 122768 280262 122802 280292
rect 122768 280190 122802 280224
rect 122768 280122 122802 280156
rect 122768 280054 122802 280084
rect 122768 279986 122802 280012
rect 122768 279919 122802 279940
rect 123010 280406 123044 280427
rect 123010 280334 123044 280360
rect 123010 280262 123044 280292
rect 123010 280190 123044 280224
rect 123010 280122 123044 280156
rect 123010 280054 123044 280084
rect 123010 279986 123044 280012
rect 123010 279919 123044 279940
rect 123468 280406 123502 280427
rect 123468 280334 123502 280360
rect 123468 280262 123502 280292
rect 123468 280190 123502 280224
rect 123468 280122 123502 280156
rect 123468 280054 123502 280084
rect 123468 279986 123502 280012
rect 123468 279919 123502 279940
rect 123604 280382 123638 280416
rect 123604 280314 123638 280348
rect 123604 280246 123638 280280
rect 123604 280178 123638 280212
rect 123604 280110 123638 280144
rect 123604 280042 123638 280076
rect 123604 279974 123638 280008
rect 121694 279910 122310 279919
rect 121728 279906 122310 279910
rect 121728 279886 122178 279906
rect 121728 279876 121859 279886
rect 121694 279842 121859 279876
rect 122212 279872 122310 279906
rect 123604 279906 123638 279940
rect 121728 279808 121859 279842
rect 122181 279838 122310 279872
rect 122356 279842 122395 279876
rect 122437 279842 122467 279876
rect 122505 279842 122539 279876
rect 122573 279842 122607 279876
rect 122645 279842 122675 279876
rect 122717 279842 122756 279876
rect 123056 279842 123095 279876
rect 123137 279842 123167 279876
rect 123205 279842 123239 279876
rect 123273 279842 123307 279876
rect 123345 279842 123375 279876
rect 123417 279842 123456 279876
rect 121694 279774 121859 279808
rect 122212 279804 122310 279838
rect 120271 279740 120395 279749
rect 120237 279706 120395 279740
rect 121728 279740 121859 279774
rect 122181 279770 122310 279804
rect 121694 279706 121859 279740
rect 122212 279736 122310 279770
rect 120271 279672 120395 279706
rect 120429 279672 120468 279706
rect 120510 279672 120540 279706
rect 120578 279672 120612 279706
rect 120646 279672 120680 279706
rect 120718 279672 120748 279706
rect 120790 279672 120829 279706
rect 121129 279672 121168 279706
rect 121210 279672 121240 279706
rect 121278 279672 121312 279706
rect 121346 279672 121380 279706
rect 121418 279672 121448 279706
rect 121490 279672 121529 279706
rect 121728 279672 121859 279706
rect 122181 279702 122310 279736
rect 123604 279838 123638 279872
rect 123604 279770 123638 279804
rect 120237 279638 120395 279672
rect 120271 279604 120395 279638
rect 120237 279570 120395 279604
rect 120271 279536 120395 279570
rect 121694 279638 121859 279672
rect 122212 279668 122310 279702
rect 122356 279686 122395 279720
rect 122437 279686 122467 279720
rect 122505 279686 122539 279720
rect 122573 279686 122607 279720
rect 122645 279686 122675 279720
rect 122717 279686 122756 279720
rect 123056 279686 123095 279720
rect 123137 279686 123167 279720
rect 123205 279686 123239 279720
rect 123273 279686 123307 279720
rect 123345 279686 123375 279720
rect 123417 279686 123456 279720
rect 123604 279702 123638 279736
rect 121728 279604 121859 279638
rect 122181 279643 122310 279668
rect 122181 279634 122344 279643
rect 121694 279570 121859 279604
rect 122212 279622 122344 279634
rect 122212 279600 122310 279622
rect 120237 279502 120395 279536
rect 120429 279516 120468 279550
rect 120510 279516 120540 279550
rect 120578 279516 120612 279550
rect 120646 279516 120680 279550
rect 120718 279516 120748 279550
rect 120790 279516 120829 279550
rect 121129 279516 121168 279550
rect 121210 279516 121240 279550
rect 121278 279516 121312 279550
rect 121346 279516 121380 279550
rect 121418 279516 121448 279550
rect 121490 279516 121529 279550
rect 121728 279536 121859 279570
rect 122181 279576 122310 279600
rect 122181 279566 122344 279576
rect 120271 279473 120395 279502
rect 121694 279502 121859 279536
rect 122212 279550 122344 279566
rect 122212 279532 122310 279550
rect 120271 279468 120417 279473
rect 120237 279452 120417 279468
rect 120237 279434 120383 279452
rect 120271 279406 120383 279434
rect 120271 279400 120417 279406
rect 120237 279380 120417 279400
rect 120237 279366 120383 279380
rect 120271 279338 120383 279366
rect 120271 279332 120417 279338
rect 120237 279308 120417 279332
rect 120237 279298 120383 279308
rect 120271 279270 120383 279298
rect 120271 279264 120417 279270
rect 120237 279236 120417 279264
rect 120237 279230 120383 279236
rect 120271 279202 120383 279230
rect 120271 279196 120417 279202
rect 120237 279168 120417 279196
rect 120237 279162 120383 279168
rect 120271 279130 120383 279162
rect 120271 279128 120417 279130
rect 120237 279100 120417 279128
rect 120237 279094 120383 279100
rect 120271 279060 120383 279094
rect 120237 279058 120383 279060
rect 120237 279032 120417 279058
rect 120237 279026 120383 279032
rect 120271 278992 120383 279026
rect 120237 278986 120383 278992
rect 120237 278965 120417 278986
rect 120841 279452 120875 279473
rect 120841 279380 120875 279406
rect 120841 279308 120875 279338
rect 120841 279236 120875 279270
rect 120841 279168 120875 279202
rect 120841 279100 120875 279130
rect 120841 279032 120875 279058
rect 120841 278965 120875 278986
rect 121083 279452 121117 279473
rect 121083 279380 121117 279406
rect 121083 279308 121117 279338
rect 121083 279236 121117 279270
rect 121083 279168 121117 279202
rect 121083 279100 121117 279130
rect 121083 279032 121117 279058
rect 121083 278965 121117 278986
rect 121541 279452 121575 279473
rect 121541 279380 121575 279406
rect 121541 279308 121575 279338
rect 121541 279236 121575 279270
rect 121541 279168 121575 279202
rect 121541 279100 121575 279130
rect 121541 279032 121575 279058
rect 121541 278965 121575 278986
rect 121728 279468 121859 279502
rect 122181 279508 122310 279532
rect 122181 279498 122344 279508
rect 121694 279434 121859 279468
rect 122212 279478 122344 279498
rect 122212 279464 122310 279478
rect 121728 279400 121859 279434
rect 122181 279440 122310 279464
rect 122181 279430 122344 279440
rect 121694 279366 121859 279400
rect 122212 279406 122344 279430
rect 122212 279396 122310 279406
rect 121728 279332 121859 279366
rect 122181 279372 122310 279396
rect 122181 279362 122344 279372
rect 121694 279298 121859 279332
rect 122212 279338 122344 279362
rect 122212 279328 122310 279338
rect 121728 279276 121859 279298
rect 122181 279300 122310 279328
rect 122181 279294 122344 279300
rect 121728 279264 122178 279276
rect 121694 279260 122178 279264
rect 122212 279270 122344 279294
rect 122212 279260 122310 279270
rect 121694 279230 122310 279260
rect 121728 279228 122310 279230
rect 121728 279226 122344 279228
rect 121728 279196 122178 279226
rect 121694 279192 122178 279196
rect 122212 279202 122344 279226
rect 122212 279192 122310 279202
rect 121694 279162 122310 279192
rect 121728 279158 122310 279162
rect 121728 279128 122178 279158
rect 121694 279124 122178 279128
rect 122212 279156 122310 279158
rect 122212 279135 122344 279156
rect 122768 279622 122802 279643
rect 122768 279550 122802 279576
rect 122768 279478 122802 279508
rect 122768 279406 122802 279440
rect 122768 279338 122802 279372
rect 122768 279270 122802 279300
rect 122768 279202 122802 279228
rect 122768 279135 122802 279156
rect 123010 279622 123044 279643
rect 123010 279550 123044 279576
rect 123010 279478 123044 279508
rect 123010 279406 123044 279440
rect 123010 279338 123044 279372
rect 123010 279270 123044 279300
rect 123010 279202 123044 279228
rect 123010 279135 123044 279156
rect 123468 279622 123502 279643
rect 123468 279550 123502 279576
rect 123468 279478 123502 279508
rect 123468 279406 123502 279440
rect 123468 279338 123502 279372
rect 123468 279270 123502 279300
rect 123468 279202 123502 279228
rect 123468 279135 123502 279156
rect 123604 279634 123638 279668
rect 123604 279566 123638 279600
rect 123604 279498 123638 279532
rect 123604 279430 123638 279464
rect 123604 279362 123638 279396
rect 123604 279294 123638 279328
rect 123604 279226 123638 279260
rect 123604 279158 123638 279192
rect 121694 279094 122212 279124
rect 121728 279090 122212 279094
rect 121728 279060 122178 279090
rect 121694 279056 122178 279060
rect 122356 279058 122395 279092
rect 122437 279058 122467 279092
rect 122505 279058 122539 279092
rect 122573 279058 122607 279092
rect 122645 279058 122675 279092
rect 122717 279058 122756 279092
rect 123056 279058 123095 279092
rect 123137 279058 123167 279092
rect 123205 279058 123239 279092
rect 123273 279058 123307 279092
rect 123345 279058 123375 279092
rect 123417 279058 123456 279092
rect 123604 279090 123638 279124
rect 121694 279026 122212 279056
rect 121728 279000 122212 279026
rect 123604 279000 123638 279056
rect 121728 278992 122245 279000
rect 121694 278966 122245 278992
rect 122279 278966 122313 279000
rect 122347 278966 122381 279000
rect 122415 278966 122449 279000
rect 122483 278966 122517 279000
rect 122551 278966 122585 279000
rect 122619 278966 122653 279000
rect 122687 278966 122721 279000
rect 122755 278966 122789 279000
rect 122823 278966 122857 279000
rect 122891 278966 122925 279000
rect 122959 278966 122993 279000
rect 123027 278966 123061 279000
rect 123095 278966 123129 279000
rect 123163 278966 123197 279000
rect 123231 278966 123265 279000
rect 123299 278966 123333 279000
rect 123367 278966 123401 279000
rect 123435 278966 123469 279000
rect 123503 278966 123537 279000
rect 123571 278966 123638 279000
rect 120237 278958 120395 278965
rect 120271 278924 120395 278958
rect 120237 278890 120395 278924
rect 121694 278958 123358 278966
rect 121728 278924 123358 278958
rect 120271 278856 120395 278890
rect 120429 278888 120468 278922
rect 120510 278888 120540 278922
rect 120578 278888 120612 278922
rect 120646 278888 120680 278922
rect 120718 278888 120748 278922
rect 120790 278888 120829 278922
rect 121129 278888 121168 278922
rect 121210 278888 121240 278922
rect 121278 278888 121312 278922
rect 121346 278888 121380 278922
rect 121418 278888 121448 278922
rect 121490 278888 121529 278922
rect 121694 278890 123358 278924
rect 120237 278822 120395 278856
rect 120271 278788 120395 278822
rect 120237 278754 120395 278788
rect 121728 278870 123358 278890
rect 121728 278856 121809 278870
rect 121694 278822 121809 278856
rect 121728 278788 121809 278822
rect 120271 278720 120395 278754
rect 120429 278732 120468 278766
rect 120510 278732 120540 278766
rect 120578 278732 120612 278766
rect 120646 278732 120680 278766
rect 120718 278732 120748 278766
rect 120790 278732 120829 278766
rect 121129 278732 121168 278766
rect 121210 278732 121240 278766
rect 121278 278732 121312 278766
rect 121346 278732 121380 278766
rect 121418 278732 121448 278766
rect 121490 278732 121529 278766
rect 121694 278754 121809 278788
rect 120237 278689 120395 278720
rect 121728 278720 121809 278754
rect 120237 278686 120417 278689
rect 120271 278668 120417 278686
rect 120271 278652 120383 278668
rect 120237 278622 120383 278652
rect 120237 278618 120417 278622
rect 120271 278596 120417 278618
rect 120271 278584 120383 278596
rect 120237 278554 120383 278584
rect 120237 278550 120417 278554
rect 120271 278524 120417 278550
rect 120271 278516 120383 278524
rect 120237 278486 120383 278516
rect 120237 278482 120417 278486
rect 120271 278452 120417 278482
rect 120271 278448 120383 278452
rect 120237 278418 120383 278448
rect 120237 278414 120417 278418
rect 120271 278384 120417 278414
rect 120271 278380 120383 278384
rect 120237 278346 120383 278380
rect 120271 278316 120417 278346
rect 120271 278312 120383 278316
rect 120237 278278 120383 278312
rect 120271 278274 120383 278278
rect 120271 278248 120417 278274
rect 120271 278244 120383 278248
rect 120237 278210 120383 278244
rect 120271 278202 120383 278210
rect 120271 278181 120417 278202
rect 120841 278668 120875 278689
rect 120841 278596 120875 278622
rect 120841 278524 120875 278554
rect 120841 278452 120875 278486
rect 120841 278384 120875 278418
rect 120841 278316 120875 278346
rect 120841 278248 120875 278274
rect 120841 278181 120875 278202
rect 121083 278668 121117 278689
rect 121083 278596 121117 278622
rect 121083 278524 121117 278554
rect 121083 278452 121117 278486
rect 121083 278384 121117 278418
rect 121083 278316 121117 278346
rect 121083 278248 121117 278274
rect 121083 278181 121117 278202
rect 121541 278668 121575 278689
rect 121541 278596 121575 278622
rect 121541 278524 121575 278554
rect 121541 278452 121575 278486
rect 121541 278384 121575 278418
rect 121541 278316 121575 278346
rect 121541 278248 121575 278274
rect 121541 278181 121575 278202
rect 121694 278686 121809 278720
rect 121728 278652 121809 278686
rect 121694 278618 121809 278652
rect 121728 278584 121809 278618
rect 121694 278550 121809 278584
rect 121728 278516 121809 278550
rect 121694 278482 121809 278516
rect 121728 278448 121809 278482
rect 121694 278414 121809 278448
rect 121728 278380 121809 278414
rect 121694 278346 121809 278380
rect 121728 278312 121809 278346
rect 121694 278278 121809 278312
rect 121728 278244 121809 278278
rect 121694 278210 121809 278244
rect 120271 278176 120395 278181
rect 120237 278142 120395 278176
rect 120271 278108 120395 278142
rect 121728 278176 121809 278210
rect 121694 278142 121809 278176
rect 120237 278074 120395 278108
rect 120429 278104 120468 278138
rect 120510 278104 120540 278138
rect 120578 278104 120612 278138
rect 120646 278104 120680 278138
rect 120718 278104 120748 278138
rect 120790 278104 120829 278138
rect 121129 278104 121168 278138
rect 121210 278104 121240 278138
rect 121278 278104 121312 278138
rect 121346 278104 121380 278138
rect 121418 278104 121448 278138
rect 121490 278104 121529 278138
rect 121728 278108 121809 278142
rect 120271 278040 120395 278074
rect 120237 278006 120395 278040
rect 120271 277972 120395 278006
rect 121694 278074 121809 278108
rect 121728 278040 121809 278074
rect 121694 278006 121809 278040
rect 120237 277938 120395 277972
rect 120429 277948 120468 277982
rect 120510 277948 120540 277982
rect 120578 277948 120612 277982
rect 120646 277948 120680 277982
rect 120718 277948 120748 277982
rect 120790 277948 120829 277982
rect 121129 277948 121168 277982
rect 121210 277948 121240 277982
rect 121278 277948 121312 277982
rect 121346 277948 121380 277982
rect 121418 277948 121448 277982
rect 121490 277948 121529 277982
rect 121728 277972 121809 278006
rect 120271 277905 120395 277938
rect 121694 277938 121809 277972
rect 120271 277904 120417 277905
rect 120237 277884 120417 277904
rect 120237 277870 120383 277884
rect 120271 277838 120383 277870
rect 120271 277836 120417 277838
rect 120237 277812 120417 277836
rect 120237 277802 120383 277812
rect 120271 277770 120383 277802
rect 120271 277768 120417 277770
rect 120237 277740 120417 277768
rect 120237 277734 120383 277740
rect 120271 277702 120383 277734
rect 120271 277700 120417 277702
rect 120237 277668 120417 277700
rect 120237 277666 120383 277668
rect 120271 277634 120383 277666
rect 120271 277632 120417 277634
rect 120237 277600 120417 277632
rect 120237 277598 120383 277600
rect 120271 277564 120383 277598
rect 120237 277562 120383 277564
rect 120237 277532 120417 277562
rect 120237 277530 120383 277532
rect 120271 277496 120383 277530
rect 120237 277490 120383 277496
rect 120237 277464 120417 277490
rect 120237 277462 120383 277464
rect 120271 277428 120383 277462
rect 120237 277418 120383 277428
rect 120237 277397 120417 277418
rect 120841 277884 120875 277905
rect 120841 277812 120875 277838
rect 120841 277740 120875 277770
rect 120841 277668 120875 277702
rect 120841 277600 120875 277634
rect 120841 277532 120875 277562
rect 120841 277464 120875 277490
rect 120841 277397 120875 277418
rect 121083 277884 121117 277905
rect 121083 277812 121117 277838
rect 121083 277740 121117 277770
rect 121083 277668 121117 277702
rect 121083 277600 121117 277634
rect 121083 277532 121117 277562
rect 121083 277464 121117 277490
rect 121083 277397 121117 277418
rect 121541 277884 121575 277905
rect 121541 277812 121575 277838
rect 121541 277740 121575 277770
rect 121541 277668 121575 277702
rect 121541 277600 121575 277634
rect 121541 277532 121575 277562
rect 121541 277464 121575 277490
rect 121541 277397 121575 277418
rect 121728 277904 121809 277938
rect 121694 277870 121809 277904
rect 121728 277836 121809 277870
rect 121694 277802 121809 277836
rect 121728 277768 121809 277802
rect 121694 277734 121809 277768
rect 121728 277700 121809 277734
rect 121694 277666 121809 277700
rect 121728 277632 121809 277666
rect 121694 277598 121809 277632
rect 121728 277564 121809 277598
rect 121694 277530 121809 277564
rect 121728 277496 121809 277530
rect 121694 277462 121809 277496
rect 121728 277428 121809 277462
rect 120237 277394 120395 277397
rect 120271 277360 120395 277394
rect 120237 277326 120395 277360
rect 121694 277394 121809 277428
rect 121728 277360 121809 277394
rect 120271 277292 120395 277326
rect 120429 277320 120468 277354
rect 120510 277320 120540 277354
rect 120578 277320 120612 277354
rect 120646 277320 120680 277354
rect 120718 277320 120748 277354
rect 120790 277320 120829 277354
rect 121129 277320 121168 277354
rect 121210 277320 121240 277354
rect 121278 277320 121312 277354
rect 121346 277320 121380 277354
rect 121418 277320 121448 277354
rect 121490 277320 121529 277354
rect 121694 277326 121809 277360
rect 120237 277258 120395 277292
rect 120271 277224 120395 277258
rect 120237 277190 120395 277224
rect 121728 277292 121809 277326
rect 121694 277258 121809 277292
rect 121728 277224 121809 277258
rect 120271 277156 120395 277190
rect 120429 277164 120468 277198
rect 120510 277164 120540 277198
rect 120578 277164 120612 277198
rect 120646 277164 120680 277198
rect 120718 277164 120748 277198
rect 120790 277164 120829 277198
rect 121129 277164 121168 277198
rect 121210 277164 121240 277198
rect 121278 277164 121312 277198
rect 121346 277164 121380 277198
rect 121418 277164 121448 277198
rect 121490 277164 121529 277198
rect 121694 277190 121809 277224
rect 120237 277122 120395 277156
rect 120271 277121 120395 277122
rect 121728 277156 121809 277190
rect 121694 277122 121809 277156
rect 120271 277100 120417 277121
rect 120271 277088 120383 277100
rect 120237 277054 120383 277088
rect 120271 277028 120417 277054
rect 120271 277020 120383 277028
rect 120237 276986 120383 277020
rect 120271 276956 120417 276986
rect 120271 276952 120383 276956
rect 120237 276918 120383 276952
rect 120271 276884 120417 276918
rect 120237 276850 120383 276884
rect 120271 276816 120417 276850
rect 120237 276782 120383 276816
rect 120271 276778 120383 276782
rect 120271 276748 120417 276778
rect 120237 276714 120383 276748
rect 120271 276706 120383 276714
rect 120271 276680 120417 276706
rect 120237 276646 120383 276680
rect 120271 276634 120383 276646
rect 120271 276613 120417 276634
rect 120841 277100 120875 277121
rect 120841 277028 120875 277054
rect 120841 276956 120875 276986
rect 120841 276884 120875 276918
rect 120841 276816 120875 276850
rect 120841 276748 120875 276778
rect 120841 276680 120875 276706
rect 120841 276613 120875 276634
rect 121083 277100 121117 277121
rect 121083 277028 121117 277054
rect 121083 276956 121117 276986
rect 121083 276884 121117 276918
rect 121083 276816 121117 276850
rect 121083 276748 121117 276778
rect 121083 276680 121117 276706
rect 121083 276613 121117 276634
rect 121541 277100 121575 277121
rect 121541 277028 121575 277054
rect 121541 276956 121575 276986
rect 121541 276884 121575 276918
rect 121541 276816 121575 276850
rect 121541 276748 121575 276778
rect 121541 276680 121575 276706
rect 121541 276613 121575 276634
rect 121728 277088 121809 277122
rect 121694 277054 121809 277088
rect 121728 277020 121809 277054
rect 121694 276986 121809 277020
rect 121728 276952 121809 276986
rect 121694 276918 121809 276952
rect 121728 276884 121809 276918
rect 121694 276850 121809 276884
rect 121728 276816 121809 276850
rect 121694 276782 121809 276816
rect 121728 276748 121809 276782
rect 121694 276714 121809 276748
rect 121728 276680 121809 276714
rect 121694 276646 121809 276680
rect 120271 276612 120395 276613
rect 120237 276578 120395 276612
rect 120271 276544 120395 276578
rect 121728 276612 121809 276646
rect 121694 276578 121809 276612
rect 120237 276510 120395 276544
rect 120429 276536 120468 276570
rect 120510 276536 120540 276570
rect 120578 276536 120612 276570
rect 120646 276536 120680 276570
rect 120718 276536 120748 276570
rect 120790 276536 120829 276570
rect 121129 276536 121168 276570
rect 121210 276536 121240 276570
rect 121278 276536 121312 276570
rect 121346 276536 121380 276570
rect 121418 276536 121448 276570
rect 121490 276536 121529 276570
rect 121728 276544 121809 276578
rect 120271 276476 120395 276510
rect 120237 276442 120395 276476
rect 120271 276408 120395 276442
rect 121694 276510 121809 276544
rect 121728 276476 121809 276510
rect 121694 276442 121809 276476
rect 120237 276374 120395 276408
rect 120429 276380 120468 276414
rect 120510 276380 120540 276414
rect 120578 276380 120612 276414
rect 120646 276380 120680 276414
rect 120718 276380 120748 276414
rect 120790 276380 120829 276414
rect 121129 276380 121168 276414
rect 121210 276380 121240 276414
rect 121278 276380 121312 276414
rect 121346 276380 121380 276414
rect 121418 276380 121448 276414
rect 121490 276380 121529 276414
rect 121728 276408 121809 276442
rect 120271 276340 120395 276374
rect 120237 276337 120395 276340
rect 121694 276374 121809 276408
rect 121728 276340 121809 276374
rect 120237 276316 120417 276337
rect 120237 276306 120383 276316
rect 120271 276272 120383 276306
rect 120237 276270 120383 276272
rect 120237 276244 120417 276270
rect 120237 276238 120383 276244
rect 120271 276204 120383 276238
rect 120237 276202 120383 276204
rect 120237 276172 120417 276202
rect 120237 276170 120383 276172
rect 120271 276136 120383 276170
rect 120237 276134 120383 276136
rect 120237 276102 120417 276134
rect 120271 276100 120417 276102
rect 120271 276068 120383 276100
rect 120237 276066 120383 276068
rect 120237 276034 120417 276066
rect 120271 276032 120417 276034
rect 120271 276000 120383 276032
rect 120237 275994 120383 276000
rect 120237 275966 120417 275994
rect 120271 275964 120417 275966
rect 120271 275932 120383 275964
rect 120237 275922 120383 275932
rect 120237 275898 120417 275922
rect 120271 275896 120417 275898
rect 120271 275864 120383 275896
rect 120237 275850 120383 275864
rect 120237 275830 120417 275850
rect 120271 275829 120417 275830
rect 120841 276316 120875 276337
rect 120841 276244 120875 276270
rect 120841 276172 120875 276202
rect 121083 276316 121117 276337
rect 121083 276244 121117 276270
rect 121083 276172 121117 276202
rect 120875 276134 121083 276139
rect 120841 276103 121117 276134
rect 120841 276100 120969 276103
rect 120875 276069 120969 276100
rect 121003 276100 121117 276103
rect 121003 276069 121083 276100
rect 120875 276066 121083 276069
rect 120841 276032 121117 276066
rect 120841 275964 120875 275994
rect 120841 275896 120875 275922
rect 120841 275829 120875 275850
rect 121083 275964 121117 275994
rect 121083 275896 121117 275922
rect 121083 275829 121117 275850
rect 121541 276316 121575 276337
rect 121541 276244 121575 276270
rect 121541 276172 121575 276202
rect 121541 276100 121575 276134
rect 121541 276032 121575 276066
rect 121541 275964 121575 275994
rect 121541 275896 121575 275922
rect 121541 275829 121575 275850
rect 121694 276306 121809 276340
rect 121728 276272 121809 276306
rect 121694 276238 121809 276272
rect 121728 276204 121809 276238
rect 122027 278588 122144 278635
rect 122027 276225 122034 278588
rect 121694 276170 121809 276204
rect 121728 276136 121809 276170
rect 121694 276102 121809 276136
rect 121728 276068 121809 276102
rect 121694 276034 121809 276068
rect 122022 276038 122034 276225
rect 121728 276000 121809 276034
rect 121694 275966 121809 276000
rect 121728 275932 121809 275966
rect 121694 275898 121809 275932
rect 121728 275864 121809 275898
rect 121694 275830 121809 275864
rect 120271 275796 120395 275829
rect 120237 275762 120395 275796
rect 121728 275796 121809 275830
rect 120271 275728 120395 275762
rect 120429 275752 120468 275786
rect 120510 275752 120540 275786
rect 120578 275752 120612 275786
rect 120646 275752 120680 275786
rect 120718 275752 120748 275786
rect 120790 275752 120829 275786
rect 121129 275752 121168 275786
rect 121210 275752 121240 275786
rect 121278 275752 121312 275786
rect 121346 275752 121380 275786
rect 121418 275752 121448 275786
rect 121490 275752 121529 275786
rect 121694 275762 121809 275796
rect 120237 275694 120395 275728
rect 120271 275660 120395 275694
rect 120237 275626 120395 275660
rect 121728 275728 121809 275762
rect 121694 275694 121809 275728
rect 121728 275660 121809 275694
rect 120271 275592 120395 275626
rect 120429 275596 120468 275630
rect 120510 275596 120540 275630
rect 120578 275596 120612 275630
rect 120646 275596 120680 275630
rect 120718 275596 120748 275630
rect 120790 275596 120829 275630
rect 121129 275596 121168 275630
rect 121210 275596 121240 275630
rect 121278 275596 121312 275630
rect 121346 275596 121380 275630
rect 121418 275596 121448 275630
rect 121490 275596 121529 275630
rect 121694 275626 121809 275660
rect 120237 275558 120395 275592
rect 120271 275553 120395 275558
rect 121728 275592 121809 275626
rect 121694 275558 121809 275592
rect 120271 275532 120417 275553
rect 120271 275524 120383 275532
rect 120237 275490 120383 275524
rect 120271 275486 120383 275490
rect 120271 275460 120417 275486
rect 120271 275456 120383 275460
rect 120237 275422 120383 275456
rect 120271 275418 120383 275422
rect 120271 275388 120417 275418
rect 120237 275354 120383 275388
rect 120271 275350 120383 275354
rect 120271 275320 120417 275350
rect 120237 275316 120417 275320
rect 120237 275286 120383 275316
rect 120271 275282 120383 275286
rect 120271 275252 120417 275282
rect 120237 275248 120417 275252
rect 120237 275218 120383 275248
rect 120271 275210 120383 275218
rect 120271 275184 120417 275210
rect 120237 275180 120417 275184
rect 120237 275150 120383 275180
rect 120271 275138 120383 275150
rect 120271 275116 120417 275138
rect 120237 275112 120417 275116
rect 120237 275082 120383 275112
rect 120271 275066 120383 275082
rect 120271 275048 120417 275066
rect 120237 275045 120417 275048
rect 120841 275532 120875 275553
rect 120841 275460 120875 275486
rect 120841 275388 120875 275418
rect 121083 275532 121117 275553
rect 121083 275460 121117 275486
rect 121083 275388 121117 275418
rect 120875 275350 121083 275353
rect 120841 275316 121117 275350
rect 120875 275282 121083 275316
rect 120841 275248 121117 275282
rect 120875 275246 121083 275248
rect 120841 275180 120875 275210
rect 120841 275112 120875 275138
rect 120841 275045 120875 275066
rect 120237 275014 120395 275045
rect 120271 274980 120395 275014
rect 120237 274946 120395 274980
rect 120429 274968 120468 275002
rect 120510 274968 120540 275002
rect 120578 274968 120612 275002
rect 120646 274968 120680 275002
rect 120718 274968 120748 275002
rect 120790 274968 120829 275002
rect 120271 274912 120395 274946
rect 120237 274878 120395 274912
rect 120271 274844 120395 274878
rect 120237 274810 120395 274844
rect 120429 274812 120468 274846
rect 120510 274812 120540 274846
rect 120578 274812 120612 274846
rect 120646 274812 120680 274846
rect 120718 274812 120748 274846
rect 120790 274812 120829 274846
rect 120271 274776 120395 274810
rect 120237 274769 120395 274776
rect 120237 274748 120417 274769
rect 120237 274742 120383 274748
rect 120271 274708 120383 274742
rect 120237 274702 120383 274708
rect 120237 274676 120417 274702
rect 120237 274674 120383 274676
rect 120271 274640 120383 274674
rect 120237 274634 120383 274640
rect 120237 274606 120417 274634
rect 120271 274604 120417 274606
rect 120271 274572 120383 274604
rect 120237 274566 120383 274572
rect 120237 274538 120417 274566
rect 120271 274532 120417 274538
rect 120271 274504 120383 274532
rect 120237 274498 120383 274504
rect 120237 274470 120417 274498
rect 120271 274464 120417 274470
rect 120271 274436 120383 274464
rect 120237 274426 120383 274436
rect 120237 274402 120417 274426
rect 120271 274396 120417 274402
rect 120271 274368 120383 274396
rect 120237 274354 120383 274368
rect 120237 274334 120417 274354
rect 120271 274328 120417 274334
rect 120271 274300 120383 274328
rect 120237 274282 120383 274300
rect 120237 274266 120417 274282
rect 120271 274261 120417 274266
rect 120841 274748 120875 274769
rect 120841 274676 120875 274702
rect 120841 274604 120875 274634
rect 120943 274579 121039 275246
rect 121083 275180 121117 275210
rect 121083 275112 121117 275138
rect 121083 275045 121117 275066
rect 121541 275532 121575 275553
rect 121541 275460 121575 275486
rect 121541 275388 121575 275418
rect 121541 275316 121575 275350
rect 121541 275248 121575 275282
rect 121541 275180 121575 275210
rect 121541 275112 121575 275138
rect 121541 275045 121575 275066
rect 121728 275524 121809 275558
rect 121694 275490 121809 275524
rect 122027 275562 122034 276038
rect 122136 276225 122144 278588
rect 122260 278482 123358 278870
rect 122254 278448 122343 278482
rect 122377 278448 122411 278482
rect 122445 278448 122479 278482
rect 122513 278448 122547 278482
rect 122581 278448 122615 278482
rect 122649 278448 122683 278482
rect 122717 278448 122751 278482
rect 122785 278448 122819 278482
rect 122853 278448 122887 278482
rect 122921 278448 122955 278482
rect 122989 278448 123023 278482
rect 123057 278448 123091 278482
rect 123125 278448 123159 278482
rect 123193 278448 123227 278482
rect 123261 278448 123295 278482
rect 123329 278448 123363 278482
rect 123397 278448 123431 278482
rect 123465 278448 123499 278482
rect 123533 278448 123567 278482
rect 123601 278448 123635 278482
rect 123669 278448 123703 278482
rect 123737 278448 123771 278482
rect 123805 278448 123839 278482
rect 123873 278448 123907 278482
rect 123941 278448 123975 278482
rect 124009 278448 124043 278482
rect 124077 278448 124111 278482
rect 124145 278448 124179 278482
rect 124213 278448 124247 278482
rect 124281 278448 124370 278482
rect 122254 278395 122374 278448
rect 122288 278361 122374 278395
rect 122254 278327 122374 278361
rect 124336 278395 124370 278448
rect 122288 278293 122374 278327
rect 122414 278313 122439 278347
rect 122495 278313 122511 278347
rect 122563 278313 122583 278347
rect 122631 278313 122655 278347
rect 122699 278313 122727 278347
rect 122767 278313 122799 278347
rect 122835 278313 122869 278347
rect 122905 278313 122937 278347
rect 122977 278313 123005 278347
rect 123049 278313 123073 278347
rect 123121 278313 123141 278347
rect 123193 278313 123209 278347
rect 123265 278313 123290 278347
rect 124336 278327 124370 278361
rect 122254 278270 122374 278293
rect 122254 278259 122402 278270
rect 122288 278250 122402 278259
rect 122288 278225 122368 278250
rect 122254 278192 122368 278225
rect 122254 278191 122402 278192
rect 122288 278182 122402 278191
rect 122288 278157 122368 278182
rect 122254 278123 122368 278157
rect 122288 278120 122368 278123
rect 122288 278114 122402 278120
rect 122288 278089 122368 278114
rect 122254 278055 122368 278089
rect 122288 278048 122368 278055
rect 122288 278046 122402 278048
rect 122288 278021 122368 278046
rect 122254 278012 122368 278021
rect 122254 278010 122402 278012
rect 122254 277987 122368 278010
rect 122288 277953 122368 277987
rect 122254 277944 122368 277953
rect 122254 277938 122402 277944
rect 122254 277919 122368 277938
rect 122288 277885 122368 277919
rect 122254 277876 122368 277885
rect 122254 277866 122402 277876
rect 122254 277851 122368 277866
rect 122288 277817 122368 277851
rect 122254 277808 122368 277817
rect 122254 277788 122402 277808
rect 123302 278250 123336 278270
rect 124336 278259 124370 278293
rect 123336 278192 124210 278193
rect 123302 278182 124210 278192
rect 123336 278161 124210 278182
rect 123336 278154 123678 278161
rect 123302 278114 123336 278120
rect 123302 278046 123336 278048
rect 123302 278010 123336 278012
rect 123302 277938 123336 277944
rect 123302 277866 123336 277876
rect 123302 277788 123336 277808
rect 122254 277783 122374 277788
rect 122288 277749 122374 277783
rect 122254 277715 122374 277749
rect 122288 277681 122374 277715
rect 122414 277711 122439 277745
rect 122495 277711 122511 277745
rect 122563 277711 122583 277745
rect 122631 277711 122655 277745
rect 122699 277711 122727 277745
rect 122767 277711 122799 277745
rect 122835 277711 122869 277745
rect 122905 277711 122937 277745
rect 122977 277711 123005 277745
rect 123049 277711 123073 277745
rect 123121 277711 123141 277745
rect 123193 277711 123209 277745
rect 123265 277711 123290 277745
rect 122254 277647 122374 277681
rect 122288 277613 122374 277647
rect 122254 277579 122374 277613
rect 122288 277545 122374 277579
rect 122416 277547 122439 277581
rect 122493 277547 122511 277581
rect 122561 277547 122583 277581
rect 122629 277547 122655 277581
rect 122697 277547 122727 277581
rect 122765 277547 122799 277581
rect 122833 277547 122867 277581
rect 122905 277547 122935 277581
rect 122977 277547 123003 277581
rect 123049 277547 123071 277581
rect 123121 277547 123139 277581
rect 123193 277547 123216 277581
rect 122254 277511 122374 277545
rect 122288 277504 122374 277511
rect 122288 277477 122404 277504
rect 122254 277467 122404 277477
rect 122254 277443 122370 277467
rect 122288 277433 122370 277443
rect 122288 277409 122404 277433
rect 122254 277396 122404 277409
rect 123228 277467 123262 277504
rect 123228 277396 123262 277433
rect 122254 277375 122374 277396
rect 122288 277341 122374 277375
rect 122254 277307 122374 277341
rect 122416 277319 122439 277353
rect 122493 277319 122511 277353
rect 122561 277319 122583 277353
rect 122629 277319 122655 277353
rect 122697 277319 122727 277353
rect 122765 277319 122799 277353
rect 122833 277319 122867 277353
rect 122905 277319 122935 277353
rect 122977 277319 123003 277353
rect 123049 277319 123071 277353
rect 123121 277319 123139 277353
rect 123193 277319 123216 277353
rect 123494 277330 123535 278154
rect 123656 278127 123678 278154
rect 123734 278127 123746 278161
rect 123806 278127 123814 278161
rect 123878 278127 123882 278161
rect 123984 278127 123988 278161
rect 124052 278127 124060 278161
rect 124120 278127 124132 278161
rect 124188 278127 124210 278161
rect 124336 278191 124370 278225
rect 124336 278123 124370 278157
rect 123610 278060 123644 278084
rect 123610 277992 123644 278008
rect 123610 277924 123644 277936
rect 123610 277856 123644 277864
rect 123610 277788 123644 277792
rect 123610 277682 123644 277686
rect 123610 277610 123644 277618
rect 123610 277538 123644 277550
rect 123610 277466 123644 277482
rect 123610 277390 123644 277414
rect 124222 278060 124256 278084
rect 124222 277992 124256 278008
rect 124222 277924 124256 277936
rect 124222 277856 124256 277864
rect 124222 277788 124256 277792
rect 124222 277682 124256 277686
rect 124222 277610 124256 277618
rect 124222 277538 124256 277550
rect 124222 277466 124256 277482
rect 124222 277390 124256 277414
rect 124336 278055 124370 278089
rect 124336 277987 124370 278021
rect 124336 277919 124370 277953
rect 124336 277851 124370 277885
rect 124336 277783 124370 277817
rect 124336 277715 124370 277749
rect 124336 277647 124370 277681
rect 124336 277579 124370 277613
rect 124336 277511 124370 277545
rect 124336 277443 124370 277477
rect 124336 277375 124370 277409
rect 123656 277330 123678 277347
rect 122288 277273 122374 277307
rect 123494 277313 123678 277330
rect 123734 277313 123746 277347
rect 123806 277313 123814 277347
rect 123878 277313 123882 277347
rect 123984 277313 123988 277347
rect 124052 277313 124060 277347
rect 124120 277313 124132 277347
rect 124188 277313 124210 277347
rect 123494 277290 124210 277313
rect 124336 277307 124370 277341
rect 122254 277221 122374 277273
rect 124336 277221 124370 277273
rect 122254 277187 122343 277221
rect 122377 277187 122411 277221
rect 122445 277187 122479 277221
rect 122513 277187 122547 277221
rect 122581 277187 122615 277221
rect 122649 277187 122683 277221
rect 122717 277187 122751 277221
rect 122785 277187 122819 277221
rect 122853 277187 122887 277221
rect 122921 277187 122955 277221
rect 122989 277187 123023 277221
rect 123057 277187 123091 277221
rect 123125 277187 123159 277221
rect 123193 277187 123227 277221
rect 123261 277187 123295 277221
rect 123329 277187 123363 277221
rect 123397 277187 123431 277221
rect 123465 277187 123499 277221
rect 123533 277187 123567 277221
rect 123601 277187 123635 277221
rect 123669 277187 123703 277221
rect 123737 277187 123771 277221
rect 123805 277187 123839 277221
rect 123873 277187 123907 277221
rect 123941 277187 123975 277221
rect 124009 277187 124043 277221
rect 124077 277187 124111 277221
rect 124145 277187 124179 277221
rect 124213 277187 124247 277221
rect 124281 277187 124370 277221
rect 123686 277010 123945 277076
rect 123686 276904 123771 277010
rect 123877 276904 123945 277010
rect 123686 276851 123945 276904
rect 122278 276817 122404 276851
rect 122438 276817 122472 276851
rect 122506 276817 122540 276851
rect 122574 276817 122608 276851
rect 122642 276817 122676 276851
rect 122710 276817 122744 276851
rect 122778 276817 122812 276851
rect 122846 276817 122880 276851
rect 122914 276817 122948 276851
rect 122982 276817 123016 276851
rect 123050 276817 123084 276851
rect 123118 276817 123152 276851
rect 123186 276817 123220 276851
rect 123254 276817 123288 276851
rect 123322 276817 123356 276851
rect 123390 276817 123424 276851
rect 123458 276817 123492 276851
rect 123526 276817 123560 276851
rect 123594 276817 123628 276851
rect 123662 276817 123696 276851
rect 123730 276817 123764 276851
rect 123798 276817 123832 276851
rect 123866 276817 123992 276851
rect 122278 276749 123860 276817
rect 122278 276733 122470 276749
rect 122312 276715 122470 276733
rect 122506 276715 122540 276749
rect 122576 276715 122608 276749
rect 122648 276715 122676 276749
rect 122720 276715 122744 276749
rect 122792 276715 122812 276749
rect 122864 276715 122880 276749
rect 122936 276715 122948 276749
rect 123008 276715 123016 276749
rect 123080 276715 123084 276749
rect 123186 276715 123190 276749
rect 123254 276715 123262 276749
rect 123322 276715 123334 276749
rect 123390 276715 123406 276749
rect 123458 276715 123478 276749
rect 123526 276715 123550 276749
rect 123594 276715 123622 276749
rect 123662 276715 123694 276749
rect 123730 276715 123764 276749
rect 123800 276740 123860 276749
rect 123800 276715 123832 276740
rect 123958 276733 123992 276817
rect 125047 276742 125058 280856
rect 122312 276699 122426 276715
rect 122278 276665 122426 276699
rect 122312 276633 122426 276665
rect 122312 276631 122392 276633
rect 122278 276597 122392 276631
rect 122312 276563 122426 276597
rect 122278 276529 122392 276563
rect 122312 276527 122392 276529
rect 122312 276495 122426 276527
rect 122278 276461 122426 276495
rect 123844 276633 123878 276672
rect 123844 276563 123878 276597
rect 123844 276488 123878 276527
rect 123958 276665 123992 276699
rect 123958 276597 123992 276631
rect 123958 276529 123992 276563
rect 122312 276445 122426 276461
rect 123958 276461 123992 276495
rect 122312 276427 122470 276445
rect 122278 276411 122470 276427
rect 122506 276411 122540 276445
rect 122576 276411 122608 276445
rect 122648 276411 122676 276445
rect 122720 276411 122744 276445
rect 122792 276411 122812 276445
rect 122864 276411 122880 276445
rect 122936 276411 122948 276445
rect 123008 276411 123016 276445
rect 123080 276411 123084 276445
rect 123186 276411 123190 276445
rect 123254 276411 123262 276445
rect 123322 276411 123334 276445
rect 123390 276411 123406 276445
rect 123458 276411 123478 276445
rect 123526 276411 123550 276445
rect 123594 276411 123622 276445
rect 123662 276411 123694 276445
rect 123730 276411 123764 276445
rect 123800 276419 123832 276445
rect 123800 276411 123862 276419
rect 122278 276343 123862 276411
rect 123958 276343 123992 276427
rect 122278 276309 122404 276343
rect 122438 276309 122472 276343
rect 122506 276309 122540 276343
rect 122574 276309 122608 276343
rect 122642 276309 122676 276343
rect 122710 276309 122744 276343
rect 122778 276309 122812 276343
rect 122846 276309 122880 276343
rect 122914 276309 122948 276343
rect 122982 276309 123016 276343
rect 123050 276309 123084 276343
rect 123118 276309 123152 276343
rect 123186 276309 123220 276343
rect 123254 276309 123288 276343
rect 123322 276309 123356 276343
rect 123390 276309 123424 276343
rect 123458 276309 123492 276343
rect 123526 276309 123560 276343
rect 123594 276309 123628 276343
rect 123662 276309 123696 276343
rect 123730 276309 123764 276343
rect 123798 276309 123832 276343
rect 123866 276309 123992 276343
rect 124173 276382 125058 276742
rect 122136 276212 122552 276225
rect 124173 276212 124291 276382
rect 122136 276205 124313 276212
rect 122136 276112 122531 276205
rect 122136 276078 122137 276112
rect 122171 276078 122209 276112
rect 122243 276078 122281 276112
rect 122315 276078 122353 276112
rect 122387 276103 122531 276112
rect 124265 276103 124313 276205
rect 122387 276097 124313 276103
rect 122387 276078 122552 276097
rect 122136 276038 122552 276078
rect 124445 276049 124567 276110
rect 122136 276035 122427 276038
rect 122136 275562 122144 276035
rect 124445 276015 124490 276049
rect 124524 276015 124567 276049
rect 124445 275971 124567 276015
rect 122027 275515 122144 275562
rect 122283 275937 122379 275971
rect 122413 275937 122447 275971
rect 122481 275937 122515 275971
rect 122549 275937 122583 275971
rect 122617 275937 122651 275971
rect 122685 275937 122719 275971
rect 122753 275937 122787 275971
rect 122821 275937 122855 275971
rect 122889 275937 122923 275971
rect 122957 275937 122991 275971
rect 123025 275937 123059 275971
rect 123093 275937 123127 275971
rect 123161 275937 123195 275971
rect 123229 275937 123263 275971
rect 123297 275937 123331 275971
rect 123365 275937 123399 275971
rect 123433 275937 123467 275971
rect 123501 275937 123535 275971
rect 123569 275937 123603 275971
rect 123637 275937 123671 275971
rect 123705 275937 123739 275971
rect 123773 275937 123807 275971
rect 123841 275937 123875 275971
rect 123909 275937 123943 275971
rect 123977 275937 124011 275971
rect 124045 275937 124079 275971
rect 124113 275937 124147 275971
rect 124181 275937 124215 275971
rect 124249 275937 124283 275971
rect 124317 275937 124351 275971
rect 124385 275937 124419 275971
rect 124453 275937 124487 275971
rect 124521 275937 124555 275971
rect 124589 275937 124623 275971
rect 124657 275937 124691 275971
rect 124725 275937 124759 275971
rect 124793 275937 124827 275971
rect 124861 275937 124957 275971
rect 122283 275846 122317 275937
rect 122462 275823 122479 275857
rect 122539 275823 122547 275857
rect 122611 275823 122615 275857
rect 122717 275823 122721 275857
rect 122785 275823 122793 275857
rect 122853 275823 122870 275857
rect 123098 275823 123115 275857
rect 123175 275823 123183 275857
rect 123247 275823 123251 275857
rect 123353 275823 123357 275857
rect 123421 275823 123429 275857
rect 123489 275823 123506 275857
rect 123734 275823 123751 275857
rect 123811 275823 123819 275857
rect 123883 275823 123887 275857
rect 123989 275823 123993 275857
rect 124057 275823 124065 275857
rect 124125 275823 124142 275857
rect 124370 275823 124387 275857
rect 124447 275823 124455 275857
rect 124519 275823 124523 275857
rect 124625 275823 124629 275857
rect 124693 275823 124701 275857
rect 124761 275823 124778 275857
rect 124923 275846 124957 275937
rect 122283 275778 122317 275812
rect 122283 275710 122317 275744
rect 122385 275778 122419 275811
rect 122385 275711 122419 275744
rect 122913 275778 122947 275811
rect 122913 275711 122947 275744
rect 123021 275778 123055 275811
rect 123021 275711 123055 275744
rect 123549 275778 123583 275811
rect 123549 275711 123583 275744
rect 123657 275778 123691 275811
rect 123657 275711 123691 275744
rect 124185 275778 124219 275811
rect 124185 275711 124219 275744
rect 124293 275778 124327 275811
rect 124293 275711 124327 275744
rect 124821 275778 124855 275811
rect 124821 275711 124855 275744
rect 124923 275778 124957 275812
rect 124923 275710 124957 275744
rect 122283 275585 122317 275676
rect 122462 275665 122479 275699
rect 122539 275665 122547 275699
rect 122611 275665 122615 275699
rect 122717 275665 122721 275699
rect 122785 275665 122793 275699
rect 122853 275665 122870 275699
rect 122462 275585 122870 275665
rect 123098 275665 123115 275699
rect 123175 275665 123183 275699
rect 123247 275665 123251 275699
rect 123353 275665 123357 275699
rect 123421 275665 123429 275699
rect 123489 275665 123506 275699
rect 123098 275585 123506 275665
rect 123734 275665 123751 275699
rect 123811 275665 123819 275699
rect 123883 275665 123887 275699
rect 123989 275665 123993 275699
rect 124057 275665 124065 275699
rect 124125 275665 124142 275699
rect 123734 275585 124142 275665
rect 124370 275665 124387 275699
rect 124447 275665 124455 275699
rect 124519 275665 124523 275699
rect 124625 275665 124629 275699
rect 124693 275665 124701 275699
rect 124761 275665 124778 275699
rect 124370 275585 124778 275665
rect 124923 275585 124957 275676
rect 122283 275551 122379 275585
rect 122413 275551 122447 275585
rect 122481 275551 122515 275585
rect 122549 275551 122583 275585
rect 122617 275551 122651 275585
rect 122685 275551 122719 275585
rect 122753 275551 122787 275585
rect 122821 275551 122855 275585
rect 122889 275551 122923 275585
rect 122957 275551 122991 275585
rect 123025 275551 123059 275585
rect 123093 275551 123127 275585
rect 123161 275551 123195 275585
rect 123229 275551 123263 275585
rect 123297 275551 123331 275585
rect 123365 275551 123399 275585
rect 123433 275551 123467 275585
rect 123501 275551 123535 275585
rect 123569 275551 123603 275585
rect 123637 275551 123671 275585
rect 123705 275551 123739 275585
rect 123773 275551 123807 275585
rect 123841 275551 123875 275585
rect 123909 275551 123943 275585
rect 123977 275551 124011 275585
rect 124045 275551 124079 275585
rect 124113 275551 124147 275585
rect 124181 275551 124215 275585
rect 124249 275551 124283 275585
rect 124317 275551 124351 275585
rect 124385 275551 124419 275585
rect 124453 275551 124487 275585
rect 124521 275551 124555 275585
rect 124589 275551 124623 275585
rect 124657 275551 124691 275585
rect 124725 275551 124759 275585
rect 124793 275551 124827 275585
rect 124861 275551 124957 275585
rect 121728 275456 121809 275490
rect 121694 275422 121809 275456
rect 123246 275431 123421 275551
rect 121728 275388 121809 275422
rect 121694 275354 121809 275388
rect 121728 275320 121809 275354
rect 121694 275286 121809 275320
rect 121728 275252 121809 275286
rect 121694 275218 121809 275252
rect 121728 275184 121809 275218
rect 121694 275150 121809 275184
rect 121728 275116 121809 275150
rect 123213 275368 123457 275431
rect 123213 275190 123246 275368
rect 123424 275190 123457 275368
rect 123213 275140 123457 275190
rect 121694 275082 121809 275116
rect 121728 275048 121809 275082
rect 121694 275014 121809 275048
rect 121129 274968 121168 275002
rect 121210 274968 121240 275002
rect 121278 274968 121312 275002
rect 121346 274968 121380 275002
rect 121418 274968 121448 275002
rect 121490 274968 121529 275002
rect 121728 274980 121809 275014
rect 121694 274946 121809 274980
rect 121728 274912 121809 274946
rect 121694 274878 121809 274912
rect 121129 274812 121168 274846
rect 121210 274812 121240 274846
rect 121278 274812 121312 274846
rect 121346 274812 121380 274846
rect 121418 274812 121448 274846
rect 121490 274812 121529 274846
rect 121728 274844 121809 274878
rect 121694 274810 121809 274844
rect 121728 274776 121809 274810
rect 121083 274748 121117 274769
rect 121083 274676 121117 274702
rect 121083 274604 121117 274634
rect 120875 274566 121083 274579
rect 120841 274532 121117 274566
rect 120875 274498 121083 274532
rect 120841 274472 121117 274498
rect 120841 274464 120875 274472
rect 120841 274396 120875 274426
rect 120841 274328 120875 274354
rect 120841 274261 120875 274282
rect 121083 274464 121117 274472
rect 121083 274396 121117 274426
rect 121083 274328 121117 274354
rect 121083 274261 121117 274282
rect 121541 274748 121575 274769
rect 121541 274676 121575 274702
rect 121541 274604 121575 274634
rect 121541 274532 121575 274566
rect 121541 274464 121575 274498
rect 121541 274396 121575 274426
rect 121541 274328 121575 274354
rect 121541 274261 121575 274282
rect 121694 274742 121809 274776
rect 121728 274708 121809 274742
rect 121694 274674 121809 274708
rect 121728 274640 121809 274674
rect 121694 274606 121809 274640
rect 121728 274572 121809 274606
rect 121694 274538 121809 274572
rect 122792 275002 122891 275036
rect 122925 275002 122959 275036
rect 122993 275002 123027 275036
rect 123061 275002 123095 275036
rect 123129 275002 123163 275036
rect 123197 275002 123231 275036
rect 123265 275002 123299 275036
rect 123333 275002 123367 275036
rect 123401 275002 123435 275036
rect 123469 275002 123503 275036
rect 123537 275002 123571 275036
rect 123605 275002 123639 275036
rect 123673 275002 123707 275036
rect 123741 275002 123775 275036
rect 123809 275002 123843 275036
rect 123877 275002 123911 275036
rect 123945 275002 123979 275036
rect 124013 275002 124112 275036
rect 122792 274915 122826 275002
rect 122952 274900 122993 274934
rect 123037 274900 123061 274934
rect 123109 274900 123129 274934
rect 123181 274900 123197 274934
rect 123253 274900 123265 274934
rect 123325 274900 123333 274934
rect 123397 274900 123401 274934
rect 123503 274900 123507 274934
rect 123571 274900 123579 274934
rect 123639 274900 123651 274934
rect 123707 274900 123723 274934
rect 123775 274900 123795 274934
rect 123843 274900 123867 274934
rect 123911 274900 123952 274934
rect 124078 274915 124112 275002
rect 122792 274847 122826 274881
rect 122792 274779 122826 274813
rect 122792 274711 122826 274745
rect 122792 274643 122826 274677
rect 122906 274847 122940 274866
rect 122906 274779 122940 274781
rect 122906 274743 122940 274745
rect 122906 274658 122940 274677
rect 123964 274847 123998 274866
rect 124078 274847 124112 274881
rect 123998 274813 124078 274816
rect 123998 274781 124112 274813
rect 123964 274779 124112 274781
rect 123998 274745 124078 274779
rect 123964 274743 124112 274745
rect 123998 274715 124112 274743
rect 123964 274658 123998 274677
rect 124078 274711 124112 274715
rect 124078 274643 124112 274677
rect 122792 274562 122826 274609
rect 122952 274590 122993 274624
rect 123037 274590 123061 274624
rect 123109 274590 123129 274624
rect 123181 274590 123197 274624
rect 123253 274590 123265 274624
rect 123325 274590 123333 274624
rect 123397 274590 123401 274624
rect 123503 274590 123507 274624
rect 123571 274590 123579 274624
rect 123639 274590 123651 274624
rect 123707 274590 123723 274624
rect 123775 274590 123795 274624
rect 123843 274590 123867 274624
rect 123911 274590 123952 274624
rect 121728 274504 121809 274538
rect 121694 274470 121809 274504
rect 121728 274436 121809 274470
rect 121694 274402 121809 274436
rect 121728 274368 121809 274402
rect 121694 274334 121809 274368
rect 122060 274541 122826 274562
rect 122060 274507 122110 274541
rect 122144 274507 122178 274541
rect 122212 274507 122246 274541
rect 122280 274507 122314 274541
rect 122348 274507 122382 274541
rect 122416 274507 122450 274541
rect 122484 274507 122518 274541
rect 122552 274507 122586 274541
rect 122620 274507 122654 274541
rect 122688 274522 122826 274541
rect 124078 274537 124112 274609
rect 124202 274555 124840 274582
rect 125047 274555 125058 276382
rect 124202 274552 125058 274555
rect 124202 274537 124232 274552
rect 124078 274522 124232 274537
rect 122688 274507 122891 274522
rect 122060 274488 122891 274507
rect 122925 274488 122959 274522
rect 122993 274488 123027 274522
rect 123061 274488 123095 274522
rect 123129 274488 123163 274522
rect 123197 274488 123231 274522
rect 123265 274488 123299 274522
rect 123333 274488 123367 274522
rect 123401 274488 123435 274522
rect 123469 274488 123503 274522
rect 123537 274488 123571 274522
rect 123605 274488 123639 274522
rect 123673 274488 123707 274522
rect 123741 274488 123775 274522
rect 123809 274488 123843 274522
rect 123877 274488 123911 274522
rect 123945 274488 123979 274522
rect 124013 274518 124232 274522
rect 124266 274518 124300 274552
rect 124334 274518 124368 274552
rect 124402 274518 124436 274552
rect 124470 274518 124504 274552
rect 124538 274518 124572 274552
rect 124606 274518 124640 274552
rect 124674 274518 124708 274552
rect 124742 274518 124776 274552
rect 124810 274518 125058 274552
rect 124013 274488 125058 274518
rect 122060 274486 122730 274488
rect 122060 274354 122253 274486
rect 122523 274354 122558 274392
rect 121728 274300 121809 274334
rect 121694 274266 121809 274300
rect 122061 274350 122558 274354
rect 122061 274316 122324 274350
rect 122360 274316 122394 274350
rect 122430 274316 122558 274350
rect 122693 274316 122740 274350
rect 122776 274316 122810 274350
rect 122846 274316 122893 274350
rect 122061 274282 122558 274316
rect 122939 274282 122974 274488
rect 123497 274443 123670 274452
rect 123497 274437 123534 274443
rect 123354 274409 123534 274437
rect 123568 274409 123606 274443
rect 123640 274437 123670 274443
rect 123640 274409 123806 274437
rect 123354 274399 123806 274409
rect 123354 274387 123390 274399
rect 123109 274316 123156 274350
rect 123192 274316 123226 274350
rect 123262 274316 123309 274350
rect 123355 274282 123390 274387
rect 123525 274316 123572 274350
rect 123608 274316 123642 274350
rect 123678 274316 123725 274350
rect 123771 274282 123806 274399
rect 123941 274316 123988 274350
rect 124024 274316 124058 274350
rect 124094 274316 124141 274350
rect 124187 274282 124222 274488
rect 124603 274354 124638 274392
rect 124726 274354 125058 274488
rect 120271 274232 120395 274261
rect 120237 274198 120395 274232
rect 121728 274232 121809 274266
rect 120271 274164 120395 274198
rect 120429 274184 120468 274218
rect 120510 274184 120540 274218
rect 120578 274184 120612 274218
rect 120646 274184 120680 274218
rect 120718 274184 120748 274218
rect 120790 274184 120829 274218
rect 121129 274184 121168 274218
rect 121210 274184 121240 274218
rect 121278 274184 121312 274218
rect 121346 274184 121380 274218
rect 121418 274184 121448 274218
rect 121490 274184 121529 274218
rect 121694 274198 121809 274232
rect 120237 274130 120395 274164
rect 120271 274096 120395 274130
rect 120237 274062 120395 274096
rect 121728 274164 121809 274198
rect 121694 274130 121809 274164
rect 121728 274096 121809 274130
rect 121694 274062 121809 274096
rect 120271 274028 120395 274062
rect 120429 274028 120468 274062
rect 120510 274028 120540 274062
rect 120578 274028 120612 274062
rect 120646 274028 120680 274062
rect 120718 274028 120748 274062
rect 120790 274028 120829 274062
rect 121129 274028 121168 274062
rect 121210 274028 121240 274062
rect 121278 274028 121312 274062
rect 121346 274028 121380 274062
rect 121418 274028 121448 274062
rect 121490 274028 121529 274062
rect 121728 274028 121809 274062
rect 120237 273994 120395 274028
rect 120271 273985 120395 273994
rect 121694 273994 121809 274028
rect 120271 273964 120417 273985
rect 120271 273960 120383 273964
rect 120237 273926 120383 273960
rect 120271 273918 120383 273926
rect 120271 273892 120417 273918
rect 120237 273858 120383 273892
rect 120271 273850 120383 273858
rect 120271 273824 120417 273850
rect 120237 273820 120417 273824
rect 120237 273790 120383 273820
rect 120271 273782 120383 273790
rect 120271 273756 120417 273782
rect 120237 273748 120417 273756
rect 120237 273722 120383 273748
rect 120271 273714 120383 273722
rect 120271 273688 120417 273714
rect 120237 273680 120417 273688
rect 120237 273654 120383 273680
rect 120271 273642 120383 273654
rect 120271 273620 120417 273642
rect 120237 273612 120417 273620
rect 120237 273586 120383 273612
rect 120271 273570 120383 273586
rect 120271 273552 120417 273570
rect 120237 273544 120417 273552
rect 120237 273518 120383 273544
rect 120271 273498 120383 273518
rect 120271 273484 120417 273498
rect 120237 273477 120417 273484
rect 120841 273964 120875 273985
rect 120841 273892 120875 273918
rect 120841 273820 120875 273850
rect 120841 273778 120875 273782
rect 121083 273964 121117 273985
rect 121083 273892 121117 273918
rect 121083 273820 121117 273850
rect 121083 273778 121117 273782
rect 120841 273748 121117 273778
rect 120875 273741 121083 273748
rect 120875 273714 120972 273741
rect 120841 273707 120972 273714
rect 121006 273714 121083 273741
rect 121006 273707 121117 273714
rect 120841 273680 121117 273707
rect 120875 273671 121083 273680
rect 120841 273612 120875 273642
rect 120841 273544 120875 273570
rect 120841 273477 120875 273498
rect 121083 273612 121117 273642
rect 121083 273544 121117 273570
rect 121083 273477 121117 273498
rect 121541 273964 121575 273985
rect 121541 273892 121575 273918
rect 121541 273820 121575 273850
rect 121541 273748 121575 273782
rect 121541 273680 121575 273714
rect 121541 273612 121575 273642
rect 121541 273544 121575 273570
rect 121541 273477 121575 273498
rect 121728 273960 121809 273994
rect 121694 273926 121809 273960
rect 121728 273892 121809 273926
rect 121694 273858 121809 273892
rect 121728 273824 121809 273858
rect 121694 273790 121809 273824
rect 121728 273756 121809 273790
rect 121694 273722 121809 273756
rect 121728 273688 121809 273722
rect 121694 273654 121809 273688
rect 121728 273620 121809 273654
rect 121694 273586 121809 273620
rect 121728 273552 121809 273586
rect 121694 273518 121809 273552
rect 122062 274281 122265 274282
rect 122062 274247 122089 274281
rect 122123 274261 122265 274281
rect 122123 274247 122231 274261
rect 122062 274215 122231 274247
rect 122062 274213 122265 274215
rect 122062 274179 122089 274213
rect 122123 274189 122265 274213
rect 122123 274179 122231 274189
rect 122062 274147 122231 274179
rect 122062 274145 122265 274147
rect 122062 274111 122089 274145
rect 122123 274117 122265 274145
rect 122123 274111 122231 274117
rect 122062 274079 122231 274111
rect 122062 274077 122265 274079
rect 122062 274043 122089 274077
rect 122123 274045 122265 274077
rect 122123 274043 122231 274045
rect 122062 274011 122231 274043
rect 122062 274009 122265 274011
rect 122062 273975 122089 274009
rect 122123 273977 122265 274009
rect 122123 273975 122231 273977
rect 122062 273941 122231 273975
rect 122062 273907 122089 273941
rect 122123 273939 122231 273941
rect 122123 273909 122265 273939
rect 122123 273907 122231 273909
rect 122062 273873 122231 273907
rect 122062 273839 122089 273873
rect 122123 273867 122231 273873
rect 122123 273841 122265 273867
rect 122123 273839 122231 273841
rect 122062 273805 122231 273839
rect 122062 273771 122089 273805
rect 122123 273795 122231 273805
rect 122123 273774 122265 273795
rect 122489 274261 122558 274282
rect 122523 274215 122558 274261
rect 122489 274189 122558 274215
rect 122523 274147 122558 274189
rect 122489 274117 122558 274147
rect 122523 274079 122558 274117
rect 122489 274045 122558 274079
rect 122523 274011 122558 274045
rect 122489 273977 122558 274011
rect 122523 273939 122558 273977
rect 122489 273909 122558 273939
rect 122523 273867 122558 273909
rect 122489 273841 122558 273867
rect 122523 273795 122558 273841
rect 122489 273774 122558 273795
rect 122647 274261 122681 274282
rect 122647 274189 122681 274215
rect 122647 274117 122681 274147
rect 122647 274045 122681 274079
rect 122647 273977 122681 274011
rect 122647 273909 122681 273939
rect 122647 273841 122681 273867
rect 122647 273774 122681 273795
rect 122905 274261 122974 274282
rect 122939 274215 122974 274261
rect 122905 274189 122974 274215
rect 122939 274147 122974 274189
rect 122905 274117 122974 274147
rect 122939 274079 122974 274117
rect 122905 274045 122974 274079
rect 122939 274011 122974 274045
rect 122905 273977 122974 274011
rect 122939 273939 122974 273977
rect 122905 273909 122974 273939
rect 122939 273867 122974 273909
rect 122905 273841 122974 273867
rect 122939 273795 122974 273841
rect 122905 273774 122974 273795
rect 123063 274261 123097 274282
rect 123063 274189 123097 274215
rect 123063 274117 123097 274147
rect 123063 274045 123097 274079
rect 123063 273977 123097 274011
rect 123063 273909 123097 273939
rect 123063 273841 123097 273867
rect 123063 273774 123097 273795
rect 123321 274261 123390 274282
rect 123355 274215 123390 274261
rect 123321 274189 123390 274215
rect 123355 274147 123390 274189
rect 123321 274117 123390 274147
rect 123355 274079 123390 274117
rect 123321 274045 123390 274079
rect 123355 274011 123390 274045
rect 123321 273977 123390 274011
rect 123355 273939 123390 273977
rect 123321 273909 123390 273939
rect 123355 273867 123390 273909
rect 123321 273841 123390 273867
rect 123355 273795 123390 273841
rect 123321 273774 123390 273795
rect 123479 274261 123513 274282
rect 123479 274189 123513 274215
rect 123479 274117 123513 274147
rect 123479 274045 123513 274079
rect 123479 273977 123513 274011
rect 123479 273909 123513 273939
rect 123479 273841 123513 273867
rect 123479 273774 123513 273795
rect 123737 274261 123806 274282
rect 123771 274215 123806 274261
rect 123737 274189 123806 274215
rect 123771 274147 123806 274189
rect 123737 274117 123806 274147
rect 123771 274079 123806 274117
rect 123737 274045 123806 274079
rect 123771 274011 123806 274045
rect 123737 273977 123806 274011
rect 123771 273939 123806 273977
rect 123737 273909 123806 273939
rect 123771 273867 123806 273909
rect 123737 273841 123806 273867
rect 123771 273795 123806 273841
rect 123737 273774 123806 273795
rect 123895 274261 123929 274282
rect 123895 274189 123929 274215
rect 123895 274117 123929 274147
rect 123895 274045 123929 274079
rect 123895 273977 123929 274011
rect 123895 273909 123929 273939
rect 123895 273841 123929 273867
rect 123895 273774 123929 273795
rect 124153 274261 124222 274282
rect 124187 274215 124222 274261
rect 124153 274189 124222 274215
rect 124187 274147 124222 274189
rect 124153 274117 124222 274147
rect 124187 274079 124222 274117
rect 124153 274045 124222 274079
rect 124187 274011 124222 274045
rect 124153 273977 124222 274011
rect 124187 273939 124222 273977
rect 124153 273909 124222 273939
rect 124187 273867 124222 273909
rect 124153 273841 124222 273867
rect 124187 273795 124222 273841
rect 124153 273774 124222 273795
rect 124311 274350 125058 274354
rect 124311 274316 124404 274350
rect 124440 274316 124474 274350
rect 124510 274316 125058 274350
rect 124311 274297 125058 274316
rect 124311 274282 124753 274297
rect 124311 274261 124345 274282
rect 124311 274189 124345 274215
rect 124311 274117 124345 274147
rect 124311 274045 124345 274079
rect 124311 273977 124345 274011
rect 124311 273909 124345 273939
rect 124311 273841 124345 273867
rect 124311 273774 124345 273795
rect 124569 274263 124753 274282
rect 124787 274263 125058 274297
rect 124569 274261 125058 274263
rect 124603 274229 125058 274261
rect 124603 274215 124753 274229
rect 124569 274195 124753 274215
rect 124787 274195 125058 274229
rect 124569 274189 125058 274195
rect 124603 274161 125058 274189
rect 124603 274147 124753 274161
rect 124569 274127 124753 274147
rect 124787 274127 125058 274161
rect 124569 274117 125058 274127
rect 124603 274093 125058 274117
rect 124603 274079 124753 274093
rect 124569 274059 124753 274079
rect 124787 274059 125058 274093
rect 124569 274045 125058 274059
rect 124603 274025 125058 274045
rect 124603 274011 124753 274025
rect 124569 273991 124753 274011
rect 124787 273991 125058 274025
rect 124569 273977 125058 273991
rect 124603 273957 125058 273977
rect 124603 273939 124753 273957
rect 124569 273923 124753 273939
rect 124787 273923 125058 273957
rect 124569 273909 125058 273923
rect 124603 273889 125058 273909
rect 124603 273867 124753 273889
rect 124569 273855 124753 273867
rect 124787 273855 125058 273889
rect 124569 273841 125058 273855
rect 124603 273821 125058 273841
rect 124603 273795 124753 273821
rect 124569 273787 124753 273795
rect 124787 273787 125058 273821
rect 124569 273774 125058 273787
rect 122123 273771 122558 273774
rect 122062 273740 122558 273771
rect 124311 273753 125058 273774
rect 124311 273740 124753 273753
rect 122062 273737 122324 273740
rect 122062 273703 122089 273737
rect 122123 273706 122324 273737
rect 122360 273706 122394 273740
rect 122430 273706 122558 273740
rect 122693 273706 122740 273740
rect 122776 273706 122810 273740
rect 122846 273706 122893 273740
rect 123109 273706 123156 273740
rect 123192 273706 123226 273740
rect 123262 273706 123309 273740
rect 123525 273706 123572 273740
rect 123608 273706 123642 273740
rect 123678 273706 123725 273740
rect 123941 273706 123988 273740
rect 124024 273706 124058 273740
rect 124094 273706 124141 273740
rect 124311 273706 124404 273740
rect 124440 273706 124474 273740
rect 124510 273719 124753 273740
rect 124787 273719 125058 273753
rect 124510 273706 125058 273719
rect 122123 273703 122558 273706
rect 122062 273702 122558 273703
rect 124311 273702 125058 273706
rect 122062 273669 122253 273702
rect 122062 273635 122089 273669
rect 122123 273635 122253 273669
rect 122062 273618 122253 273635
rect 124610 273685 125058 273702
rect 124610 273651 124753 273685
rect 124787 273651 125058 273685
rect 124610 273618 125058 273651
rect 122062 273598 125058 273618
rect 122062 273564 122243 273598
rect 122277 273564 122311 273598
rect 122345 273564 122379 273598
rect 122413 273564 122447 273598
rect 122481 273564 122515 273598
rect 122549 273564 122583 273598
rect 122617 273564 122651 273598
rect 122685 273564 122719 273598
rect 122753 273564 122787 273598
rect 122821 273564 122855 273598
rect 122889 273564 122923 273598
rect 122957 273564 122991 273598
rect 123025 273564 123059 273598
rect 123093 273564 123127 273598
rect 123161 273564 123195 273598
rect 123229 273564 123263 273598
rect 123297 273564 123331 273598
rect 123365 273564 123399 273598
rect 123433 273564 123467 273598
rect 123501 273564 123535 273598
rect 123569 273564 123603 273598
rect 123637 273564 123671 273598
rect 123705 273564 123739 273598
rect 123773 273564 123807 273598
rect 123841 273564 123875 273598
rect 123909 273564 123943 273598
rect 123977 273564 124011 273598
rect 124045 273564 124079 273598
rect 124113 273564 124147 273598
rect 124181 273564 124215 273598
rect 124249 273564 124283 273598
rect 124317 273564 124351 273598
rect 124385 273564 124419 273598
rect 124453 273564 124487 273598
rect 124521 273564 124555 273598
rect 124589 273564 125058 273598
rect 122062 273545 125058 273564
rect 121728 273484 121809 273518
rect 120237 273450 120395 273477
rect 120271 273416 120395 273450
rect 121694 273450 121809 273484
rect 120237 273382 120395 273416
rect 120429 273400 120468 273434
rect 120510 273400 120540 273434
rect 120578 273400 120612 273434
rect 120646 273400 120680 273434
rect 120718 273400 120748 273434
rect 120790 273400 120829 273434
rect 121129 273400 121168 273434
rect 121210 273400 121240 273434
rect 121278 273400 121312 273434
rect 121346 273400 121380 273434
rect 121418 273400 121448 273434
rect 121490 273400 121529 273434
rect 121728 273416 121809 273450
rect 120271 273348 120395 273382
rect 120237 273314 120395 273348
rect 120271 273280 120395 273314
rect 120237 273246 120395 273280
rect 121694 273382 121809 273416
rect 121728 273348 121809 273382
rect 121694 273314 121809 273348
rect 121728 273280 121809 273314
rect 120271 273212 120395 273246
rect 120429 273244 120468 273278
rect 120510 273244 120540 273278
rect 120578 273244 120612 273278
rect 120646 273244 120680 273278
rect 120718 273244 120748 273278
rect 120790 273244 120829 273278
rect 121129 273244 121168 273278
rect 121210 273244 121240 273278
rect 121278 273244 121312 273278
rect 121346 273244 121380 273278
rect 121418 273244 121448 273278
rect 121490 273244 121529 273278
rect 121694 273246 121809 273280
rect 120237 273201 120395 273212
rect 121728 273212 121809 273246
rect 120237 273180 120417 273201
rect 120237 273178 120383 273180
rect 120271 273144 120383 273178
rect 120237 273134 120383 273144
rect 120237 273110 120417 273134
rect 120271 273108 120417 273110
rect 120271 273076 120383 273108
rect 120237 273066 120383 273076
rect 120237 273042 120417 273066
rect 120271 273036 120417 273042
rect 120271 273008 120383 273036
rect 120237 272998 120383 273008
rect 120237 272974 120417 272998
rect 120271 272964 120417 272974
rect 120271 272940 120383 272964
rect 120237 272930 120383 272940
rect 120237 272906 120417 272930
rect 120271 272896 120417 272906
rect 120271 272872 120383 272896
rect 120237 272858 120383 272872
rect 120237 272838 120417 272858
rect 120271 272828 120417 272838
rect 120271 272804 120383 272828
rect 120237 272786 120383 272804
rect 120237 272770 120417 272786
rect 120271 272760 120417 272770
rect 120271 272736 120383 272760
rect 120237 272714 120383 272736
rect 120237 272702 120417 272714
rect 120271 272693 120417 272702
rect 120841 273180 120875 273201
rect 120841 273108 120875 273134
rect 120841 273036 120875 273066
rect 120841 272964 120875 272998
rect 120841 272896 120875 272930
rect 120841 272828 120875 272858
rect 120841 272760 120875 272786
rect 120841 272693 120875 272714
rect 121083 273180 121117 273201
rect 121083 273108 121117 273134
rect 121083 273036 121117 273066
rect 121083 272964 121117 272998
rect 121083 272896 121117 272930
rect 121083 272828 121117 272858
rect 121083 272760 121117 272786
rect 121083 272693 121117 272714
rect 121541 273180 121575 273201
rect 121541 273108 121575 273134
rect 121541 273036 121575 273066
rect 121541 272964 121575 272998
rect 121541 272896 121575 272930
rect 121541 272828 121575 272858
rect 121541 272760 121575 272786
rect 121541 272693 121575 272714
rect 121694 273178 121809 273212
rect 121728 273144 121809 273178
rect 121694 273110 121809 273144
rect 121728 273076 121809 273110
rect 121694 273057 121809 273076
rect 121694 273042 123538 273057
rect 121728 273008 123538 273042
rect 121694 272998 123538 273008
rect 121694 272974 122006 272998
rect 121728 272964 122006 272974
rect 122040 272964 122074 272998
rect 122108 272964 122142 272998
rect 122176 272964 122210 272998
rect 122244 272964 122278 272998
rect 122312 272964 122346 272998
rect 122380 272964 122414 272998
rect 122448 272964 122482 272998
rect 122516 272964 122550 272998
rect 122584 272964 122618 272998
rect 122652 272964 122686 272998
rect 122720 272964 122754 272998
rect 122788 272964 122822 272998
rect 122856 272964 122890 272998
rect 122924 272964 122958 272998
rect 122992 272964 123026 272998
rect 123060 272964 123094 272998
rect 123128 272964 123162 272998
rect 123196 272964 123230 272998
rect 123264 272964 123298 272998
rect 123332 272964 123366 272998
rect 123400 272964 123434 272998
rect 123468 272964 123554 272998
rect 121728 272954 123554 272964
rect 121728 272940 121954 272954
rect 121694 272917 121954 272940
rect 121694 272906 121920 272917
rect 121728 272883 121920 272906
rect 121728 272872 121954 272883
rect 121694 272849 121954 272872
rect 121694 272838 121920 272849
rect 121728 272815 121920 272838
rect 121728 272804 121954 272815
rect 121694 272781 121954 272804
rect 121694 272770 121920 272781
rect 121728 272747 121920 272770
rect 121728 272736 121954 272747
rect 121694 272713 121954 272736
rect 121694 272702 121920 272713
rect 120271 272668 120395 272693
rect 120237 272634 120395 272668
rect 121728 272679 121920 272702
rect 121728 272668 121954 272679
rect 120271 272600 120395 272634
rect 120429 272616 120468 272650
rect 120510 272616 120540 272650
rect 120578 272616 120612 272650
rect 120646 272616 120680 272650
rect 120718 272616 120748 272650
rect 120790 272616 120829 272650
rect 121129 272616 121168 272650
rect 121210 272616 121240 272650
rect 121278 272616 121312 272650
rect 121346 272616 121380 272650
rect 121418 272616 121448 272650
rect 121490 272616 121529 272650
rect 121694 272645 121954 272668
rect 121694 272634 121920 272645
rect 120237 272566 120395 272600
rect 120271 272532 120395 272566
rect 120237 272498 120395 272532
rect 120271 272464 120395 272498
rect 121728 272611 121920 272634
rect 122079 272894 122571 272954
rect 122079 272860 122164 272894
rect 122206 272860 122236 272894
rect 122274 272860 122308 272894
rect 122342 272860 122376 272894
rect 122414 272860 122444 272894
rect 122486 272860 122571 272894
rect 122079 272780 122125 272860
rect 122113 272746 122125 272780
rect 122079 272666 122125 272746
rect 122525 272780 122571 272860
rect 122525 272746 122537 272780
rect 122525 272666 122571 272746
rect 122079 272632 122164 272666
rect 122206 272632 122236 272666
rect 122274 272632 122308 272666
rect 122342 272632 122376 272666
rect 122414 272632 122444 272666
rect 122486 272632 122571 272666
rect 122779 272894 123271 272954
rect 122779 272860 122864 272894
rect 122906 272860 122936 272894
rect 122974 272860 123008 272894
rect 123042 272860 123076 272894
rect 123114 272860 123144 272894
rect 123186 272860 123271 272894
rect 122779 272780 122825 272860
rect 122813 272746 122825 272780
rect 122779 272666 122825 272746
rect 123225 272780 123271 272860
rect 123225 272746 123237 272780
rect 123225 272666 123271 272746
rect 122779 272632 122864 272666
rect 122906 272632 122936 272666
rect 122974 272632 123008 272666
rect 123042 272632 123076 272666
rect 123114 272632 123144 272666
rect 123186 272632 123271 272666
rect 123520 272917 123554 272954
rect 123520 272849 123554 272883
rect 123520 272781 123554 272815
rect 123520 272713 123554 272747
rect 121728 272600 121954 272611
rect 121694 272577 121954 272600
rect 121694 272566 121920 272577
rect 121728 272543 121920 272566
rect 121728 272532 121954 272543
rect 121694 272509 121954 272532
rect 123333 272625 123462 272656
rect 123333 272591 123382 272625
rect 123416 272591 123462 272625
rect 123333 272553 123462 272591
rect 123333 272519 123382 272553
rect 123416 272519 123462 272553
rect 123333 272510 123462 272519
rect 121694 272498 121920 272509
rect 120237 272430 120395 272464
rect 120429 272460 120468 272494
rect 120510 272460 120540 272494
rect 120578 272460 120612 272494
rect 120646 272460 120680 272494
rect 120718 272460 120748 272494
rect 120790 272460 120829 272494
rect 121129 272460 121168 272494
rect 121210 272460 121240 272494
rect 121278 272460 121312 272494
rect 121346 272460 121380 272494
rect 121418 272460 121448 272494
rect 121490 272460 121529 272494
rect 121728 272475 121920 272498
rect 122125 272476 122164 272510
rect 122206 272476 122236 272510
rect 122274 272476 122308 272510
rect 122342 272476 122376 272510
rect 122414 272476 122444 272510
rect 122486 272476 122525 272510
rect 122825 272476 122864 272510
rect 122906 272476 122936 272510
rect 122974 272476 123008 272510
rect 123042 272476 123076 272510
rect 123114 272476 123144 272510
rect 123186 272481 123462 272510
rect 123186 272476 123382 272481
rect 121728 272464 121954 272475
rect 120271 272417 120395 272430
rect 121694 272441 121954 272464
rect 121694 272430 121920 272441
rect 120271 272396 120417 272417
rect 120237 272362 120383 272396
rect 120271 272350 120383 272362
rect 120271 272328 120417 272350
rect 120237 272324 120417 272328
rect 120237 272294 120383 272324
rect 120271 272282 120383 272294
rect 120271 272260 120417 272282
rect 120237 272252 120417 272260
rect 120237 272226 120383 272252
rect 120271 272214 120383 272226
rect 120271 272192 120417 272214
rect 120237 272180 120417 272192
rect 120237 272158 120383 272180
rect 120271 272146 120383 272158
rect 120271 272124 120417 272146
rect 120237 272112 120417 272124
rect 120237 272090 120383 272112
rect 120271 272074 120383 272090
rect 120271 272056 120417 272074
rect 120237 272044 120417 272056
rect 120237 272022 120383 272044
rect 120271 272002 120383 272022
rect 120271 271988 120417 272002
rect 120237 271976 120417 271988
rect 120237 271954 120383 271976
rect 120271 271930 120383 271954
rect 120271 271920 120417 271930
rect 120237 271909 120417 271920
rect 120841 272396 120875 272417
rect 120841 272324 120875 272350
rect 120841 272252 120875 272282
rect 120841 272180 120875 272214
rect 120841 272112 120875 272146
rect 120841 272044 120875 272074
rect 120841 271976 120875 272002
rect 120841 271909 120875 271930
rect 121083 272396 121117 272417
rect 121083 272324 121117 272350
rect 121083 272252 121117 272282
rect 121083 272180 121117 272214
rect 121083 272112 121117 272146
rect 121083 272044 121117 272074
rect 121083 271976 121117 272002
rect 121083 271909 121117 271930
rect 121541 272396 121575 272417
rect 121541 272324 121575 272350
rect 121541 272252 121575 272282
rect 121541 272180 121575 272214
rect 121541 272112 121575 272146
rect 121541 272044 121575 272074
rect 121541 271976 121575 272002
rect 121541 271909 121575 271930
rect 121728 272407 121920 272430
rect 123333 272447 123382 272476
rect 123416 272447 123462 272481
rect 121728 272396 121954 272407
rect 121694 272373 121954 272396
rect 121694 272362 121920 272373
rect 121728 272339 121920 272362
rect 121728 272328 121954 272339
rect 121694 272305 121954 272328
rect 121694 272294 121920 272305
rect 121728 272271 121920 272294
rect 121728 272260 121954 272271
rect 121694 272248 121954 272260
rect 122079 272412 122113 272433
rect 122079 272340 122113 272366
rect 122079 272268 122113 272298
rect 121694 272237 122079 272248
rect 121694 272226 121920 272237
rect 121728 272203 121920 272226
rect 121954 272230 122079 272237
rect 121954 272203 122113 272230
rect 121728 272196 122113 272203
rect 121728 272192 122079 272196
rect 121694 272169 122079 272192
rect 121694 272158 121920 272169
rect 121728 272135 121920 272158
rect 121954 272162 122079 272169
rect 121954 272135 122113 272162
rect 121728 272128 122113 272135
rect 121728 272124 122079 272128
rect 121694 272123 122079 272124
rect 121694 272101 121954 272123
rect 121694 272090 121920 272101
rect 121728 272067 121920 272090
rect 121728 272056 121954 272067
rect 121694 272033 121954 272056
rect 121694 272022 121920 272033
rect 121728 271999 121920 272022
rect 121728 271988 121954 271999
rect 121694 271965 121954 271988
rect 121694 271954 121920 271965
rect 121728 271931 121920 271954
rect 121728 271920 121954 271931
rect 122079 272060 122113 272090
rect 122079 271992 122113 272018
rect 122079 271925 122113 271946
rect 122537 272412 122571 272433
rect 122537 272340 122571 272366
rect 122537 272268 122571 272298
rect 122779 272412 122813 272433
rect 122779 272340 122813 272366
rect 122779 272268 122813 272298
rect 122571 272230 122779 272235
rect 122537 272199 122813 272230
rect 122537 272196 122665 272199
rect 122571 272165 122665 272196
rect 122699 272196 122813 272199
rect 122699 272165 122779 272196
rect 122571 272162 122779 272165
rect 122537 272128 122813 272162
rect 122537 272060 122571 272090
rect 122537 271992 122571 272018
rect 122537 271925 122571 271946
rect 122779 272060 122813 272090
rect 122779 271992 122813 272018
rect 122779 271925 122813 271946
rect 123237 272412 123271 272433
rect 123237 272340 123271 272366
rect 123237 272268 123271 272298
rect 123237 272196 123271 272230
rect 123237 272128 123271 272162
rect 123237 272060 123271 272090
rect 123237 271992 123271 272018
rect 123237 271925 123271 271946
rect 123333 272427 123462 272447
rect 123520 272645 123554 272679
rect 123520 272577 123554 272611
rect 123520 272509 123554 272543
rect 123520 272441 123554 272475
rect 120237 271886 120395 271909
rect 120271 271852 120395 271886
rect 121694 271897 121954 271920
rect 121694 271886 121920 271897
rect 120237 271818 120395 271852
rect 120429 271832 120468 271866
rect 120510 271832 120540 271866
rect 120578 271832 120612 271866
rect 120646 271832 120680 271866
rect 120718 271832 120748 271866
rect 120790 271832 120829 271866
rect 121129 271832 121168 271866
rect 121210 271832 121240 271866
rect 121278 271832 121312 271866
rect 121346 271832 121380 271866
rect 121418 271832 121448 271866
rect 121490 271832 121529 271866
rect 121728 271863 121920 271886
rect 123333 271882 123367 272427
rect 121728 271852 121954 271863
rect 120271 271784 120395 271818
rect 120237 271750 120395 271784
rect 120271 271716 120395 271750
rect 120237 271682 120395 271716
rect 121694 271829 121954 271852
rect 122125 271848 122164 271882
rect 122206 271848 122236 271882
rect 122274 271848 122308 271882
rect 122342 271848 122376 271882
rect 122414 271848 122444 271882
rect 122486 271848 122525 271882
rect 122825 271848 122864 271882
rect 122906 271848 122936 271882
rect 122974 271848 123008 271882
rect 123042 271848 123076 271882
rect 123114 271848 123144 271882
rect 123186 271848 123367 271882
rect 123520 272373 123554 272407
rect 123520 272305 123554 272339
rect 123520 272237 123554 272271
rect 123520 272169 123554 272203
rect 123520 272101 123554 272135
rect 123520 272033 123554 272067
rect 123520 271965 123554 271999
rect 123520 271897 123554 271931
rect 121694 271818 121920 271829
rect 121728 271795 121920 271818
rect 121728 271784 121954 271795
rect 121694 271761 121954 271784
rect 121694 271750 121920 271761
rect 121728 271727 121920 271750
rect 121728 271716 121954 271727
rect 123520 271829 123554 271863
rect 123520 271761 123554 271795
rect 120271 271648 120395 271682
rect 120429 271676 120468 271710
rect 120510 271676 120540 271710
rect 120578 271676 120612 271710
rect 120646 271676 120680 271710
rect 120718 271676 120748 271710
rect 120790 271676 120829 271710
rect 121129 271676 121168 271710
rect 121210 271676 121240 271710
rect 121278 271676 121312 271710
rect 121346 271676 121380 271710
rect 121418 271676 121448 271710
rect 121490 271676 121529 271710
rect 121694 271693 121954 271716
rect 121694 271682 121920 271693
rect 120237 271633 120395 271648
rect 121728 271659 121920 271682
rect 122125 271692 122164 271726
rect 122206 271692 122236 271726
rect 122274 271692 122308 271726
rect 122342 271692 122376 271726
rect 122414 271692 122444 271726
rect 122486 271692 122525 271726
rect 122825 271692 122864 271726
rect 122906 271692 122936 271726
rect 122974 271692 123008 271726
rect 123042 271692 123076 271726
rect 123114 271692 123144 271726
rect 123186 271692 123225 271726
rect 123520 271693 123554 271727
rect 121728 271648 121954 271659
rect 120237 271614 120417 271633
rect 120271 271612 120417 271614
rect 120271 271580 120383 271612
rect 120237 271566 120383 271580
rect 120237 271546 120417 271566
rect 120271 271540 120417 271546
rect 120271 271512 120383 271540
rect 120237 271498 120383 271512
rect 120237 271478 120417 271498
rect 120271 271468 120417 271478
rect 120271 271444 120383 271468
rect 120237 271430 120383 271444
rect 120237 271410 120417 271430
rect 120271 271396 120417 271410
rect 120271 271376 120383 271396
rect 120237 271362 120383 271376
rect 120237 271342 120417 271362
rect 120271 271328 120417 271342
rect 120271 271308 120383 271328
rect 120237 271290 120383 271308
rect 120237 271274 120417 271290
rect 120271 271260 120417 271274
rect 120271 271240 120383 271260
rect 120237 271218 120383 271240
rect 120237 271206 120417 271218
rect 120271 271192 120417 271206
rect 120271 271172 120383 271192
rect 120237 271146 120383 271172
rect 120237 271138 120417 271146
rect 120271 271125 120417 271138
rect 120841 271612 120875 271633
rect 120841 271540 120875 271566
rect 120841 271468 120875 271498
rect 120841 271396 120875 271430
rect 120841 271328 120875 271362
rect 120841 271260 120875 271290
rect 120841 271192 120875 271218
rect 120841 271125 120875 271146
rect 121083 271612 121117 271633
rect 121083 271540 121117 271566
rect 121083 271468 121117 271498
rect 121083 271396 121117 271430
rect 121083 271328 121117 271362
rect 121083 271260 121117 271290
rect 121083 271192 121117 271218
rect 121083 271125 121117 271146
rect 121541 271612 121575 271633
rect 121541 271540 121575 271566
rect 121541 271468 121575 271498
rect 121541 271396 121575 271430
rect 121541 271328 121575 271362
rect 121541 271260 121575 271290
rect 121541 271192 121575 271218
rect 121541 271125 121575 271146
rect 121694 271625 121954 271648
rect 121694 271614 121920 271625
rect 121728 271591 121920 271614
rect 121728 271580 121954 271591
rect 121694 271557 121954 271580
rect 121694 271546 121920 271557
rect 121728 271523 121920 271546
rect 121728 271512 121954 271523
rect 121694 271489 121954 271512
rect 121694 271478 121920 271489
rect 121728 271455 121920 271478
rect 122079 271628 122113 271649
rect 122079 271556 122113 271582
rect 122079 271484 122113 271514
rect 121954 271455 122079 271456
rect 121728 271446 122079 271455
rect 121728 271444 122113 271446
rect 121694 271421 122113 271444
rect 121694 271410 121920 271421
rect 121728 271387 121920 271410
rect 121954 271412 122113 271421
rect 121954 271387 122079 271412
rect 121728 271378 122079 271387
rect 121728 271376 122113 271378
rect 121694 271353 122113 271376
rect 121694 271342 121920 271353
rect 121728 271319 121920 271342
rect 121954 271344 122113 271353
rect 121954 271331 122079 271344
rect 121728 271308 121954 271319
rect 121694 271285 121954 271308
rect 121694 271274 121920 271285
rect 121728 271251 121920 271274
rect 121728 271240 121954 271251
rect 121694 271217 121954 271240
rect 121694 271206 121920 271217
rect 121728 271183 121920 271206
rect 121728 271172 121954 271183
rect 121694 271149 121954 271172
rect 121694 271138 121920 271149
rect 120271 271104 120395 271125
rect 120237 271070 120395 271104
rect 121728 271115 121920 271138
rect 122079 271276 122113 271306
rect 122079 271208 122113 271234
rect 122079 271141 122113 271162
rect 122537 271628 122571 271649
rect 122537 271556 122571 271582
rect 122537 271484 122571 271514
rect 122779 271628 122813 271649
rect 122779 271556 122813 271582
rect 122779 271484 122813 271514
rect 122571 271446 122779 271449
rect 122537 271412 122813 271446
rect 122571 271378 122779 271412
rect 122537 271344 122813 271378
rect 122571 271342 122779 271344
rect 122537 271276 122571 271306
rect 122537 271208 122571 271234
rect 122537 271141 122571 271162
rect 121728 271104 121954 271115
rect 120271 271036 120395 271070
rect 120429 271048 120468 271082
rect 120510 271048 120540 271082
rect 120578 271048 120612 271082
rect 120646 271048 120680 271082
rect 120718 271048 120748 271082
rect 120790 271048 120829 271082
rect 121129 271048 121168 271082
rect 121210 271048 121240 271082
rect 121278 271048 121312 271082
rect 121346 271048 121380 271082
rect 121418 271048 121448 271082
rect 121490 271048 121529 271082
rect 121694 271081 121954 271104
rect 121694 271070 121920 271081
rect 120237 271002 120395 271036
rect 120271 270968 120395 271002
rect 120237 270934 120395 270968
rect 120271 270900 120395 270934
rect 121728 271047 121920 271070
rect 122125 271064 122164 271098
rect 122206 271064 122236 271098
rect 122274 271064 122308 271098
rect 122342 271064 122376 271098
rect 122414 271064 122444 271098
rect 122486 271064 122525 271098
rect 121728 271036 121954 271047
rect 121694 271013 121954 271036
rect 121694 271002 121920 271013
rect 121728 270979 121920 271002
rect 121728 270968 121954 270979
rect 121694 270945 121954 270968
rect 121694 270934 121920 270945
rect 120237 270866 120395 270900
rect 120429 270892 120468 270926
rect 120510 270892 120540 270926
rect 120578 270892 120612 270926
rect 120646 270892 120680 270926
rect 120718 270892 120748 270926
rect 120790 270892 120829 270926
rect 121129 270892 121168 270926
rect 121210 270892 121240 270926
rect 121278 270892 121312 270926
rect 121346 270892 121380 270926
rect 121418 270892 121448 270926
rect 121490 270892 121529 270926
rect 121728 270911 121920 270934
rect 121728 270900 121954 270911
rect 122125 270908 122164 270942
rect 122206 270908 122236 270942
rect 122274 270908 122308 270942
rect 122342 270908 122376 270942
rect 122414 270908 122444 270942
rect 122486 270908 122525 270942
rect 120271 270849 120395 270866
rect 121694 270877 121954 270900
rect 121694 270866 121920 270877
rect 120271 270832 120417 270849
rect 120237 270828 120417 270832
rect 120237 270798 120383 270828
rect 120271 270782 120383 270798
rect 120271 270764 120417 270782
rect 120237 270756 120417 270764
rect 120237 270730 120383 270756
rect 120271 270714 120383 270730
rect 120271 270696 120417 270714
rect 120237 270684 120417 270696
rect 120237 270662 120383 270684
rect 120271 270646 120383 270662
rect 120271 270628 120417 270646
rect 120237 270612 120417 270628
rect 120237 270594 120383 270612
rect 120271 270578 120383 270594
rect 120271 270560 120417 270578
rect 120237 270544 120417 270560
rect 120237 270526 120383 270544
rect 120271 270506 120383 270526
rect 120271 270492 120417 270506
rect 120237 270476 120417 270492
rect 120237 270458 120383 270476
rect 120271 270434 120383 270458
rect 120271 270424 120417 270434
rect 120237 270408 120417 270424
rect 120237 270390 120383 270408
rect 120271 270362 120383 270390
rect 120271 270356 120417 270362
rect 120237 270341 120417 270356
rect 120841 270828 120875 270849
rect 120841 270756 120875 270782
rect 120841 270684 120875 270714
rect 120841 270612 120875 270646
rect 120841 270544 120875 270578
rect 120841 270476 120875 270506
rect 120841 270408 120875 270434
rect 120841 270341 120875 270362
rect 121083 270828 121117 270849
rect 121083 270756 121117 270782
rect 121083 270684 121117 270714
rect 121083 270612 121117 270646
rect 121083 270544 121117 270578
rect 121083 270476 121117 270506
rect 121083 270408 121117 270434
rect 121083 270341 121117 270362
rect 121541 270828 121575 270849
rect 121541 270756 121575 270782
rect 121541 270684 121575 270714
rect 121541 270612 121575 270646
rect 121541 270544 121575 270578
rect 121541 270476 121575 270506
rect 121541 270408 121575 270434
rect 121541 270341 121575 270362
rect 121728 270843 121920 270866
rect 121728 270832 121954 270843
rect 121694 270809 121954 270832
rect 121694 270798 121920 270809
rect 121728 270775 121920 270798
rect 121728 270764 121954 270775
rect 121694 270741 121954 270764
rect 121694 270730 121920 270741
rect 121728 270707 121920 270730
rect 121728 270696 121954 270707
rect 121694 270673 121954 270696
rect 121694 270662 121920 270673
rect 121728 270639 121920 270662
rect 122079 270844 122113 270865
rect 122079 270772 122113 270798
rect 122079 270700 122113 270730
rect 121954 270662 122079 270672
rect 121954 270639 122113 270662
rect 121728 270628 122113 270639
rect 121694 270605 122079 270628
rect 121694 270594 121920 270605
rect 121728 270571 121920 270594
rect 121954 270594 122079 270605
rect 121954 270571 122113 270594
rect 121728 270560 122113 270571
rect 121694 270547 122079 270560
rect 121694 270537 121954 270547
rect 121694 270526 121920 270537
rect 121728 270503 121920 270526
rect 121728 270492 121954 270503
rect 121694 270469 121954 270492
rect 121694 270458 121920 270469
rect 121728 270435 121920 270458
rect 121728 270424 121954 270435
rect 121694 270401 121954 270424
rect 121694 270390 121920 270401
rect 121728 270367 121920 270390
rect 121728 270356 121954 270367
rect 122079 270492 122113 270522
rect 122079 270424 122113 270450
rect 122079 270357 122113 270378
rect 122537 270844 122571 270865
rect 122537 270772 122571 270798
rect 122537 270700 122571 270730
rect 122639 270675 122735 271342
rect 122779 271276 122813 271306
rect 122779 271208 122813 271234
rect 122779 271141 122813 271162
rect 123237 271628 123271 271649
rect 123237 271556 123271 271582
rect 123237 271484 123271 271514
rect 123237 271412 123271 271446
rect 123237 271344 123271 271378
rect 123237 271276 123271 271306
rect 123237 271208 123271 271234
rect 123237 271141 123271 271162
rect 123520 271625 123554 271659
rect 123520 271557 123554 271591
rect 123520 271489 123554 271523
rect 123520 271421 123554 271455
rect 123520 271353 123554 271387
rect 123520 271285 123554 271319
rect 123520 271217 123554 271251
rect 123520 271149 123554 271183
rect 122825 271064 122864 271098
rect 122906 271064 122936 271098
rect 122974 271064 123008 271098
rect 123042 271064 123076 271098
rect 123114 271064 123144 271098
rect 123186 271064 123225 271098
rect 123520 271081 123554 271115
rect 123520 271013 123554 271047
rect 123520 270945 123554 270979
rect 122825 270908 122864 270942
rect 122906 270908 122936 270942
rect 122974 270908 123008 270942
rect 123042 270908 123076 270942
rect 123114 270908 123144 270942
rect 123186 270908 123225 270942
rect 123520 270877 123554 270911
rect 122779 270844 122813 270865
rect 122779 270772 122813 270798
rect 122779 270700 122813 270730
rect 122571 270662 122779 270675
rect 122537 270628 122813 270662
rect 122571 270594 122779 270628
rect 122537 270568 122813 270594
rect 122537 270560 122571 270568
rect 122537 270492 122571 270522
rect 122537 270424 122571 270450
rect 122537 270357 122571 270378
rect 122779 270560 122813 270568
rect 122779 270492 122813 270522
rect 122779 270424 122813 270450
rect 122779 270357 122813 270378
rect 123237 270844 123271 270865
rect 123237 270772 123271 270798
rect 123237 270700 123271 270730
rect 123237 270628 123271 270662
rect 123237 270560 123271 270594
rect 123237 270492 123271 270522
rect 123237 270424 123271 270450
rect 123237 270357 123271 270378
rect 123520 270809 123554 270843
rect 123520 270741 123554 270775
rect 123520 270673 123554 270707
rect 123520 270605 123554 270639
rect 123520 270537 123554 270571
rect 123520 270469 123554 270503
rect 123520 270401 123554 270435
rect 120237 270322 120395 270341
rect 120271 270288 120395 270322
rect 121694 270333 121954 270356
rect 121694 270322 121920 270333
rect 120237 270254 120395 270288
rect 120429 270264 120468 270298
rect 120510 270264 120540 270298
rect 120578 270264 120612 270298
rect 120646 270264 120680 270298
rect 120718 270264 120748 270298
rect 120790 270264 120829 270298
rect 121129 270264 121168 270298
rect 121210 270264 121240 270298
rect 121278 270264 121312 270298
rect 121346 270264 121380 270298
rect 121418 270264 121448 270298
rect 121490 270264 121529 270298
rect 121728 270299 121920 270322
rect 123520 270333 123554 270367
rect 121728 270288 121954 270299
rect 121694 270265 121954 270288
rect 122125 270280 122164 270314
rect 122206 270280 122236 270314
rect 122274 270280 122308 270314
rect 122342 270280 122376 270314
rect 122414 270280 122444 270314
rect 122486 270280 122525 270314
rect 122825 270280 122864 270314
rect 122906 270280 122936 270314
rect 122974 270280 123008 270314
rect 123042 270280 123076 270314
rect 123114 270280 123144 270314
rect 123186 270280 123225 270314
rect 120271 270220 120395 270254
rect 120237 270186 120395 270220
rect 120271 270152 120395 270186
rect 120237 270118 120395 270152
rect 121694 270254 121920 270265
rect 121728 270231 121920 270254
rect 121728 270220 121954 270231
rect 121694 270197 121954 270220
rect 121694 270186 121920 270197
rect 121728 270163 121920 270186
rect 121728 270152 121954 270163
rect 123520 270265 123554 270299
rect 123520 270197 123554 270231
rect 120271 270084 120395 270118
rect 120429 270108 120468 270142
rect 120510 270108 120540 270142
rect 120578 270108 120612 270142
rect 120646 270108 120680 270142
rect 120718 270108 120748 270142
rect 120790 270108 120829 270142
rect 121129 270108 121168 270142
rect 121210 270108 121240 270142
rect 121278 270108 121312 270142
rect 121346 270108 121380 270142
rect 121418 270108 121448 270142
rect 121490 270108 121529 270142
rect 121694 270129 121954 270152
rect 121694 270118 121920 270129
rect 120237 270065 120395 270084
rect 121728 270095 121920 270118
rect 122125 270124 122164 270158
rect 122206 270124 122236 270158
rect 122274 270124 122308 270158
rect 122342 270124 122376 270158
rect 122414 270124 122444 270158
rect 122486 270124 122525 270158
rect 122825 270124 122864 270158
rect 122906 270124 122936 270158
rect 122974 270124 123008 270158
rect 123042 270124 123076 270158
rect 123114 270124 123144 270158
rect 123186 270124 123351 270158
rect 121728 270084 121954 270095
rect 120237 270050 120417 270065
rect 120271 270044 120417 270050
rect 120271 270016 120383 270044
rect 120237 269998 120383 270016
rect 120237 269982 120417 269998
rect 120271 269972 120417 269982
rect 120271 269948 120383 269972
rect 120237 269930 120383 269948
rect 120237 269914 120417 269930
rect 120271 269900 120417 269914
rect 120271 269880 120383 269900
rect 120237 269862 120383 269880
rect 120237 269846 120417 269862
rect 120271 269828 120417 269846
rect 120271 269812 120383 269828
rect 120237 269794 120383 269812
rect 120237 269778 120417 269794
rect 120271 269760 120417 269778
rect 120271 269744 120383 269760
rect 120237 269722 120383 269744
rect 120237 269710 120417 269722
rect 120271 269692 120417 269710
rect 120271 269676 120383 269692
rect 120237 269650 120383 269676
rect 120237 269642 120417 269650
rect 120271 269624 120417 269642
rect 120271 269608 120383 269624
rect 120237 269578 120383 269608
rect 120237 269574 120417 269578
rect 120271 269557 120417 269574
rect 120841 270044 120875 270065
rect 120841 269972 120875 269998
rect 120841 269900 120875 269930
rect 120841 269828 120875 269862
rect 120841 269760 120875 269794
rect 120841 269692 120875 269722
rect 120841 269624 120875 269650
rect 120841 269557 120875 269578
rect 121083 270044 121117 270065
rect 121083 269972 121117 269998
rect 121083 269900 121117 269930
rect 121083 269828 121117 269862
rect 121083 269760 121117 269794
rect 121083 269692 121117 269722
rect 121083 269624 121117 269650
rect 121083 269557 121117 269578
rect 121541 270044 121575 270065
rect 121541 269972 121575 269998
rect 121541 269900 121575 269930
rect 121541 269828 121575 269862
rect 121541 269760 121575 269794
rect 121541 269692 121575 269722
rect 121541 269624 121575 269650
rect 121541 269557 121575 269578
rect 121694 270061 121954 270084
rect 121694 270050 121920 270061
rect 121728 270027 121920 270050
rect 121728 270016 121954 270027
rect 121694 269993 121954 270016
rect 121694 269982 121920 269993
rect 121728 269959 121920 269982
rect 121728 269948 121954 269959
rect 121694 269925 121954 269948
rect 121694 269914 121920 269925
rect 121728 269891 121920 269914
rect 121728 269882 121954 269891
rect 122079 270060 122113 270081
rect 122079 269988 122113 270014
rect 122079 269916 122113 269946
rect 121728 269880 122079 269882
rect 121694 269878 122079 269880
rect 121694 269857 122113 269878
rect 121694 269846 121920 269857
rect 121728 269823 121920 269846
rect 121954 269844 122113 269857
rect 121954 269823 122079 269844
rect 121728 269812 122079 269823
rect 121694 269810 122079 269812
rect 121694 269789 122113 269810
rect 121694 269778 121920 269789
rect 121728 269755 121920 269778
rect 121954 269776 122113 269789
rect 121954 269757 122079 269776
rect 121728 269744 121954 269755
rect 121694 269721 121954 269744
rect 121694 269710 121920 269721
rect 121728 269687 121920 269710
rect 121728 269676 121954 269687
rect 121694 269653 121954 269676
rect 121694 269642 121920 269653
rect 121728 269619 121920 269642
rect 121728 269608 121954 269619
rect 121694 269585 121954 269608
rect 121694 269574 121920 269585
rect 120271 269540 120395 269557
rect 120237 269506 120395 269540
rect 121728 269551 121920 269574
rect 122079 269708 122113 269738
rect 122079 269640 122113 269666
rect 122079 269573 122113 269594
rect 122537 270060 122571 270081
rect 122537 269988 122571 270014
rect 122537 269916 122571 269946
rect 122537 269874 122571 269878
rect 122779 270060 122813 270081
rect 122779 269988 122813 270014
rect 122779 269916 122813 269946
rect 122779 269874 122813 269878
rect 122537 269844 122813 269874
rect 122571 269837 122779 269844
rect 122571 269810 122668 269837
rect 122537 269803 122668 269810
rect 122702 269810 122779 269837
rect 122702 269803 122813 269810
rect 122537 269776 122813 269803
rect 122571 269767 122779 269776
rect 122537 269708 122571 269738
rect 122537 269640 122571 269666
rect 122537 269573 122571 269594
rect 122779 269708 122813 269738
rect 122779 269640 122813 269666
rect 122779 269573 122813 269594
rect 123237 270060 123271 270081
rect 123237 269988 123271 270014
rect 123237 269916 123271 269946
rect 123237 269844 123271 269878
rect 123237 269776 123271 269810
rect 123237 269708 123271 269738
rect 123237 269640 123271 269666
rect 123237 269573 123271 269594
rect 121728 269540 121954 269551
rect 121694 269517 121954 269540
rect 123317 269530 123351 270124
rect 120271 269472 120395 269506
rect 120429 269480 120468 269514
rect 120510 269480 120540 269514
rect 120578 269480 120612 269514
rect 120646 269480 120680 269514
rect 120718 269480 120748 269514
rect 120790 269480 120829 269514
rect 121129 269480 121168 269514
rect 121210 269480 121240 269514
rect 121278 269480 121312 269514
rect 121346 269480 121380 269514
rect 121418 269480 121448 269514
rect 121490 269480 121529 269514
rect 121694 269506 121920 269517
rect 120237 269438 120395 269472
rect 120271 269404 120395 269438
rect 120237 269370 120395 269404
rect 120271 269336 120395 269370
rect 121728 269483 121920 269506
rect 122125 269496 122164 269530
rect 122206 269496 122236 269530
rect 122274 269496 122308 269530
rect 122342 269496 122376 269530
rect 122414 269496 122444 269530
rect 122486 269496 122525 269530
rect 122825 269496 122864 269530
rect 122906 269496 122936 269530
rect 122974 269496 123008 269530
rect 123042 269496 123076 269530
rect 123114 269496 123144 269530
rect 123186 269496 123351 269530
rect 123520 270129 123554 270163
rect 123520 270061 123554 270095
rect 123520 269993 123554 270027
rect 123520 269925 123554 269959
rect 123520 269857 123554 269891
rect 123520 269789 123554 269823
rect 123520 269721 123554 269755
rect 123520 269653 123554 269687
rect 123520 269585 123554 269619
rect 123520 269517 123554 269551
rect 121728 269472 121954 269483
rect 121694 269449 121954 269472
rect 121694 269438 121920 269449
rect 121728 269415 121920 269438
rect 121728 269404 121954 269415
rect 121694 269381 121954 269404
rect 121694 269370 121920 269381
rect 120237 269302 120395 269336
rect 120429 269324 120468 269358
rect 120510 269324 120540 269358
rect 120578 269324 120612 269358
rect 120646 269324 120680 269358
rect 120718 269324 120748 269358
rect 120790 269324 120829 269358
rect 121129 269324 121168 269358
rect 121210 269324 121240 269358
rect 121278 269324 121312 269358
rect 121346 269324 121380 269358
rect 121418 269324 121448 269358
rect 121490 269324 121529 269358
rect 121728 269347 121920 269370
rect 123520 269449 123554 269483
rect 123520 269381 123554 269415
rect 121728 269336 121954 269347
rect 120271 269281 120395 269302
rect 121694 269313 121954 269336
rect 121694 269302 121920 269313
rect 120271 269268 120417 269281
rect 120237 269244 120417 269268
rect 120237 269234 120383 269244
rect 120271 269210 120383 269234
rect 120271 269200 120417 269210
rect 120237 269173 120417 269200
rect 120841 269244 120875 269281
rect 120841 269173 120875 269210
rect 120237 269166 120429 269173
rect 120271 269132 120429 269166
rect 120237 269130 120429 269132
rect 120829 269130 120875 269173
rect 120237 269098 120468 269130
rect 120271 269096 120468 269098
rect 120510 269096 120540 269130
rect 120578 269096 120612 269130
rect 120646 269096 120680 269130
rect 120718 269096 120748 269130
rect 120790 269114 120875 269130
rect 121083 269244 121117 269281
rect 121083 269173 121117 269210
rect 121541 269244 121575 269281
rect 121541 269173 121575 269210
rect 121083 269130 121129 269173
rect 121529 269130 121575 269173
rect 121083 269114 121168 269130
rect 120790 269096 121168 269114
rect 121210 269096 121240 269130
rect 121278 269096 121312 269130
rect 121346 269096 121380 269130
rect 121418 269096 121448 269130
rect 121490 269114 121575 269130
rect 121728 269279 121920 269302
rect 121728 269268 121954 269279
rect 121694 269245 121954 269268
rect 121694 269234 121920 269245
rect 121728 269211 121920 269234
rect 121728 269200 121954 269211
rect 121694 269177 121954 269200
rect 121694 269166 121920 269177
rect 121728 269143 121920 269166
rect 121728 269132 121954 269143
rect 121694 269114 121954 269132
rect 121490 269109 121954 269114
rect 121490 269098 121920 269109
rect 121490 269096 121694 269098
rect 120271 269064 121694 269096
rect 121728 269075 121920 269098
rect 121728 269066 121954 269075
rect 122079 269340 122164 269374
rect 122206 269340 122236 269374
rect 122274 269340 122308 269374
rect 122342 269340 122376 269374
rect 122414 269340 122444 269374
rect 122486 269340 122571 269374
rect 122079 269260 122125 269340
rect 122113 269226 122125 269260
rect 122079 269146 122125 269226
rect 122525 269260 122571 269340
rect 122525 269226 122537 269260
rect 122525 269146 122571 269226
rect 122079 269112 122164 269146
rect 122206 269112 122236 269146
rect 122274 269112 122308 269146
rect 122342 269112 122376 269146
rect 122414 269112 122444 269146
rect 122486 269112 122571 269146
rect 122079 269066 122571 269112
rect 122779 269340 122864 269374
rect 122906 269340 122936 269374
rect 122974 269340 123008 269374
rect 123042 269340 123076 269374
rect 123114 269340 123144 269374
rect 123186 269340 123271 269374
rect 122779 269260 122825 269340
rect 122813 269226 122825 269260
rect 122779 269146 122825 269226
rect 123225 269260 123271 269340
rect 123225 269226 123237 269260
rect 123225 269146 123271 269226
rect 122779 269112 122864 269146
rect 122906 269112 122936 269146
rect 122974 269112 123008 269146
rect 123042 269112 123076 269146
rect 123114 269112 123144 269146
rect 123186 269112 123271 269146
rect 122779 269066 123271 269112
rect 123520 269313 123554 269347
rect 123520 269245 123554 269279
rect 123520 269177 123554 269211
rect 123520 269109 123554 269143
rect 123520 269066 123554 269075
rect 121728 269064 123554 269066
rect 120237 269028 123554 269064
rect 120237 269012 122006 269028
rect 120237 268978 120319 269012
rect 120353 268978 120387 269012
rect 120421 268978 120455 269012
rect 120489 268978 120523 269012
rect 120557 268978 120591 269012
rect 120625 268978 120659 269012
rect 120693 268978 120727 269012
rect 120761 268978 120795 269012
rect 120829 268978 120863 269012
rect 120897 268978 120931 269012
rect 120965 268978 120999 269012
rect 121033 268978 121067 269012
rect 121101 268978 121135 269012
rect 121169 268978 121203 269012
rect 121237 268978 121271 269012
rect 121305 268978 121339 269012
rect 121373 268978 121407 269012
rect 121441 268978 121475 269012
rect 121509 268978 121543 269012
rect 121577 268978 121611 269012
rect 121645 268994 122006 269012
rect 122040 268994 122074 269028
rect 122108 268994 122142 269028
rect 122176 268994 122210 269028
rect 122244 268994 122278 269028
rect 122312 268994 122346 269028
rect 122380 268994 122414 269028
rect 122448 268994 122482 269028
rect 122516 268994 122550 269028
rect 122584 268994 122618 269028
rect 122652 268994 122686 269028
rect 122720 268994 122754 269028
rect 122788 268994 122822 269028
rect 122856 268994 122890 269028
rect 122924 268994 122958 269028
rect 122992 268994 123026 269028
rect 123060 268994 123094 269028
rect 123128 268994 123162 269028
rect 123196 268994 123230 269028
rect 123264 268994 123298 269028
rect 123332 268994 123366 269028
rect 123400 268994 123434 269028
rect 123468 268994 123554 269028
rect 123827 272777 124279 273545
rect 123827 272770 124768 272777
rect 125047 272770 125058 273545
rect 123827 272750 125058 272770
rect 123827 272716 124065 272750
rect 124099 272716 124133 272750
rect 124167 272716 124201 272750
rect 124235 272716 124269 272750
rect 124303 272716 124337 272750
rect 124371 272716 124405 272750
rect 124439 272716 124473 272750
rect 124507 272716 124541 272750
rect 124575 272716 124609 272750
rect 124643 272716 124677 272750
rect 124711 272716 125058 272750
rect 123827 272689 125058 272716
rect 123827 272592 124029 272689
rect 123827 272558 123986 272592
rect 124020 272558 124029 272592
rect 123827 272524 124029 272558
rect 123827 272490 123986 272524
rect 124020 272490 124029 272524
rect 123827 272456 124029 272490
rect 123827 272422 123986 272456
rect 124020 272422 124029 272456
rect 123827 272388 124029 272422
rect 123827 272354 123986 272388
rect 124020 272354 124029 272388
rect 123827 272320 124029 272354
rect 123827 272286 123986 272320
rect 124020 272286 124029 272320
rect 123827 272252 124029 272286
rect 124116 272601 124188 272689
rect 124696 272687 125058 272689
rect 124696 272653 124828 272687
rect 124862 272653 125058 272687
rect 124696 272619 125058 272653
rect 124696 272601 124828 272619
rect 124116 272585 124828 272601
rect 124862 272585 125058 272619
rect 124116 272580 125058 272585
rect 124116 272566 124880 272580
rect 124116 272532 124209 272566
rect 124255 272532 124281 272566
rect 124323 272532 124353 272566
rect 124391 272532 124425 272566
rect 124459 272532 124493 272566
rect 124531 272532 124561 272566
rect 124603 272532 124629 272566
rect 124675 272532 124768 272566
rect 124116 272473 124188 272532
rect 124116 272437 124120 272473
rect 124154 272437 124188 272473
rect 124116 272403 124188 272437
rect 124116 272367 124120 272403
rect 124154 272367 124188 272403
rect 124116 272308 124188 272367
rect 124696 272473 124768 272532
rect 124696 272437 124730 272473
rect 124764 272437 124768 272473
rect 124696 272403 124768 272437
rect 124696 272367 124730 272403
rect 124764 272367 124768 272403
rect 124696 272308 124768 272367
rect 124116 272274 124209 272308
rect 124255 272274 124281 272308
rect 124323 272274 124353 272308
rect 124391 272274 124425 272308
rect 124459 272274 124493 272308
rect 124531 272274 124561 272308
rect 124603 272274 124629 272308
rect 124675 272274 124768 272308
rect 124811 272551 124880 272566
rect 124811 272517 124828 272551
rect 124862 272517 124880 272551
rect 124811 272483 124880 272517
rect 124811 272449 124828 272483
rect 124862 272449 124880 272483
rect 124811 272415 124880 272449
rect 124811 272381 124828 272415
rect 124862 272381 124880 272415
rect 124811 272347 124880 272381
rect 124811 272313 124828 272347
rect 124862 272313 124880 272347
rect 124811 272279 124880 272313
rect 123827 272218 123986 272252
rect 124020 272218 124029 272252
rect 123827 272184 124029 272218
rect 124811 272245 124828 272279
rect 124862 272245 124880 272279
rect 124811 272211 124880 272245
rect 124811 272185 124828 272211
rect 123827 272150 123986 272184
rect 124020 272150 124029 272184
rect 123827 272116 124029 272150
rect 124188 272177 124828 272185
rect 124862 272177 124880 272211
rect 124188 272150 124880 272177
rect 124188 272116 124209 272150
rect 124255 272116 124281 272150
rect 124323 272116 124353 272150
rect 124391 272116 124425 272150
rect 124459 272116 124493 272150
rect 124531 272116 124561 272150
rect 124603 272116 124629 272150
rect 124675 272116 124696 272150
rect 124811 272143 124880 272150
rect 123827 272082 123986 272116
rect 124020 272082 124029 272116
rect 124811 272109 124828 272143
rect 124862 272109 124880 272143
rect 123827 272048 124029 272082
rect 123827 272014 123986 272048
rect 124020 272014 124029 272048
rect 123827 271980 124029 272014
rect 123827 271946 123986 271980
rect 124020 271946 124029 271980
rect 123827 271912 124029 271946
rect 123827 271878 123986 271912
rect 124020 271878 124029 271912
rect 123827 271844 124029 271878
rect 123827 271810 123986 271844
rect 124020 271810 124029 271844
rect 123827 271776 124029 271810
rect 123827 271742 123986 271776
rect 124020 271742 124029 271776
rect 123827 271708 124029 271742
rect 123827 271674 123986 271708
rect 124020 271674 124029 271708
rect 123827 271640 124029 271674
rect 123827 271606 123986 271640
rect 124020 271606 124029 271640
rect 123827 271572 124029 271606
rect 123827 271538 123986 271572
rect 124020 271538 124029 271572
rect 123827 271504 124029 271538
rect 123827 271470 123986 271504
rect 124020 271470 124029 271504
rect 123827 271436 124029 271470
rect 123827 271402 123986 271436
rect 124020 271402 124029 271436
rect 123827 271368 124029 271402
rect 123827 271334 123986 271368
rect 124020 271334 124029 271368
rect 123827 271300 124029 271334
rect 123827 271266 123986 271300
rect 124020 271266 124029 271300
rect 123827 271232 124029 271266
rect 123827 271198 123986 271232
rect 124020 271198 124029 271232
rect 123827 271164 124029 271198
rect 123827 271130 123986 271164
rect 124020 271130 124029 271164
rect 123827 271096 124029 271130
rect 123827 271062 123986 271096
rect 124020 271062 124029 271096
rect 123827 271028 124029 271062
rect 123827 270994 123986 271028
rect 124020 270994 124029 271028
rect 123827 270960 124029 270994
rect 123827 270926 123986 270960
rect 124020 270926 124029 270960
rect 123827 270892 124029 270926
rect 123827 270858 123986 270892
rect 124020 270858 124029 270892
rect 123827 270824 124029 270858
rect 123827 270790 123986 270824
rect 124020 270790 124029 270824
rect 123827 270756 124029 270790
rect 123827 270722 123986 270756
rect 124020 270722 124029 270756
rect 123827 270688 124029 270722
rect 123827 270654 123986 270688
rect 124020 270654 124029 270688
rect 123827 270620 124029 270654
rect 123827 270586 123986 270620
rect 124020 270586 124029 270620
rect 123827 270552 124029 270586
rect 123827 270518 123986 270552
rect 124020 270518 124029 270552
rect 123827 270484 124029 270518
rect 123827 270450 123986 270484
rect 124020 270450 124029 270484
rect 123827 270416 124029 270450
rect 123827 270382 123986 270416
rect 124020 270382 124029 270416
rect 123827 270348 124029 270382
rect 123827 270314 123986 270348
rect 124020 270314 124029 270348
rect 123827 270280 124029 270314
rect 123827 270246 123986 270280
rect 124020 270246 124029 270280
rect 123827 270212 124029 270246
rect 123827 270178 123986 270212
rect 124020 270178 124029 270212
rect 123827 270144 124029 270178
rect 123827 270110 123986 270144
rect 124020 270110 124029 270144
rect 123827 270076 124029 270110
rect 123827 270042 123986 270076
rect 124020 270042 124029 270076
rect 123827 270008 124029 270042
rect 123827 269974 123986 270008
rect 124020 269974 124029 270008
rect 123827 269940 124029 269974
rect 123827 269906 123986 269940
rect 124020 269906 124029 269940
rect 123827 269872 124029 269906
rect 123827 269838 123986 269872
rect 124020 269838 124029 269872
rect 123827 269804 124029 269838
rect 124084 272057 124154 272104
rect 124084 272021 124120 272057
rect 124084 271987 124154 272021
rect 124084 271951 124120 271987
rect 124084 271904 124154 271951
rect 124730 272057 124764 272104
rect 124730 271987 124764 272021
rect 124730 271904 124764 271951
rect 124811 272075 124880 272109
rect 124811 272041 124828 272075
rect 124862 272041 124880 272075
rect 124811 272007 124880 272041
rect 124811 271973 124828 272007
rect 124862 271973 124880 272007
rect 124811 271939 124880 271973
rect 124811 271905 124828 271939
rect 124862 271905 124880 271939
rect 124084 271688 124120 271904
rect 124188 271858 124209 271892
rect 124255 271858 124281 271892
rect 124323 271858 124353 271892
rect 124391 271858 124425 271892
rect 124459 271858 124493 271892
rect 124531 271858 124561 271892
rect 124603 271858 124629 271892
rect 124675 271858 124696 271892
rect 124811 271871 124880 271905
rect 124811 271837 124828 271871
rect 124862 271837 124880 271871
rect 124811 271803 124880 271837
rect 124811 271769 124828 271803
rect 124862 271769 124880 271803
rect 124188 271735 124880 271769
rect 124188 271734 124828 271735
rect 124188 271700 124209 271734
rect 124255 271700 124281 271734
rect 124323 271700 124353 271734
rect 124391 271700 124425 271734
rect 124459 271700 124493 271734
rect 124531 271700 124561 271734
rect 124603 271700 124629 271734
rect 124675 271700 124696 271734
rect 124811 271701 124828 271734
rect 124862 271701 124880 271735
rect 124084 271641 124154 271688
rect 124084 271605 124120 271641
rect 124084 271571 124154 271605
rect 124084 271535 124120 271571
rect 124084 271488 124154 271535
rect 124730 271641 124764 271688
rect 124730 271571 124764 271605
rect 124730 271488 124764 271535
rect 124811 271667 124880 271701
rect 124811 271633 124828 271667
rect 124862 271633 124880 271667
rect 124811 271599 124880 271633
rect 124811 271565 124828 271599
rect 124862 271565 124880 271599
rect 124811 271531 124880 271565
rect 124811 271497 124828 271531
rect 124862 271497 124880 271531
rect 124084 271272 124120 271488
rect 124188 271442 124209 271476
rect 124255 271442 124281 271476
rect 124323 271442 124353 271476
rect 124391 271442 124425 271476
rect 124459 271442 124493 271476
rect 124531 271442 124561 271476
rect 124603 271442 124629 271476
rect 124675 271442 124696 271476
rect 124811 271463 124880 271497
rect 124811 271429 124828 271463
rect 124862 271429 124880 271463
rect 124811 271395 124880 271429
rect 124811 271361 124828 271395
rect 124862 271361 124880 271395
rect 124811 271353 124880 271361
rect 124188 271327 124880 271353
rect 124188 271318 124828 271327
rect 124188 271284 124209 271318
rect 124255 271284 124281 271318
rect 124323 271284 124353 271318
rect 124391 271284 124425 271318
rect 124459 271284 124493 271318
rect 124531 271284 124561 271318
rect 124603 271284 124629 271318
rect 124675 271284 124696 271318
rect 124811 271293 124828 271318
rect 124862 271293 124880 271327
rect 124084 271225 124154 271272
rect 124084 271189 124120 271225
rect 124084 271155 124154 271189
rect 124084 271119 124120 271155
rect 124084 271072 124154 271119
rect 124730 271225 124764 271272
rect 124730 271155 124764 271189
rect 124730 271072 124764 271119
rect 124811 271259 124880 271293
rect 124811 271225 124828 271259
rect 124862 271225 124880 271259
rect 124811 271191 124880 271225
rect 124811 271157 124828 271191
rect 124862 271157 124880 271191
rect 124811 271123 124880 271157
rect 124811 271089 124828 271123
rect 124862 271089 124880 271123
rect 124084 270856 124120 271072
rect 124188 271026 124209 271060
rect 124255 271026 124281 271060
rect 124323 271026 124353 271060
rect 124391 271026 124425 271060
rect 124459 271026 124493 271060
rect 124531 271026 124561 271060
rect 124603 271026 124629 271060
rect 124675 271026 124696 271060
rect 124811 271055 124880 271089
rect 124811 271021 124828 271055
rect 124862 271021 124880 271055
rect 124811 270987 124880 271021
rect 124811 270953 124828 270987
rect 124862 270953 124880 270987
rect 124811 270937 124880 270953
rect 124188 270919 124880 270937
rect 124188 270902 124828 270919
rect 124188 270868 124209 270902
rect 124255 270868 124281 270902
rect 124323 270868 124353 270902
rect 124391 270868 124425 270902
rect 124459 270868 124493 270902
rect 124531 270868 124561 270902
rect 124603 270868 124629 270902
rect 124675 270868 124696 270902
rect 124811 270885 124828 270902
rect 124862 270885 124880 270919
rect 124084 270809 124154 270856
rect 124084 270773 124120 270809
rect 124084 270739 124154 270773
rect 124084 270703 124120 270739
rect 124084 270656 124154 270703
rect 124730 270809 124764 270856
rect 124730 270739 124764 270773
rect 124730 270656 124764 270703
rect 124811 270851 124880 270885
rect 124811 270817 124828 270851
rect 124862 270817 124880 270851
rect 124811 270783 124880 270817
rect 124811 270749 124828 270783
rect 124862 270749 124880 270783
rect 124811 270715 124880 270749
rect 124811 270681 124828 270715
rect 124862 270681 124880 270715
rect 124084 270440 124120 270656
rect 124811 270647 124880 270681
rect 124188 270610 124209 270644
rect 124255 270610 124281 270644
rect 124323 270610 124353 270644
rect 124391 270610 124425 270644
rect 124459 270610 124493 270644
rect 124531 270610 124561 270644
rect 124603 270610 124629 270644
rect 124675 270610 124696 270644
rect 124811 270613 124828 270647
rect 124862 270613 124880 270647
rect 124811 270579 124880 270613
rect 124811 270545 124828 270579
rect 124862 270545 124880 270579
rect 124811 270521 124880 270545
rect 124188 270511 124880 270521
rect 124188 270486 124828 270511
rect 124188 270452 124209 270486
rect 124255 270452 124281 270486
rect 124323 270452 124353 270486
rect 124391 270452 124425 270486
rect 124459 270452 124493 270486
rect 124531 270452 124561 270486
rect 124603 270452 124629 270486
rect 124675 270452 124696 270486
rect 124811 270477 124828 270486
rect 124862 270477 124880 270511
rect 124811 270443 124880 270477
rect 124084 270393 124154 270440
rect 124084 270357 124120 270393
rect 124084 270323 124154 270357
rect 124084 270287 124120 270323
rect 124084 270240 124154 270287
rect 124730 270393 124764 270440
rect 124730 270323 124764 270357
rect 124730 270240 124764 270287
rect 124811 270409 124828 270443
rect 124862 270409 124880 270443
rect 124811 270375 124880 270409
rect 124811 270341 124828 270375
rect 124862 270341 124880 270375
rect 124811 270307 124880 270341
rect 124811 270273 124828 270307
rect 124862 270273 124880 270307
rect 124084 270024 124120 270240
rect 124811 270239 124880 270273
rect 124188 270194 124209 270228
rect 124255 270194 124281 270228
rect 124323 270194 124353 270228
rect 124391 270194 124425 270228
rect 124459 270194 124493 270228
rect 124531 270194 124561 270228
rect 124603 270194 124629 270228
rect 124675 270194 124696 270228
rect 124811 270205 124828 270239
rect 124862 270205 124880 270239
rect 124811 270171 124880 270205
rect 124811 270137 124828 270171
rect 124862 270137 124880 270171
rect 124811 270105 124880 270137
rect 124188 270103 124880 270105
rect 124188 270070 124828 270103
rect 124188 270036 124209 270070
rect 124255 270036 124281 270070
rect 124323 270036 124353 270070
rect 124391 270036 124425 270070
rect 124459 270036 124493 270070
rect 124531 270036 124561 270070
rect 124603 270036 124629 270070
rect 124675 270036 124696 270070
rect 124811 270069 124828 270070
rect 124862 270069 124880 270103
rect 124811 270035 124880 270069
rect 124084 269977 124154 270024
rect 124084 269941 124120 269977
rect 124084 269907 124154 269941
rect 124084 269871 124120 269907
rect 124084 269824 124154 269871
rect 124730 269977 124764 270024
rect 124730 269907 124764 269941
rect 124730 269824 124764 269871
rect 124811 270001 124828 270035
rect 124862 270001 124880 270035
rect 124811 269967 124880 270001
rect 124811 269933 124828 269967
rect 124862 269933 124880 269967
rect 124811 269899 124880 269933
rect 124811 269865 124828 269899
rect 124862 269865 124880 269899
rect 124811 269831 124880 269865
rect 123827 269770 123986 269804
rect 124020 269770 124029 269804
rect 124188 269778 124209 269812
rect 124255 269778 124281 269812
rect 124323 269778 124353 269812
rect 124391 269778 124425 269812
rect 124459 269778 124493 269812
rect 124531 269778 124561 269812
rect 124603 269778 124629 269812
rect 124675 269778 124696 269812
rect 124811 269797 124828 269831
rect 124862 269797 124880 269831
rect 123827 269736 124029 269770
rect 123827 269702 123986 269736
rect 124020 269702 124029 269736
rect 123827 269668 124029 269702
rect 124811 269763 124880 269797
rect 124811 269729 124828 269763
rect 124862 269729 124880 269763
rect 124811 269695 124880 269729
rect 124811 269689 124828 269695
rect 123827 269634 123986 269668
rect 124020 269634 124029 269668
rect 123827 269600 124029 269634
rect 123827 269566 123986 269600
rect 124020 269566 124029 269600
rect 123827 269532 124029 269566
rect 123827 269498 123986 269532
rect 124020 269498 124029 269532
rect 123827 269464 124029 269498
rect 123827 269430 123986 269464
rect 124020 269430 124029 269464
rect 123827 269396 124029 269430
rect 123827 269362 123986 269396
rect 124020 269362 124029 269396
rect 123827 269281 124029 269362
rect 124116 269661 124828 269689
rect 124862 269668 124880 269695
rect 125047 269668 125058 272580
rect 124862 269661 125058 269668
rect 124116 269654 125058 269661
rect 124116 269620 124209 269654
rect 124255 269620 124281 269654
rect 124323 269620 124353 269654
rect 124391 269620 124425 269654
rect 124459 269620 124493 269654
rect 124531 269620 124561 269654
rect 124603 269620 124629 269654
rect 124675 269627 125058 269654
rect 124675 269620 124828 269627
rect 124116 269561 124188 269620
rect 124116 269525 124120 269561
rect 124154 269525 124188 269561
rect 124116 269491 124188 269525
rect 124116 269455 124120 269491
rect 124154 269455 124188 269491
rect 124116 269396 124188 269455
rect 124696 269593 124828 269620
rect 124862 269593 125058 269627
rect 124696 269561 125058 269593
rect 124696 269525 124730 269561
rect 124764 269559 125058 269561
rect 124764 269525 124828 269559
rect 124862 269525 125058 269559
rect 124696 269491 125058 269525
rect 124696 269455 124730 269491
rect 124764 269457 124828 269491
rect 124862 269457 125058 269491
rect 124764 269455 125058 269457
rect 124696 269423 125058 269455
rect 124696 269396 124828 269423
rect 124116 269362 124209 269396
rect 124255 269362 124281 269396
rect 124323 269362 124353 269396
rect 124391 269362 124425 269396
rect 124459 269362 124493 269396
rect 124531 269362 124561 269396
rect 124603 269362 124629 269396
rect 124675 269389 124828 269396
rect 124862 269389 125058 269423
rect 124675 269362 125058 269389
rect 124116 269281 124188 269362
rect 124696 269355 125058 269362
rect 124696 269321 124828 269355
rect 124862 269321 125058 269355
rect 124696 269281 125058 269321
rect 123827 269254 125058 269281
rect 123827 269220 124049 269254
rect 124083 269220 124117 269254
rect 124151 269220 124185 269254
rect 124219 269220 124253 269254
rect 124287 269220 124321 269254
rect 124355 269220 124389 269254
rect 124423 269220 124457 269254
rect 124491 269220 124525 269254
rect 124559 269220 124593 269254
rect 124627 269220 124661 269254
rect 124695 269220 125058 269254
rect 121645 268978 123550 268994
rect 120307 268946 123550 268978
rect 121789 268938 123550 268946
rect 123827 268990 125058 269220
rect 125160 275523 125658 280856
rect 125160 275151 128452 275523
rect 125160 268990 125825 275151
rect 123827 268861 125825 268990
rect 120072 268835 125825 268861
rect 120072 268785 120283 268835
rect 119938 268733 120283 268785
rect 125145 268733 125825 268835
rect 119938 268708 125825 268733
rect 111939 268659 119151 268677
rect 112005 268607 119104 268659
rect 123847 268607 125825 268708
rect 105957 268349 125825 268607
rect 128019 268349 128452 275151
rect 105957 268022 128452 268349
rect 105957 268007 125658 268022
<< viali >>
rect 106406 280851 106440 280885
rect 106806 280851 106840 280885
rect 107206 280851 107240 280885
rect 107606 280851 107640 280885
rect 108006 280851 108040 280885
rect 108406 280851 108440 280885
rect 108806 280851 108840 280885
rect 109206 280851 109240 280885
rect 109606 280851 109640 280885
rect 110006 280851 110040 280885
rect 106311 280762 106345 280788
rect 106311 280754 106345 280762
rect 106311 280694 106345 280716
rect 106311 280682 106345 280694
rect 106311 280626 106345 280644
rect 106311 280610 106345 280626
rect 106311 280558 106345 280572
rect 106311 280538 106345 280558
rect 106311 280490 106345 280500
rect 106311 280466 106345 280490
rect 106311 280422 106345 280428
rect 106311 280394 106345 280422
rect 106311 280354 106345 280356
rect 106311 280322 106345 280354
rect 106311 280252 106345 280284
rect 106311 280250 106345 280252
rect 106311 280184 106345 280212
rect 106311 280178 106345 280184
rect 106311 280116 106345 280140
rect 106311 280106 106345 280116
rect 106311 280048 106345 280068
rect 106311 280034 106345 280048
rect 106311 279980 106345 279996
rect 106311 279962 106345 279980
rect 106311 279912 106345 279924
rect 106311 279890 106345 279912
rect 106311 279844 106345 279852
rect 106311 279818 106345 279844
rect 106501 280762 106535 280788
rect 106501 280754 106535 280762
rect 106501 280694 106535 280716
rect 106501 280682 106535 280694
rect 106501 280626 106535 280644
rect 106501 280610 106535 280626
rect 106501 280558 106535 280572
rect 106501 280538 106535 280558
rect 106501 280490 106535 280500
rect 106501 280466 106535 280490
rect 106501 280422 106535 280428
rect 106501 280394 106535 280422
rect 106501 280354 106535 280356
rect 106501 280322 106535 280354
rect 106501 280252 106535 280284
rect 106501 280250 106535 280252
rect 106501 280184 106535 280212
rect 106501 280178 106535 280184
rect 106501 280116 106535 280140
rect 106501 280106 106535 280116
rect 106501 280048 106535 280068
rect 106501 280034 106535 280048
rect 106501 279980 106535 279996
rect 106501 279962 106535 279980
rect 106501 279912 106535 279924
rect 106501 279890 106535 279912
rect 106501 279844 106535 279852
rect 106501 279818 106535 279844
rect 106711 280762 106745 280788
rect 106711 280754 106745 280762
rect 106711 280694 106745 280716
rect 106711 280682 106745 280694
rect 106711 280626 106745 280644
rect 106711 280610 106745 280626
rect 106711 280558 106745 280572
rect 106711 280538 106745 280558
rect 106711 280490 106745 280500
rect 106711 280466 106745 280490
rect 106711 280422 106745 280428
rect 106711 280394 106745 280422
rect 106711 280354 106745 280356
rect 106711 280322 106745 280354
rect 106711 280252 106745 280284
rect 106711 280250 106745 280252
rect 106711 280184 106745 280212
rect 106711 280178 106745 280184
rect 106711 280116 106745 280140
rect 106711 280106 106745 280116
rect 106711 280048 106745 280068
rect 106711 280034 106745 280048
rect 106711 279980 106745 279996
rect 106711 279962 106745 279980
rect 106711 279912 106745 279924
rect 106711 279890 106745 279912
rect 106711 279844 106745 279852
rect 106711 279818 106745 279844
rect 106901 280762 106935 280788
rect 106901 280754 106935 280762
rect 106901 280694 106935 280716
rect 106901 280682 106935 280694
rect 106901 280626 106935 280644
rect 106901 280610 106935 280626
rect 106901 280558 106935 280572
rect 106901 280538 106935 280558
rect 106901 280490 106935 280500
rect 106901 280466 106935 280490
rect 106901 280422 106935 280428
rect 106901 280394 106935 280422
rect 106901 280354 106935 280356
rect 106901 280322 106935 280354
rect 106901 280252 106935 280284
rect 106901 280250 106935 280252
rect 106901 280184 106935 280212
rect 106901 280178 106935 280184
rect 106901 280116 106935 280140
rect 106901 280106 106935 280116
rect 106901 280048 106935 280068
rect 106901 280034 106935 280048
rect 106901 279980 106935 279996
rect 106901 279962 106935 279980
rect 106901 279912 106935 279924
rect 106901 279890 106935 279912
rect 106901 279844 106935 279852
rect 106901 279818 106935 279844
rect 107111 280762 107145 280788
rect 107111 280754 107145 280762
rect 107111 280694 107145 280716
rect 107111 280682 107145 280694
rect 107111 280626 107145 280644
rect 107111 280610 107145 280626
rect 107111 280558 107145 280572
rect 107111 280538 107145 280558
rect 107111 280490 107145 280500
rect 107111 280466 107145 280490
rect 107111 280422 107145 280428
rect 107111 280394 107145 280422
rect 107111 280354 107145 280356
rect 107111 280322 107145 280354
rect 107111 280252 107145 280284
rect 107111 280250 107145 280252
rect 107111 280184 107145 280212
rect 107111 280178 107145 280184
rect 107111 280116 107145 280140
rect 107111 280106 107145 280116
rect 107111 280048 107145 280068
rect 107111 280034 107145 280048
rect 107111 279980 107145 279996
rect 107111 279962 107145 279980
rect 107111 279912 107145 279924
rect 107111 279890 107145 279912
rect 107111 279844 107145 279852
rect 107111 279818 107145 279844
rect 107301 280762 107335 280788
rect 107301 280754 107335 280762
rect 107301 280694 107335 280716
rect 107301 280682 107335 280694
rect 107301 280626 107335 280644
rect 107301 280610 107335 280626
rect 107301 280558 107335 280572
rect 107301 280538 107335 280558
rect 107301 280490 107335 280500
rect 107301 280466 107335 280490
rect 107301 280422 107335 280428
rect 107301 280394 107335 280422
rect 107301 280354 107335 280356
rect 107301 280322 107335 280354
rect 107301 280252 107335 280284
rect 107301 280250 107335 280252
rect 107301 280184 107335 280212
rect 107301 280178 107335 280184
rect 107301 280116 107335 280140
rect 107301 280106 107335 280116
rect 107301 280048 107335 280068
rect 107301 280034 107335 280048
rect 107301 279980 107335 279996
rect 107301 279962 107335 279980
rect 107301 279912 107335 279924
rect 107301 279890 107335 279912
rect 107301 279844 107335 279852
rect 107301 279818 107335 279844
rect 107511 280762 107545 280788
rect 107511 280754 107545 280762
rect 107511 280694 107545 280716
rect 107511 280682 107545 280694
rect 107511 280626 107545 280644
rect 107511 280610 107545 280626
rect 107511 280558 107545 280572
rect 107511 280538 107545 280558
rect 107511 280490 107545 280500
rect 107511 280466 107545 280490
rect 107511 280422 107545 280428
rect 107511 280394 107545 280422
rect 107511 280354 107545 280356
rect 107511 280322 107545 280354
rect 107511 280252 107545 280284
rect 107511 280250 107545 280252
rect 107511 280184 107545 280212
rect 107511 280178 107545 280184
rect 107511 280116 107545 280140
rect 107511 280106 107545 280116
rect 107511 280048 107545 280068
rect 107511 280034 107545 280048
rect 107511 279980 107545 279996
rect 107511 279962 107545 279980
rect 107511 279912 107545 279924
rect 107511 279890 107545 279912
rect 107511 279844 107545 279852
rect 107511 279818 107545 279844
rect 107701 280762 107735 280788
rect 107701 280754 107735 280762
rect 107701 280694 107735 280716
rect 107701 280682 107735 280694
rect 107701 280626 107735 280644
rect 107701 280610 107735 280626
rect 107701 280558 107735 280572
rect 107701 280538 107735 280558
rect 107701 280490 107735 280500
rect 107701 280466 107735 280490
rect 107701 280422 107735 280428
rect 107701 280394 107735 280422
rect 107701 280354 107735 280356
rect 107701 280322 107735 280354
rect 107701 280252 107735 280284
rect 107701 280250 107735 280252
rect 107701 280184 107735 280212
rect 107701 280178 107735 280184
rect 107701 280116 107735 280140
rect 107701 280106 107735 280116
rect 107701 280048 107735 280068
rect 107701 280034 107735 280048
rect 107701 279980 107735 279996
rect 107701 279962 107735 279980
rect 107701 279912 107735 279924
rect 107701 279890 107735 279912
rect 107701 279844 107735 279852
rect 107701 279818 107735 279844
rect 107911 280762 107945 280788
rect 107911 280754 107945 280762
rect 107911 280694 107945 280716
rect 107911 280682 107945 280694
rect 107911 280626 107945 280644
rect 107911 280610 107945 280626
rect 107911 280558 107945 280572
rect 107911 280538 107945 280558
rect 107911 280490 107945 280500
rect 107911 280466 107945 280490
rect 107911 280422 107945 280428
rect 107911 280394 107945 280422
rect 107911 280354 107945 280356
rect 107911 280322 107945 280354
rect 107911 280252 107945 280284
rect 107911 280250 107945 280252
rect 107911 280184 107945 280212
rect 107911 280178 107945 280184
rect 107911 280116 107945 280140
rect 107911 280106 107945 280116
rect 107911 280048 107945 280068
rect 107911 280034 107945 280048
rect 107911 279980 107945 279996
rect 107911 279962 107945 279980
rect 107911 279912 107945 279924
rect 107911 279890 107945 279912
rect 107911 279844 107945 279852
rect 107911 279818 107945 279844
rect 108101 280762 108135 280788
rect 108101 280754 108135 280762
rect 108101 280694 108135 280716
rect 108101 280682 108135 280694
rect 108101 280626 108135 280644
rect 108101 280610 108135 280626
rect 108101 280558 108135 280572
rect 108101 280538 108135 280558
rect 108101 280490 108135 280500
rect 108101 280466 108135 280490
rect 108101 280422 108135 280428
rect 108101 280394 108135 280422
rect 108101 280354 108135 280356
rect 108101 280322 108135 280354
rect 108101 280252 108135 280284
rect 108101 280250 108135 280252
rect 108101 280184 108135 280212
rect 108101 280178 108135 280184
rect 108101 280116 108135 280140
rect 108101 280106 108135 280116
rect 108101 280048 108135 280068
rect 108101 280034 108135 280048
rect 108101 279980 108135 279996
rect 108101 279962 108135 279980
rect 108101 279912 108135 279924
rect 108101 279890 108135 279912
rect 108101 279844 108135 279852
rect 108101 279818 108135 279844
rect 108311 280762 108345 280788
rect 108311 280754 108345 280762
rect 108311 280694 108345 280716
rect 108311 280682 108345 280694
rect 108311 280626 108345 280644
rect 108311 280610 108345 280626
rect 108311 280558 108345 280572
rect 108311 280538 108345 280558
rect 108311 280490 108345 280500
rect 108311 280466 108345 280490
rect 108311 280422 108345 280428
rect 108311 280394 108345 280422
rect 108311 280354 108345 280356
rect 108311 280322 108345 280354
rect 108311 280252 108345 280284
rect 108311 280250 108345 280252
rect 108311 280184 108345 280212
rect 108311 280178 108345 280184
rect 108311 280116 108345 280140
rect 108311 280106 108345 280116
rect 108311 280048 108345 280068
rect 108311 280034 108345 280048
rect 108311 279980 108345 279996
rect 108311 279962 108345 279980
rect 108311 279912 108345 279924
rect 108311 279890 108345 279912
rect 108311 279844 108345 279852
rect 108311 279818 108345 279844
rect 108501 280762 108535 280788
rect 108501 280754 108535 280762
rect 108501 280694 108535 280716
rect 108501 280682 108535 280694
rect 108501 280626 108535 280644
rect 108501 280610 108535 280626
rect 108501 280558 108535 280572
rect 108501 280538 108535 280558
rect 108501 280490 108535 280500
rect 108501 280466 108535 280490
rect 108501 280422 108535 280428
rect 108501 280394 108535 280422
rect 108501 280354 108535 280356
rect 108501 280322 108535 280354
rect 108501 280252 108535 280284
rect 108501 280250 108535 280252
rect 108501 280184 108535 280212
rect 108501 280178 108535 280184
rect 108501 280116 108535 280140
rect 108501 280106 108535 280116
rect 108501 280048 108535 280068
rect 108501 280034 108535 280048
rect 108501 279980 108535 279996
rect 108501 279962 108535 279980
rect 108501 279912 108535 279924
rect 108501 279890 108535 279912
rect 108501 279844 108535 279852
rect 108501 279818 108535 279844
rect 108711 280762 108745 280788
rect 108711 280754 108745 280762
rect 108711 280694 108745 280716
rect 108711 280682 108745 280694
rect 108711 280626 108745 280644
rect 108711 280610 108745 280626
rect 108711 280558 108745 280572
rect 108711 280538 108745 280558
rect 108711 280490 108745 280500
rect 108711 280466 108745 280490
rect 108711 280422 108745 280428
rect 108711 280394 108745 280422
rect 108711 280354 108745 280356
rect 108711 280322 108745 280354
rect 108711 280252 108745 280284
rect 108711 280250 108745 280252
rect 108711 280184 108745 280212
rect 108711 280178 108745 280184
rect 108711 280116 108745 280140
rect 108711 280106 108745 280116
rect 108711 280048 108745 280068
rect 108711 280034 108745 280048
rect 108711 279980 108745 279996
rect 108711 279962 108745 279980
rect 108711 279912 108745 279924
rect 108711 279890 108745 279912
rect 108711 279844 108745 279852
rect 108711 279818 108745 279844
rect 108901 280762 108935 280788
rect 108901 280754 108935 280762
rect 108901 280694 108935 280716
rect 108901 280682 108935 280694
rect 108901 280626 108935 280644
rect 108901 280610 108935 280626
rect 108901 280558 108935 280572
rect 108901 280538 108935 280558
rect 108901 280490 108935 280500
rect 108901 280466 108935 280490
rect 108901 280422 108935 280428
rect 108901 280394 108935 280422
rect 108901 280354 108935 280356
rect 108901 280322 108935 280354
rect 108901 280252 108935 280284
rect 108901 280250 108935 280252
rect 108901 280184 108935 280212
rect 108901 280178 108935 280184
rect 108901 280116 108935 280140
rect 108901 280106 108935 280116
rect 108901 280048 108935 280068
rect 108901 280034 108935 280048
rect 108901 279980 108935 279996
rect 108901 279962 108935 279980
rect 108901 279912 108935 279924
rect 108901 279890 108935 279912
rect 108901 279844 108935 279852
rect 108901 279818 108935 279844
rect 109111 280762 109145 280788
rect 109111 280754 109145 280762
rect 109111 280694 109145 280716
rect 109111 280682 109145 280694
rect 109111 280626 109145 280644
rect 109111 280610 109145 280626
rect 109111 280558 109145 280572
rect 109111 280538 109145 280558
rect 109111 280490 109145 280500
rect 109111 280466 109145 280490
rect 109111 280422 109145 280428
rect 109111 280394 109145 280422
rect 109111 280354 109145 280356
rect 109111 280322 109145 280354
rect 109111 280252 109145 280284
rect 109111 280250 109145 280252
rect 109111 280184 109145 280212
rect 109111 280178 109145 280184
rect 109111 280116 109145 280140
rect 109111 280106 109145 280116
rect 109111 280048 109145 280068
rect 109111 280034 109145 280048
rect 109111 279980 109145 279996
rect 109111 279962 109145 279980
rect 109111 279912 109145 279924
rect 109111 279890 109145 279912
rect 109111 279844 109145 279852
rect 109111 279818 109145 279844
rect 109301 280762 109335 280788
rect 109301 280754 109335 280762
rect 109301 280694 109335 280716
rect 109301 280682 109335 280694
rect 109301 280626 109335 280644
rect 109301 280610 109335 280626
rect 109301 280558 109335 280572
rect 109301 280538 109335 280558
rect 109301 280490 109335 280500
rect 109301 280466 109335 280490
rect 109301 280422 109335 280428
rect 109301 280394 109335 280422
rect 109301 280354 109335 280356
rect 109301 280322 109335 280354
rect 109301 280252 109335 280284
rect 109301 280250 109335 280252
rect 109301 280184 109335 280212
rect 109301 280178 109335 280184
rect 109301 280116 109335 280140
rect 109301 280106 109335 280116
rect 109301 280048 109335 280068
rect 109301 280034 109335 280048
rect 109301 279980 109335 279996
rect 109301 279962 109335 279980
rect 109301 279912 109335 279924
rect 109301 279890 109335 279912
rect 109301 279844 109335 279852
rect 109301 279818 109335 279844
rect 109511 280762 109545 280788
rect 109511 280754 109545 280762
rect 109511 280694 109545 280716
rect 109511 280682 109545 280694
rect 109511 280626 109545 280644
rect 109511 280610 109545 280626
rect 109511 280558 109545 280572
rect 109511 280538 109545 280558
rect 109511 280490 109545 280500
rect 109511 280466 109545 280490
rect 109511 280422 109545 280428
rect 109511 280394 109545 280422
rect 109511 280354 109545 280356
rect 109511 280322 109545 280354
rect 109511 280252 109545 280284
rect 109511 280250 109545 280252
rect 109511 280184 109545 280212
rect 109511 280178 109545 280184
rect 109511 280116 109545 280140
rect 109511 280106 109545 280116
rect 109511 280048 109545 280068
rect 109511 280034 109545 280048
rect 109511 279980 109545 279996
rect 109511 279962 109545 279980
rect 109511 279912 109545 279924
rect 109511 279890 109545 279912
rect 109511 279844 109545 279852
rect 109511 279818 109545 279844
rect 109701 280762 109735 280788
rect 109701 280754 109735 280762
rect 109701 280694 109735 280716
rect 109701 280682 109735 280694
rect 109701 280626 109735 280644
rect 109701 280610 109735 280626
rect 109701 280558 109735 280572
rect 109701 280538 109735 280558
rect 109701 280490 109735 280500
rect 109701 280466 109735 280490
rect 109701 280422 109735 280428
rect 109701 280394 109735 280422
rect 109701 280354 109735 280356
rect 109701 280322 109735 280354
rect 109701 280252 109735 280284
rect 109701 280250 109735 280252
rect 109701 280184 109735 280212
rect 109701 280178 109735 280184
rect 109701 280116 109735 280140
rect 109701 280106 109735 280116
rect 109701 280048 109735 280068
rect 109701 280034 109735 280048
rect 109701 279980 109735 279996
rect 109701 279962 109735 279980
rect 109701 279912 109735 279924
rect 109701 279890 109735 279912
rect 109701 279844 109735 279852
rect 109701 279818 109735 279844
rect 109911 280762 109945 280788
rect 109911 280754 109945 280762
rect 109911 280694 109945 280716
rect 109911 280682 109945 280694
rect 109911 280626 109945 280644
rect 109911 280610 109945 280626
rect 109911 280558 109945 280572
rect 109911 280538 109945 280558
rect 109911 280490 109945 280500
rect 109911 280466 109945 280490
rect 109911 280422 109945 280428
rect 109911 280394 109945 280422
rect 109911 280354 109945 280356
rect 109911 280322 109945 280354
rect 109911 280252 109945 280284
rect 109911 280250 109945 280252
rect 109911 280184 109945 280212
rect 109911 280178 109945 280184
rect 109911 280116 109945 280140
rect 109911 280106 109945 280116
rect 109911 280048 109945 280068
rect 109911 280034 109945 280048
rect 109911 279980 109945 279996
rect 109911 279962 109945 279980
rect 109911 279912 109945 279924
rect 109911 279890 109945 279912
rect 109911 279844 109945 279852
rect 109911 279818 109945 279844
rect 110101 280762 110135 280788
rect 110101 280754 110135 280762
rect 110101 280694 110135 280716
rect 110101 280682 110135 280694
rect 110101 280626 110135 280644
rect 110101 280610 110135 280626
rect 110101 280558 110135 280572
rect 110101 280538 110135 280558
rect 110101 280490 110135 280500
rect 110101 280466 110135 280490
rect 110101 280422 110135 280428
rect 110101 280394 110135 280422
rect 110101 280354 110135 280356
rect 110101 280322 110135 280354
rect 110101 280252 110135 280284
rect 110101 280250 110135 280252
rect 110101 280184 110135 280212
rect 110101 280178 110135 280184
rect 110101 280116 110135 280140
rect 110101 280106 110135 280116
rect 110101 280048 110135 280068
rect 110101 280034 110135 280048
rect 110101 279980 110135 279996
rect 110101 279962 110135 279980
rect 110101 279912 110135 279924
rect 110101 279890 110135 279912
rect 110101 279844 110135 279852
rect 110101 279818 110135 279844
rect 106406 279721 106440 279755
rect 106806 279721 106840 279755
rect 107206 279721 107240 279755
rect 107606 279721 107640 279755
rect 108006 279721 108040 279755
rect 108406 279721 108440 279755
rect 108806 279721 108840 279755
rect 109206 279721 109240 279755
rect 109606 279721 109640 279755
rect 110006 279721 110040 279755
rect 106382 279023 106414 279057
rect 106414 279023 106416 279057
rect 106454 279023 106482 279057
rect 106482 279023 106488 279057
rect 106526 279023 106550 279057
rect 106550 279023 106560 279057
rect 106598 279023 106618 279057
rect 106618 279023 106632 279057
rect 106670 279023 106686 279057
rect 106686 279023 106704 279057
rect 106742 279023 106754 279057
rect 106754 279023 106776 279057
rect 106814 279023 106822 279057
rect 106822 279023 106848 279057
rect 106886 279023 106890 279057
rect 106890 279023 106920 279057
rect 106958 279023 106992 279057
rect 107030 279023 107060 279057
rect 107060 279023 107064 279057
rect 107102 279023 107128 279057
rect 107128 279023 107136 279057
rect 107174 279023 107196 279057
rect 107196 279023 107208 279057
rect 107246 279023 107264 279057
rect 107264 279023 107280 279057
rect 107318 279023 107332 279057
rect 107332 279023 107352 279057
rect 107390 279023 107400 279057
rect 107400 279023 107424 279057
rect 107462 279023 107468 279057
rect 107468 279023 107496 279057
rect 107534 279023 107536 279057
rect 107536 279023 107568 279057
rect 106287 278969 106321 278973
rect 106287 278939 106321 278969
rect 106287 278867 106321 278901
rect 106287 278799 106321 278829
rect 106287 278795 106321 278799
rect 107629 278969 107663 278973
rect 107629 278939 107663 278969
rect 107629 278867 107663 278901
rect 107629 278799 107663 278829
rect 107629 278795 107663 278799
rect 106382 278711 106414 278745
rect 106414 278711 106416 278745
rect 106454 278711 106482 278745
rect 106482 278711 106488 278745
rect 106526 278711 106550 278745
rect 106550 278711 106560 278745
rect 106598 278711 106618 278745
rect 106618 278711 106632 278745
rect 106670 278711 106686 278745
rect 106686 278711 106704 278745
rect 106742 278711 106754 278745
rect 106754 278711 106776 278745
rect 106814 278711 106822 278745
rect 106822 278711 106848 278745
rect 106886 278711 106890 278745
rect 106890 278711 106920 278745
rect 106958 278711 106992 278745
rect 107030 278711 107060 278745
rect 107060 278711 107064 278745
rect 107102 278711 107128 278745
rect 107128 278711 107136 278745
rect 107174 278711 107196 278745
rect 107196 278711 107208 278745
rect 107246 278711 107264 278745
rect 107264 278711 107280 278745
rect 107318 278711 107332 278745
rect 107332 278711 107352 278745
rect 107390 278711 107400 278745
rect 107400 278711 107424 278745
rect 107462 278711 107468 278745
rect 107468 278711 107496 278745
rect 107534 278711 107536 278745
rect 107536 278711 107568 278745
rect 106382 278423 106414 278457
rect 106414 278423 106416 278457
rect 106454 278423 106482 278457
rect 106482 278423 106488 278457
rect 106526 278423 106550 278457
rect 106550 278423 106560 278457
rect 106598 278423 106618 278457
rect 106618 278423 106632 278457
rect 106670 278423 106686 278457
rect 106686 278423 106704 278457
rect 106742 278423 106754 278457
rect 106754 278423 106776 278457
rect 106814 278423 106822 278457
rect 106822 278423 106848 278457
rect 106886 278423 106890 278457
rect 106890 278423 106920 278457
rect 106958 278423 106992 278457
rect 107030 278423 107060 278457
rect 107060 278423 107064 278457
rect 107102 278423 107128 278457
rect 107128 278423 107136 278457
rect 107174 278423 107196 278457
rect 107196 278423 107208 278457
rect 107246 278423 107264 278457
rect 107264 278423 107280 278457
rect 107318 278423 107332 278457
rect 107332 278423 107352 278457
rect 107390 278423 107400 278457
rect 107400 278423 107424 278457
rect 107462 278423 107468 278457
rect 107468 278423 107496 278457
rect 107534 278423 107536 278457
rect 107536 278423 107568 278457
rect 106287 278369 106321 278373
rect 106287 278339 106321 278369
rect 106287 278267 106321 278301
rect 106287 278199 106321 278229
rect 106287 278195 106321 278199
rect 107629 278369 107663 278373
rect 107629 278339 107663 278369
rect 107629 278267 107663 278301
rect 107629 278199 107663 278229
rect 107629 278195 107663 278199
rect 106382 278111 106414 278145
rect 106414 278111 106416 278145
rect 106454 278111 106482 278145
rect 106482 278111 106488 278145
rect 106526 278111 106550 278145
rect 106550 278111 106560 278145
rect 106598 278111 106618 278145
rect 106618 278111 106632 278145
rect 106670 278111 106686 278145
rect 106686 278111 106704 278145
rect 106742 278111 106754 278145
rect 106754 278111 106776 278145
rect 106814 278111 106822 278145
rect 106822 278111 106848 278145
rect 106886 278111 106890 278145
rect 106890 278111 106920 278145
rect 106958 278111 106992 278145
rect 107030 278111 107060 278145
rect 107060 278111 107064 278145
rect 107102 278111 107128 278145
rect 107128 278111 107136 278145
rect 107174 278111 107196 278145
rect 107196 278111 107208 278145
rect 107246 278111 107264 278145
rect 107264 278111 107280 278145
rect 107318 278111 107332 278145
rect 107332 278111 107352 278145
rect 107390 278111 107400 278145
rect 107400 278111 107424 278145
rect 107462 278111 107468 278145
rect 107468 278111 107496 278145
rect 107534 278111 107536 278145
rect 107536 278111 107568 278145
rect 106966 277984 107072 278053
rect 106966 277950 106985 277984
rect 106985 277950 107019 277984
rect 107019 277950 107053 277984
rect 107053 277950 107072 277984
rect 109795 279049 109801 279083
rect 109801 279049 109829 279083
rect 109867 279049 109869 279083
rect 109869 279049 109901 279083
rect 109939 279049 109971 279083
rect 109971 279049 109973 279083
rect 110011 279049 110039 279083
rect 110039 279049 110045 279083
rect 106966 277803 107072 277950
rect 109731 278951 109765 278977
rect 109731 278943 109765 278951
rect 109731 278883 109765 278905
rect 109731 278871 109765 278883
rect 109731 278815 109765 278833
rect 109731 278799 109765 278815
rect 109731 278747 109765 278761
rect 109731 278727 109765 278747
rect 109731 278679 109765 278689
rect 109731 278655 109765 278679
rect 109731 278611 109765 278617
rect 109731 278583 109765 278611
rect 109731 278543 109765 278545
rect 109731 278511 109765 278543
rect 109731 278441 109765 278473
rect 109731 278439 109765 278441
rect 109731 278373 109765 278401
rect 109731 278367 109765 278373
rect 109731 278305 109765 278329
rect 109731 278295 109765 278305
rect 109731 278237 109765 278257
rect 109731 278223 109765 278237
rect 109731 278169 109765 278185
rect 109731 278151 109765 278169
rect 109731 278101 109765 278113
rect 109731 278079 109765 278101
rect 109731 278033 109765 278041
rect 109731 278007 109765 278033
rect 110075 278951 110109 278977
rect 110075 278943 110109 278951
rect 110075 278883 110109 278905
rect 110075 278871 110109 278883
rect 110075 278815 110109 278833
rect 110075 278799 110109 278815
rect 110075 278747 110109 278761
rect 110075 278727 110109 278747
rect 110075 278679 110109 278689
rect 110075 278655 110109 278679
rect 110075 278611 110109 278617
rect 110075 278583 110109 278611
rect 110075 278543 110109 278545
rect 110075 278511 110109 278543
rect 110075 278441 110109 278473
rect 110075 278439 110109 278441
rect 110075 278373 110109 278401
rect 110075 278367 110109 278373
rect 110075 278305 110109 278329
rect 110075 278295 110109 278305
rect 110075 278237 110109 278257
rect 110075 278223 110109 278237
rect 110075 278169 110109 278185
rect 110075 278151 110109 278169
rect 110075 278101 110109 278113
rect 110075 278079 110109 278101
rect 110075 278033 110109 278041
rect 110075 278007 110109 278033
rect 109795 277901 109801 277935
rect 109801 277901 109829 277935
rect 109867 277901 109869 277935
rect 109869 277901 109901 277935
rect 109939 277901 109971 277935
rect 109971 277901 109973 277935
rect 110011 277901 110039 277935
rect 110039 277901 110045 277935
rect 109795 277793 109801 277827
rect 109801 277793 109829 277827
rect 109867 277793 109869 277827
rect 109869 277793 109901 277827
rect 109939 277793 109971 277827
rect 109971 277793 109973 277827
rect 110011 277793 110039 277827
rect 110039 277793 110045 277827
rect 106523 277176 106549 277210
rect 106549 277176 106557 277210
rect 106595 277176 106617 277210
rect 106617 277176 106629 277210
rect 106667 277176 106685 277210
rect 106685 277176 106701 277210
rect 106739 277176 106753 277210
rect 106753 277176 106773 277210
rect 106811 277176 106821 277210
rect 106821 277176 106845 277210
rect 106883 277176 106889 277210
rect 106889 277176 106917 277210
rect 106955 277176 106957 277210
rect 106957 277176 106989 277210
rect 107027 277176 107059 277210
rect 107059 277176 107061 277210
rect 107099 277176 107127 277210
rect 107127 277176 107133 277210
rect 107171 277176 107195 277210
rect 107195 277176 107205 277210
rect 107243 277176 107263 277210
rect 107263 277176 107277 277210
rect 107315 277176 107331 277210
rect 107331 277176 107349 277210
rect 107387 277176 107399 277210
rect 107399 277176 107421 277210
rect 107459 277176 107467 277210
rect 107467 277176 107493 277210
rect 106410 277110 106444 277144
rect 107572 277110 107606 277144
rect 106523 277044 106549 277078
rect 106549 277044 106557 277078
rect 106595 277044 106617 277078
rect 106617 277044 106629 277078
rect 106667 277044 106685 277078
rect 106685 277044 106701 277078
rect 106739 277044 106753 277078
rect 106753 277044 106773 277078
rect 106811 277044 106821 277078
rect 106821 277044 106845 277078
rect 106883 277044 106889 277078
rect 106889 277044 106917 277078
rect 106955 277044 106957 277078
rect 106957 277044 106989 277078
rect 107027 277044 107059 277078
rect 107059 277044 107061 277078
rect 107099 277044 107127 277078
rect 107127 277044 107133 277078
rect 107171 277044 107195 277078
rect 107195 277044 107205 277078
rect 107243 277044 107263 277078
rect 107263 277044 107277 277078
rect 107315 277044 107331 277078
rect 107331 277044 107349 277078
rect 107387 277044 107399 277078
rect 107399 277044 107421 277078
rect 107459 277044 107467 277078
rect 107467 277044 107493 277078
rect 109731 277695 109765 277721
rect 109731 277687 109765 277695
rect 109731 277627 109765 277649
rect 109731 277615 109765 277627
rect 109731 277559 109765 277577
rect 109731 277543 109765 277559
rect 109731 277491 109765 277505
rect 109731 277471 109765 277491
rect 109731 277423 109765 277433
rect 109731 277399 109765 277423
rect 109731 277355 109765 277361
rect 109731 277327 109765 277355
rect 109731 277287 109765 277289
rect 109731 277255 109765 277287
rect 109731 277185 109765 277217
rect 109731 277183 109765 277185
rect 109731 277117 109765 277145
rect 109731 277111 109765 277117
rect 109731 277049 109765 277073
rect 109731 277039 109765 277049
rect 109731 276981 109765 277001
rect 109731 276967 109765 276981
rect 109731 276913 109765 276929
rect 109731 276895 109765 276913
rect 109731 276845 109765 276857
rect 109731 276823 109765 276845
rect 109731 276777 109765 276785
rect 109731 276751 109765 276777
rect 110075 277695 110109 277721
rect 110075 277687 110109 277695
rect 110075 277627 110109 277649
rect 110075 277615 110109 277627
rect 110075 277559 110109 277577
rect 110075 277543 110109 277559
rect 110075 277491 110109 277505
rect 110075 277471 110109 277491
rect 110075 277423 110109 277433
rect 110075 277399 110109 277423
rect 110075 277355 110109 277361
rect 110075 277327 110109 277355
rect 110075 277287 110109 277289
rect 110075 277255 110109 277287
rect 110075 277185 110109 277217
rect 110075 277183 110109 277185
rect 110075 277117 110109 277145
rect 110075 277111 110109 277117
rect 110075 277049 110109 277073
rect 110075 277039 110109 277049
rect 110075 276981 110109 277001
rect 110075 276967 110109 276981
rect 110075 276913 110109 276929
rect 110075 276895 110109 276913
rect 110075 276845 110109 276857
rect 110075 276823 110109 276845
rect 110075 276777 110109 276785
rect 110075 276751 110109 276777
rect 109795 276645 109801 276679
rect 109801 276645 109829 276679
rect 109867 276645 109869 276679
rect 109869 276645 109901 276679
rect 109939 276645 109971 276679
rect 109971 276645 109973 276679
rect 110011 276645 110039 276679
rect 110039 276645 110045 276679
rect 106409 274870 106515 276272
rect 106987 275725 106989 275759
rect 106989 275725 107021 275759
rect 107059 275725 107091 275759
rect 107091 275725 107093 275759
rect 107487 275725 107489 275759
rect 107489 275725 107521 275759
rect 107559 275725 107591 275759
rect 107591 275725 107593 275759
rect 107987 275725 107989 275759
rect 107989 275725 108021 275759
rect 108059 275725 108091 275759
rect 108091 275725 108093 275759
rect 108487 275725 108489 275759
rect 108489 275725 108521 275759
rect 108559 275725 108591 275759
rect 108591 275725 108593 275759
rect 108987 275725 108989 275759
rect 108989 275725 109021 275759
rect 109059 275725 109091 275759
rect 109091 275725 109093 275759
rect 109487 275725 109489 275759
rect 109489 275725 109521 275759
rect 109559 275725 109591 275759
rect 109591 275725 109593 275759
rect 106870 275647 106904 275665
rect 106870 275631 106904 275647
rect 106870 275579 106904 275593
rect 106870 275559 106904 275579
rect 106870 275511 106904 275521
rect 106870 275487 106904 275511
rect 106870 275443 106904 275449
rect 106870 275415 106904 275443
rect 106870 275375 106904 275377
rect 106870 275343 106904 275375
rect 106870 275273 106904 275305
rect 106870 275271 106904 275273
rect 106870 275205 106904 275233
rect 106870 275199 106904 275205
rect 106870 275137 106904 275161
rect 106870 275127 106904 275137
rect 106870 275069 106904 275089
rect 106870 275055 106904 275069
rect 106870 275001 106904 275017
rect 106870 274983 106904 275001
rect 107176 275647 107210 275665
rect 107176 275631 107210 275647
rect 107176 275579 107210 275593
rect 107176 275559 107210 275579
rect 107176 275511 107210 275521
rect 107176 275487 107210 275511
rect 107176 275443 107210 275449
rect 107176 275415 107210 275443
rect 107176 275375 107210 275377
rect 107176 275343 107210 275375
rect 107176 275273 107210 275305
rect 107176 275271 107210 275273
rect 107176 275205 107210 275233
rect 107176 275199 107210 275205
rect 107176 275137 107210 275161
rect 107176 275127 107210 275137
rect 107176 275069 107210 275089
rect 107176 275055 107210 275069
rect 107176 275001 107210 275017
rect 107176 274983 107210 275001
rect 107370 275647 107404 275665
rect 107370 275631 107404 275647
rect 107370 275579 107404 275593
rect 107370 275559 107404 275579
rect 107370 275511 107404 275521
rect 107370 275487 107404 275511
rect 107370 275443 107404 275449
rect 107370 275415 107404 275443
rect 107370 275375 107404 275377
rect 107370 275343 107404 275375
rect 107370 275273 107404 275305
rect 107370 275271 107404 275273
rect 107370 275205 107404 275233
rect 107370 275199 107404 275205
rect 107370 275137 107404 275161
rect 107370 275127 107404 275137
rect 107370 275069 107404 275089
rect 107370 275055 107404 275069
rect 107370 275001 107404 275017
rect 107370 274983 107404 275001
rect 107676 275647 107710 275665
rect 107676 275631 107710 275647
rect 107676 275579 107710 275593
rect 107676 275559 107710 275579
rect 107676 275511 107710 275521
rect 107676 275487 107710 275511
rect 107676 275443 107710 275449
rect 107676 275415 107710 275443
rect 107676 275375 107710 275377
rect 107676 275343 107710 275375
rect 107676 275273 107710 275305
rect 107676 275271 107710 275273
rect 107676 275205 107710 275233
rect 107676 275199 107710 275205
rect 107676 275137 107710 275161
rect 107676 275127 107710 275137
rect 107676 275069 107710 275089
rect 107676 275055 107710 275069
rect 107676 275001 107710 275017
rect 107676 274983 107710 275001
rect 107870 275647 107904 275665
rect 107870 275631 107904 275647
rect 107870 275579 107904 275593
rect 107870 275559 107904 275579
rect 107870 275511 107904 275521
rect 107870 275487 107904 275511
rect 107870 275443 107904 275449
rect 107870 275415 107904 275443
rect 107870 275375 107904 275377
rect 107870 275343 107904 275375
rect 107870 275273 107904 275305
rect 107870 275271 107904 275273
rect 107870 275205 107904 275233
rect 107870 275199 107904 275205
rect 107870 275137 107904 275161
rect 107870 275127 107904 275137
rect 107870 275069 107904 275089
rect 107870 275055 107904 275069
rect 107870 275001 107904 275017
rect 107870 274983 107904 275001
rect 108176 275647 108210 275665
rect 108176 275631 108210 275647
rect 108176 275579 108210 275593
rect 108176 275559 108210 275579
rect 108176 275511 108210 275521
rect 108176 275487 108210 275511
rect 108176 275443 108210 275449
rect 108176 275415 108210 275443
rect 108176 275375 108210 275377
rect 108176 275343 108210 275375
rect 108176 275273 108210 275305
rect 108176 275271 108210 275273
rect 108176 275205 108210 275233
rect 108176 275199 108210 275205
rect 108176 275137 108210 275161
rect 108176 275127 108210 275137
rect 108176 275069 108210 275089
rect 108176 275055 108210 275069
rect 108176 275001 108210 275017
rect 108176 274983 108210 275001
rect 108370 275647 108404 275665
rect 108370 275631 108404 275647
rect 108370 275579 108404 275593
rect 108370 275559 108404 275579
rect 108370 275511 108404 275521
rect 108370 275487 108404 275511
rect 108370 275443 108404 275449
rect 108370 275415 108404 275443
rect 108370 275375 108404 275377
rect 108370 275343 108404 275375
rect 108370 275273 108404 275305
rect 108370 275271 108404 275273
rect 108370 275205 108404 275233
rect 108370 275199 108404 275205
rect 108370 275137 108404 275161
rect 108370 275127 108404 275137
rect 108370 275069 108404 275089
rect 108370 275055 108404 275069
rect 108370 275001 108404 275017
rect 108370 274983 108404 275001
rect 108676 275647 108710 275665
rect 108676 275631 108710 275647
rect 108676 275579 108710 275593
rect 108676 275559 108710 275579
rect 108676 275511 108710 275521
rect 108676 275487 108710 275511
rect 108676 275443 108710 275449
rect 108676 275415 108710 275443
rect 108676 275375 108710 275377
rect 108676 275343 108710 275375
rect 108676 275273 108710 275305
rect 108676 275271 108710 275273
rect 108676 275205 108710 275233
rect 108676 275199 108710 275205
rect 108676 275137 108710 275161
rect 108676 275127 108710 275137
rect 108676 275069 108710 275089
rect 108676 275055 108710 275069
rect 108676 275001 108710 275017
rect 108676 274983 108710 275001
rect 108870 275647 108904 275665
rect 108870 275631 108904 275647
rect 108870 275579 108904 275593
rect 108870 275559 108904 275579
rect 108870 275511 108904 275521
rect 108870 275487 108904 275511
rect 108870 275443 108904 275449
rect 108870 275415 108904 275443
rect 108870 275375 108904 275377
rect 108870 275343 108904 275375
rect 108870 275273 108904 275305
rect 108870 275271 108904 275273
rect 108870 275205 108904 275233
rect 108870 275199 108904 275205
rect 108870 275137 108904 275161
rect 108870 275127 108904 275137
rect 108870 275069 108904 275089
rect 108870 275055 108904 275069
rect 108870 275001 108904 275017
rect 108870 274983 108904 275001
rect 109176 275647 109210 275665
rect 109176 275631 109210 275647
rect 109176 275579 109210 275593
rect 109176 275559 109210 275579
rect 109176 275511 109210 275521
rect 109176 275487 109210 275511
rect 109176 275443 109210 275449
rect 109176 275415 109210 275443
rect 109176 275375 109210 275377
rect 109176 275343 109210 275375
rect 109176 275273 109210 275305
rect 109176 275271 109210 275273
rect 109176 275205 109210 275233
rect 109176 275199 109210 275205
rect 109176 275137 109210 275161
rect 109176 275127 109210 275137
rect 109176 275069 109210 275089
rect 109176 275055 109210 275069
rect 109176 275001 109210 275017
rect 109176 274983 109210 275001
rect 109370 275647 109404 275665
rect 109370 275631 109404 275647
rect 109370 275579 109404 275593
rect 109370 275559 109404 275579
rect 109370 275511 109404 275521
rect 109370 275487 109404 275511
rect 109370 275443 109404 275449
rect 109370 275415 109404 275443
rect 109370 275375 109404 275377
rect 109370 275343 109404 275375
rect 109370 275273 109404 275305
rect 109370 275271 109404 275273
rect 109370 275205 109404 275233
rect 109370 275199 109404 275205
rect 109370 275137 109404 275161
rect 109370 275127 109404 275137
rect 109370 275069 109404 275089
rect 109370 275055 109404 275069
rect 109370 275001 109404 275017
rect 109370 274983 109404 275001
rect 109676 275647 109710 275665
rect 109676 275631 109710 275647
rect 109676 275579 109710 275593
rect 109676 275559 109710 275579
rect 109676 275511 109710 275521
rect 109676 275487 109710 275511
rect 109676 275443 109710 275449
rect 109676 275415 109710 275443
rect 109676 275375 109710 275377
rect 109676 275343 109710 275375
rect 109676 275273 109710 275305
rect 109676 275271 109710 275273
rect 109676 275205 109710 275233
rect 109676 275199 109710 275205
rect 109676 275137 109710 275161
rect 109676 275127 109710 275137
rect 109676 275069 109710 275089
rect 109676 275055 109710 275069
rect 109676 275001 109710 275017
rect 109676 274983 109710 275001
rect 106987 274889 106989 274923
rect 106989 274889 107021 274923
rect 107059 274889 107091 274923
rect 107091 274889 107093 274923
rect 107487 274889 107489 274923
rect 107489 274889 107521 274923
rect 107559 274889 107591 274923
rect 107591 274889 107593 274923
rect 107987 274889 107989 274923
rect 107989 274889 108021 274923
rect 108059 274889 108091 274923
rect 108091 274889 108093 274923
rect 108487 274889 108489 274923
rect 108489 274889 108521 274923
rect 108559 274889 108591 274923
rect 108591 274889 108593 274923
rect 108987 274889 108989 274923
rect 108989 274889 109021 274923
rect 109059 274889 109091 274923
rect 109091 274889 109093 274923
rect 109487 274889 109489 274923
rect 109489 274889 109521 274923
rect 109559 274889 109591 274923
rect 109591 274889 109593 274923
rect 107500 272117 107514 272151
rect 107514 272117 107534 272151
rect 107572 272117 107582 272151
rect 107582 272117 107606 272151
rect 107644 272117 107650 272151
rect 107650 272117 107678 272151
rect 107716 272117 107718 272151
rect 107718 272117 107750 272151
rect 107788 272117 107820 272151
rect 107820 272117 107822 272151
rect 107860 272117 107888 272151
rect 107888 272117 107894 272151
rect 107932 272117 107956 272151
rect 107956 272117 107966 272151
rect 108004 272117 108024 272151
rect 108024 272117 108038 272151
rect 106997 272009 107001 272043
rect 107001 272009 107031 272043
rect 107069 272009 107103 272043
rect 107141 272009 107171 272043
rect 107171 272009 107175 272043
rect 107413 272026 107447 272032
rect 107413 271998 107447 272026
rect 106935 271940 106969 271942
rect 106935 271908 106969 271940
rect 106935 271838 106969 271870
rect 106935 271836 106969 271838
rect 107203 271940 107237 271942
rect 107203 271908 107237 271940
rect 107203 271838 107237 271870
rect 107203 271836 107237 271838
rect 107413 271958 107447 271960
rect 107413 271926 107447 271958
rect 107413 271856 107447 271888
rect 107413 271854 107447 271856
rect 107413 271788 107447 271816
rect 107413 271782 107447 271788
rect 106997 271735 107001 271769
rect 107001 271735 107031 271769
rect 107069 271735 107103 271769
rect 107141 271735 107171 271769
rect 107171 271735 107175 271769
rect 108091 272026 108125 272032
rect 108091 271998 108125 272026
rect 108091 271958 108125 271960
rect 108091 271926 108125 271958
rect 108091 271856 108125 271888
rect 108091 271854 108125 271856
rect 108091 271788 108125 271816
rect 108091 271782 108125 271788
rect 107500 271663 107514 271697
rect 107514 271663 107534 271697
rect 107572 271663 107582 271697
rect 107582 271663 107606 271697
rect 107644 271663 107650 271697
rect 107650 271663 107678 271697
rect 107716 271663 107718 271697
rect 107718 271663 107750 271697
rect 107788 271663 107820 271697
rect 107820 271663 107822 271697
rect 107860 271663 107888 271697
rect 107888 271663 107894 271697
rect 107932 271663 107956 271697
rect 107956 271663 107966 271697
rect 108004 271663 108024 271697
rect 108024 271663 108038 271697
rect 107216 271501 107246 271535
rect 107246 271501 107250 271535
rect 107288 271501 107314 271535
rect 107314 271501 107322 271535
rect 107360 271501 107382 271535
rect 107382 271501 107394 271535
rect 107432 271501 107450 271535
rect 107450 271501 107466 271535
rect 107504 271501 107518 271535
rect 107518 271501 107538 271535
rect 107576 271501 107586 271535
rect 107586 271501 107610 271535
rect 107648 271501 107654 271535
rect 107654 271501 107682 271535
rect 107720 271501 107722 271535
rect 107722 271501 107754 271535
rect 107792 271501 107824 271535
rect 107824 271501 107826 271535
rect 107864 271501 107892 271535
rect 107892 271501 107898 271535
rect 107936 271501 107960 271535
rect 107960 271501 107970 271535
rect 108008 271501 108028 271535
rect 108028 271501 108042 271535
rect 108080 271501 108096 271535
rect 108096 271501 108114 271535
rect 108152 271501 108164 271535
rect 108164 271501 108186 271535
rect 108224 271501 108232 271535
rect 108232 271501 108258 271535
rect 108296 271501 108300 271535
rect 108300 271501 108330 271535
rect 107101 271451 107135 271453
rect 107101 271419 107135 271451
rect 107101 271349 107135 271381
rect 107101 271347 107135 271349
rect 108411 271451 108445 271453
rect 108411 271419 108445 271451
rect 108411 271349 108445 271381
rect 108411 271347 108445 271349
rect 107216 271265 107246 271299
rect 107246 271265 107250 271299
rect 107288 271265 107314 271299
rect 107314 271265 107322 271299
rect 107360 271265 107382 271299
rect 107382 271265 107394 271299
rect 107432 271265 107450 271299
rect 107450 271265 107466 271299
rect 107504 271265 107518 271299
rect 107518 271265 107538 271299
rect 107576 271265 107586 271299
rect 107586 271265 107610 271299
rect 107648 271265 107654 271299
rect 107654 271265 107682 271299
rect 107720 271265 107722 271299
rect 107722 271265 107754 271299
rect 107792 271265 107824 271299
rect 107824 271265 107826 271299
rect 107864 271265 107892 271299
rect 107892 271265 107898 271299
rect 107936 271265 107960 271299
rect 107960 271265 107970 271299
rect 108008 271265 108028 271299
rect 108028 271265 108042 271299
rect 108080 271265 108096 271299
rect 108096 271265 108114 271299
rect 108152 271265 108164 271299
rect 108164 271265 108186 271299
rect 108224 271265 108232 271299
rect 108232 271265 108258 271299
rect 108296 271265 108300 271299
rect 108300 271265 108330 271299
rect 107216 271131 107246 271165
rect 107246 271131 107250 271165
rect 107288 271131 107314 271165
rect 107314 271131 107322 271165
rect 107360 271131 107382 271165
rect 107382 271131 107394 271165
rect 107432 271131 107450 271165
rect 107450 271131 107466 271165
rect 107504 271131 107518 271165
rect 107518 271131 107538 271165
rect 107576 271131 107586 271165
rect 107586 271131 107610 271165
rect 107648 271131 107654 271165
rect 107654 271131 107682 271165
rect 107720 271131 107722 271165
rect 107722 271131 107754 271165
rect 107792 271131 107824 271165
rect 107824 271131 107826 271165
rect 107864 271131 107892 271165
rect 107892 271131 107898 271165
rect 107936 271131 107960 271165
rect 107960 271131 107970 271165
rect 108008 271131 108028 271165
rect 108028 271131 108042 271165
rect 108080 271131 108096 271165
rect 108096 271131 108114 271165
rect 108152 271131 108164 271165
rect 108164 271131 108186 271165
rect 108224 271131 108232 271165
rect 108232 271131 108258 271165
rect 108296 271131 108300 271165
rect 108300 271131 108330 271165
rect 107101 271081 107135 271083
rect 107101 271049 107135 271081
rect 107101 270979 107135 271011
rect 107101 270977 107135 270979
rect 108411 271081 108445 271083
rect 108411 271049 108445 271081
rect 108411 270979 108445 271011
rect 108411 270977 108445 270979
rect 107216 270895 107246 270929
rect 107246 270895 107250 270929
rect 107288 270895 107314 270929
rect 107314 270895 107322 270929
rect 107360 270895 107382 270929
rect 107382 270895 107394 270929
rect 107432 270895 107450 270929
rect 107450 270895 107466 270929
rect 107504 270895 107518 270929
rect 107518 270895 107538 270929
rect 107576 270895 107586 270929
rect 107586 270895 107610 270929
rect 107648 270895 107654 270929
rect 107654 270895 107682 270929
rect 107720 270895 107722 270929
rect 107722 270895 107754 270929
rect 107792 270895 107824 270929
rect 107824 270895 107826 270929
rect 107864 270895 107892 270929
rect 107892 270895 107898 270929
rect 107936 270895 107960 270929
rect 107960 270895 107970 270929
rect 108008 270895 108028 270929
rect 108028 270895 108042 270929
rect 108080 270895 108096 270929
rect 108096 270895 108114 270929
rect 108152 270895 108164 270929
rect 108164 270895 108186 270929
rect 108224 270895 108232 270929
rect 108232 270895 108258 270929
rect 108296 270895 108300 270929
rect 108300 270895 108330 270929
rect 109009 270940 109043 270974
rect 109009 270868 109043 270902
rect 109458 272473 109492 272507
rect 109394 272399 109428 272411
rect 109394 272377 109428 272399
rect 109394 272331 109428 272339
rect 109394 272305 109428 272331
rect 109394 272263 109428 272267
rect 109394 272233 109428 272263
rect 109394 272161 109428 272195
rect 109394 272093 109428 272123
rect 109394 272089 109428 272093
rect 109394 272025 109428 272051
rect 109394 272017 109428 272025
rect 109394 271957 109428 271979
rect 109394 271945 109428 271957
rect 109394 271889 109428 271907
rect 109394 271873 109428 271889
rect 109394 271821 109428 271835
rect 109394 271801 109428 271821
rect 109394 271753 109428 271763
rect 109394 271729 109428 271753
rect 109394 271685 109428 271691
rect 109394 271657 109428 271685
rect 109394 271617 109428 271619
rect 109394 271585 109428 271617
rect 109394 271515 109428 271547
rect 109394 271513 109428 271515
rect 109394 271447 109428 271475
rect 109394 271441 109428 271447
rect 109394 271379 109428 271403
rect 109394 271369 109428 271379
rect 109394 271311 109428 271331
rect 109394 271297 109428 271311
rect 109394 271243 109428 271259
rect 109394 271225 109428 271243
rect 109394 271175 109428 271187
rect 109394 271153 109428 271175
rect 109394 271107 109428 271115
rect 109394 271081 109428 271107
rect 109394 271039 109428 271043
rect 109394 271009 109428 271039
rect 109394 270937 109428 270971
rect 109394 270869 109428 270899
rect 109394 270865 109428 270869
rect 109394 270801 109428 270827
rect 109394 270793 109428 270801
rect 109394 270733 109428 270755
rect 109394 270721 109428 270733
rect 109522 272399 109556 272411
rect 109522 272377 109556 272399
rect 109522 272331 109556 272339
rect 109522 272305 109556 272331
rect 109522 272263 109556 272267
rect 109522 272233 109556 272263
rect 109522 272161 109556 272195
rect 109522 272093 109556 272123
rect 109522 272089 109556 272093
rect 109522 272025 109556 272051
rect 109522 272017 109556 272025
rect 109522 271957 109556 271979
rect 109522 271945 109556 271957
rect 109522 271889 109556 271907
rect 109522 271873 109556 271889
rect 109522 271821 109556 271835
rect 109522 271801 109556 271821
rect 109522 271753 109556 271763
rect 109522 271729 109556 271753
rect 109522 271685 109556 271691
rect 109522 271657 109556 271685
rect 109522 271617 109556 271619
rect 109522 271585 109556 271617
rect 109522 271515 109556 271547
rect 109522 271513 109556 271515
rect 109522 271447 109556 271475
rect 109522 271441 109556 271447
rect 109522 271379 109556 271403
rect 109522 271369 109556 271379
rect 109522 271311 109556 271331
rect 109522 271297 109556 271311
rect 109522 271243 109556 271259
rect 109522 271225 109556 271243
rect 109522 271175 109556 271187
rect 109522 271153 109556 271175
rect 109522 271107 109556 271115
rect 109522 271081 109556 271107
rect 109522 271039 109556 271043
rect 109522 271009 109556 271039
rect 109522 270937 109556 270971
rect 109522 270869 109556 270899
rect 109522 270865 109556 270869
rect 109522 270801 109556 270827
rect 109522 270793 109556 270801
rect 109522 270733 109556 270755
rect 109522 270721 109556 270733
rect 109458 270625 109492 270659
rect 111553 280832 111581 280866
rect 111581 280832 111587 280866
rect 111625 280832 111649 280866
rect 111649 280832 111659 280866
rect 111697 280832 111717 280866
rect 111717 280832 111731 280866
rect 111769 280832 111785 280866
rect 111785 280832 111803 280866
rect 111841 280832 111853 280866
rect 111853 280832 111875 280866
rect 111913 280832 111921 280866
rect 111921 280832 111947 280866
rect 111985 280832 111989 280866
rect 111989 280832 112019 280866
rect 112057 280832 112091 280866
rect 112129 280832 112159 280866
rect 112159 280832 112163 280866
rect 112201 280832 112227 280866
rect 112227 280832 112235 280866
rect 112273 280832 112295 280866
rect 112295 280832 112307 280866
rect 112345 280832 112363 280866
rect 112363 280832 112379 280866
rect 112417 280832 112431 280866
rect 112431 280832 112451 280866
rect 112489 280832 112499 280866
rect 112499 280832 112523 280866
rect 112561 280832 112567 280866
rect 112567 280832 112595 280866
rect 111452 280791 111486 280793
rect 111452 280759 111486 280791
rect 111452 280689 111486 280721
rect 111452 280687 111486 280689
rect 112662 280791 112696 280793
rect 112662 280759 112696 280791
rect 112662 280689 112696 280721
rect 112662 280687 112696 280689
rect 111553 280614 111581 280648
rect 111581 280614 111587 280648
rect 111625 280614 111649 280648
rect 111649 280614 111659 280648
rect 111697 280614 111717 280648
rect 111717 280614 111731 280648
rect 111769 280614 111785 280648
rect 111785 280614 111803 280648
rect 111841 280614 111853 280648
rect 111853 280614 111875 280648
rect 111913 280614 111921 280648
rect 111921 280614 111947 280648
rect 111985 280614 111989 280648
rect 111989 280614 112019 280648
rect 112057 280614 112091 280648
rect 112129 280614 112159 280648
rect 112159 280614 112163 280648
rect 112201 280614 112227 280648
rect 112227 280614 112235 280648
rect 112273 280614 112295 280648
rect 112295 280614 112307 280648
rect 112345 280614 112363 280648
rect 112363 280614 112379 280648
rect 112417 280614 112431 280648
rect 112431 280614 112451 280648
rect 112489 280614 112499 280648
rect 112499 280614 112523 280648
rect 112561 280614 112567 280648
rect 112567 280614 112595 280648
rect 112999 280840 113027 280874
rect 113027 280840 113033 280874
rect 113071 280840 113095 280874
rect 113095 280840 113105 280874
rect 113143 280840 113163 280874
rect 113163 280840 113177 280874
rect 113215 280840 113231 280874
rect 113231 280840 113249 280874
rect 113287 280840 113299 280874
rect 113299 280840 113321 280874
rect 113359 280840 113367 280874
rect 113367 280840 113393 280874
rect 113431 280840 113435 280874
rect 113435 280840 113465 280874
rect 113503 280840 113537 280874
rect 113575 280840 113605 280874
rect 113605 280840 113609 280874
rect 113647 280840 113673 280874
rect 113673 280840 113681 280874
rect 113719 280840 113741 280874
rect 113741 280840 113753 280874
rect 113791 280840 113809 280874
rect 113809 280840 113825 280874
rect 113863 280840 113877 280874
rect 113877 280840 113897 280874
rect 113935 280840 113945 280874
rect 113945 280840 113969 280874
rect 114007 280840 114013 280874
rect 114013 280840 114041 280874
rect 112898 280779 112932 280781
rect 112898 280747 112932 280779
rect 112898 280677 112932 280709
rect 112898 280675 112932 280677
rect 114108 280779 114142 280781
rect 114108 280747 114142 280779
rect 114108 280677 114142 280709
rect 114108 280675 114142 280677
rect 114704 280815 114706 280849
rect 114706 280815 114738 280849
rect 114776 280815 114808 280849
rect 114808 280815 114810 280849
rect 112999 280582 113027 280616
rect 113027 280582 113033 280616
rect 113071 280582 113095 280616
rect 113095 280582 113105 280616
rect 113143 280582 113163 280616
rect 113163 280582 113177 280616
rect 113215 280582 113231 280616
rect 113231 280582 113249 280616
rect 113287 280582 113299 280616
rect 113299 280582 113321 280616
rect 113359 280582 113367 280616
rect 113367 280582 113393 280616
rect 113431 280582 113435 280616
rect 113435 280582 113465 280616
rect 113503 280582 113537 280616
rect 113575 280582 113605 280616
rect 113605 280582 113609 280616
rect 113647 280582 113673 280616
rect 113673 280582 113681 280616
rect 113719 280582 113741 280616
rect 113741 280582 113753 280616
rect 113791 280582 113809 280616
rect 113809 280582 113825 280616
rect 113863 280582 113877 280616
rect 113877 280582 113897 280616
rect 113935 280582 113945 280616
rect 113945 280582 113969 280616
rect 114007 280582 114013 280616
rect 114013 280582 114041 280616
rect 111553 280472 111581 280506
rect 111581 280472 111587 280506
rect 111625 280472 111649 280506
rect 111649 280472 111659 280506
rect 111697 280472 111717 280506
rect 111717 280472 111731 280506
rect 111769 280472 111785 280506
rect 111785 280472 111803 280506
rect 111841 280472 111853 280506
rect 111853 280472 111875 280506
rect 111913 280472 111921 280506
rect 111921 280472 111947 280506
rect 111985 280472 111989 280506
rect 111989 280472 112019 280506
rect 112057 280472 112091 280506
rect 112129 280472 112159 280506
rect 112159 280472 112163 280506
rect 112201 280472 112227 280506
rect 112227 280472 112235 280506
rect 112273 280472 112295 280506
rect 112295 280472 112307 280506
rect 112345 280472 112363 280506
rect 112363 280472 112379 280506
rect 112417 280472 112431 280506
rect 112431 280472 112451 280506
rect 112489 280472 112499 280506
rect 112499 280472 112523 280506
rect 112561 280472 112567 280506
rect 112567 280472 112595 280506
rect 111452 280431 111486 280433
rect 111452 280399 111486 280431
rect 111452 280329 111486 280361
rect 111452 280327 111486 280329
rect 112662 280431 112696 280433
rect 112662 280399 112696 280431
rect 112662 280329 112696 280361
rect 112662 280327 112696 280329
rect 111553 280254 111581 280288
rect 111581 280254 111587 280288
rect 111625 280254 111649 280288
rect 111649 280254 111659 280288
rect 111697 280254 111717 280288
rect 111717 280254 111731 280288
rect 111769 280254 111785 280288
rect 111785 280254 111803 280288
rect 111841 280254 111853 280288
rect 111853 280254 111875 280288
rect 111913 280254 111921 280288
rect 111921 280254 111947 280288
rect 111985 280254 111989 280288
rect 111989 280254 112019 280288
rect 112057 280254 112091 280288
rect 112129 280254 112159 280288
rect 112159 280254 112163 280288
rect 112201 280254 112227 280288
rect 112227 280254 112235 280288
rect 112273 280254 112295 280288
rect 112295 280254 112307 280288
rect 112345 280254 112363 280288
rect 112363 280254 112379 280288
rect 112417 280254 112431 280288
rect 112431 280254 112451 280288
rect 112489 280254 112499 280288
rect 112499 280254 112523 280288
rect 112561 280254 112567 280288
rect 112567 280254 112595 280288
rect 112999 280416 113027 280450
rect 113027 280416 113033 280450
rect 113071 280416 113095 280450
rect 113095 280416 113105 280450
rect 113143 280416 113163 280450
rect 113163 280416 113177 280450
rect 113215 280416 113231 280450
rect 113231 280416 113249 280450
rect 113287 280416 113299 280450
rect 113299 280416 113321 280450
rect 113359 280416 113367 280450
rect 113367 280416 113393 280450
rect 113431 280416 113435 280450
rect 113435 280416 113465 280450
rect 113503 280416 113537 280450
rect 113575 280416 113605 280450
rect 113605 280416 113609 280450
rect 113647 280416 113673 280450
rect 113673 280416 113681 280450
rect 113719 280416 113741 280450
rect 113741 280416 113753 280450
rect 113791 280416 113809 280450
rect 113809 280416 113825 280450
rect 113863 280416 113877 280450
rect 113877 280416 113897 280450
rect 113935 280416 113945 280450
rect 113945 280416 113969 280450
rect 114007 280416 114013 280450
rect 114013 280416 114041 280450
rect 112898 280355 112932 280357
rect 112898 280323 112932 280355
rect 112898 280253 112932 280285
rect 112898 280251 112932 280253
rect 114108 280355 114142 280357
rect 114108 280323 114142 280355
rect 114108 280253 114142 280285
rect 114108 280251 114142 280253
rect 112999 280158 113027 280192
rect 113027 280158 113033 280192
rect 113071 280158 113095 280192
rect 113095 280158 113105 280192
rect 113143 280158 113163 280192
rect 113163 280158 113177 280192
rect 113215 280158 113231 280192
rect 113231 280158 113249 280192
rect 113287 280158 113299 280192
rect 113299 280158 113321 280192
rect 113359 280158 113367 280192
rect 113367 280158 113393 280192
rect 113431 280158 113435 280192
rect 113435 280158 113465 280192
rect 113503 280158 113537 280192
rect 113575 280158 113605 280192
rect 113605 280158 113609 280192
rect 113647 280158 113673 280192
rect 113673 280158 113681 280192
rect 113719 280158 113741 280192
rect 113741 280158 113753 280192
rect 113791 280158 113809 280192
rect 113809 280158 113825 280192
rect 113863 280158 113877 280192
rect 113877 280158 113897 280192
rect 113935 280158 113945 280192
rect 113945 280158 113969 280192
rect 114007 280158 114013 280192
rect 114013 280158 114041 280192
rect 111553 280112 111581 280146
rect 111581 280112 111587 280146
rect 111625 280112 111649 280146
rect 111649 280112 111659 280146
rect 111697 280112 111717 280146
rect 111717 280112 111731 280146
rect 111769 280112 111785 280146
rect 111785 280112 111803 280146
rect 111841 280112 111853 280146
rect 111853 280112 111875 280146
rect 111913 280112 111921 280146
rect 111921 280112 111947 280146
rect 111985 280112 111989 280146
rect 111989 280112 112019 280146
rect 112057 280112 112091 280146
rect 112129 280112 112159 280146
rect 112159 280112 112163 280146
rect 112201 280112 112227 280146
rect 112227 280112 112235 280146
rect 112273 280112 112295 280146
rect 112295 280112 112307 280146
rect 112345 280112 112363 280146
rect 112363 280112 112379 280146
rect 112417 280112 112431 280146
rect 112431 280112 112451 280146
rect 112489 280112 112499 280146
rect 112499 280112 112523 280146
rect 112561 280112 112567 280146
rect 112567 280112 112595 280146
rect 111452 280071 111486 280073
rect 111452 280039 111486 280071
rect 111452 279969 111486 280001
rect 111452 279967 111486 279969
rect 112662 280071 112696 280073
rect 112662 280039 112696 280071
rect 112662 279969 112696 280001
rect 112662 279967 112696 279969
rect 111553 279894 111581 279928
rect 111581 279894 111587 279928
rect 111625 279894 111649 279928
rect 111649 279894 111659 279928
rect 111697 279894 111717 279928
rect 111717 279894 111731 279928
rect 111769 279894 111785 279928
rect 111785 279894 111803 279928
rect 111841 279894 111853 279928
rect 111853 279894 111875 279928
rect 111913 279894 111921 279928
rect 111921 279894 111947 279928
rect 111985 279894 111989 279928
rect 111989 279894 112019 279928
rect 112057 279894 112091 279928
rect 112129 279894 112159 279928
rect 112159 279894 112163 279928
rect 112201 279894 112227 279928
rect 112227 279894 112235 279928
rect 112273 279894 112295 279928
rect 112295 279894 112307 279928
rect 112345 279894 112363 279928
rect 112363 279894 112379 279928
rect 112417 279894 112431 279928
rect 112431 279894 112451 279928
rect 112489 279894 112499 279928
rect 112499 279894 112523 279928
rect 112561 279894 112567 279928
rect 112567 279894 112595 279928
rect 113029 280014 113057 280048
rect 113057 280014 113063 280048
rect 113101 280014 113125 280048
rect 113125 280014 113135 280048
rect 113173 280014 113193 280048
rect 113193 280014 113207 280048
rect 113245 280014 113261 280048
rect 113261 280014 113279 280048
rect 113317 280014 113329 280048
rect 113329 280014 113351 280048
rect 113389 280014 113397 280048
rect 113397 280014 113423 280048
rect 113461 280014 113465 280048
rect 113465 280014 113495 280048
rect 113533 280014 113567 280048
rect 113605 280014 113635 280048
rect 113635 280014 113639 280048
rect 113677 280014 113703 280048
rect 113703 280014 113711 280048
rect 113749 280014 113771 280048
rect 113771 280014 113783 280048
rect 113821 280014 113839 280048
rect 113839 280014 113855 280048
rect 113893 280014 113907 280048
rect 113907 280014 113927 280048
rect 113965 280014 113975 280048
rect 113975 280014 113999 280048
rect 114037 280014 114043 280048
rect 114043 280014 114071 280048
rect 112928 279945 112962 279979
rect 114138 279945 114172 279979
rect 114342 279917 114376 279951
rect 113029 279876 113057 279910
rect 113057 279876 113063 279910
rect 113101 279876 113125 279910
rect 113125 279876 113135 279910
rect 113173 279876 113193 279910
rect 113193 279876 113207 279910
rect 113245 279876 113261 279910
rect 113261 279876 113279 279910
rect 113317 279876 113329 279910
rect 113329 279876 113351 279910
rect 113389 279876 113397 279910
rect 113397 279876 113423 279910
rect 113461 279876 113465 279910
rect 113465 279876 113495 279910
rect 113533 279876 113567 279910
rect 113605 279876 113635 279910
rect 113635 279876 113639 279910
rect 113677 279876 113703 279910
rect 113703 279876 113711 279910
rect 113749 279876 113771 279910
rect 113771 279876 113783 279910
rect 113821 279876 113839 279910
rect 113839 279876 113855 279910
rect 113893 279876 113907 279910
rect 113907 279876 113927 279910
rect 113965 279876 113975 279910
rect 113975 279876 113999 279910
rect 114037 279876 114043 279910
rect 114043 279876 114071 279910
rect 114576 280756 114610 280764
rect 114576 280730 114610 280756
rect 114576 280688 114610 280692
rect 114576 280658 114610 280688
rect 114576 280586 114610 280620
rect 114576 280518 114610 280548
rect 114576 280514 114610 280518
rect 114576 280450 114610 280476
rect 114576 280442 114610 280450
rect 114904 280756 114938 280764
rect 114904 280730 114938 280756
rect 114904 280688 114938 280692
rect 114904 280658 114938 280688
rect 114904 280586 114938 280620
rect 114904 280518 114938 280548
rect 114904 280514 114938 280518
rect 114904 280450 114938 280476
rect 114904 280442 114938 280450
rect 114704 280357 114706 280391
rect 114706 280357 114738 280391
rect 114776 280357 114808 280391
rect 114808 280357 114810 280391
rect 115395 280815 115397 280849
rect 115397 280815 115429 280849
rect 115467 280815 115499 280849
rect 115499 280815 115501 280849
rect 114899 280243 114933 280277
rect 115267 280756 115301 280764
rect 115267 280730 115301 280756
rect 115267 280688 115301 280692
rect 115267 280658 115301 280688
rect 115267 280586 115301 280620
rect 115267 280518 115301 280548
rect 115267 280514 115301 280518
rect 115267 280450 115301 280476
rect 115267 280442 115301 280450
rect 115595 280756 115629 280764
rect 115595 280730 115629 280756
rect 115595 280688 115629 280692
rect 115595 280658 115629 280688
rect 115595 280586 115629 280620
rect 115595 280518 115629 280548
rect 115595 280514 115629 280518
rect 115595 280450 115629 280476
rect 115595 280442 115629 280450
rect 115395 280357 115397 280391
rect 115397 280357 115429 280391
rect 115467 280357 115499 280391
rect 115499 280357 115501 280391
rect 114704 280129 114706 280163
rect 114706 280129 114738 280163
rect 114776 280129 114808 280163
rect 114808 280129 114810 280163
rect 114576 280088 114610 280090
rect 114576 280056 114610 280088
rect 114576 279986 114610 280018
rect 114576 279984 114610 279986
rect 114904 280088 114938 280090
rect 114904 280056 114938 280088
rect 114904 279986 114938 280018
rect 114904 279984 114938 279986
rect 115271 280243 115305 280277
rect 115395 280129 115397 280163
rect 115397 280129 115429 280163
rect 115467 280129 115499 280163
rect 115499 280129 115501 280163
rect 115267 280088 115301 280090
rect 115267 280056 115301 280088
rect 115267 279986 115301 280018
rect 115267 279984 115301 279986
rect 115595 280088 115629 280090
rect 115595 280056 115629 280088
rect 115595 279986 115629 280018
rect 115595 279984 115629 279986
rect 116164 280840 116192 280874
rect 116192 280840 116198 280874
rect 116236 280840 116260 280874
rect 116260 280840 116270 280874
rect 116308 280840 116328 280874
rect 116328 280840 116342 280874
rect 116380 280840 116396 280874
rect 116396 280840 116414 280874
rect 116452 280840 116464 280874
rect 116464 280840 116486 280874
rect 116524 280840 116532 280874
rect 116532 280840 116558 280874
rect 116596 280840 116600 280874
rect 116600 280840 116630 280874
rect 116668 280840 116702 280874
rect 116740 280840 116770 280874
rect 116770 280840 116774 280874
rect 116812 280840 116838 280874
rect 116838 280840 116846 280874
rect 116884 280840 116906 280874
rect 116906 280840 116918 280874
rect 116956 280840 116974 280874
rect 116974 280840 116990 280874
rect 117028 280840 117042 280874
rect 117042 280840 117062 280874
rect 117100 280840 117110 280874
rect 117110 280840 117134 280874
rect 117172 280840 117178 280874
rect 117178 280840 117206 280874
rect 116063 280779 116097 280781
rect 116063 280747 116097 280779
rect 116063 280677 116097 280709
rect 116063 280675 116097 280677
rect 117273 280779 117307 280781
rect 117273 280747 117307 280779
rect 117273 280677 117307 280709
rect 117273 280675 117307 280677
rect 116164 280582 116192 280616
rect 116192 280582 116198 280616
rect 116236 280582 116260 280616
rect 116260 280582 116270 280616
rect 116308 280582 116328 280616
rect 116328 280582 116342 280616
rect 116380 280582 116396 280616
rect 116396 280582 116414 280616
rect 116452 280582 116464 280616
rect 116464 280582 116486 280616
rect 116524 280582 116532 280616
rect 116532 280582 116558 280616
rect 116596 280582 116600 280616
rect 116600 280582 116630 280616
rect 116668 280582 116702 280616
rect 116740 280582 116770 280616
rect 116770 280582 116774 280616
rect 116812 280582 116838 280616
rect 116838 280582 116846 280616
rect 116884 280582 116906 280616
rect 116906 280582 116918 280616
rect 116956 280582 116974 280616
rect 116974 280582 116990 280616
rect 117028 280582 117042 280616
rect 117042 280582 117062 280616
rect 117100 280582 117110 280616
rect 117110 280582 117134 280616
rect 117172 280582 117178 280616
rect 117178 280582 117206 280616
rect 117610 280832 117638 280866
rect 117638 280832 117644 280866
rect 117682 280832 117706 280866
rect 117706 280832 117716 280866
rect 117754 280832 117774 280866
rect 117774 280832 117788 280866
rect 117826 280832 117842 280866
rect 117842 280832 117860 280866
rect 117898 280832 117910 280866
rect 117910 280832 117932 280866
rect 117970 280832 117978 280866
rect 117978 280832 118004 280866
rect 118042 280832 118046 280866
rect 118046 280832 118076 280866
rect 118114 280832 118148 280866
rect 118186 280832 118216 280866
rect 118216 280832 118220 280866
rect 118258 280832 118284 280866
rect 118284 280832 118292 280866
rect 118330 280832 118352 280866
rect 118352 280832 118364 280866
rect 118402 280832 118420 280866
rect 118420 280832 118436 280866
rect 118474 280832 118488 280866
rect 118488 280832 118508 280866
rect 118546 280832 118556 280866
rect 118556 280832 118580 280866
rect 118618 280832 118624 280866
rect 118624 280832 118652 280866
rect 117509 280791 117543 280793
rect 117509 280759 117543 280791
rect 117509 280689 117543 280721
rect 117509 280687 117543 280689
rect 118719 280791 118753 280793
rect 118719 280759 118753 280791
rect 118719 280689 118753 280721
rect 118719 280687 118753 280689
rect 117610 280614 117638 280648
rect 117638 280614 117644 280648
rect 117682 280614 117706 280648
rect 117706 280614 117716 280648
rect 117754 280614 117774 280648
rect 117774 280614 117788 280648
rect 117826 280614 117842 280648
rect 117842 280614 117860 280648
rect 117898 280614 117910 280648
rect 117910 280614 117932 280648
rect 117970 280614 117978 280648
rect 117978 280614 118004 280648
rect 118042 280614 118046 280648
rect 118046 280614 118076 280648
rect 118114 280614 118148 280648
rect 118186 280614 118216 280648
rect 118216 280614 118220 280648
rect 118258 280614 118284 280648
rect 118284 280614 118292 280648
rect 118330 280614 118352 280648
rect 118352 280614 118364 280648
rect 118402 280614 118420 280648
rect 118420 280614 118436 280648
rect 118474 280614 118488 280648
rect 118488 280614 118508 280648
rect 118546 280614 118556 280648
rect 118556 280614 118580 280648
rect 118618 280614 118624 280648
rect 118624 280614 118652 280648
rect 116164 280416 116192 280450
rect 116192 280416 116198 280450
rect 116236 280416 116260 280450
rect 116260 280416 116270 280450
rect 116308 280416 116328 280450
rect 116328 280416 116342 280450
rect 116380 280416 116396 280450
rect 116396 280416 116414 280450
rect 116452 280416 116464 280450
rect 116464 280416 116486 280450
rect 116524 280416 116532 280450
rect 116532 280416 116558 280450
rect 116596 280416 116600 280450
rect 116600 280416 116630 280450
rect 116668 280416 116702 280450
rect 116740 280416 116770 280450
rect 116770 280416 116774 280450
rect 116812 280416 116838 280450
rect 116838 280416 116846 280450
rect 116884 280416 116906 280450
rect 116906 280416 116918 280450
rect 116956 280416 116974 280450
rect 116974 280416 116990 280450
rect 117028 280416 117042 280450
rect 117042 280416 117062 280450
rect 117100 280416 117110 280450
rect 117110 280416 117134 280450
rect 117172 280416 117178 280450
rect 117178 280416 117206 280450
rect 116063 280355 116097 280357
rect 116063 280323 116097 280355
rect 116063 280253 116097 280285
rect 116063 280251 116097 280253
rect 117273 280355 117307 280357
rect 117273 280323 117307 280355
rect 117273 280253 117307 280285
rect 117273 280251 117307 280253
rect 116164 280158 116192 280192
rect 116192 280158 116198 280192
rect 116236 280158 116260 280192
rect 116260 280158 116270 280192
rect 116308 280158 116328 280192
rect 116328 280158 116342 280192
rect 116380 280158 116396 280192
rect 116396 280158 116414 280192
rect 116452 280158 116464 280192
rect 116464 280158 116486 280192
rect 116524 280158 116532 280192
rect 116532 280158 116558 280192
rect 116596 280158 116600 280192
rect 116600 280158 116630 280192
rect 116668 280158 116702 280192
rect 116740 280158 116770 280192
rect 116770 280158 116774 280192
rect 116812 280158 116838 280192
rect 116838 280158 116846 280192
rect 116884 280158 116906 280192
rect 116906 280158 116918 280192
rect 116956 280158 116974 280192
rect 116974 280158 116990 280192
rect 117028 280158 117042 280192
rect 117042 280158 117062 280192
rect 117100 280158 117110 280192
rect 117110 280158 117134 280192
rect 117172 280158 117178 280192
rect 117178 280158 117206 280192
rect 117610 280472 117638 280506
rect 117638 280472 117644 280506
rect 117682 280472 117706 280506
rect 117706 280472 117716 280506
rect 117754 280472 117774 280506
rect 117774 280472 117788 280506
rect 117826 280472 117842 280506
rect 117842 280472 117860 280506
rect 117898 280472 117910 280506
rect 117910 280472 117932 280506
rect 117970 280472 117978 280506
rect 117978 280472 118004 280506
rect 118042 280472 118046 280506
rect 118046 280472 118076 280506
rect 118114 280472 118148 280506
rect 118186 280472 118216 280506
rect 118216 280472 118220 280506
rect 118258 280472 118284 280506
rect 118284 280472 118292 280506
rect 118330 280472 118352 280506
rect 118352 280472 118364 280506
rect 118402 280472 118420 280506
rect 118420 280472 118436 280506
rect 118474 280472 118488 280506
rect 118488 280472 118508 280506
rect 118546 280472 118556 280506
rect 118556 280472 118580 280506
rect 118618 280472 118624 280506
rect 118624 280472 118652 280506
rect 117509 280431 117543 280433
rect 117509 280399 117543 280431
rect 117509 280329 117543 280361
rect 117509 280327 117543 280329
rect 118719 280431 118753 280433
rect 118719 280399 118753 280431
rect 118719 280329 118753 280361
rect 118719 280327 118753 280329
rect 117610 280254 117638 280288
rect 117638 280254 117644 280288
rect 117682 280254 117706 280288
rect 117706 280254 117716 280288
rect 117754 280254 117774 280288
rect 117774 280254 117788 280288
rect 117826 280254 117842 280288
rect 117842 280254 117860 280288
rect 117898 280254 117910 280288
rect 117910 280254 117932 280288
rect 117970 280254 117978 280288
rect 117978 280254 118004 280288
rect 118042 280254 118046 280288
rect 118046 280254 118076 280288
rect 118114 280254 118148 280288
rect 118186 280254 118216 280288
rect 118216 280254 118220 280288
rect 118258 280254 118284 280288
rect 118284 280254 118292 280288
rect 118330 280254 118352 280288
rect 118352 280254 118364 280288
rect 118402 280254 118420 280288
rect 118420 280254 118436 280288
rect 118474 280254 118488 280288
rect 118488 280254 118508 280288
rect 118546 280254 118556 280288
rect 118556 280254 118580 280288
rect 118618 280254 118624 280288
rect 118624 280254 118652 280288
rect 111553 279752 111581 279786
rect 111581 279752 111587 279786
rect 111625 279752 111649 279786
rect 111649 279752 111659 279786
rect 111697 279752 111717 279786
rect 111717 279752 111731 279786
rect 111769 279752 111785 279786
rect 111785 279752 111803 279786
rect 111841 279752 111853 279786
rect 111853 279752 111875 279786
rect 111913 279752 111921 279786
rect 111921 279752 111947 279786
rect 111985 279752 111989 279786
rect 111989 279752 112019 279786
rect 112057 279752 112091 279786
rect 112129 279752 112159 279786
rect 112159 279752 112163 279786
rect 112201 279752 112227 279786
rect 112227 279752 112235 279786
rect 112273 279752 112295 279786
rect 112295 279752 112307 279786
rect 112345 279752 112363 279786
rect 112363 279752 112379 279786
rect 112417 279752 112431 279786
rect 112431 279752 112451 279786
rect 112489 279752 112499 279786
rect 112499 279752 112523 279786
rect 112561 279752 112567 279786
rect 112567 279752 112595 279786
rect 111452 279711 111486 279713
rect 111452 279679 111486 279711
rect 111452 279609 111486 279641
rect 111452 279607 111486 279609
rect 113029 279716 113057 279750
rect 113057 279716 113063 279750
rect 113101 279716 113125 279750
rect 113125 279716 113135 279750
rect 113173 279716 113193 279750
rect 113193 279716 113207 279750
rect 113245 279716 113261 279750
rect 113261 279716 113279 279750
rect 113317 279716 113329 279750
rect 113329 279716 113351 279750
rect 113389 279716 113397 279750
rect 113397 279716 113423 279750
rect 113461 279716 113465 279750
rect 113465 279716 113495 279750
rect 113533 279716 113567 279750
rect 113605 279716 113635 279750
rect 113635 279716 113639 279750
rect 113677 279716 113703 279750
rect 113703 279716 113711 279750
rect 113749 279716 113771 279750
rect 113771 279716 113783 279750
rect 113821 279716 113839 279750
rect 113839 279716 113855 279750
rect 113893 279716 113907 279750
rect 113907 279716 113927 279750
rect 113965 279716 113975 279750
rect 113975 279716 113999 279750
rect 114037 279716 114043 279750
rect 114043 279716 114071 279750
rect 112662 279711 112696 279713
rect 112662 279679 112696 279711
rect 112662 279609 112696 279641
rect 112928 279647 112962 279681
rect 114138 279647 114172 279681
rect 112662 279607 112696 279609
rect 113029 279578 113057 279612
rect 113057 279578 113063 279612
rect 113101 279578 113125 279612
rect 113125 279578 113135 279612
rect 113173 279578 113193 279612
rect 113193 279578 113207 279612
rect 113245 279578 113261 279612
rect 113261 279578 113279 279612
rect 113317 279578 113329 279612
rect 113329 279578 113351 279612
rect 113389 279578 113397 279612
rect 113397 279578 113423 279612
rect 113461 279578 113465 279612
rect 113465 279578 113495 279612
rect 113533 279578 113567 279612
rect 113605 279578 113635 279612
rect 113635 279578 113639 279612
rect 113677 279578 113703 279612
rect 113703 279578 113711 279612
rect 113749 279578 113771 279612
rect 113771 279578 113783 279612
rect 113821 279578 113839 279612
rect 113839 279578 113855 279612
rect 113893 279578 113907 279612
rect 113907 279578 113927 279612
rect 113965 279578 113975 279612
rect 113975 279578 113999 279612
rect 114037 279578 114043 279612
rect 114043 279578 114071 279612
rect 114704 279911 114706 279945
rect 114706 279911 114738 279945
rect 114776 279911 114808 279945
rect 114808 279911 114810 279945
rect 111553 279534 111581 279568
rect 111581 279534 111587 279568
rect 111625 279534 111649 279568
rect 111649 279534 111659 279568
rect 111697 279534 111717 279568
rect 111717 279534 111731 279568
rect 111769 279534 111785 279568
rect 111785 279534 111803 279568
rect 111841 279534 111853 279568
rect 111853 279534 111875 279568
rect 111913 279534 111921 279568
rect 111921 279534 111947 279568
rect 111985 279534 111989 279568
rect 111989 279534 112019 279568
rect 112057 279534 112091 279568
rect 112129 279534 112159 279568
rect 112159 279534 112163 279568
rect 112201 279534 112227 279568
rect 112227 279534 112235 279568
rect 112273 279534 112295 279568
rect 112295 279534 112307 279568
rect 112345 279534 112363 279568
rect 112363 279534 112379 279568
rect 112417 279534 112431 279568
rect 112431 279534 112451 279568
rect 112489 279534 112499 279568
rect 112499 279534 112523 279568
rect 112561 279534 112567 279568
rect 112567 279534 112595 279568
rect 114899 279820 114933 279854
rect 115395 279911 115397 279945
rect 115397 279911 115429 279945
rect 115467 279911 115499 279945
rect 115499 279911 115501 279945
rect 114704 279721 114706 279755
rect 114706 279721 114738 279755
rect 114776 279721 114808 279755
rect 114808 279721 114810 279755
rect 114576 279680 114610 279682
rect 114576 279648 114610 279680
rect 114576 279578 114610 279610
rect 114576 279576 114610 279578
rect 114904 279680 114938 279682
rect 114904 279648 114938 279680
rect 114904 279578 114938 279610
rect 114904 279576 114938 279578
rect 115271 279820 115305 279854
rect 115395 279721 115397 279755
rect 115397 279721 115429 279755
rect 115467 279721 115499 279755
rect 115499 279721 115501 279755
rect 115267 279680 115301 279682
rect 115267 279648 115301 279680
rect 115267 279578 115301 279610
rect 115267 279576 115301 279578
rect 115595 279680 115629 279682
rect 115595 279648 115629 279680
rect 115595 279578 115629 279610
rect 115595 279576 115629 279578
rect 116134 280014 116162 280048
rect 116162 280014 116168 280048
rect 116206 280014 116230 280048
rect 116230 280014 116240 280048
rect 116278 280014 116298 280048
rect 116298 280014 116312 280048
rect 116350 280014 116366 280048
rect 116366 280014 116384 280048
rect 116422 280014 116434 280048
rect 116434 280014 116456 280048
rect 116494 280014 116502 280048
rect 116502 280014 116528 280048
rect 116566 280014 116570 280048
rect 116570 280014 116600 280048
rect 116638 280014 116672 280048
rect 116710 280014 116740 280048
rect 116740 280014 116744 280048
rect 116782 280014 116808 280048
rect 116808 280014 116816 280048
rect 116854 280014 116876 280048
rect 116876 280014 116888 280048
rect 116926 280014 116944 280048
rect 116944 280014 116960 280048
rect 116998 280014 117012 280048
rect 117012 280014 117032 280048
rect 117070 280014 117080 280048
rect 117080 280014 117104 280048
rect 117142 280014 117148 280048
rect 117148 280014 117176 280048
rect 115828 279917 115862 279951
rect 116033 279945 116067 279979
rect 117243 279945 117277 279979
rect 116134 279876 116162 279910
rect 116162 279876 116168 279910
rect 116206 279876 116230 279910
rect 116230 279876 116240 279910
rect 116278 279876 116298 279910
rect 116298 279876 116312 279910
rect 116350 279876 116366 279910
rect 116366 279876 116384 279910
rect 116422 279876 116434 279910
rect 116434 279876 116456 279910
rect 116494 279876 116502 279910
rect 116502 279876 116528 279910
rect 116566 279876 116570 279910
rect 116570 279876 116600 279910
rect 116638 279876 116672 279910
rect 116710 279876 116740 279910
rect 116740 279876 116744 279910
rect 116782 279876 116808 279910
rect 116808 279876 116816 279910
rect 116854 279876 116876 279910
rect 116876 279876 116888 279910
rect 116926 279876 116944 279910
rect 116944 279876 116960 279910
rect 116998 279876 117012 279910
rect 117012 279876 117032 279910
rect 117070 279876 117080 279910
rect 117080 279876 117104 279910
rect 117142 279876 117148 279910
rect 117148 279876 117176 279910
rect 117610 280112 117638 280146
rect 117638 280112 117644 280146
rect 117682 280112 117706 280146
rect 117706 280112 117716 280146
rect 117754 280112 117774 280146
rect 117774 280112 117788 280146
rect 117826 280112 117842 280146
rect 117842 280112 117860 280146
rect 117898 280112 117910 280146
rect 117910 280112 117932 280146
rect 117970 280112 117978 280146
rect 117978 280112 118004 280146
rect 118042 280112 118046 280146
rect 118046 280112 118076 280146
rect 118114 280112 118148 280146
rect 118186 280112 118216 280146
rect 118216 280112 118220 280146
rect 118258 280112 118284 280146
rect 118284 280112 118292 280146
rect 118330 280112 118352 280146
rect 118352 280112 118364 280146
rect 118402 280112 118420 280146
rect 118420 280112 118436 280146
rect 118474 280112 118488 280146
rect 118488 280112 118508 280146
rect 118546 280112 118556 280146
rect 118556 280112 118580 280146
rect 118618 280112 118624 280146
rect 118624 280112 118652 280146
rect 117509 280071 117543 280073
rect 117509 280039 117543 280071
rect 117509 279969 117543 280001
rect 117509 279967 117543 279969
rect 118719 280071 118753 280073
rect 118719 280039 118753 280071
rect 118719 279969 118753 280001
rect 118719 279967 118753 279969
rect 117610 279894 117638 279928
rect 117638 279894 117644 279928
rect 117682 279894 117706 279928
rect 117706 279894 117716 279928
rect 117754 279894 117774 279928
rect 117774 279894 117788 279928
rect 117826 279894 117842 279928
rect 117842 279894 117860 279928
rect 117898 279894 117910 279928
rect 117910 279894 117932 279928
rect 117970 279894 117978 279928
rect 117978 279894 118004 279928
rect 118042 279894 118046 279928
rect 118046 279894 118076 279928
rect 118114 279894 118148 279928
rect 118186 279894 118216 279928
rect 118216 279894 118220 279928
rect 118258 279894 118284 279928
rect 118284 279894 118292 279928
rect 118330 279894 118352 279928
rect 118352 279894 118364 279928
rect 118402 279894 118420 279928
rect 118420 279894 118436 279928
rect 118474 279894 118488 279928
rect 118488 279894 118508 279928
rect 118546 279894 118556 279928
rect 118556 279894 118580 279928
rect 118618 279894 118624 279928
rect 118624 279894 118652 279928
rect 117610 279752 117638 279786
rect 117638 279752 117644 279786
rect 117682 279752 117706 279786
rect 117706 279752 117716 279786
rect 117754 279752 117774 279786
rect 117774 279752 117788 279786
rect 117826 279752 117842 279786
rect 117842 279752 117860 279786
rect 117898 279752 117910 279786
rect 117910 279752 117932 279786
rect 117970 279752 117978 279786
rect 117978 279752 118004 279786
rect 118042 279752 118046 279786
rect 118046 279752 118076 279786
rect 118114 279752 118148 279786
rect 118186 279752 118216 279786
rect 118216 279752 118220 279786
rect 118258 279752 118284 279786
rect 118284 279752 118292 279786
rect 118330 279752 118352 279786
rect 118352 279752 118364 279786
rect 118402 279752 118420 279786
rect 118420 279752 118436 279786
rect 118474 279752 118488 279786
rect 118488 279752 118508 279786
rect 118546 279752 118556 279786
rect 118556 279752 118580 279786
rect 118618 279752 118624 279786
rect 118624 279752 118652 279786
rect 116134 279716 116162 279750
rect 116162 279716 116168 279750
rect 116206 279716 116230 279750
rect 116230 279716 116240 279750
rect 116278 279716 116298 279750
rect 116298 279716 116312 279750
rect 116350 279716 116366 279750
rect 116366 279716 116384 279750
rect 116422 279716 116434 279750
rect 116434 279716 116456 279750
rect 116494 279716 116502 279750
rect 116502 279716 116528 279750
rect 116566 279716 116570 279750
rect 116570 279716 116600 279750
rect 116638 279716 116672 279750
rect 116710 279716 116740 279750
rect 116740 279716 116744 279750
rect 116782 279716 116808 279750
rect 116808 279716 116816 279750
rect 116854 279716 116876 279750
rect 116876 279716 116888 279750
rect 116926 279716 116944 279750
rect 116944 279716 116960 279750
rect 116998 279716 117012 279750
rect 117012 279716 117032 279750
rect 117070 279716 117080 279750
rect 117080 279716 117104 279750
rect 117142 279716 117148 279750
rect 117148 279716 117176 279750
rect 117509 279711 117543 279713
rect 116033 279647 116067 279681
rect 117243 279647 117277 279681
rect 117509 279679 117543 279711
rect 116134 279578 116162 279612
rect 116162 279578 116168 279612
rect 116206 279578 116230 279612
rect 116230 279578 116240 279612
rect 116278 279578 116298 279612
rect 116298 279578 116312 279612
rect 116350 279578 116366 279612
rect 116366 279578 116384 279612
rect 116422 279578 116434 279612
rect 116434 279578 116456 279612
rect 116494 279578 116502 279612
rect 116502 279578 116528 279612
rect 116566 279578 116570 279612
rect 116570 279578 116600 279612
rect 116638 279578 116672 279612
rect 116710 279578 116740 279612
rect 116740 279578 116744 279612
rect 116782 279578 116808 279612
rect 116808 279578 116816 279612
rect 116854 279578 116876 279612
rect 116876 279578 116888 279612
rect 116926 279578 116944 279612
rect 116944 279578 116960 279612
rect 116998 279578 117012 279612
rect 117012 279578 117032 279612
rect 117070 279578 117080 279612
rect 117080 279578 117104 279612
rect 117142 279578 117148 279612
rect 117148 279578 117176 279612
rect 117509 279609 117543 279641
rect 117509 279607 117543 279609
rect 118719 279711 118753 279713
rect 118719 279679 118753 279711
rect 118719 279609 118753 279641
rect 118719 279607 118753 279609
rect 114704 279503 114706 279537
rect 114706 279503 114738 279537
rect 114776 279503 114808 279537
rect 114808 279503 114810 279537
rect 115395 279503 115397 279537
rect 115397 279503 115429 279537
rect 115467 279503 115499 279537
rect 115499 279503 115501 279537
rect 117610 279534 117638 279568
rect 117638 279534 117644 279568
rect 117682 279534 117706 279568
rect 117706 279534 117716 279568
rect 117754 279534 117774 279568
rect 117774 279534 117788 279568
rect 117826 279534 117842 279568
rect 117842 279534 117860 279568
rect 117898 279534 117910 279568
rect 117910 279534 117932 279568
rect 117970 279534 117978 279568
rect 117978 279534 118004 279568
rect 118042 279534 118046 279568
rect 118046 279534 118076 279568
rect 118114 279534 118148 279568
rect 118186 279534 118216 279568
rect 118216 279534 118220 279568
rect 118258 279534 118284 279568
rect 118284 279534 118292 279568
rect 118330 279534 118352 279568
rect 118352 279534 118364 279568
rect 118402 279534 118420 279568
rect 118420 279534 118436 279568
rect 118474 279534 118488 279568
rect 118488 279534 118508 279568
rect 118546 279534 118556 279568
rect 118556 279534 118580 279568
rect 118618 279534 118624 279568
rect 118624 279534 118652 279568
rect 114034 279397 114068 279399
rect 114106 279397 114140 279399
rect 114178 279397 114212 279399
rect 114034 279365 114060 279397
rect 114060 279365 114068 279397
rect 114106 279365 114128 279397
rect 114128 279365 114140 279397
rect 114178 279365 114196 279397
rect 114196 279365 114212 279397
rect 115992 279397 116026 279399
rect 116064 279397 116098 279399
rect 116136 279397 116170 279399
rect 115992 279365 116009 279397
rect 116009 279365 116026 279397
rect 116064 279365 116077 279397
rect 116077 279365 116098 279397
rect 116136 279365 116145 279397
rect 116145 279365 116170 279397
rect 111553 279166 111581 279200
rect 111581 279166 111587 279200
rect 111625 279166 111649 279200
rect 111649 279166 111659 279200
rect 111697 279166 111717 279200
rect 111717 279166 111731 279200
rect 111769 279166 111785 279200
rect 111785 279166 111803 279200
rect 111841 279166 111853 279200
rect 111853 279166 111875 279200
rect 111913 279166 111921 279200
rect 111921 279166 111947 279200
rect 111985 279166 111989 279200
rect 111989 279166 112019 279200
rect 112057 279166 112091 279200
rect 112129 279166 112159 279200
rect 112159 279166 112163 279200
rect 112201 279166 112227 279200
rect 112227 279166 112235 279200
rect 112273 279166 112295 279200
rect 112295 279166 112307 279200
rect 112345 279166 112363 279200
rect 112363 279166 112379 279200
rect 112417 279166 112431 279200
rect 112431 279166 112451 279200
rect 112489 279166 112499 279200
rect 112499 279166 112523 279200
rect 112561 279166 112567 279200
rect 112567 279166 112595 279200
rect 111452 279125 111486 279127
rect 111452 279093 111486 279125
rect 111452 279023 111486 279055
rect 111452 279021 111486 279023
rect 112662 279125 112696 279127
rect 112662 279093 112696 279125
rect 112662 279023 112696 279055
rect 112662 279021 112696 279023
rect 111553 278948 111581 278982
rect 111581 278948 111587 278982
rect 111625 278948 111649 278982
rect 111649 278948 111659 278982
rect 111697 278948 111717 278982
rect 111717 278948 111731 278982
rect 111769 278948 111785 278982
rect 111785 278948 111803 278982
rect 111841 278948 111853 278982
rect 111853 278948 111875 278982
rect 111913 278948 111921 278982
rect 111921 278948 111947 278982
rect 111985 278948 111989 278982
rect 111989 278948 112019 278982
rect 112057 278948 112091 278982
rect 112129 278948 112159 278982
rect 112159 278948 112163 278982
rect 112201 278948 112227 278982
rect 112227 278948 112235 278982
rect 112273 278948 112295 278982
rect 112295 278948 112307 278982
rect 112345 278948 112363 278982
rect 112363 278948 112379 278982
rect 112417 278948 112431 278982
rect 112431 278948 112451 278982
rect 112489 278948 112499 278982
rect 112499 278948 112523 278982
rect 112561 278948 112567 278982
rect 112567 278948 112595 278982
rect 112999 279174 113027 279208
rect 113027 279174 113033 279208
rect 113071 279174 113095 279208
rect 113095 279174 113105 279208
rect 113143 279174 113163 279208
rect 113163 279174 113177 279208
rect 113215 279174 113231 279208
rect 113231 279174 113249 279208
rect 113287 279174 113299 279208
rect 113299 279174 113321 279208
rect 113359 279174 113367 279208
rect 113367 279174 113393 279208
rect 113431 279174 113435 279208
rect 113435 279174 113465 279208
rect 113503 279174 113537 279208
rect 113575 279174 113605 279208
rect 113605 279174 113609 279208
rect 113647 279174 113673 279208
rect 113673 279174 113681 279208
rect 113719 279174 113741 279208
rect 113741 279174 113753 279208
rect 113791 279174 113809 279208
rect 113809 279174 113825 279208
rect 113863 279174 113877 279208
rect 113877 279174 113897 279208
rect 113935 279174 113945 279208
rect 113945 279174 113969 279208
rect 114007 279174 114013 279208
rect 114013 279174 114041 279208
rect 112898 279113 112932 279115
rect 112898 279081 112932 279113
rect 112898 279011 112932 279043
rect 112898 279009 112932 279011
rect 114108 279113 114142 279115
rect 114108 279081 114142 279113
rect 114108 279011 114142 279043
rect 114108 279009 114142 279011
rect 114704 279149 114706 279183
rect 114706 279149 114738 279183
rect 114776 279149 114808 279183
rect 114808 279149 114810 279183
rect 112999 278916 113027 278950
rect 113027 278916 113033 278950
rect 113071 278916 113095 278950
rect 113095 278916 113105 278950
rect 113143 278916 113163 278950
rect 113163 278916 113177 278950
rect 113215 278916 113231 278950
rect 113231 278916 113249 278950
rect 113287 278916 113299 278950
rect 113299 278916 113321 278950
rect 113359 278916 113367 278950
rect 113367 278916 113393 278950
rect 113431 278916 113435 278950
rect 113435 278916 113465 278950
rect 113503 278916 113537 278950
rect 113575 278916 113605 278950
rect 113605 278916 113609 278950
rect 113647 278916 113673 278950
rect 113673 278916 113681 278950
rect 113719 278916 113741 278950
rect 113741 278916 113753 278950
rect 113791 278916 113809 278950
rect 113809 278916 113825 278950
rect 113863 278916 113877 278950
rect 113877 278916 113897 278950
rect 113935 278916 113945 278950
rect 113945 278916 113969 278950
rect 114007 278916 114013 278950
rect 114013 278916 114041 278950
rect 111553 278806 111581 278840
rect 111581 278806 111587 278840
rect 111625 278806 111649 278840
rect 111649 278806 111659 278840
rect 111697 278806 111717 278840
rect 111717 278806 111731 278840
rect 111769 278806 111785 278840
rect 111785 278806 111803 278840
rect 111841 278806 111853 278840
rect 111853 278806 111875 278840
rect 111913 278806 111921 278840
rect 111921 278806 111947 278840
rect 111985 278806 111989 278840
rect 111989 278806 112019 278840
rect 112057 278806 112091 278840
rect 112129 278806 112159 278840
rect 112159 278806 112163 278840
rect 112201 278806 112227 278840
rect 112227 278806 112235 278840
rect 112273 278806 112295 278840
rect 112295 278806 112307 278840
rect 112345 278806 112363 278840
rect 112363 278806 112379 278840
rect 112417 278806 112431 278840
rect 112431 278806 112451 278840
rect 112489 278806 112499 278840
rect 112499 278806 112523 278840
rect 112561 278806 112567 278840
rect 112567 278806 112595 278840
rect 111452 278765 111486 278767
rect 111452 278733 111486 278765
rect 111452 278663 111486 278695
rect 111452 278661 111486 278663
rect 112662 278765 112696 278767
rect 112662 278733 112696 278765
rect 112662 278663 112696 278695
rect 112662 278661 112696 278663
rect 111553 278588 111581 278622
rect 111581 278588 111587 278622
rect 111625 278588 111649 278622
rect 111649 278588 111659 278622
rect 111697 278588 111717 278622
rect 111717 278588 111731 278622
rect 111769 278588 111785 278622
rect 111785 278588 111803 278622
rect 111841 278588 111853 278622
rect 111853 278588 111875 278622
rect 111913 278588 111921 278622
rect 111921 278588 111947 278622
rect 111985 278588 111989 278622
rect 111989 278588 112019 278622
rect 112057 278588 112091 278622
rect 112129 278588 112159 278622
rect 112159 278588 112163 278622
rect 112201 278588 112227 278622
rect 112227 278588 112235 278622
rect 112273 278588 112295 278622
rect 112295 278588 112307 278622
rect 112345 278588 112363 278622
rect 112363 278588 112379 278622
rect 112417 278588 112431 278622
rect 112431 278588 112451 278622
rect 112489 278588 112499 278622
rect 112499 278588 112523 278622
rect 112561 278588 112567 278622
rect 112567 278588 112595 278622
rect 112999 278750 113027 278784
rect 113027 278750 113033 278784
rect 113071 278750 113095 278784
rect 113095 278750 113105 278784
rect 113143 278750 113163 278784
rect 113163 278750 113177 278784
rect 113215 278750 113231 278784
rect 113231 278750 113249 278784
rect 113287 278750 113299 278784
rect 113299 278750 113321 278784
rect 113359 278750 113367 278784
rect 113367 278750 113393 278784
rect 113431 278750 113435 278784
rect 113435 278750 113465 278784
rect 113503 278750 113537 278784
rect 113575 278750 113605 278784
rect 113605 278750 113609 278784
rect 113647 278750 113673 278784
rect 113673 278750 113681 278784
rect 113719 278750 113741 278784
rect 113741 278750 113753 278784
rect 113791 278750 113809 278784
rect 113809 278750 113825 278784
rect 113863 278750 113877 278784
rect 113877 278750 113897 278784
rect 113935 278750 113945 278784
rect 113945 278750 113969 278784
rect 114007 278750 114013 278784
rect 114013 278750 114041 278784
rect 112898 278689 112932 278691
rect 112898 278657 112932 278689
rect 112898 278587 112932 278619
rect 112898 278585 112932 278587
rect 114108 278689 114142 278691
rect 114108 278657 114142 278689
rect 114108 278587 114142 278619
rect 114108 278585 114142 278587
rect 112999 278492 113027 278526
rect 113027 278492 113033 278526
rect 113071 278492 113095 278526
rect 113095 278492 113105 278526
rect 113143 278492 113163 278526
rect 113163 278492 113177 278526
rect 113215 278492 113231 278526
rect 113231 278492 113249 278526
rect 113287 278492 113299 278526
rect 113299 278492 113321 278526
rect 113359 278492 113367 278526
rect 113367 278492 113393 278526
rect 113431 278492 113435 278526
rect 113435 278492 113465 278526
rect 113503 278492 113537 278526
rect 113575 278492 113605 278526
rect 113605 278492 113609 278526
rect 113647 278492 113673 278526
rect 113673 278492 113681 278526
rect 113719 278492 113741 278526
rect 113741 278492 113753 278526
rect 113791 278492 113809 278526
rect 113809 278492 113825 278526
rect 113863 278492 113877 278526
rect 113877 278492 113897 278526
rect 113935 278492 113945 278526
rect 113945 278492 113969 278526
rect 114007 278492 114013 278526
rect 114013 278492 114041 278526
rect 111553 278446 111581 278480
rect 111581 278446 111587 278480
rect 111625 278446 111649 278480
rect 111649 278446 111659 278480
rect 111697 278446 111717 278480
rect 111717 278446 111731 278480
rect 111769 278446 111785 278480
rect 111785 278446 111803 278480
rect 111841 278446 111853 278480
rect 111853 278446 111875 278480
rect 111913 278446 111921 278480
rect 111921 278446 111947 278480
rect 111985 278446 111989 278480
rect 111989 278446 112019 278480
rect 112057 278446 112091 278480
rect 112129 278446 112159 278480
rect 112159 278446 112163 278480
rect 112201 278446 112227 278480
rect 112227 278446 112235 278480
rect 112273 278446 112295 278480
rect 112295 278446 112307 278480
rect 112345 278446 112363 278480
rect 112363 278446 112379 278480
rect 112417 278446 112431 278480
rect 112431 278446 112451 278480
rect 112489 278446 112499 278480
rect 112499 278446 112523 278480
rect 112561 278446 112567 278480
rect 112567 278446 112595 278480
rect 111452 278405 111486 278407
rect 111452 278373 111486 278405
rect 111452 278303 111486 278335
rect 111452 278301 111486 278303
rect 112662 278405 112696 278407
rect 112662 278373 112696 278405
rect 112662 278303 112696 278335
rect 112662 278301 112696 278303
rect 111553 278228 111581 278262
rect 111581 278228 111587 278262
rect 111625 278228 111649 278262
rect 111649 278228 111659 278262
rect 111697 278228 111717 278262
rect 111717 278228 111731 278262
rect 111769 278228 111785 278262
rect 111785 278228 111803 278262
rect 111841 278228 111853 278262
rect 111853 278228 111875 278262
rect 111913 278228 111921 278262
rect 111921 278228 111947 278262
rect 111985 278228 111989 278262
rect 111989 278228 112019 278262
rect 112057 278228 112091 278262
rect 112129 278228 112159 278262
rect 112159 278228 112163 278262
rect 112201 278228 112227 278262
rect 112227 278228 112235 278262
rect 112273 278228 112295 278262
rect 112295 278228 112307 278262
rect 112345 278228 112363 278262
rect 112363 278228 112379 278262
rect 112417 278228 112431 278262
rect 112431 278228 112451 278262
rect 112489 278228 112499 278262
rect 112499 278228 112523 278262
rect 112561 278228 112567 278262
rect 112567 278228 112595 278262
rect 113029 278348 113057 278382
rect 113057 278348 113063 278382
rect 113101 278348 113125 278382
rect 113125 278348 113135 278382
rect 113173 278348 113193 278382
rect 113193 278348 113207 278382
rect 113245 278348 113261 278382
rect 113261 278348 113279 278382
rect 113317 278348 113329 278382
rect 113329 278348 113351 278382
rect 113389 278348 113397 278382
rect 113397 278348 113423 278382
rect 113461 278348 113465 278382
rect 113465 278348 113495 278382
rect 113533 278348 113567 278382
rect 113605 278348 113635 278382
rect 113635 278348 113639 278382
rect 113677 278348 113703 278382
rect 113703 278348 113711 278382
rect 113749 278348 113771 278382
rect 113771 278348 113783 278382
rect 113821 278348 113839 278382
rect 113839 278348 113855 278382
rect 113893 278348 113907 278382
rect 113907 278348 113927 278382
rect 113965 278348 113975 278382
rect 113975 278348 113999 278382
rect 114037 278348 114043 278382
rect 114043 278348 114071 278382
rect 112928 278279 112962 278313
rect 114138 278279 114172 278313
rect 114342 278251 114376 278285
rect 113029 278210 113057 278244
rect 113057 278210 113063 278244
rect 113101 278210 113125 278244
rect 113125 278210 113135 278244
rect 113173 278210 113193 278244
rect 113193 278210 113207 278244
rect 113245 278210 113261 278244
rect 113261 278210 113279 278244
rect 113317 278210 113329 278244
rect 113329 278210 113351 278244
rect 113389 278210 113397 278244
rect 113397 278210 113423 278244
rect 113461 278210 113465 278244
rect 113465 278210 113495 278244
rect 113533 278210 113567 278244
rect 113605 278210 113635 278244
rect 113635 278210 113639 278244
rect 113677 278210 113703 278244
rect 113703 278210 113711 278244
rect 113749 278210 113771 278244
rect 113771 278210 113783 278244
rect 113821 278210 113839 278244
rect 113839 278210 113855 278244
rect 113893 278210 113907 278244
rect 113907 278210 113927 278244
rect 113965 278210 113975 278244
rect 113975 278210 113999 278244
rect 114037 278210 114043 278244
rect 114043 278210 114071 278244
rect 114576 279090 114610 279098
rect 114576 279064 114610 279090
rect 114576 279022 114610 279026
rect 114576 278992 114610 279022
rect 114576 278920 114610 278954
rect 114576 278852 114610 278882
rect 114576 278848 114610 278852
rect 114576 278784 114610 278810
rect 114576 278776 114610 278784
rect 114904 279090 114938 279098
rect 114904 279064 114938 279090
rect 114904 279022 114938 279026
rect 114904 278992 114938 279022
rect 114904 278920 114938 278954
rect 114904 278852 114938 278882
rect 114904 278848 114938 278852
rect 114904 278784 114938 278810
rect 114904 278776 114938 278784
rect 114704 278691 114706 278725
rect 114706 278691 114738 278725
rect 114776 278691 114808 278725
rect 114808 278691 114810 278725
rect 115395 279149 115397 279183
rect 115397 279149 115429 279183
rect 115467 279149 115499 279183
rect 115499 279149 115501 279183
rect 114899 278577 114933 278611
rect 115267 279090 115301 279098
rect 115267 279064 115301 279090
rect 115267 279022 115301 279026
rect 115267 278992 115301 279022
rect 115267 278920 115301 278954
rect 115267 278852 115301 278882
rect 115267 278848 115301 278852
rect 115267 278784 115301 278810
rect 115267 278776 115301 278784
rect 115595 279090 115629 279098
rect 115595 279064 115629 279090
rect 115595 279022 115629 279026
rect 115595 278992 115629 279022
rect 115595 278920 115629 278954
rect 115595 278852 115629 278882
rect 115595 278848 115629 278852
rect 115595 278784 115629 278810
rect 115595 278776 115629 278784
rect 115395 278691 115397 278725
rect 115397 278691 115429 278725
rect 115467 278691 115499 278725
rect 115499 278691 115501 278725
rect 114704 278463 114706 278497
rect 114706 278463 114738 278497
rect 114776 278463 114808 278497
rect 114808 278463 114810 278497
rect 114576 278422 114610 278424
rect 114576 278390 114610 278422
rect 114576 278320 114610 278352
rect 114576 278318 114610 278320
rect 114904 278422 114938 278424
rect 114904 278390 114938 278422
rect 114904 278320 114938 278352
rect 114904 278318 114938 278320
rect 115271 278577 115305 278611
rect 115395 278463 115397 278497
rect 115397 278463 115429 278497
rect 115467 278463 115499 278497
rect 115499 278463 115501 278497
rect 115267 278422 115301 278424
rect 115267 278390 115301 278422
rect 115267 278320 115301 278352
rect 115267 278318 115301 278320
rect 115595 278422 115629 278424
rect 115595 278390 115629 278422
rect 115595 278320 115629 278352
rect 115595 278318 115629 278320
rect 116164 279174 116192 279208
rect 116192 279174 116198 279208
rect 116236 279174 116260 279208
rect 116260 279174 116270 279208
rect 116308 279174 116328 279208
rect 116328 279174 116342 279208
rect 116380 279174 116396 279208
rect 116396 279174 116414 279208
rect 116452 279174 116464 279208
rect 116464 279174 116486 279208
rect 116524 279174 116532 279208
rect 116532 279174 116558 279208
rect 116596 279174 116600 279208
rect 116600 279174 116630 279208
rect 116668 279174 116702 279208
rect 116740 279174 116770 279208
rect 116770 279174 116774 279208
rect 116812 279174 116838 279208
rect 116838 279174 116846 279208
rect 116884 279174 116906 279208
rect 116906 279174 116918 279208
rect 116956 279174 116974 279208
rect 116974 279174 116990 279208
rect 117028 279174 117042 279208
rect 117042 279174 117062 279208
rect 117100 279174 117110 279208
rect 117110 279174 117134 279208
rect 117172 279174 117178 279208
rect 117178 279174 117206 279208
rect 116063 279113 116097 279115
rect 116063 279081 116097 279113
rect 116063 279011 116097 279043
rect 116063 279009 116097 279011
rect 117273 279113 117307 279115
rect 117273 279081 117307 279113
rect 117273 279011 117307 279043
rect 117273 279009 117307 279011
rect 116164 278916 116192 278950
rect 116192 278916 116198 278950
rect 116236 278916 116260 278950
rect 116260 278916 116270 278950
rect 116308 278916 116328 278950
rect 116328 278916 116342 278950
rect 116380 278916 116396 278950
rect 116396 278916 116414 278950
rect 116452 278916 116464 278950
rect 116464 278916 116486 278950
rect 116524 278916 116532 278950
rect 116532 278916 116558 278950
rect 116596 278916 116600 278950
rect 116600 278916 116630 278950
rect 116668 278916 116702 278950
rect 116740 278916 116770 278950
rect 116770 278916 116774 278950
rect 116812 278916 116838 278950
rect 116838 278916 116846 278950
rect 116884 278916 116906 278950
rect 116906 278916 116918 278950
rect 116956 278916 116974 278950
rect 116974 278916 116990 278950
rect 117028 278916 117042 278950
rect 117042 278916 117062 278950
rect 117100 278916 117110 278950
rect 117110 278916 117134 278950
rect 117172 278916 117178 278950
rect 117178 278916 117206 278950
rect 117610 279166 117638 279200
rect 117638 279166 117644 279200
rect 117682 279166 117706 279200
rect 117706 279166 117716 279200
rect 117754 279166 117774 279200
rect 117774 279166 117788 279200
rect 117826 279166 117842 279200
rect 117842 279166 117860 279200
rect 117898 279166 117910 279200
rect 117910 279166 117932 279200
rect 117970 279166 117978 279200
rect 117978 279166 118004 279200
rect 118042 279166 118046 279200
rect 118046 279166 118076 279200
rect 118114 279166 118148 279200
rect 118186 279166 118216 279200
rect 118216 279166 118220 279200
rect 118258 279166 118284 279200
rect 118284 279166 118292 279200
rect 118330 279166 118352 279200
rect 118352 279166 118364 279200
rect 118402 279166 118420 279200
rect 118420 279166 118436 279200
rect 118474 279166 118488 279200
rect 118488 279166 118508 279200
rect 118546 279166 118556 279200
rect 118556 279166 118580 279200
rect 118618 279166 118624 279200
rect 118624 279166 118652 279200
rect 117509 279125 117543 279127
rect 117509 279093 117543 279125
rect 117509 279023 117543 279055
rect 117509 279021 117543 279023
rect 118719 279125 118753 279127
rect 118719 279093 118753 279125
rect 118719 279023 118753 279055
rect 118719 279021 118753 279023
rect 117610 278948 117638 278982
rect 117638 278948 117644 278982
rect 117682 278948 117706 278982
rect 117706 278948 117716 278982
rect 117754 278948 117774 278982
rect 117774 278948 117788 278982
rect 117826 278948 117842 278982
rect 117842 278948 117860 278982
rect 117898 278948 117910 278982
rect 117910 278948 117932 278982
rect 117970 278948 117978 278982
rect 117978 278948 118004 278982
rect 118042 278948 118046 278982
rect 118046 278948 118076 278982
rect 118114 278948 118148 278982
rect 118186 278948 118216 278982
rect 118216 278948 118220 278982
rect 118258 278948 118284 278982
rect 118284 278948 118292 278982
rect 118330 278948 118352 278982
rect 118352 278948 118364 278982
rect 118402 278948 118420 278982
rect 118420 278948 118436 278982
rect 118474 278948 118488 278982
rect 118488 278948 118508 278982
rect 118546 278948 118556 278982
rect 118556 278948 118580 278982
rect 118618 278948 118624 278982
rect 118624 278948 118652 278982
rect 116164 278750 116192 278784
rect 116192 278750 116198 278784
rect 116236 278750 116260 278784
rect 116260 278750 116270 278784
rect 116308 278750 116328 278784
rect 116328 278750 116342 278784
rect 116380 278750 116396 278784
rect 116396 278750 116414 278784
rect 116452 278750 116464 278784
rect 116464 278750 116486 278784
rect 116524 278750 116532 278784
rect 116532 278750 116558 278784
rect 116596 278750 116600 278784
rect 116600 278750 116630 278784
rect 116668 278750 116702 278784
rect 116740 278750 116770 278784
rect 116770 278750 116774 278784
rect 116812 278750 116838 278784
rect 116838 278750 116846 278784
rect 116884 278750 116906 278784
rect 116906 278750 116918 278784
rect 116956 278750 116974 278784
rect 116974 278750 116990 278784
rect 117028 278750 117042 278784
rect 117042 278750 117062 278784
rect 117100 278750 117110 278784
rect 117110 278750 117134 278784
rect 117172 278750 117178 278784
rect 117178 278750 117206 278784
rect 116063 278689 116097 278691
rect 116063 278657 116097 278689
rect 116063 278587 116097 278619
rect 116063 278585 116097 278587
rect 117273 278689 117307 278691
rect 117273 278657 117307 278689
rect 117273 278587 117307 278619
rect 117273 278585 117307 278587
rect 116164 278492 116192 278526
rect 116192 278492 116198 278526
rect 116236 278492 116260 278526
rect 116260 278492 116270 278526
rect 116308 278492 116328 278526
rect 116328 278492 116342 278526
rect 116380 278492 116396 278526
rect 116396 278492 116414 278526
rect 116452 278492 116464 278526
rect 116464 278492 116486 278526
rect 116524 278492 116532 278526
rect 116532 278492 116558 278526
rect 116596 278492 116600 278526
rect 116600 278492 116630 278526
rect 116668 278492 116702 278526
rect 116740 278492 116770 278526
rect 116770 278492 116774 278526
rect 116812 278492 116838 278526
rect 116838 278492 116846 278526
rect 116884 278492 116906 278526
rect 116906 278492 116918 278526
rect 116956 278492 116974 278526
rect 116974 278492 116990 278526
rect 117028 278492 117042 278526
rect 117042 278492 117062 278526
rect 117100 278492 117110 278526
rect 117110 278492 117134 278526
rect 117172 278492 117178 278526
rect 117178 278492 117206 278526
rect 117610 278806 117638 278840
rect 117638 278806 117644 278840
rect 117682 278806 117706 278840
rect 117706 278806 117716 278840
rect 117754 278806 117774 278840
rect 117774 278806 117788 278840
rect 117826 278806 117842 278840
rect 117842 278806 117860 278840
rect 117898 278806 117910 278840
rect 117910 278806 117932 278840
rect 117970 278806 117978 278840
rect 117978 278806 118004 278840
rect 118042 278806 118046 278840
rect 118046 278806 118076 278840
rect 118114 278806 118148 278840
rect 118186 278806 118216 278840
rect 118216 278806 118220 278840
rect 118258 278806 118284 278840
rect 118284 278806 118292 278840
rect 118330 278806 118352 278840
rect 118352 278806 118364 278840
rect 118402 278806 118420 278840
rect 118420 278806 118436 278840
rect 118474 278806 118488 278840
rect 118488 278806 118508 278840
rect 118546 278806 118556 278840
rect 118556 278806 118580 278840
rect 118618 278806 118624 278840
rect 118624 278806 118652 278840
rect 117509 278765 117543 278767
rect 117509 278733 117543 278765
rect 117509 278663 117543 278695
rect 117509 278661 117543 278663
rect 118719 278765 118753 278767
rect 118719 278733 118753 278765
rect 118719 278663 118753 278695
rect 118719 278661 118753 278663
rect 117610 278588 117638 278622
rect 117638 278588 117644 278622
rect 117682 278588 117706 278622
rect 117706 278588 117716 278622
rect 117754 278588 117774 278622
rect 117774 278588 117788 278622
rect 117826 278588 117842 278622
rect 117842 278588 117860 278622
rect 117898 278588 117910 278622
rect 117910 278588 117932 278622
rect 117970 278588 117978 278622
rect 117978 278588 118004 278622
rect 118042 278588 118046 278622
rect 118046 278588 118076 278622
rect 118114 278588 118148 278622
rect 118186 278588 118216 278622
rect 118216 278588 118220 278622
rect 118258 278588 118284 278622
rect 118284 278588 118292 278622
rect 118330 278588 118352 278622
rect 118352 278588 118364 278622
rect 118402 278588 118420 278622
rect 118420 278588 118436 278622
rect 118474 278588 118488 278622
rect 118488 278588 118508 278622
rect 118546 278588 118556 278622
rect 118556 278588 118580 278622
rect 118618 278588 118624 278622
rect 118624 278588 118652 278622
rect 111553 278086 111581 278120
rect 111581 278086 111587 278120
rect 111625 278086 111649 278120
rect 111649 278086 111659 278120
rect 111697 278086 111717 278120
rect 111717 278086 111731 278120
rect 111769 278086 111785 278120
rect 111785 278086 111803 278120
rect 111841 278086 111853 278120
rect 111853 278086 111875 278120
rect 111913 278086 111921 278120
rect 111921 278086 111947 278120
rect 111985 278086 111989 278120
rect 111989 278086 112019 278120
rect 112057 278086 112091 278120
rect 112129 278086 112159 278120
rect 112159 278086 112163 278120
rect 112201 278086 112227 278120
rect 112227 278086 112235 278120
rect 112273 278086 112295 278120
rect 112295 278086 112307 278120
rect 112345 278086 112363 278120
rect 112363 278086 112379 278120
rect 112417 278086 112431 278120
rect 112431 278086 112451 278120
rect 112489 278086 112499 278120
rect 112499 278086 112523 278120
rect 112561 278086 112567 278120
rect 112567 278086 112595 278120
rect 111452 278045 111486 278047
rect 111452 278013 111486 278045
rect 111452 277943 111486 277975
rect 111452 277941 111486 277943
rect 113029 278050 113057 278084
rect 113057 278050 113063 278084
rect 113101 278050 113125 278084
rect 113125 278050 113135 278084
rect 113173 278050 113193 278084
rect 113193 278050 113207 278084
rect 113245 278050 113261 278084
rect 113261 278050 113279 278084
rect 113317 278050 113329 278084
rect 113329 278050 113351 278084
rect 113389 278050 113397 278084
rect 113397 278050 113423 278084
rect 113461 278050 113465 278084
rect 113465 278050 113495 278084
rect 113533 278050 113567 278084
rect 113605 278050 113635 278084
rect 113635 278050 113639 278084
rect 113677 278050 113703 278084
rect 113703 278050 113711 278084
rect 113749 278050 113771 278084
rect 113771 278050 113783 278084
rect 113821 278050 113839 278084
rect 113839 278050 113855 278084
rect 113893 278050 113907 278084
rect 113907 278050 113927 278084
rect 113965 278050 113975 278084
rect 113975 278050 113999 278084
rect 114037 278050 114043 278084
rect 114043 278050 114071 278084
rect 112662 278045 112696 278047
rect 112662 278013 112696 278045
rect 112662 277943 112696 277975
rect 112928 277981 112962 278015
rect 114138 277981 114172 278015
rect 112662 277941 112696 277943
rect 113029 277912 113057 277946
rect 113057 277912 113063 277946
rect 113101 277912 113125 277946
rect 113125 277912 113135 277946
rect 113173 277912 113193 277946
rect 113193 277912 113207 277946
rect 113245 277912 113261 277946
rect 113261 277912 113279 277946
rect 113317 277912 113329 277946
rect 113329 277912 113351 277946
rect 113389 277912 113397 277946
rect 113397 277912 113423 277946
rect 113461 277912 113465 277946
rect 113465 277912 113495 277946
rect 113533 277912 113567 277946
rect 113605 277912 113635 277946
rect 113635 277912 113639 277946
rect 113677 277912 113703 277946
rect 113703 277912 113711 277946
rect 113749 277912 113771 277946
rect 113771 277912 113783 277946
rect 113821 277912 113839 277946
rect 113839 277912 113855 277946
rect 113893 277912 113907 277946
rect 113907 277912 113927 277946
rect 113965 277912 113975 277946
rect 113975 277912 113999 277946
rect 114037 277912 114043 277946
rect 114043 277912 114071 277946
rect 114704 278245 114706 278279
rect 114706 278245 114738 278279
rect 114776 278245 114808 278279
rect 114808 278245 114810 278279
rect 111553 277868 111581 277902
rect 111581 277868 111587 277902
rect 111625 277868 111649 277902
rect 111649 277868 111659 277902
rect 111697 277868 111717 277902
rect 111717 277868 111731 277902
rect 111769 277868 111785 277902
rect 111785 277868 111803 277902
rect 111841 277868 111853 277902
rect 111853 277868 111875 277902
rect 111913 277868 111921 277902
rect 111921 277868 111947 277902
rect 111985 277868 111989 277902
rect 111989 277868 112019 277902
rect 112057 277868 112091 277902
rect 112129 277868 112159 277902
rect 112159 277868 112163 277902
rect 112201 277868 112227 277902
rect 112227 277868 112235 277902
rect 112273 277868 112295 277902
rect 112295 277868 112307 277902
rect 112345 277868 112363 277902
rect 112363 277868 112379 277902
rect 112417 277868 112431 277902
rect 112431 277868 112451 277902
rect 112489 277868 112499 277902
rect 112499 277868 112523 277902
rect 112561 277868 112567 277902
rect 112567 277868 112595 277902
rect 114899 278154 114933 278188
rect 115395 278245 115397 278279
rect 115397 278245 115429 278279
rect 115467 278245 115499 278279
rect 115499 278245 115501 278279
rect 114704 278055 114706 278089
rect 114706 278055 114738 278089
rect 114776 278055 114808 278089
rect 114808 278055 114810 278089
rect 114576 278014 114610 278016
rect 114576 277982 114610 278014
rect 114576 277912 114610 277944
rect 114576 277910 114610 277912
rect 114904 278014 114938 278016
rect 114904 277982 114938 278014
rect 114904 277912 114938 277944
rect 114904 277910 114938 277912
rect 115271 278154 115305 278188
rect 115395 278055 115397 278089
rect 115397 278055 115429 278089
rect 115467 278055 115499 278089
rect 115499 278055 115501 278089
rect 115267 278014 115301 278016
rect 115267 277982 115301 278014
rect 115267 277912 115301 277944
rect 115267 277910 115301 277912
rect 115595 278014 115629 278016
rect 115595 277982 115629 278014
rect 115595 277912 115629 277944
rect 115595 277910 115629 277912
rect 116134 278348 116162 278382
rect 116162 278348 116168 278382
rect 116206 278348 116230 278382
rect 116230 278348 116240 278382
rect 116278 278348 116298 278382
rect 116298 278348 116312 278382
rect 116350 278348 116366 278382
rect 116366 278348 116384 278382
rect 116422 278348 116434 278382
rect 116434 278348 116456 278382
rect 116494 278348 116502 278382
rect 116502 278348 116528 278382
rect 116566 278348 116570 278382
rect 116570 278348 116600 278382
rect 116638 278348 116672 278382
rect 116710 278348 116740 278382
rect 116740 278348 116744 278382
rect 116782 278348 116808 278382
rect 116808 278348 116816 278382
rect 116854 278348 116876 278382
rect 116876 278348 116888 278382
rect 116926 278348 116944 278382
rect 116944 278348 116960 278382
rect 116998 278348 117012 278382
rect 117012 278348 117032 278382
rect 117070 278348 117080 278382
rect 117080 278348 117104 278382
rect 117142 278348 117148 278382
rect 117148 278348 117176 278382
rect 115828 278251 115862 278285
rect 116033 278279 116067 278313
rect 117243 278279 117277 278313
rect 116134 278210 116162 278244
rect 116162 278210 116168 278244
rect 116206 278210 116230 278244
rect 116230 278210 116240 278244
rect 116278 278210 116298 278244
rect 116298 278210 116312 278244
rect 116350 278210 116366 278244
rect 116366 278210 116384 278244
rect 116422 278210 116434 278244
rect 116434 278210 116456 278244
rect 116494 278210 116502 278244
rect 116502 278210 116528 278244
rect 116566 278210 116570 278244
rect 116570 278210 116600 278244
rect 116638 278210 116672 278244
rect 116710 278210 116740 278244
rect 116740 278210 116744 278244
rect 116782 278210 116808 278244
rect 116808 278210 116816 278244
rect 116854 278210 116876 278244
rect 116876 278210 116888 278244
rect 116926 278210 116944 278244
rect 116944 278210 116960 278244
rect 116998 278210 117012 278244
rect 117012 278210 117032 278244
rect 117070 278210 117080 278244
rect 117080 278210 117104 278244
rect 117142 278210 117148 278244
rect 117148 278210 117176 278244
rect 117610 278446 117638 278480
rect 117638 278446 117644 278480
rect 117682 278446 117706 278480
rect 117706 278446 117716 278480
rect 117754 278446 117774 278480
rect 117774 278446 117788 278480
rect 117826 278446 117842 278480
rect 117842 278446 117860 278480
rect 117898 278446 117910 278480
rect 117910 278446 117932 278480
rect 117970 278446 117978 278480
rect 117978 278446 118004 278480
rect 118042 278446 118046 278480
rect 118046 278446 118076 278480
rect 118114 278446 118148 278480
rect 118186 278446 118216 278480
rect 118216 278446 118220 278480
rect 118258 278446 118284 278480
rect 118284 278446 118292 278480
rect 118330 278446 118352 278480
rect 118352 278446 118364 278480
rect 118402 278446 118420 278480
rect 118420 278446 118436 278480
rect 118474 278446 118488 278480
rect 118488 278446 118508 278480
rect 118546 278446 118556 278480
rect 118556 278446 118580 278480
rect 118618 278446 118624 278480
rect 118624 278446 118652 278480
rect 117509 278405 117543 278407
rect 117509 278373 117543 278405
rect 117509 278303 117543 278335
rect 117509 278301 117543 278303
rect 118719 278405 118753 278407
rect 118719 278373 118753 278405
rect 118719 278303 118753 278335
rect 118719 278301 118753 278303
rect 117610 278228 117638 278262
rect 117638 278228 117644 278262
rect 117682 278228 117706 278262
rect 117706 278228 117716 278262
rect 117754 278228 117774 278262
rect 117774 278228 117788 278262
rect 117826 278228 117842 278262
rect 117842 278228 117860 278262
rect 117898 278228 117910 278262
rect 117910 278228 117932 278262
rect 117970 278228 117978 278262
rect 117978 278228 118004 278262
rect 118042 278228 118046 278262
rect 118046 278228 118076 278262
rect 118114 278228 118148 278262
rect 118186 278228 118216 278262
rect 118216 278228 118220 278262
rect 118258 278228 118284 278262
rect 118284 278228 118292 278262
rect 118330 278228 118352 278262
rect 118352 278228 118364 278262
rect 118402 278228 118420 278262
rect 118420 278228 118436 278262
rect 118474 278228 118488 278262
rect 118488 278228 118508 278262
rect 118546 278228 118556 278262
rect 118556 278228 118580 278262
rect 118618 278228 118624 278262
rect 118624 278228 118652 278262
rect 117610 278086 117638 278120
rect 117638 278086 117644 278120
rect 117682 278086 117706 278120
rect 117706 278086 117716 278120
rect 117754 278086 117774 278120
rect 117774 278086 117788 278120
rect 117826 278086 117842 278120
rect 117842 278086 117860 278120
rect 117898 278086 117910 278120
rect 117910 278086 117932 278120
rect 117970 278086 117978 278120
rect 117978 278086 118004 278120
rect 118042 278086 118046 278120
rect 118046 278086 118076 278120
rect 118114 278086 118148 278120
rect 118186 278086 118216 278120
rect 118216 278086 118220 278120
rect 118258 278086 118284 278120
rect 118284 278086 118292 278120
rect 118330 278086 118352 278120
rect 118352 278086 118364 278120
rect 118402 278086 118420 278120
rect 118420 278086 118436 278120
rect 118474 278086 118488 278120
rect 118488 278086 118508 278120
rect 118546 278086 118556 278120
rect 118556 278086 118580 278120
rect 118618 278086 118624 278120
rect 118624 278086 118652 278120
rect 116134 278050 116162 278084
rect 116162 278050 116168 278084
rect 116206 278050 116230 278084
rect 116230 278050 116240 278084
rect 116278 278050 116298 278084
rect 116298 278050 116312 278084
rect 116350 278050 116366 278084
rect 116366 278050 116384 278084
rect 116422 278050 116434 278084
rect 116434 278050 116456 278084
rect 116494 278050 116502 278084
rect 116502 278050 116528 278084
rect 116566 278050 116570 278084
rect 116570 278050 116600 278084
rect 116638 278050 116672 278084
rect 116710 278050 116740 278084
rect 116740 278050 116744 278084
rect 116782 278050 116808 278084
rect 116808 278050 116816 278084
rect 116854 278050 116876 278084
rect 116876 278050 116888 278084
rect 116926 278050 116944 278084
rect 116944 278050 116960 278084
rect 116998 278050 117012 278084
rect 117012 278050 117032 278084
rect 117070 278050 117080 278084
rect 117080 278050 117104 278084
rect 117142 278050 117148 278084
rect 117148 278050 117176 278084
rect 117509 278045 117543 278047
rect 116033 277981 116067 278015
rect 117243 277981 117277 278015
rect 117509 278013 117543 278045
rect 116134 277912 116162 277946
rect 116162 277912 116168 277946
rect 116206 277912 116230 277946
rect 116230 277912 116240 277946
rect 116278 277912 116298 277946
rect 116298 277912 116312 277946
rect 116350 277912 116366 277946
rect 116366 277912 116384 277946
rect 116422 277912 116434 277946
rect 116434 277912 116456 277946
rect 116494 277912 116502 277946
rect 116502 277912 116528 277946
rect 116566 277912 116570 277946
rect 116570 277912 116600 277946
rect 116638 277912 116672 277946
rect 116710 277912 116740 277946
rect 116740 277912 116744 277946
rect 116782 277912 116808 277946
rect 116808 277912 116816 277946
rect 116854 277912 116876 277946
rect 116876 277912 116888 277946
rect 116926 277912 116944 277946
rect 116944 277912 116960 277946
rect 116998 277912 117012 277946
rect 117012 277912 117032 277946
rect 117070 277912 117080 277946
rect 117080 277912 117104 277946
rect 117142 277912 117148 277946
rect 117148 277912 117176 277946
rect 117509 277943 117543 277975
rect 117509 277941 117543 277943
rect 118719 278045 118753 278047
rect 118719 278013 118753 278045
rect 118719 277943 118753 277975
rect 118719 277941 118753 277943
rect 114704 277837 114706 277871
rect 114706 277837 114738 277871
rect 114776 277837 114808 277871
rect 114808 277837 114810 277871
rect 115395 277837 115397 277871
rect 115397 277837 115429 277871
rect 115467 277837 115499 277871
rect 115499 277837 115501 277871
rect 117610 277868 117638 277902
rect 117638 277868 117644 277902
rect 117682 277868 117706 277902
rect 117706 277868 117716 277902
rect 117754 277868 117774 277902
rect 117774 277868 117788 277902
rect 117826 277868 117842 277902
rect 117842 277868 117860 277902
rect 117898 277868 117910 277902
rect 117910 277868 117932 277902
rect 117970 277868 117978 277902
rect 117978 277868 118004 277902
rect 118042 277868 118046 277902
rect 118046 277868 118076 277902
rect 118114 277868 118148 277902
rect 118186 277868 118216 277902
rect 118216 277868 118220 277902
rect 118258 277868 118284 277902
rect 118284 277868 118292 277902
rect 118330 277868 118352 277902
rect 118352 277868 118364 277902
rect 118402 277868 118420 277902
rect 118420 277868 118436 277902
rect 118474 277868 118488 277902
rect 118488 277868 118508 277902
rect 118546 277868 118556 277902
rect 118556 277868 118580 277902
rect 118618 277868 118624 277902
rect 118624 277868 118652 277902
rect 114034 277731 114068 277733
rect 114106 277731 114140 277733
rect 114178 277731 114212 277733
rect 114034 277699 114060 277731
rect 114060 277699 114068 277731
rect 114106 277699 114128 277731
rect 114128 277699 114140 277731
rect 114178 277699 114196 277731
rect 114196 277699 114212 277731
rect 115992 277731 116026 277733
rect 116064 277731 116098 277733
rect 116136 277731 116170 277733
rect 115992 277699 116009 277731
rect 116009 277699 116026 277731
rect 116064 277699 116077 277731
rect 116077 277699 116098 277731
rect 116136 277699 116145 277731
rect 116145 277699 116170 277731
rect 111553 277500 111581 277534
rect 111581 277500 111587 277534
rect 111625 277500 111649 277534
rect 111649 277500 111659 277534
rect 111697 277500 111717 277534
rect 111717 277500 111731 277534
rect 111769 277500 111785 277534
rect 111785 277500 111803 277534
rect 111841 277500 111853 277534
rect 111853 277500 111875 277534
rect 111913 277500 111921 277534
rect 111921 277500 111947 277534
rect 111985 277500 111989 277534
rect 111989 277500 112019 277534
rect 112057 277500 112091 277534
rect 112129 277500 112159 277534
rect 112159 277500 112163 277534
rect 112201 277500 112227 277534
rect 112227 277500 112235 277534
rect 112273 277500 112295 277534
rect 112295 277500 112307 277534
rect 112345 277500 112363 277534
rect 112363 277500 112379 277534
rect 112417 277500 112431 277534
rect 112431 277500 112451 277534
rect 112489 277500 112499 277534
rect 112499 277500 112523 277534
rect 112561 277500 112567 277534
rect 112567 277500 112595 277534
rect 111452 277459 111486 277461
rect 111452 277427 111486 277459
rect 111452 277357 111486 277389
rect 111452 277355 111486 277357
rect 112662 277459 112696 277461
rect 112662 277427 112696 277459
rect 112662 277357 112696 277389
rect 112662 277355 112696 277357
rect 111553 277282 111581 277316
rect 111581 277282 111587 277316
rect 111625 277282 111649 277316
rect 111649 277282 111659 277316
rect 111697 277282 111717 277316
rect 111717 277282 111731 277316
rect 111769 277282 111785 277316
rect 111785 277282 111803 277316
rect 111841 277282 111853 277316
rect 111853 277282 111875 277316
rect 111913 277282 111921 277316
rect 111921 277282 111947 277316
rect 111985 277282 111989 277316
rect 111989 277282 112019 277316
rect 112057 277282 112091 277316
rect 112129 277282 112159 277316
rect 112159 277282 112163 277316
rect 112201 277282 112227 277316
rect 112227 277282 112235 277316
rect 112273 277282 112295 277316
rect 112295 277282 112307 277316
rect 112345 277282 112363 277316
rect 112363 277282 112379 277316
rect 112417 277282 112431 277316
rect 112431 277282 112451 277316
rect 112489 277282 112499 277316
rect 112499 277282 112523 277316
rect 112561 277282 112567 277316
rect 112567 277282 112595 277316
rect 112999 277508 113027 277542
rect 113027 277508 113033 277542
rect 113071 277508 113095 277542
rect 113095 277508 113105 277542
rect 113143 277508 113163 277542
rect 113163 277508 113177 277542
rect 113215 277508 113231 277542
rect 113231 277508 113249 277542
rect 113287 277508 113299 277542
rect 113299 277508 113321 277542
rect 113359 277508 113367 277542
rect 113367 277508 113393 277542
rect 113431 277508 113435 277542
rect 113435 277508 113465 277542
rect 113503 277508 113537 277542
rect 113575 277508 113605 277542
rect 113605 277508 113609 277542
rect 113647 277508 113673 277542
rect 113673 277508 113681 277542
rect 113719 277508 113741 277542
rect 113741 277508 113753 277542
rect 113791 277508 113809 277542
rect 113809 277508 113825 277542
rect 113863 277508 113877 277542
rect 113877 277508 113897 277542
rect 113935 277508 113945 277542
rect 113945 277508 113969 277542
rect 114007 277508 114013 277542
rect 114013 277508 114041 277542
rect 112898 277447 112932 277449
rect 112898 277415 112932 277447
rect 112898 277345 112932 277377
rect 112898 277343 112932 277345
rect 114108 277447 114142 277449
rect 114108 277415 114142 277447
rect 114108 277345 114142 277377
rect 114108 277343 114142 277345
rect 114704 277483 114706 277517
rect 114706 277483 114738 277517
rect 114776 277483 114808 277517
rect 114808 277483 114810 277517
rect 112999 277250 113027 277284
rect 113027 277250 113033 277284
rect 113071 277250 113095 277284
rect 113095 277250 113105 277284
rect 113143 277250 113163 277284
rect 113163 277250 113177 277284
rect 113215 277250 113231 277284
rect 113231 277250 113249 277284
rect 113287 277250 113299 277284
rect 113299 277250 113321 277284
rect 113359 277250 113367 277284
rect 113367 277250 113393 277284
rect 113431 277250 113435 277284
rect 113435 277250 113465 277284
rect 113503 277250 113537 277284
rect 113575 277250 113605 277284
rect 113605 277250 113609 277284
rect 113647 277250 113673 277284
rect 113673 277250 113681 277284
rect 113719 277250 113741 277284
rect 113741 277250 113753 277284
rect 113791 277250 113809 277284
rect 113809 277250 113825 277284
rect 113863 277250 113877 277284
rect 113877 277250 113897 277284
rect 113935 277250 113945 277284
rect 113945 277250 113969 277284
rect 114007 277250 114013 277284
rect 114013 277250 114041 277284
rect 111553 277140 111581 277174
rect 111581 277140 111587 277174
rect 111625 277140 111649 277174
rect 111649 277140 111659 277174
rect 111697 277140 111717 277174
rect 111717 277140 111731 277174
rect 111769 277140 111785 277174
rect 111785 277140 111803 277174
rect 111841 277140 111853 277174
rect 111853 277140 111875 277174
rect 111913 277140 111921 277174
rect 111921 277140 111947 277174
rect 111985 277140 111989 277174
rect 111989 277140 112019 277174
rect 112057 277140 112091 277174
rect 112129 277140 112159 277174
rect 112159 277140 112163 277174
rect 112201 277140 112227 277174
rect 112227 277140 112235 277174
rect 112273 277140 112295 277174
rect 112295 277140 112307 277174
rect 112345 277140 112363 277174
rect 112363 277140 112379 277174
rect 112417 277140 112431 277174
rect 112431 277140 112451 277174
rect 112489 277140 112499 277174
rect 112499 277140 112523 277174
rect 112561 277140 112567 277174
rect 112567 277140 112595 277174
rect 111452 277099 111486 277101
rect 111452 277067 111486 277099
rect 111452 276997 111486 277029
rect 111452 276995 111486 276997
rect 112662 277099 112696 277101
rect 112662 277067 112696 277099
rect 112662 276997 112696 277029
rect 112662 276995 112696 276997
rect 111553 276922 111581 276956
rect 111581 276922 111587 276956
rect 111625 276922 111649 276956
rect 111649 276922 111659 276956
rect 111697 276922 111717 276956
rect 111717 276922 111731 276956
rect 111769 276922 111785 276956
rect 111785 276922 111803 276956
rect 111841 276922 111853 276956
rect 111853 276922 111875 276956
rect 111913 276922 111921 276956
rect 111921 276922 111947 276956
rect 111985 276922 111989 276956
rect 111989 276922 112019 276956
rect 112057 276922 112091 276956
rect 112129 276922 112159 276956
rect 112159 276922 112163 276956
rect 112201 276922 112227 276956
rect 112227 276922 112235 276956
rect 112273 276922 112295 276956
rect 112295 276922 112307 276956
rect 112345 276922 112363 276956
rect 112363 276922 112379 276956
rect 112417 276922 112431 276956
rect 112431 276922 112451 276956
rect 112489 276922 112499 276956
rect 112499 276922 112523 276956
rect 112561 276922 112567 276956
rect 112567 276922 112595 276956
rect 112999 277084 113027 277118
rect 113027 277084 113033 277118
rect 113071 277084 113095 277118
rect 113095 277084 113105 277118
rect 113143 277084 113163 277118
rect 113163 277084 113177 277118
rect 113215 277084 113231 277118
rect 113231 277084 113249 277118
rect 113287 277084 113299 277118
rect 113299 277084 113321 277118
rect 113359 277084 113367 277118
rect 113367 277084 113393 277118
rect 113431 277084 113435 277118
rect 113435 277084 113465 277118
rect 113503 277084 113537 277118
rect 113575 277084 113605 277118
rect 113605 277084 113609 277118
rect 113647 277084 113673 277118
rect 113673 277084 113681 277118
rect 113719 277084 113741 277118
rect 113741 277084 113753 277118
rect 113791 277084 113809 277118
rect 113809 277084 113825 277118
rect 113863 277084 113877 277118
rect 113877 277084 113897 277118
rect 113935 277084 113945 277118
rect 113945 277084 113969 277118
rect 114007 277084 114013 277118
rect 114013 277084 114041 277118
rect 112898 277023 112932 277025
rect 112898 276991 112932 277023
rect 112898 276921 112932 276953
rect 112898 276919 112932 276921
rect 114108 277023 114142 277025
rect 114108 276991 114142 277023
rect 114108 276921 114142 276953
rect 114108 276919 114142 276921
rect 112999 276826 113027 276860
rect 113027 276826 113033 276860
rect 113071 276826 113095 276860
rect 113095 276826 113105 276860
rect 113143 276826 113163 276860
rect 113163 276826 113177 276860
rect 113215 276826 113231 276860
rect 113231 276826 113249 276860
rect 113287 276826 113299 276860
rect 113299 276826 113321 276860
rect 113359 276826 113367 276860
rect 113367 276826 113393 276860
rect 113431 276826 113435 276860
rect 113435 276826 113465 276860
rect 113503 276826 113537 276860
rect 113575 276826 113605 276860
rect 113605 276826 113609 276860
rect 113647 276826 113673 276860
rect 113673 276826 113681 276860
rect 113719 276826 113741 276860
rect 113741 276826 113753 276860
rect 113791 276826 113809 276860
rect 113809 276826 113825 276860
rect 113863 276826 113877 276860
rect 113877 276826 113897 276860
rect 113935 276826 113945 276860
rect 113945 276826 113969 276860
rect 114007 276826 114013 276860
rect 114013 276826 114041 276860
rect 111553 276780 111581 276814
rect 111581 276780 111587 276814
rect 111625 276780 111649 276814
rect 111649 276780 111659 276814
rect 111697 276780 111717 276814
rect 111717 276780 111731 276814
rect 111769 276780 111785 276814
rect 111785 276780 111803 276814
rect 111841 276780 111853 276814
rect 111853 276780 111875 276814
rect 111913 276780 111921 276814
rect 111921 276780 111947 276814
rect 111985 276780 111989 276814
rect 111989 276780 112019 276814
rect 112057 276780 112091 276814
rect 112129 276780 112159 276814
rect 112159 276780 112163 276814
rect 112201 276780 112227 276814
rect 112227 276780 112235 276814
rect 112273 276780 112295 276814
rect 112295 276780 112307 276814
rect 112345 276780 112363 276814
rect 112363 276780 112379 276814
rect 112417 276780 112431 276814
rect 112431 276780 112451 276814
rect 112489 276780 112499 276814
rect 112499 276780 112523 276814
rect 112561 276780 112567 276814
rect 112567 276780 112595 276814
rect 111452 276739 111486 276741
rect 111452 276707 111486 276739
rect 111452 276637 111486 276669
rect 111452 276635 111486 276637
rect 112662 276739 112696 276741
rect 112662 276707 112696 276739
rect 112662 276637 112696 276669
rect 112662 276635 112696 276637
rect 111553 276562 111581 276596
rect 111581 276562 111587 276596
rect 111625 276562 111649 276596
rect 111649 276562 111659 276596
rect 111697 276562 111717 276596
rect 111717 276562 111731 276596
rect 111769 276562 111785 276596
rect 111785 276562 111803 276596
rect 111841 276562 111853 276596
rect 111853 276562 111875 276596
rect 111913 276562 111921 276596
rect 111921 276562 111947 276596
rect 111985 276562 111989 276596
rect 111989 276562 112019 276596
rect 112057 276562 112091 276596
rect 112129 276562 112159 276596
rect 112159 276562 112163 276596
rect 112201 276562 112227 276596
rect 112227 276562 112235 276596
rect 112273 276562 112295 276596
rect 112295 276562 112307 276596
rect 112345 276562 112363 276596
rect 112363 276562 112379 276596
rect 112417 276562 112431 276596
rect 112431 276562 112451 276596
rect 112489 276562 112499 276596
rect 112499 276562 112523 276596
rect 112561 276562 112567 276596
rect 112567 276562 112595 276596
rect 113029 276682 113057 276716
rect 113057 276682 113063 276716
rect 113101 276682 113125 276716
rect 113125 276682 113135 276716
rect 113173 276682 113193 276716
rect 113193 276682 113207 276716
rect 113245 276682 113261 276716
rect 113261 276682 113279 276716
rect 113317 276682 113329 276716
rect 113329 276682 113351 276716
rect 113389 276682 113397 276716
rect 113397 276682 113423 276716
rect 113461 276682 113465 276716
rect 113465 276682 113495 276716
rect 113533 276682 113567 276716
rect 113605 276682 113635 276716
rect 113635 276682 113639 276716
rect 113677 276682 113703 276716
rect 113703 276682 113711 276716
rect 113749 276682 113771 276716
rect 113771 276682 113783 276716
rect 113821 276682 113839 276716
rect 113839 276682 113855 276716
rect 113893 276682 113907 276716
rect 113907 276682 113927 276716
rect 113965 276682 113975 276716
rect 113975 276682 113999 276716
rect 114037 276682 114043 276716
rect 114043 276682 114071 276716
rect 112928 276613 112962 276647
rect 114138 276613 114172 276647
rect 114342 276585 114376 276619
rect 113029 276544 113057 276578
rect 113057 276544 113063 276578
rect 113101 276544 113125 276578
rect 113125 276544 113135 276578
rect 113173 276544 113193 276578
rect 113193 276544 113207 276578
rect 113245 276544 113261 276578
rect 113261 276544 113279 276578
rect 113317 276544 113329 276578
rect 113329 276544 113351 276578
rect 113389 276544 113397 276578
rect 113397 276544 113423 276578
rect 113461 276544 113465 276578
rect 113465 276544 113495 276578
rect 113533 276544 113567 276578
rect 113605 276544 113635 276578
rect 113635 276544 113639 276578
rect 113677 276544 113703 276578
rect 113703 276544 113711 276578
rect 113749 276544 113771 276578
rect 113771 276544 113783 276578
rect 113821 276544 113839 276578
rect 113839 276544 113855 276578
rect 113893 276544 113907 276578
rect 113907 276544 113927 276578
rect 113965 276544 113975 276578
rect 113975 276544 113999 276578
rect 114037 276544 114043 276578
rect 114043 276544 114071 276578
rect 114576 277424 114610 277432
rect 114576 277398 114610 277424
rect 114576 277356 114610 277360
rect 114576 277326 114610 277356
rect 114576 277254 114610 277288
rect 114576 277186 114610 277216
rect 114576 277182 114610 277186
rect 114576 277118 114610 277144
rect 114576 277110 114610 277118
rect 114904 277424 114938 277432
rect 114904 277398 114938 277424
rect 114904 277356 114938 277360
rect 114904 277326 114938 277356
rect 114904 277254 114938 277288
rect 114904 277186 114938 277216
rect 114904 277182 114938 277186
rect 114904 277118 114938 277144
rect 114904 277110 114938 277118
rect 114704 277025 114706 277059
rect 114706 277025 114738 277059
rect 114776 277025 114808 277059
rect 114808 277025 114810 277059
rect 115395 277483 115397 277517
rect 115397 277483 115429 277517
rect 115467 277483 115499 277517
rect 115499 277483 115501 277517
rect 114899 276911 114933 276945
rect 115267 277424 115301 277432
rect 115267 277398 115301 277424
rect 115267 277356 115301 277360
rect 115267 277326 115301 277356
rect 115267 277254 115301 277288
rect 115267 277186 115301 277216
rect 115267 277182 115301 277186
rect 115267 277118 115301 277144
rect 115267 277110 115301 277118
rect 115595 277424 115629 277432
rect 115595 277398 115629 277424
rect 115595 277356 115629 277360
rect 115595 277326 115629 277356
rect 115595 277254 115629 277288
rect 115595 277186 115629 277216
rect 115595 277182 115629 277186
rect 115595 277118 115629 277144
rect 115595 277110 115629 277118
rect 115395 277025 115397 277059
rect 115397 277025 115429 277059
rect 115467 277025 115499 277059
rect 115499 277025 115501 277059
rect 114704 276797 114706 276831
rect 114706 276797 114738 276831
rect 114776 276797 114808 276831
rect 114808 276797 114810 276831
rect 114576 276756 114610 276758
rect 114576 276724 114610 276756
rect 114576 276654 114610 276686
rect 114576 276652 114610 276654
rect 114904 276756 114938 276758
rect 114904 276724 114938 276756
rect 114904 276654 114938 276686
rect 114904 276652 114938 276654
rect 115271 276911 115305 276945
rect 115395 276797 115397 276831
rect 115397 276797 115429 276831
rect 115467 276797 115499 276831
rect 115499 276797 115501 276831
rect 115267 276756 115301 276758
rect 115267 276724 115301 276756
rect 115267 276654 115301 276686
rect 115267 276652 115301 276654
rect 115595 276756 115629 276758
rect 115595 276724 115629 276756
rect 115595 276654 115629 276686
rect 115595 276652 115629 276654
rect 116164 277508 116192 277542
rect 116192 277508 116198 277542
rect 116236 277508 116260 277542
rect 116260 277508 116270 277542
rect 116308 277508 116328 277542
rect 116328 277508 116342 277542
rect 116380 277508 116396 277542
rect 116396 277508 116414 277542
rect 116452 277508 116464 277542
rect 116464 277508 116486 277542
rect 116524 277508 116532 277542
rect 116532 277508 116558 277542
rect 116596 277508 116600 277542
rect 116600 277508 116630 277542
rect 116668 277508 116702 277542
rect 116740 277508 116770 277542
rect 116770 277508 116774 277542
rect 116812 277508 116838 277542
rect 116838 277508 116846 277542
rect 116884 277508 116906 277542
rect 116906 277508 116918 277542
rect 116956 277508 116974 277542
rect 116974 277508 116990 277542
rect 117028 277508 117042 277542
rect 117042 277508 117062 277542
rect 117100 277508 117110 277542
rect 117110 277508 117134 277542
rect 117172 277508 117178 277542
rect 117178 277508 117206 277542
rect 116063 277447 116097 277449
rect 116063 277415 116097 277447
rect 116063 277345 116097 277377
rect 116063 277343 116097 277345
rect 117273 277447 117307 277449
rect 117273 277415 117307 277447
rect 117273 277345 117307 277377
rect 117273 277343 117307 277345
rect 116164 277250 116192 277284
rect 116192 277250 116198 277284
rect 116236 277250 116260 277284
rect 116260 277250 116270 277284
rect 116308 277250 116328 277284
rect 116328 277250 116342 277284
rect 116380 277250 116396 277284
rect 116396 277250 116414 277284
rect 116452 277250 116464 277284
rect 116464 277250 116486 277284
rect 116524 277250 116532 277284
rect 116532 277250 116558 277284
rect 116596 277250 116600 277284
rect 116600 277250 116630 277284
rect 116668 277250 116702 277284
rect 116740 277250 116770 277284
rect 116770 277250 116774 277284
rect 116812 277250 116838 277284
rect 116838 277250 116846 277284
rect 116884 277250 116906 277284
rect 116906 277250 116918 277284
rect 116956 277250 116974 277284
rect 116974 277250 116990 277284
rect 117028 277250 117042 277284
rect 117042 277250 117062 277284
rect 117100 277250 117110 277284
rect 117110 277250 117134 277284
rect 117172 277250 117178 277284
rect 117178 277250 117206 277284
rect 117610 277500 117638 277534
rect 117638 277500 117644 277534
rect 117682 277500 117706 277534
rect 117706 277500 117716 277534
rect 117754 277500 117774 277534
rect 117774 277500 117788 277534
rect 117826 277500 117842 277534
rect 117842 277500 117860 277534
rect 117898 277500 117910 277534
rect 117910 277500 117932 277534
rect 117970 277500 117978 277534
rect 117978 277500 118004 277534
rect 118042 277500 118046 277534
rect 118046 277500 118076 277534
rect 118114 277500 118148 277534
rect 118186 277500 118216 277534
rect 118216 277500 118220 277534
rect 118258 277500 118284 277534
rect 118284 277500 118292 277534
rect 118330 277500 118352 277534
rect 118352 277500 118364 277534
rect 118402 277500 118420 277534
rect 118420 277500 118436 277534
rect 118474 277500 118488 277534
rect 118488 277500 118508 277534
rect 118546 277500 118556 277534
rect 118556 277500 118580 277534
rect 118618 277500 118624 277534
rect 118624 277500 118652 277534
rect 117509 277459 117543 277461
rect 117509 277427 117543 277459
rect 117509 277357 117543 277389
rect 117509 277355 117543 277357
rect 118719 277459 118753 277461
rect 118719 277427 118753 277459
rect 118719 277357 118753 277389
rect 118719 277355 118753 277357
rect 117610 277282 117638 277316
rect 117638 277282 117644 277316
rect 117682 277282 117706 277316
rect 117706 277282 117716 277316
rect 117754 277282 117774 277316
rect 117774 277282 117788 277316
rect 117826 277282 117842 277316
rect 117842 277282 117860 277316
rect 117898 277282 117910 277316
rect 117910 277282 117932 277316
rect 117970 277282 117978 277316
rect 117978 277282 118004 277316
rect 118042 277282 118046 277316
rect 118046 277282 118076 277316
rect 118114 277282 118148 277316
rect 118186 277282 118216 277316
rect 118216 277282 118220 277316
rect 118258 277282 118284 277316
rect 118284 277282 118292 277316
rect 118330 277282 118352 277316
rect 118352 277282 118364 277316
rect 118402 277282 118420 277316
rect 118420 277282 118436 277316
rect 118474 277282 118488 277316
rect 118488 277282 118508 277316
rect 118546 277282 118556 277316
rect 118556 277282 118580 277316
rect 118618 277282 118624 277316
rect 118624 277282 118652 277316
rect 116164 277084 116192 277118
rect 116192 277084 116198 277118
rect 116236 277084 116260 277118
rect 116260 277084 116270 277118
rect 116308 277084 116328 277118
rect 116328 277084 116342 277118
rect 116380 277084 116396 277118
rect 116396 277084 116414 277118
rect 116452 277084 116464 277118
rect 116464 277084 116486 277118
rect 116524 277084 116532 277118
rect 116532 277084 116558 277118
rect 116596 277084 116600 277118
rect 116600 277084 116630 277118
rect 116668 277084 116702 277118
rect 116740 277084 116770 277118
rect 116770 277084 116774 277118
rect 116812 277084 116838 277118
rect 116838 277084 116846 277118
rect 116884 277084 116906 277118
rect 116906 277084 116918 277118
rect 116956 277084 116974 277118
rect 116974 277084 116990 277118
rect 117028 277084 117042 277118
rect 117042 277084 117062 277118
rect 117100 277084 117110 277118
rect 117110 277084 117134 277118
rect 117172 277084 117178 277118
rect 117178 277084 117206 277118
rect 116063 277023 116097 277025
rect 116063 276991 116097 277023
rect 116063 276921 116097 276953
rect 116063 276919 116097 276921
rect 117273 277023 117307 277025
rect 117273 276991 117307 277023
rect 117273 276921 117307 276953
rect 117273 276919 117307 276921
rect 116164 276826 116192 276860
rect 116192 276826 116198 276860
rect 116236 276826 116260 276860
rect 116260 276826 116270 276860
rect 116308 276826 116328 276860
rect 116328 276826 116342 276860
rect 116380 276826 116396 276860
rect 116396 276826 116414 276860
rect 116452 276826 116464 276860
rect 116464 276826 116486 276860
rect 116524 276826 116532 276860
rect 116532 276826 116558 276860
rect 116596 276826 116600 276860
rect 116600 276826 116630 276860
rect 116668 276826 116702 276860
rect 116740 276826 116770 276860
rect 116770 276826 116774 276860
rect 116812 276826 116838 276860
rect 116838 276826 116846 276860
rect 116884 276826 116906 276860
rect 116906 276826 116918 276860
rect 116956 276826 116974 276860
rect 116974 276826 116990 276860
rect 117028 276826 117042 276860
rect 117042 276826 117062 276860
rect 117100 276826 117110 276860
rect 117110 276826 117134 276860
rect 117172 276826 117178 276860
rect 117178 276826 117206 276860
rect 117610 277140 117638 277174
rect 117638 277140 117644 277174
rect 117682 277140 117706 277174
rect 117706 277140 117716 277174
rect 117754 277140 117774 277174
rect 117774 277140 117788 277174
rect 117826 277140 117842 277174
rect 117842 277140 117860 277174
rect 117898 277140 117910 277174
rect 117910 277140 117932 277174
rect 117970 277140 117978 277174
rect 117978 277140 118004 277174
rect 118042 277140 118046 277174
rect 118046 277140 118076 277174
rect 118114 277140 118148 277174
rect 118186 277140 118216 277174
rect 118216 277140 118220 277174
rect 118258 277140 118284 277174
rect 118284 277140 118292 277174
rect 118330 277140 118352 277174
rect 118352 277140 118364 277174
rect 118402 277140 118420 277174
rect 118420 277140 118436 277174
rect 118474 277140 118488 277174
rect 118488 277140 118508 277174
rect 118546 277140 118556 277174
rect 118556 277140 118580 277174
rect 118618 277140 118624 277174
rect 118624 277140 118652 277174
rect 117509 277099 117543 277101
rect 117509 277067 117543 277099
rect 117509 276997 117543 277029
rect 117509 276995 117543 276997
rect 118719 277099 118753 277101
rect 118719 277067 118753 277099
rect 118719 276997 118753 277029
rect 118719 276995 118753 276997
rect 117610 276922 117638 276956
rect 117638 276922 117644 276956
rect 117682 276922 117706 276956
rect 117706 276922 117716 276956
rect 117754 276922 117774 276956
rect 117774 276922 117788 276956
rect 117826 276922 117842 276956
rect 117842 276922 117860 276956
rect 117898 276922 117910 276956
rect 117910 276922 117932 276956
rect 117970 276922 117978 276956
rect 117978 276922 118004 276956
rect 118042 276922 118046 276956
rect 118046 276922 118076 276956
rect 118114 276922 118148 276956
rect 118186 276922 118216 276956
rect 118216 276922 118220 276956
rect 118258 276922 118284 276956
rect 118284 276922 118292 276956
rect 118330 276922 118352 276956
rect 118352 276922 118364 276956
rect 118402 276922 118420 276956
rect 118420 276922 118436 276956
rect 118474 276922 118488 276956
rect 118488 276922 118508 276956
rect 118546 276922 118556 276956
rect 118556 276922 118580 276956
rect 118618 276922 118624 276956
rect 118624 276922 118652 276956
rect 111553 276420 111581 276454
rect 111581 276420 111587 276454
rect 111625 276420 111649 276454
rect 111649 276420 111659 276454
rect 111697 276420 111717 276454
rect 111717 276420 111731 276454
rect 111769 276420 111785 276454
rect 111785 276420 111803 276454
rect 111841 276420 111853 276454
rect 111853 276420 111875 276454
rect 111913 276420 111921 276454
rect 111921 276420 111947 276454
rect 111985 276420 111989 276454
rect 111989 276420 112019 276454
rect 112057 276420 112091 276454
rect 112129 276420 112159 276454
rect 112159 276420 112163 276454
rect 112201 276420 112227 276454
rect 112227 276420 112235 276454
rect 112273 276420 112295 276454
rect 112295 276420 112307 276454
rect 112345 276420 112363 276454
rect 112363 276420 112379 276454
rect 112417 276420 112431 276454
rect 112431 276420 112451 276454
rect 112489 276420 112499 276454
rect 112499 276420 112523 276454
rect 112561 276420 112567 276454
rect 112567 276420 112595 276454
rect 111452 276379 111486 276381
rect 111452 276347 111486 276379
rect 111452 276277 111486 276309
rect 111452 276275 111486 276277
rect 113029 276384 113057 276418
rect 113057 276384 113063 276418
rect 113101 276384 113125 276418
rect 113125 276384 113135 276418
rect 113173 276384 113193 276418
rect 113193 276384 113207 276418
rect 113245 276384 113261 276418
rect 113261 276384 113279 276418
rect 113317 276384 113329 276418
rect 113329 276384 113351 276418
rect 113389 276384 113397 276418
rect 113397 276384 113423 276418
rect 113461 276384 113465 276418
rect 113465 276384 113495 276418
rect 113533 276384 113567 276418
rect 113605 276384 113635 276418
rect 113635 276384 113639 276418
rect 113677 276384 113703 276418
rect 113703 276384 113711 276418
rect 113749 276384 113771 276418
rect 113771 276384 113783 276418
rect 113821 276384 113839 276418
rect 113839 276384 113855 276418
rect 113893 276384 113907 276418
rect 113907 276384 113927 276418
rect 113965 276384 113975 276418
rect 113975 276384 113999 276418
rect 114037 276384 114043 276418
rect 114043 276384 114071 276418
rect 112662 276379 112696 276381
rect 112662 276347 112696 276379
rect 112662 276277 112696 276309
rect 112928 276315 112962 276349
rect 114138 276315 114172 276349
rect 112662 276275 112696 276277
rect 113029 276246 113057 276280
rect 113057 276246 113063 276280
rect 113101 276246 113125 276280
rect 113125 276246 113135 276280
rect 113173 276246 113193 276280
rect 113193 276246 113207 276280
rect 113245 276246 113261 276280
rect 113261 276246 113279 276280
rect 113317 276246 113329 276280
rect 113329 276246 113351 276280
rect 113389 276246 113397 276280
rect 113397 276246 113423 276280
rect 113461 276246 113465 276280
rect 113465 276246 113495 276280
rect 113533 276246 113567 276280
rect 113605 276246 113635 276280
rect 113635 276246 113639 276280
rect 113677 276246 113703 276280
rect 113703 276246 113711 276280
rect 113749 276246 113771 276280
rect 113771 276246 113783 276280
rect 113821 276246 113839 276280
rect 113839 276246 113855 276280
rect 113893 276246 113907 276280
rect 113907 276246 113927 276280
rect 113965 276246 113975 276280
rect 113975 276246 113999 276280
rect 114037 276246 114043 276280
rect 114043 276246 114071 276280
rect 114704 276579 114706 276613
rect 114706 276579 114738 276613
rect 114776 276579 114808 276613
rect 114808 276579 114810 276613
rect 111553 276202 111581 276236
rect 111581 276202 111587 276236
rect 111625 276202 111649 276236
rect 111649 276202 111659 276236
rect 111697 276202 111717 276236
rect 111717 276202 111731 276236
rect 111769 276202 111785 276236
rect 111785 276202 111803 276236
rect 111841 276202 111853 276236
rect 111853 276202 111875 276236
rect 111913 276202 111921 276236
rect 111921 276202 111947 276236
rect 111985 276202 111989 276236
rect 111989 276202 112019 276236
rect 112057 276202 112091 276236
rect 112129 276202 112159 276236
rect 112159 276202 112163 276236
rect 112201 276202 112227 276236
rect 112227 276202 112235 276236
rect 112273 276202 112295 276236
rect 112295 276202 112307 276236
rect 112345 276202 112363 276236
rect 112363 276202 112379 276236
rect 112417 276202 112431 276236
rect 112431 276202 112451 276236
rect 112489 276202 112499 276236
rect 112499 276202 112523 276236
rect 112561 276202 112567 276236
rect 112567 276202 112595 276236
rect 114899 276488 114933 276522
rect 115395 276579 115397 276613
rect 115397 276579 115429 276613
rect 115467 276579 115499 276613
rect 115499 276579 115501 276613
rect 114704 276389 114706 276423
rect 114706 276389 114738 276423
rect 114776 276389 114808 276423
rect 114808 276389 114810 276423
rect 114576 276348 114610 276350
rect 114576 276316 114610 276348
rect 114576 276246 114610 276278
rect 114576 276244 114610 276246
rect 114904 276348 114938 276350
rect 114904 276316 114938 276348
rect 114904 276246 114938 276278
rect 114904 276244 114938 276246
rect 115271 276488 115305 276522
rect 115395 276389 115397 276423
rect 115397 276389 115429 276423
rect 115467 276389 115499 276423
rect 115499 276389 115501 276423
rect 115267 276348 115301 276350
rect 115267 276316 115301 276348
rect 115267 276246 115301 276278
rect 115267 276244 115301 276246
rect 115595 276348 115629 276350
rect 115595 276316 115629 276348
rect 115595 276246 115629 276278
rect 115595 276244 115629 276246
rect 116134 276682 116162 276716
rect 116162 276682 116168 276716
rect 116206 276682 116230 276716
rect 116230 276682 116240 276716
rect 116278 276682 116298 276716
rect 116298 276682 116312 276716
rect 116350 276682 116366 276716
rect 116366 276682 116384 276716
rect 116422 276682 116434 276716
rect 116434 276682 116456 276716
rect 116494 276682 116502 276716
rect 116502 276682 116528 276716
rect 116566 276682 116570 276716
rect 116570 276682 116600 276716
rect 116638 276682 116672 276716
rect 116710 276682 116740 276716
rect 116740 276682 116744 276716
rect 116782 276682 116808 276716
rect 116808 276682 116816 276716
rect 116854 276682 116876 276716
rect 116876 276682 116888 276716
rect 116926 276682 116944 276716
rect 116944 276682 116960 276716
rect 116998 276682 117012 276716
rect 117012 276682 117032 276716
rect 117070 276682 117080 276716
rect 117080 276682 117104 276716
rect 117142 276682 117148 276716
rect 117148 276682 117176 276716
rect 115828 276585 115862 276619
rect 116033 276613 116067 276647
rect 117243 276613 117277 276647
rect 116134 276544 116162 276578
rect 116162 276544 116168 276578
rect 116206 276544 116230 276578
rect 116230 276544 116240 276578
rect 116278 276544 116298 276578
rect 116298 276544 116312 276578
rect 116350 276544 116366 276578
rect 116366 276544 116384 276578
rect 116422 276544 116434 276578
rect 116434 276544 116456 276578
rect 116494 276544 116502 276578
rect 116502 276544 116528 276578
rect 116566 276544 116570 276578
rect 116570 276544 116600 276578
rect 116638 276544 116672 276578
rect 116710 276544 116740 276578
rect 116740 276544 116744 276578
rect 116782 276544 116808 276578
rect 116808 276544 116816 276578
rect 116854 276544 116876 276578
rect 116876 276544 116888 276578
rect 116926 276544 116944 276578
rect 116944 276544 116960 276578
rect 116998 276544 117012 276578
rect 117012 276544 117032 276578
rect 117070 276544 117080 276578
rect 117080 276544 117104 276578
rect 117142 276544 117148 276578
rect 117148 276544 117176 276578
rect 117610 276780 117638 276814
rect 117638 276780 117644 276814
rect 117682 276780 117706 276814
rect 117706 276780 117716 276814
rect 117754 276780 117774 276814
rect 117774 276780 117788 276814
rect 117826 276780 117842 276814
rect 117842 276780 117860 276814
rect 117898 276780 117910 276814
rect 117910 276780 117932 276814
rect 117970 276780 117978 276814
rect 117978 276780 118004 276814
rect 118042 276780 118046 276814
rect 118046 276780 118076 276814
rect 118114 276780 118148 276814
rect 118186 276780 118216 276814
rect 118216 276780 118220 276814
rect 118258 276780 118284 276814
rect 118284 276780 118292 276814
rect 118330 276780 118352 276814
rect 118352 276780 118364 276814
rect 118402 276780 118420 276814
rect 118420 276780 118436 276814
rect 118474 276780 118488 276814
rect 118488 276780 118508 276814
rect 118546 276780 118556 276814
rect 118556 276780 118580 276814
rect 118618 276780 118624 276814
rect 118624 276780 118652 276814
rect 117509 276739 117543 276741
rect 117509 276707 117543 276739
rect 117509 276637 117543 276669
rect 117509 276635 117543 276637
rect 118719 276739 118753 276741
rect 118719 276707 118753 276739
rect 118719 276637 118753 276669
rect 118719 276635 118753 276637
rect 117610 276562 117638 276596
rect 117638 276562 117644 276596
rect 117682 276562 117706 276596
rect 117706 276562 117716 276596
rect 117754 276562 117774 276596
rect 117774 276562 117788 276596
rect 117826 276562 117842 276596
rect 117842 276562 117860 276596
rect 117898 276562 117910 276596
rect 117910 276562 117932 276596
rect 117970 276562 117978 276596
rect 117978 276562 118004 276596
rect 118042 276562 118046 276596
rect 118046 276562 118076 276596
rect 118114 276562 118148 276596
rect 118186 276562 118216 276596
rect 118216 276562 118220 276596
rect 118258 276562 118284 276596
rect 118284 276562 118292 276596
rect 118330 276562 118352 276596
rect 118352 276562 118364 276596
rect 118402 276562 118420 276596
rect 118420 276562 118436 276596
rect 118474 276562 118488 276596
rect 118488 276562 118508 276596
rect 118546 276562 118556 276596
rect 118556 276562 118580 276596
rect 118618 276562 118624 276596
rect 118624 276562 118652 276596
rect 117610 276420 117638 276454
rect 117638 276420 117644 276454
rect 117682 276420 117706 276454
rect 117706 276420 117716 276454
rect 117754 276420 117774 276454
rect 117774 276420 117788 276454
rect 117826 276420 117842 276454
rect 117842 276420 117860 276454
rect 117898 276420 117910 276454
rect 117910 276420 117932 276454
rect 117970 276420 117978 276454
rect 117978 276420 118004 276454
rect 118042 276420 118046 276454
rect 118046 276420 118076 276454
rect 118114 276420 118148 276454
rect 118186 276420 118216 276454
rect 118216 276420 118220 276454
rect 118258 276420 118284 276454
rect 118284 276420 118292 276454
rect 118330 276420 118352 276454
rect 118352 276420 118364 276454
rect 118402 276420 118420 276454
rect 118420 276420 118436 276454
rect 118474 276420 118488 276454
rect 118488 276420 118508 276454
rect 118546 276420 118556 276454
rect 118556 276420 118580 276454
rect 118618 276420 118624 276454
rect 118624 276420 118652 276454
rect 116134 276384 116162 276418
rect 116162 276384 116168 276418
rect 116206 276384 116230 276418
rect 116230 276384 116240 276418
rect 116278 276384 116298 276418
rect 116298 276384 116312 276418
rect 116350 276384 116366 276418
rect 116366 276384 116384 276418
rect 116422 276384 116434 276418
rect 116434 276384 116456 276418
rect 116494 276384 116502 276418
rect 116502 276384 116528 276418
rect 116566 276384 116570 276418
rect 116570 276384 116600 276418
rect 116638 276384 116672 276418
rect 116710 276384 116740 276418
rect 116740 276384 116744 276418
rect 116782 276384 116808 276418
rect 116808 276384 116816 276418
rect 116854 276384 116876 276418
rect 116876 276384 116888 276418
rect 116926 276384 116944 276418
rect 116944 276384 116960 276418
rect 116998 276384 117012 276418
rect 117012 276384 117032 276418
rect 117070 276384 117080 276418
rect 117080 276384 117104 276418
rect 117142 276384 117148 276418
rect 117148 276384 117176 276418
rect 117509 276379 117543 276381
rect 116033 276315 116067 276349
rect 117243 276315 117277 276349
rect 117509 276347 117543 276379
rect 116134 276246 116162 276280
rect 116162 276246 116168 276280
rect 116206 276246 116230 276280
rect 116230 276246 116240 276280
rect 116278 276246 116298 276280
rect 116298 276246 116312 276280
rect 116350 276246 116366 276280
rect 116366 276246 116384 276280
rect 116422 276246 116434 276280
rect 116434 276246 116456 276280
rect 116494 276246 116502 276280
rect 116502 276246 116528 276280
rect 116566 276246 116570 276280
rect 116570 276246 116600 276280
rect 116638 276246 116672 276280
rect 116710 276246 116740 276280
rect 116740 276246 116744 276280
rect 116782 276246 116808 276280
rect 116808 276246 116816 276280
rect 116854 276246 116876 276280
rect 116876 276246 116888 276280
rect 116926 276246 116944 276280
rect 116944 276246 116960 276280
rect 116998 276246 117012 276280
rect 117012 276246 117032 276280
rect 117070 276246 117080 276280
rect 117080 276246 117104 276280
rect 117142 276246 117148 276280
rect 117148 276246 117176 276280
rect 117509 276277 117543 276309
rect 117509 276275 117543 276277
rect 118719 276379 118753 276381
rect 118719 276347 118753 276379
rect 118719 276277 118753 276309
rect 118719 276275 118753 276277
rect 114704 276171 114706 276205
rect 114706 276171 114738 276205
rect 114776 276171 114808 276205
rect 114808 276171 114810 276205
rect 115395 276171 115397 276205
rect 115397 276171 115429 276205
rect 115467 276171 115499 276205
rect 115499 276171 115501 276205
rect 117610 276202 117638 276236
rect 117638 276202 117644 276236
rect 117682 276202 117706 276236
rect 117706 276202 117716 276236
rect 117754 276202 117774 276236
rect 117774 276202 117788 276236
rect 117826 276202 117842 276236
rect 117842 276202 117860 276236
rect 117898 276202 117910 276236
rect 117910 276202 117932 276236
rect 117970 276202 117978 276236
rect 117978 276202 118004 276236
rect 118042 276202 118046 276236
rect 118046 276202 118076 276236
rect 118114 276202 118148 276236
rect 118186 276202 118216 276236
rect 118216 276202 118220 276236
rect 118258 276202 118284 276236
rect 118284 276202 118292 276236
rect 118330 276202 118352 276236
rect 118352 276202 118364 276236
rect 118402 276202 118420 276236
rect 118420 276202 118436 276236
rect 118474 276202 118488 276236
rect 118488 276202 118508 276236
rect 118546 276202 118556 276236
rect 118556 276202 118580 276236
rect 118618 276202 118624 276236
rect 118624 276202 118652 276236
rect 114034 276065 114068 276067
rect 114106 276065 114140 276067
rect 114178 276065 114212 276067
rect 114034 276033 114060 276065
rect 114060 276033 114068 276065
rect 114106 276033 114128 276065
rect 114128 276033 114140 276065
rect 114178 276033 114196 276065
rect 114196 276033 114212 276065
rect 115992 276065 116026 276067
rect 116064 276065 116098 276067
rect 116136 276065 116170 276067
rect 115992 276033 116009 276065
rect 116009 276033 116026 276065
rect 116064 276033 116077 276065
rect 116077 276033 116098 276065
rect 116136 276033 116145 276065
rect 116145 276033 116170 276065
rect 111553 275834 111581 275868
rect 111581 275834 111587 275868
rect 111625 275834 111649 275868
rect 111649 275834 111659 275868
rect 111697 275834 111717 275868
rect 111717 275834 111731 275868
rect 111769 275834 111785 275868
rect 111785 275834 111803 275868
rect 111841 275834 111853 275868
rect 111853 275834 111875 275868
rect 111913 275834 111921 275868
rect 111921 275834 111947 275868
rect 111985 275834 111989 275868
rect 111989 275834 112019 275868
rect 112057 275834 112091 275868
rect 112129 275834 112159 275868
rect 112159 275834 112163 275868
rect 112201 275834 112227 275868
rect 112227 275834 112235 275868
rect 112273 275834 112295 275868
rect 112295 275834 112307 275868
rect 112345 275834 112363 275868
rect 112363 275834 112379 275868
rect 112417 275834 112431 275868
rect 112431 275834 112451 275868
rect 112489 275834 112499 275868
rect 112499 275834 112523 275868
rect 112561 275834 112567 275868
rect 112567 275834 112595 275868
rect 111452 275793 111486 275795
rect 111452 275761 111486 275793
rect 111452 275691 111486 275723
rect 111452 275689 111486 275691
rect 112662 275793 112696 275795
rect 112662 275761 112696 275793
rect 112662 275691 112696 275723
rect 112662 275689 112696 275691
rect 111553 275616 111581 275650
rect 111581 275616 111587 275650
rect 111625 275616 111649 275650
rect 111649 275616 111659 275650
rect 111697 275616 111717 275650
rect 111717 275616 111731 275650
rect 111769 275616 111785 275650
rect 111785 275616 111803 275650
rect 111841 275616 111853 275650
rect 111853 275616 111875 275650
rect 111913 275616 111921 275650
rect 111921 275616 111947 275650
rect 111985 275616 111989 275650
rect 111989 275616 112019 275650
rect 112057 275616 112091 275650
rect 112129 275616 112159 275650
rect 112159 275616 112163 275650
rect 112201 275616 112227 275650
rect 112227 275616 112235 275650
rect 112273 275616 112295 275650
rect 112295 275616 112307 275650
rect 112345 275616 112363 275650
rect 112363 275616 112379 275650
rect 112417 275616 112431 275650
rect 112431 275616 112451 275650
rect 112489 275616 112499 275650
rect 112499 275616 112523 275650
rect 112561 275616 112567 275650
rect 112567 275616 112595 275650
rect 112999 275842 113027 275876
rect 113027 275842 113033 275876
rect 113071 275842 113095 275876
rect 113095 275842 113105 275876
rect 113143 275842 113163 275876
rect 113163 275842 113177 275876
rect 113215 275842 113231 275876
rect 113231 275842 113249 275876
rect 113287 275842 113299 275876
rect 113299 275842 113321 275876
rect 113359 275842 113367 275876
rect 113367 275842 113393 275876
rect 113431 275842 113435 275876
rect 113435 275842 113465 275876
rect 113503 275842 113537 275876
rect 113575 275842 113605 275876
rect 113605 275842 113609 275876
rect 113647 275842 113673 275876
rect 113673 275842 113681 275876
rect 113719 275842 113741 275876
rect 113741 275842 113753 275876
rect 113791 275842 113809 275876
rect 113809 275842 113825 275876
rect 113863 275842 113877 275876
rect 113877 275842 113897 275876
rect 113935 275842 113945 275876
rect 113945 275842 113969 275876
rect 114007 275842 114013 275876
rect 114013 275842 114041 275876
rect 112898 275781 112932 275783
rect 112898 275749 112932 275781
rect 112898 275679 112932 275711
rect 112898 275677 112932 275679
rect 114108 275781 114142 275783
rect 114108 275749 114142 275781
rect 114108 275679 114142 275711
rect 114108 275677 114142 275679
rect 114704 275817 114706 275851
rect 114706 275817 114738 275851
rect 114776 275817 114808 275851
rect 114808 275817 114810 275851
rect 112999 275584 113027 275618
rect 113027 275584 113033 275618
rect 113071 275584 113095 275618
rect 113095 275584 113105 275618
rect 113143 275584 113163 275618
rect 113163 275584 113177 275618
rect 113215 275584 113231 275618
rect 113231 275584 113249 275618
rect 113287 275584 113299 275618
rect 113299 275584 113321 275618
rect 113359 275584 113367 275618
rect 113367 275584 113393 275618
rect 113431 275584 113435 275618
rect 113435 275584 113465 275618
rect 113503 275584 113537 275618
rect 113575 275584 113605 275618
rect 113605 275584 113609 275618
rect 113647 275584 113673 275618
rect 113673 275584 113681 275618
rect 113719 275584 113741 275618
rect 113741 275584 113753 275618
rect 113791 275584 113809 275618
rect 113809 275584 113825 275618
rect 113863 275584 113877 275618
rect 113877 275584 113897 275618
rect 113935 275584 113945 275618
rect 113945 275584 113969 275618
rect 114007 275584 114013 275618
rect 114013 275584 114041 275618
rect 111553 275474 111581 275508
rect 111581 275474 111587 275508
rect 111625 275474 111649 275508
rect 111649 275474 111659 275508
rect 111697 275474 111717 275508
rect 111717 275474 111731 275508
rect 111769 275474 111785 275508
rect 111785 275474 111803 275508
rect 111841 275474 111853 275508
rect 111853 275474 111875 275508
rect 111913 275474 111921 275508
rect 111921 275474 111947 275508
rect 111985 275474 111989 275508
rect 111989 275474 112019 275508
rect 112057 275474 112091 275508
rect 112129 275474 112159 275508
rect 112159 275474 112163 275508
rect 112201 275474 112227 275508
rect 112227 275474 112235 275508
rect 112273 275474 112295 275508
rect 112295 275474 112307 275508
rect 112345 275474 112363 275508
rect 112363 275474 112379 275508
rect 112417 275474 112431 275508
rect 112431 275474 112451 275508
rect 112489 275474 112499 275508
rect 112499 275474 112523 275508
rect 112561 275474 112567 275508
rect 112567 275474 112595 275508
rect 111452 275433 111486 275435
rect 111452 275401 111486 275433
rect 111452 275331 111486 275363
rect 111452 275329 111486 275331
rect 112662 275433 112696 275435
rect 112662 275401 112696 275433
rect 112662 275331 112696 275363
rect 112662 275329 112696 275331
rect 111553 275256 111581 275290
rect 111581 275256 111587 275290
rect 111625 275256 111649 275290
rect 111649 275256 111659 275290
rect 111697 275256 111717 275290
rect 111717 275256 111731 275290
rect 111769 275256 111785 275290
rect 111785 275256 111803 275290
rect 111841 275256 111853 275290
rect 111853 275256 111875 275290
rect 111913 275256 111921 275290
rect 111921 275256 111947 275290
rect 111985 275256 111989 275290
rect 111989 275256 112019 275290
rect 112057 275256 112091 275290
rect 112129 275256 112159 275290
rect 112159 275256 112163 275290
rect 112201 275256 112227 275290
rect 112227 275256 112235 275290
rect 112273 275256 112295 275290
rect 112295 275256 112307 275290
rect 112345 275256 112363 275290
rect 112363 275256 112379 275290
rect 112417 275256 112431 275290
rect 112431 275256 112451 275290
rect 112489 275256 112499 275290
rect 112499 275256 112523 275290
rect 112561 275256 112567 275290
rect 112567 275256 112595 275290
rect 112999 275418 113027 275452
rect 113027 275418 113033 275452
rect 113071 275418 113095 275452
rect 113095 275418 113105 275452
rect 113143 275418 113163 275452
rect 113163 275418 113177 275452
rect 113215 275418 113231 275452
rect 113231 275418 113249 275452
rect 113287 275418 113299 275452
rect 113299 275418 113321 275452
rect 113359 275418 113367 275452
rect 113367 275418 113393 275452
rect 113431 275418 113435 275452
rect 113435 275418 113465 275452
rect 113503 275418 113537 275452
rect 113575 275418 113605 275452
rect 113605 275418 113609 275452
rect 113647 275418 113673 275452
rect 113673 275418 113681 275452
rect 113719 275418 113741 275452
rect 113741 275418 113753 275452
rect 113791 275418 113809 275452
rect 113809 275418 113825 275452
rect 113863 275418 113877 275452
rect 113877 275418 113897 275452
rect 113935 275418 113945 275452
rect 113945 275418 113969 275452
rect 114007 275418 114013 275452
rect 114013 275418 114041 275452
rect 112898 275357 112932 275359
rect 112898 275325 112932 275357
rect 112898 275255 112932 275287
rect 112898 275253 112932 275255
rect 114108 275357 114142 275359
rect 114108 275325 114142 275357
rect 114108 275255 114142 275287
rect 114108 275253 114142 275255
rect 112999 275160 113027 275194
rect 113027 275160 113033 275194
rect 113071 275160 113095 275194
rect 113095 275160 113105 275194
rect 113143 275160 113163 275194
rect 113163 275160 113177 275194
rect 113215 275160 113231 275194
rect 113231 275160 113249 275194
rect 113287 275160 113299 275194
rect 113299 275160 113321 275194
rect 113359 275160 113367 275194
rect 113367 275160 113393 275194
rect 113431 275160 113435 275194
rect 113435 275160 113465 275194
rect 113503 275160 113537 275194
rect 113575 275160 113605 275194
rect 113605 275160 113609 275194
rect 113647 275160 113673 275194
rect 113673 275160 113681 275194
rect 113719 275160 113741 275194
rect 113741 275160 113753 275194
rect 113791 275160 113809 275194
rect 113809 275160 113825 275194
rect 113863 275160 113877 275194
rect 113877 275160 113897 275194
rect 113935 275160 113945 275194
rect 113945 275160 113969 275194
rect 114007 275160 114013 275194
rect 114013 275160 114041 275194
rect 111553 275114 111581 275148
rect 111581 275114 111587 275148
rect 111625 275114 111649 275148
rect 111649 275114 111659 275148
rect 111697 275114 111717 275148
rect 111717 275114 111731 275148
rect 111769 275114 111785 275148
rect 111785 275114 111803 275148
rect 111841 275114 111853 275148
rect 111853 275114 111875 275148
rect 111913 275114 111921 275148
rect 111921 275114 111947 275148
rect 111985 275114 111989 275148
rect 111989 275114 112019 275148
rect 112057 275114 112091 275148
rect 112129 275114 112159 275148
rect 112159 275114 112163 275148
rect 112201 275114 112227 275148
rect 112227 275114 112235 275148
rect 112273 275114 112295 275148
rect 112295 275114 112307 275148
rect 112345 275114 112363 275148
rect 112363 275114 112379 275148
rect 112417 275114 112431 275148
rect 112431 275114 112451 275148
rect 112489 275114 112499 275148
rect 112499 275114 112523 275148
rect 112561 275114 112567 275148
rect 112567 275114 112595 275148
rect 111452 275073 111486 275075
rect 111452 275041 111486 275073
rect 111452 274971 111486 275003
rect 111452 274969 111486 274971
rect 112662 275073 112696 275075
rect 112662 275041 112696 275073
rect 112662 274971 112696 275003
rect 112662 274969 112696 274971
rect 111553 274896 111581 274930
rect 111581 274896 111587 274930
rect 111625 274896 111649 274930
rect 111649 274896 111659 274930
rect 111697 274896 111717 274930
rect 111717 274896 111731 274930
rect 111769 274896 111785 274930
rect 111785 274896 111803 274930
rect 111841 274896 111853 274930
rect 111853 274896 111875 274930
rect 111913 274896 111921 274930
rect 111921 274896 111947 274930
rect 111985 274896 111989 274930
rect 111989 274896 112019 274930
rect 112057 274896 112091 274930
rect 112129 274896 112159 274930
rect 112159 274896 112163 274930
rect 112201 274896 112227 274930
rect 112227 274896 112235 274930
rect 112273 274896 112295 274930
rect 112295 274896 112307 274930
rect 112345 274896 112363 274930
rect 112363 274896 112379 274930
rect 112417 274896 112431 274930
rect 112431 274896 112451 274930
rect 112489 274896 112499 274930
rect 112499 274896 112523 274930
rect 112561 274896 112567 274930
rect 112567 274896 112595 274930
rect 113029 275016 113057 275050
rect 113057 275016 113063 275050
rect 113101 275016 113125 275050
rect 113125 275016 113135 275050
rect 113173 275016 113193 275050
rect 113193 275016 113207 275050
rect 113245 275016 113261 275050
rect 113261 275016 113279 275050
rect 113317 275016 113329 275050
rect 113329 275016 113351 275050
rect 113389 275016 113397 275050
rect 113397 275016 113423 275050
rect 113461 275016 113465 275050
rect 113465 275016 113495 275050
rect 113533 275016 113567 275050
rect 113605 275016 113635 275050
rect 113635 275016 113639 275050
rect 113677 275016 113703 275050
rect 113703 275016 113711 275050
rect 113749 275016 113771 275050
rect 113771 275016 113783 275050
rect 113821 275016 113839 275050
rect 113839 275016 113855 275050
rect 113893 275016 113907 275050
rect 113907 275016 113927 275050
rect 113965 275016 113975 275050
rect 113975 275016 113999 275050
rect 114037 275016 114043 275050
rect 114043 275016 114071 275050
rect 112928 274947 112962 274981
rect 114138 274947 114172 274981
rect 114342 274919 114376 274953
rect 113029 274878 113057 274912
rect 113057 274878 113063 274912
rect 113101 274878 113125 274912
rect 113125 274878 113135 274912
rect 113173 274878 113193 274912
rect 113193 274878 113207 274912
rect 113245 274878 113261 274912
rect 113261 274878 113279 274912
rect 113317 274878 113329 274912
rect 113329 274878 113351 274912
rect 113389 274878 113397 274912
rect 113397 274878 113423 274912
rect 113461 274878 113465 274912
rect 113465 274878 113495 274912
rect 113533 274878 113567 274912
rect 113605 274878 113635 274912
rect 113635 274878 113639 274912
rect 113677 274878 113703 274912
rect 113703 274878 113711 274912
rect 113749 274878 113771 274912
rect 113771 274878 113783 274912
rect 113821 274878 113839 274912
rect 113839 274878 113855 274912
rect 113893 274878 113907 274912
rect 113907 274878 113927 274912
rect 113965 274878 113975 274912
rect 113975 274878 113999 274912
rect 114037 274878 114043 274912
rect 114043 274878 114071 274912
rect 114576 275758 114610 275766
rect 114576 275732 114610 275758
rect 114576 275690 114610 275694
rect 114576 275660 114610 275690
rect 114576 275588 114610 275622
rect 114576 275520 114610 275550
rect 114576 275516 114610 275520
rect 114576 275452 114610 275478
rect 114576 275444 114610 275452
rect 114904 275758 114938 275766
rect 114904 275732 114938 275758
rect 114904 275690 114938 275694
rect 114904 275660 114938 275690
rect 114904 275588 114938 275622
rect 114904 275520 114938 275550
rect 114904 275516 114938 275520
rect 114904 275452 114938 275478
rect 114904 275444 114938 275452
rect 114704 275359 114706 275393
rect 114706 275359 114738 275393
rect 114776 275359 114808 275393
rect 114808 275359 114810 275393
rect 115395 275817 115397 275851
rect 115397 275817 115429 275851
rect 115467 275817 115499 275851
rect 115499 275817 115501 275851
rect 114899 275245 114933 275279
rect 115267 275758 115301 275766
rect 115267 275732 115301 275758
rect 115267 275690 115301 275694
rect 115267 275660 115301 275690
rect 115267 275588 115301 275622
rect 115267 275520 115301 275550
rect 115267 275516 115301 275520
rect 115267 275452 115301 275478
rect 115267 275444 115301 275452
rect 115595 275758 115629 275766
rect 115595 275732 115629 275758
rect 115595 275690 115629 275694
rect 115595 275660 115629 275690
rect 115595 275588 115629 275622
rect 115595 275520 115629 275550
rect 115595 275516 115629 275520
rect 115595 275452 115629 275478
rect 115595 275444 115629 275452
rect 115395 275359 115397 275393
rect 115397 275359 115429 275393
rect 115467 275359 115499 275393
rect 115499 275359 115501 275393
rect 114704 275131 114706 275165
rect 114706 275131 114738 275165
rect 114776 275131 114808 275165
rect 114808 275131 114810 275165
rect 114576 275090 114610 275092
rect 114576 275058 114610 275090
rect 114576 274988 114610 275020
rect 114576 274986 114610 274988
rect 114904 275090 114938 275092
rect 114904 275058 114938 275090
rect 114904 274988 114938 275020
rect 114904 274986 114938 274988
rect 115271 275245 115305 275279
rect 115395 275131 115397 275165
rect 115397 275131 115429 275165
rect 115467 275131 115499 275165
rect 115499 275131 115501 275165
rect 115267 275090 115301 275092
rect 115267 275058 115301 275090
rect 115267 274988 115301 275020
rect 115267 274986 115301 274988
rect 115595 275090 115629 275092
rect 115595 275058 115629 275090
rect 115595 274988 115629 275020
rect 115595 274986 115629 274988
rect 116164 275842 116192 275876
rect 116192 275842 116198 275876
rect 116236 275842 116260 275876
rect 116260 275842 116270 275876
rect 116308 275842 116328 275876
rect 116328 275842 116342 275876
rect 116380 275842 116396 275876
rect 116396 275842 116414 275876
rect 116452 275842 116464 275876
rect 116464 275842 116486 275876
rect 116524 275842 116532 275876
rect 116532 275842 116558 275876
rect 116596 275842 116600 275876
rect 116600 275842 116630 275876
rect 116668 275842 116702 275876
rect 116740 275842 116770 275876
rect 116770 275842 116774 275876
rect 116812 275842 116838 275876
rect 116838 275842 116846 275876
rect 116884 275842 116906 275876
rect 116906 275842 116918 275876
rect 116956 275842 116974 275876
rect 116974 275842 116990 275876
rect 117028 275842 117042 275876
rect 117042 275842 117062 275876
rect 117100 275842 117110 275876
rect 117110 275842 117134 275876
rect 117172 275842 117178 275876
rect 117178 275842 117206 275876
rect 116063 275781 116097 275783
rect 116063 275749 116097 275781
rect 116063 275679 116097 275711
rect 116063 275677 116097 275679
rect 117273 275781 117307 275783
rect 117273 275749 117307 275781
rect 117273 275679 117307 275711
rect 117273 275677 117307 275679
rect 116164 275584 116192 275618
rect 116192 275584 116198 275618
rect 116236 275584 116260 275618
rect 116260 275584 116270 275618
rect 116308 275584 116328 275618
rect 116328 275584 116342 275618
rect 116380 275584 116396 275618
rect 116396 275584 116414 275618
rect 116452 275584 116464 275618
rect 116464 275584 116486 275618
rect 116524 275584 116532 275618
rect 116532 275584 116558 275618
rect 116596 275584 116600 275618
rect 116600 275584 116630 275618
rect 116668 275584 116702 275618
rect 116740 275584 116770 275618
rect 116770 275584 116774 275618
rect 116812 275584 116838 275618
rect 116838 275584 116846 275618
rect 116884 275584 116906 275618
rect 116906 275584 116918 275618
rect 116956 275584 116974 275618
rect 116974 275584 116990 275618
rect 117028 275584 117042 275618
rect 117042 275584 117062 275618
rect 117100 275584 117110 275618
rect 117110 275584 117134 275618
rect 117172 275584 117178 275618
rect 117178 275584 117206 275618
rect 117610 275834 117638 275868
rect 117638 275834 117644 275868
rect 117682 275834 117706 275868
rect 117706 275834 117716 275868
rect 117754 275834 117774 275868
rect 117774 275834 117788 275868
rect 117826 275834 117842 275868
rect 117842 275834 117860 275868
rect 117898 275834 117910 275868
rect 117910 275834 117932 275868
rect 117970 275834 117978 275868
rect 117978 275834 118004 275868
rect 118042 275834 118046 275868
rect 118046 275834 118076 275868
rect 118114 275834 118148 275868
rect 118186 275834 118216 275868
rect 118216 275834 118220 275868
rect 118258 275834 118284 275868
rect 118284 275834 118292 275868
rect 118330 275834 118352 275868
rect 118352 275834 118364 275868
rect 118402 275834 118420 275868
rect 118420 275834 118436 275868
rect 118474 275834 118488 275868
rect 118488 275834 118508 275868
rect 118546 275834 118556 275868
rect 118556 275834 118580 275868
rect 118618 275834 118624 275868
rect 118624 275834 118652 275868
rect 117509 275793 117543 275795
rect 117509 275761 117543 275793
rect 117509 275691 117543 275723
rect 117509 275689 117543 275691
rect 118719 275793 118753 275795
rect 118719 275761 118753 275793
rect 118719 275691 118753 275723
rect 118719 275689 118753 275691
rect 117610 275616 117638 275650
rect 117638 275616 117644 275650
rect 117682 275616 117706 275650
rect 117706 275616 117716 275650
rect 117754 275616 117774 275650
rect 117774 275616 117788 275650
rect 117826 275616 117842 275650
rect 117842 275616 117860 275650
rect 117898 275616 117910 275650
rect 117910 275616 117932 275650
rect 117970 275616 117978 275650
rect 117978 275616 118004 275650
rect 118042 275616 118046 275650
rect 118046 275616 118076 275650
rect 118114 275616 118148 275650
rect 118186 275616 118216 275650
rect 118216 275616 118220 275650
rect 118258 275616 118284 275650
rect 118284 275616 118292 275650
rect 118330 275616 118352 275650
rect 118352 275616 118364 275650
rect 118402 275616 118420 275650
rect 118420 275616 118436 275650
rect 118474 275616 118488 275650
rect 118488 275616 118508 275650
rect 118546 275616 118556 275650
rect 118556 275616 118580 275650
rect 118618 275616 118624 275650
rect 118624 275616 118652 275650
rect 116164 275418 116192 275452
rect 116192 275418 116198 275452
rect 116236 275418 116260 275452
rect 116260 275418 116270 275452
rect 116308 275418 116328 275452
rect 116328 275418 116342 275452
rect 116380 275418 116396 275452
rect 116396 275418 116414 275452
rect 116452 275418 116464 275452
rect 116464 275418 116486 275452
rect 116524 275418 116532 275452
rect 116532 275418 116558 275452
rect 116596 275418 116600 275452
rect 116600 275418 116630 275452
rect 116668 275418 116702 275452
rect 116740 275418 116770 275452
rect 116770 275418 116774 275452
rect 116812 275418 116838 275452
rect 116838 275418 116846 275452
rect 116884 275418 116906 275452
rect 116906 275418 116918 275452
rect 116956 275418 116974 275452
rect 116974 275418 116990 275452
rect 117028 275418 117042 275452
rect 117042 275418 117062 275452
rect 117100 275418 117110 275452
rect 117110 275418 117134 275452
rect 117172 275418 117178 275452
rect 117178 275418 117206 275452
rect 116063 275357 116097 275359
rect 116063 275325 116097 275357
rect 116063 275255 116097 275287
rect 116063 275253 116097 275255
rect 117273 275357 117307 275359
rect 117273 275325 117307 275357
rect 117273 275255 117307 275287
rect 117273 275253 117307 275255
rect 116164 275160 116192 275194
rect 116192 275160 116198 275194
rect 116236 275160 116260 275194
rect 116260 275160 116270 275194
rect 116308 275160 116328 275194
rect 116328 275160 116342 275194
rect 116380 275160 116396 275194
rect 116396 275160 116414 275194
rect 116452 275160 116464 275194
rect 116464 275160 116486 275194
rect 116524 275160 116532 275194
rect 116532 275160 116558 275194
rect 116596 275160 116600 275194
rect 116600 275160 116630 275194
rect 116668 275160 116702 275194
rect 116740 275160 116770 275194
rect 116770 275160 116774 275194
rect 116812 275160 116838 275194
rect 116838 275160 116846 275194
rect 116884 275160 116906 275194
rect 116906 275160 116918 275194
rect 116956 275160 116974 275194
rect 116974 275160 116990 275194
rect 117028 275160 117042 275194
rect 117042 275160 117062 275194
rect 117100 275160 117110 275194
rect 117110 275160 117134 275194
rect 117172 275160 117178 275194
rect 117178 275160 117206 275194
rect 117610 275474 117638 275508
rect 117638 275474 117644 275508
rect 117682 275474 117706 275508
rect 117706 275474 117716 275508
rect 117754 275474 117774 275508
rect 117774 275474 117788 275508
rect 117826 275474 117842 275508
rect 117842 275474 117860 275508
rect 117898 275474 117910 275508
rect 117910 275474 117932 275508
rect 117970 275474 117978 275508
rect 117978 275474 118004 275508
rect 118042 275474 118046 275508
rect 118046 275474 118076 275508
rect 118114 275474 118148 275508
rect 118186 275474 118216 275508
rect 118216 275474 118220 275508
rect 118258 275474 118284 275508
rect 118284 275474 118292 275508
rect 118330 275474 118352 275508
rect 118352 275474 118364 275508
rect 118402 275474 118420 275508
rect 118420 275474 118436 275508
rect 118474 275474 118488 275508
rect 118488 275474 118508 275508
rect 118546 275474 118556 275508
rect 118556 275474 118580 275508
rect 118618 275474 118624 275508
rect 118624 275474 118652 275508
rect 117509 275433 117543 275435
rect 117509 275401 117543 275433
rect 117509 275331 117543 275363
rect 117509 275329 117543 275331
rect 118719 275433 118753 275435
rect 118719 275401 118753 275433
rect 118719 275331 118753 275363
rect 118719 275329 118753 275331
rect 117610 275256 117638 275290
rect 117638 275256 117644 275290
rect 117682 275256 117706 275290
rect 117706 275256 117716 275290
rect 117754 275256 117774 275290
rect 117774 275256 117788 275290
rect 117826 275256 117842 275290
rect 117842 275256 117860 275290
rect 117898 275256 117910 275290
rect 117910 275256 117932 275290
rect 117970 275256 117978 275290
rect 117978 275256 118004 275290
rect 118042 275256 118046 275290
rect 118046 275256 118076 275290
rect 118114 275256 118148 275290
rect 118186 275256 118216 275290
rect 118216 275256 118220 275290
rect 118258 275256 118284 275290
rect 118284 275256 118292 275290
rect 118330 275256 118352 275290
rect 118352 275256 118364 275290
rect 118402 275256 118420 275290
rect 118420 275256 118436 275290
rect 118474 275256 118488 275290
rect 118488 275256 118508 275290
rect 118546 275256 118556 275290
rect 118556 275256 118580 275290
rect 118618 275256 118624 275290
rect 118624 275256 118652 275290
rect 111553 274754 111581 274788
rect 111581 274754 111587 274788
rect 111625 274754 111649 274788
rect 111649 274754 111659 274788
rect 111697 274754 111717 274788
rect 111717 274754 111731 274788
rect 111769 274754 111785 274788
rect 111785 274754 111803 274788
rect 111841 274754 111853 274788
rect 111853 274754 111875 274788
rect 111913 274754 111921 274788
rect 111921 274754 111947 274788
rect 111985 274754 111989 274788
rect 111989 274754 112019 274788
rect 112057 274754 112091 274788
rect 112129 274754 112159 274788
rect 112159 274754 112163 274788
rect 112201 274754 112227 274788
rect 112227 274754 112235 274788
rect 112273 274754 112295 274788
rect 112295 274754 112307 274788
rect 112345 274754 112363 274788
rect 112363 274754 112379 274788
rect 112417 274754 112431 274788
rect 112431 274754 112451 274788
rect 112489 274754 112499 274788
rect 112499 274754 112523 274788
rect 112561 274754 112567 274788
rect 112567 274754 112595 274788
rect 111452 274713 111486 274715
rect 111452 274681 111486 274713
rect 111452 274611 111486 274643
rect 111452 274609 111486 274611
rect 113029 274718 113057 274752
rect 113057 274718 113063 274752
rect 113101 274718 113125 274752
rect 113125 274718 113135 274752
rect 113173 274718 113193 274752
rect 113193 274718 113207 274752
rect 113245 274718 113261 274752
rect 113261 274718 113279 274752
rect 113317 274718 113329 274752
rect 113329 274718 113351 274752
rect 113389 274718 113397 274752
rect 113397 274718 113423 274752
rect 113461 274718 113465 274752
rect 113465 274718 113495 274752
rect 113533 274718 113567 274752
rect 113605 274718 113635 274752
rect 113635 274718 113639 274752
rect 113677 274718 113703 274752
rect 113703 274718 113711 274752
rect 113749 274718 113771 274752
rect 113771 274718 113783 274752
rect 113821 274718 113839 274752
rect 113839 274718 113855 274752
rect 113893 274718 113907 274752
rect 113907 274718 113927 274752
rect 113965 274718 113975 274752
rect 113975 274718 113999 274752
rect 114037 274718 114043 274752
rect 114043 274718 114071 274752
rect 112662 274713 112696 274715
rect 112662 274681 112696 274713
rect 112662 274611 112696 274643
rect 112928 274649 112962 274683
rect 114138 274649 114172 274683
rect 112662 274609 112696 274611
rect 113029 274580 113057 274614
rect 113057 274580 113063 274614
rect 113101 274580 113125 274614
rect 113125 274580 113135 274614
rect 113173 274580 113193 274614
rect 113193 274580 113207 274614
rect 113245 274580 113261 274614
rect 113261 274580 113279 274614
rect 113317 274580 113329 274614
rect 113329 274580 113351 274614
rect 113389 274580 113397 274614
rect 113397 274580 113423 274614
rect 113461 274580 113465 274614
rect 113465 274580 113495 274614
rect 113533 274580 113567 274614
rect 113605 274580 113635 274614
rect 113635 274580 113639 274614
rect 113677 274580 113703 274614
rect 113703 274580 113711 274614
rect 113749 274580 113771 274614
rect 113771 274580 113783 274614
rect 113821 274580 113839 274614
rect 113839 274580 113855 274614
rect 113893 274580 113907 274614
rect 113907 274580 113927 274614
rect 113965 274580 113975 274614
rect 113975 274580 113999 274614
rect 114037 274580 114043 274614
rect 114043 274580 114071 274614
rect 114704 274913 114706 274947
rect 114706 274913 114738 274947
rect 114776 274913 114808 274947
rect 114808 274913 114810 274947
rect 111553 274536 111581 274570
rect 111581 274536 111587 274570
rect 111625 274536 111649 274570
rect 111649 274536 111659 274570
rect 111697 274536 111717 274570
rect 111717 274536 111731 274570
rect 111769 274536 111785 274570
rect 111785 274536 111803 274570
rect 111841 274536 111853 274570
rect 111853 274536 111875 274570
rect 111913 274536 111921 274570
rect 111921 274536 111947 274570
rect 111985 274536 111989 274570
rect 111989 274536 112019 274570
rect 112057 274536 112091 274570
rect 112129 274536 112159 274570
rect 112159 274536 112163 274570
rect 112201 274536 112227 274570
rect 112227 274536 112235 274570
rect 112273 274536 112295 274570
rect 112295 274536 112307 274570
rect 112345 274536 112363 274570
rect 112363 274536 112379 274570
rect 112417 274536 112431 274570
rect 112431 274536 112451 274570
rect 112489 274536 112499 274570
rect 112499 274536 112523 274570
rect 112561 274536 112567 274570
rect 112567 274536 112595 274570
rect 114899 274822 114933 274856
rect 115395 274913 115397 274947
rect 115397 274913 115429 274947
rect 115467 274913 115499 274947
rect 115499 274913 115501 274947
rect 114704 274723 114706 274757
rect 114706 274723 114738 274757
rect 114776 274723 114808 274757
rect 114808 274723 114810 274757
rect 114576 274682 114610 274684
rect 114576 274650 114610 274682
rect 114576 274580 114610 274612
rect 114576 274578 114610 274580
rect 114904 274682 114938 274684
rect 114904 274650 114938 274682
rect 114904 274580 114938 274612
rect 114904 274578 114938 274580
rect 115271 274822 115305 274856
rect 115395 274723 115397 274757
rect 115397 274723 115429 274757
rect 115467 274723 115499 274757
rect 115499 274723 115501 274757
rect 115267 274682 115301 274684
rect 115267 274650 115301 274682
rect 115267 274580 115301 274612
rect 115267 274578 115301 274580
rect 115595 274682 115629 274684
rect 115595 274650 115629 274682
rect 115595 274580 115629 274612
rect 115595 274578 115629 274580
rect 116134 275016 116162 275050
rect 116162 275016 116168 275050
rect 116206 275016 116230 275050
rect 116230 275016 116240 275050
rect 116278 275016 116298 275050
rect 116298 275016 116312 275050
rect 116350 275016 116366 275050
rect 116366 275016 116384 275050
rect 116422 275016 116434 275050
rect 116434 275016 116456 275050
rect 116494 275016 116502 275050
rect 116502 275016 116528 275050
rect 116566 275016 116570 275050
rect 116570 275016 116600 275050
rect 116638 275016 116672 275050
rect 116710 275016 116740 275050
rect 116740 275016 116744 275050
rect 116782 275016 116808 275050
rect 116808 275016 116816 275050
rect 116854 275016 116876 275050
rect 116876 275016 116888 275050
rect 116926 275016 116944 275050
rect 116944 275016 116960 275050
rect 116998 275016 117012 275050
rect 117012 275016 117032 275050
rect 117070 275016 117080 275050
rect 117080 275016 117104 275050
rect 117142 275016 117148 275050
rect 117148 275016 117176 275050
rect 115828 274919 115862 274953
rect 116033 274947 116067 274981
rect 117243 274947 117277 274981
rect 116134 274878 116162 274912
rect 116162 274878 116168 274912
rect 116206 274878 116230 274912
rect 116230 274878 116240 274912
rect 116278 274878 116298 274912
rect 116298 274878 116312 274912
rect 116350 274878 116366 274912
rect 116366 274878 116384 274912
rect 116422 274878 116434 274912
rect 116434 274878 116456 274912
rect 116494 274878 116502 274912
rect 116502 274878 116528 274912
rect 116566 274878 116570 274912
rect 116570 274878 116600 274912
rect 116638 274878 116672 274912
rect 116710 274878 116740 274912
rect 116740 274878 116744 274912
rect 116782 274878 116808 274912
rect 116808 274878 116816 274912
rect 116854 274878 116876 274912
rect 116876 274878 116888 274912
rect 116926 274878 116944 274912
rect 116944 274878 116960 274912
rect 116998 274878 117012 274912
rect 117012 274878 117032 274912
rect 117070 274878 117080 274912
rect 117080 274878 117104 274912
rect 117142 274878 117148 274912
rect 117148 274878 117176 274912
rect 117610 275114 117638 275148
rect 117638 275114 117644 275148
rect 117682 275114 117706 275148
rect 117706 275114 117716 275148
rect 117754 275114 117774 275148
rect 117774 275114 117788 275148
rect 117826 275114 117842 275148
rect 117842 275114 117860 275148
rect 117898 275114 117910 275148
rect 117910 275114 117932 275148
rect 117970 275114 117978 275148
rect 117978 275114 118004 275148
rect 118042 275114 118046 275148
rect 118046 275114 118076 275148
rect 118114 275114 118148 275148
rect 118186 275114 118216 275148
rect 118216 275114 118220 275148
rect 118258 275114 118284 275148
rect 118284 275114 118292 275148
rect 118330 275114 118352 275148
rect 118352 275114 118364 275148
rect 118402 275114 118420 275148
rect 118420 275114 118436 275148
rect 118474 275114 118488 275148
rect 118488 275114 118508 275148
rect 118546 275114 118556 275148
rect 118556 275114 118580 275148
rect 118618 275114 118624 275148
rect 118624 275114 118652 275148
rect 117509 275073 117543 275075
rect 117509 275041 117543 275073
rect 117509 274971 117543 275003
rect 117509 274969 117543 274971
rect 118719 275073 118753 275075
rect 118719 275041 118753 275073
rect 118719 274971 118753 275003
rect 118719 274969 118753 274971
rect 117610 274896 117638 274930
rect 117638 274896 117644 274930
rect 117682 274896 117706 274930
rect 117706 274896 117716 274930
rect 117754 274896 117774 274930
rect 117774 274896 117788 274930
rect 117826 274896 117842 274930
rect 117842 274896 117860 274930
rect 117898 274896 117910 274930
rect 117910 274896 117932 274930
rect 117970 274896 117978 274930
rect 117978 274896 118004 274930
rect 118042 274896 118046 274930
rect 118046 274896 118076 274930
rect 118114 274896 118148 274930
rect 118186 274896 118216 274930
rect 118216 274896 118220 274930
rect 118258 274896 118284 274930
rect 118284 274896 118292 274930
rect 118330 274896 118352 274930
rect 118352 274896 118364 274930
rect 118402 274896 118420 274930
rect 118420 274896 118436 274930
rect 118474 274896 118488 274930
rect 118488 274896 118508 274930
rect 118546 274896 118556 274930
rect 118556 274896 118580 274930
rect 118618 274896 118624 274930
rect 118624 274896 118652 274930
rect 117610 274754 117638 274788
rect 117638 274754 117644 274788
rect 117682 274754 117706 274788
rect 117706 274754 117716 274788
rect 117754 274754 117774 274788
rect 117774 274754 117788 274788
rect 117826 274754 117842 274788
rect 117842 274754 117860 274788
rect 117898 274754 117910 274788
rect 117910 274754 117932 274788
rect 117970 274754 117978 274788
rect 117978 274754 118004 274788
rect 118042 274754 118046 274788
rect 118046 274754 118076 274788
rect 118114 274754 118148 274788
rect 118186 274754 118216 274788
rect 118216 274754 118220 274788
rect 118258 274754 118284 274788
rect 118284 274754 118292 274788
rect 118330 274754 118352 274788
rect 118352 274754 118364 274788
rect 118402 274754 118420 274788
rect 118420 274754 118436 274788
rect 118474 274754 118488 274788
rect 118488 274754 118508 274788
rect 118546 274754 118556 274788
rect 118556 274754 118580 274788
rect 118618 274754 118624 274788
rect 118624 274754 118652 274788
rect 116134 274718 116162 274752
rect 116162 274718 116168 274752
rect 116206 274718 116230 274752
rect 116230 274718 116240 274752
rect 116278 274718 116298 274752
rect 116298 274718 116312 274752
rect 116350 274718 116366 274752
rect 116366 274718 116384 274752
rect 116422 274718 116434 274752
rect 116434 274718 116456 274752
rect 116494 274718 116502 274752
rect 116502 274718 116528 274752
rect 116566 274718 116570 274752
rect 116570 274718 116600 274752
rect 116638 274718 116672 274752
rect 116710 274718 116740 274752
rect 116740 274718 116744 274752
rect 116782 274718 116808 274752
rect 116808 274718 116816 274752
rect 116854 274718 116876 274752
rect 116876 274718 116888 274752
rect 116926 274718 116944 274752
rect 116944 274718 116960 274752
rect 116998 274718 117012 274752
rect 117012 274718 117032 274752
rect 117070 274718 117080 274752
rect 117080 274718 117104 274752
rect 117142 274718 117148 274752
rect 117148 274718 117176 274752
rect 117509 274713 117543 274715
rect 116033 274649 116067 274683
rect 117243 274649 117277 274683
rect 117509 274681 117543 274713
rect 116134 274580 116162 274614
rect 116162 274580 116168 274614
rect 116206 274580 116230 274614
rect 116230 274580 116240 274614
rect 116278 274580 116298 274614
rect 116298 274580 116312 274614
rect 116350 274580 116366 274614
rect 116366 274580 116384 274614
rect 116422 274580 116434 274614
rect 116434 274580 116456 274614
rect 116494 274580 116502 274614
rect 116502 274580 116528 274614
rect 116566 274580 116570 274614
rect 116570 274580 116600 274614
rect 116638 274580 116672 274614
rect 116710 274580 116740 274614
rect 116740 274580 116744 274614
rect 116782 274580 116808 274614
rect 116808 274580 116816 274614
rect 116854 274580 116876 274614
rect 116876 274580 116888 274614
rect 116926 274580 116944 274614
rect 116944 274580 116960 274614
rect 116998 274580 117012 274614
rect 117012 274580 117032 274614
rect 117070 274580 117080 274614
rect 117080 274580 117104 274614
rect 117142 274580 117148 274614
rect 117148 274580 117176 274614
rect 117509 274611 117543 274643
rect 117509 274609 117543 274611
rect 118719 274713 118753 274715
rect 118719 274681 118753 274713
rect 118719 274611 118753 274643
rect 118719 274609 118753 274611
rect 114704 274505 114706 274539
rect 114706 274505 114738 274539
rect 114776 274505 114808 274539
rect 114808 274505 114810 274539
rect 115395 274505 115397 274539
rect 115397 274505 115429 274539
rect 115467 274505 115499 274539
rect 115499 274505 115501 274539
rect 117610 274536 117638 274570
rect 117638 274536 117644 274570
rect 117682 274536 117706 274570
rect 117706 274536 117716 274570
rect 117754 274536 117774 274570
rect 117774 274536 117788 274570
rect 117826 274536 117842 274570
rect 117842 274536 117860 274570
rect 117898 274536 117910 274570
rect 117910 274536 117932 274570
rect 117970 274536 117978 274570
rect 117978 274536 118004 274570
rect 118042 274536 118046 274570
rect 118046 274536 118076 274570
rect 118114 274536 118148 274570
rect 118186 274536 118216 274570
rect 118216 274536 118220 274570
rect 118258 274536 118284 274570
rect 118284 274536 118292 274570
rect 118330 274536 118352 274570
rect 118352 274536 118364 274570
rect 118402 274536 118420 274570
rect 118420 274536 118436 274570
rect 118474 274536 118488 274570
rect 118488 274536 118508 274570
rect 118546 274536 118556 274570
rect 118556 274536 118580 274570
rect 118618 274536 118624 274570
rect 118624 274536 118652 274570
rect 114034 274399 114068 274401
rect 114106 274399 114140 274401
rect 114178 274399 114212 274401
rect 114034 274367 114060 274399
rect 114060 274367 114068 274399
rect 114106 274367 114128 274399
rect 114128 274367 114140 274399
rect 114178 274367 114196 274399
rect 114196 274367 114212 274399
rect 115992 274399 116026 274401
rect 116064 274399 116098 274401
rect 116136 274399 116170 274401
rect 115992 274367 116009 274399
rect 116009 274367 116026 274399
rect 116064 274367 116077 274399
rect 116077 274367 116098 274399
rect 116136 274367 116145 274399
rect 116145 274367 116170 274399
rect 111553 274168 111581 274202
rect 111581 274168 111587 274202
rect 111625 274168 111649 274202
rect 111649 274168 111659 274202
rect 111697 274168 111717 274202
rect 111717 274168 111731 274202
rect 111769 274168 111785 274202
rect 111785 274168 111803 274202
rect 111841 274168 111853 274202
rect 111853 274168 111875 274202
rect 111913 274168 111921 274202
rect 111921 274168 111947 274202
rect 111985 274168 111989 274202
rect 111989 274168 112019 274202
rect 112057 274168 112091 274202
rect 112129 274168 112159 274202
rect 112159 274168 112163 274202
rect 112201 274168 112227 274202
rect 112227 274168 112235 274202
rect 112273 274168 112295 274202
rect 112295 274168 112307 274202
rect 112345 274168 112363 274202
rect 112363 274168 112379 274202
rect 112417 274168 112431 274202
rect 112431 274168 112451 274202
rect 112489 274168 112499 274202
rect 112499 274168 112523 274202
rect 112561 274168 112567 274202
rect 112567 274168 112595 274202
rect 111452 274127 111486 274129
rect 111452 274095 111486 274127
rect 111452 274025 111486 274057
rect 111452 274023 111486 274025
rect 112662 274127 112696 274129
rect 112662 274095 112696 274127
rect 112662 274025 112696 274057
rect 112662 274023 112696 274025
rect 111553 273950 111581 273984
rect 111581 273950 111587 273984
rect 111625 273950 111649 273984
rect 111649 273950 111659 273984
rect 111697 273950 111717 273984
rect 111717 273950 111731 273984
rect 111769 273950 111785 273984
rect 111785 273950 111803 273984
rect 111841 273950 111853 273984
rect 111853 273950 111875 273984
rect 111913 273950 111921 273984
rect 111921 273950 111947 273984
rect 111985 273950 111989 273984
rect 111989 273950 112019 273984
rect 112057 273950 112091 273984
rect 112129 273950 112159 273984
rect 112159 273950 112163 273984
rect 112201 273950 112227 273984
rect 112227 273950 112235 273984
rect 112273 273950 112295 273984
rect 112295 273950 112307 273984
rect 112345 273950 112363 273984
rect 112363 273950 112379 273984
rect 112417 273950 112431 273984
rect 112431 273950 112451 273984
rect 112489 273950 112499 273984
rect 112499 273950 112523 273984
rect 112561 273950 112567 273984
rect 112567 273950 112595 273984
rect 112999 274176 113027 274210
rect 113027 274176 113033 274210
rect 113071 274176 113095 274210
rect 113095 274176 113105 274210
rect 113143 274176 113163 274210
rect 113163 274176 113177 274210
rect 113215 274176 113231 274210
rect 113231 274176 113249 274210
rect 113287 274176 113299 274210
rect 113299 274176 113321 274210
rect 113359 274176 113367 274210
rect 113367 274176 113393 274210
rect 113431 274176 113435 274210
rect 113435 274176 113465 274210
rect 113503 274176 113537 274210
rect 113575 274176 113605 274210
rect 113605 274176 113609 274210
rect 113647 274176 113673 274210
rect 113673 274176 113681 274210
rect 113719 274176 113741 274210
rect 113741 274176 113753 274210
rect 113791 274176 113809 274210
rect 113809 274176 113825 274210
rect 113863 274176 113877 274210
rect 113877 274176 113897 274210
rect 113935 274176 113945 274210
rect 113945 274176 113969 274210
rect 114007 274176 114013 274210
rect 114013 274176 114041 274210
rect 112898 274115 112932 274117
rect 112898 274083 112932 274115
rect 112898 274013 112932 274045
rect 112898 274011 112932 274013
rect 114108 274115 114142 274117
rect 114108 274083 114142 274115
rect 114108 274013 114142 274045
rect 114108 274011 114142 274013
rect 114704 274151 114706 274185
rect 114706 274151 114738 274185
rect 114776 274151 114808 274185
rect 114808 274151 114810 274185
rect 112999 273918 113027 273952
rect 113027 273918 113033 273952
rect 113071 273918 113095 273952
rect 113095 273918 113105 273952
rect 113143 273918 113163 273952
rect 113163 273918 113177 273952
rect 113215 273918 113231 273952
rect 113231 273918 113249 273952
rect 113287 273918 113299 273952
rect 113299 273918 113321 273952
rect 113359 273918 113367 273952
rect 113367 273918 113393 273952
rect 113431 273918 113435 273952
rect 113435 273918 113465 273952
rect 113503 273918 113537 273952
rect 113575 273918 113605 273952
rect 113605 273918 113609 273952
rect 113647 273918 113673 273952
rect 113673 273918 113681 273952
rect 113719 273918 113741 273952
rect 113741 273918 113753 273952
rect 113791 273918 113809 273952
rect 113809 273918 113825 273952
rect 113863 273918 113877 273952
rect 113877 273918 113897 273952
rect 113935 273918 113945 273952
rect 113945 273918 113969 273952
rect 114007 273918 114013 273952
rect 114013 273918 114041 273952
rect 111553 273808 111581 273842
rect 111581 273808 111587 273842
rect 111625 273808 111649 273842
rect 111649 273808 111659 273842
rect 111697 273808 111717 273842
rect 111717 273808 111731 273842
rect 111769 273808 111785 273842
rect 111785 273808 111803 273842
rect 111841 273808 111853 273842
rect 111853 273808 111875 273842
rect 111913 273808 111921 273842
rect 111921 273808 111947 273842
rect 111985 273808 111989 273842
rect 111989 273808 112019 273842
rect 112057 273808 112091 273842
rect 112129 273808 112159 273842
rect 112159 273808 112163 273842
rect 112201 273808 112227 273842
rect 112227 273808 112235 273842
rect 112273 273808 112295 273842
rect 112295 273808 112307 273842
rect 112345 273808 112363 273842
rect 112363 273808 112379 273842
rect 112417 273808 112431 273842
rect 112431 273808 112451 273842
rect 112489 273808 112499 273842
rect 112499 273808 112523 273842
rect 112561 273808 112567 273842
rect 112567 273808 112595 273842
rect 111452 273767 111486 273769
rect 111452 273735 111486 273767
rect 111452 273665 111486 273697
rect 111452 273663 111486 273665
rect 112662 273767 112696 273769
rect 112662 273735 112696 273767
rect 112662 273665 112696 273697
rect 112662 273663 112696 273665
rect 111553 273590 111581 273624
rect 111581 273590 111587 273624
rect 111625 273590 111649 273624
rect 111649 273590 111659 273624
rect 111697 273590 111717 273624
rect 111717 273590 111731 273624
rect 111769 273590 111785 273624
rect 111785 273590 111803 273624
rect 111841 273590 111853 273624
rect 111853 273590 111875 273624
rect 111913 273590 111921 273624
rect 111921 273590 111947 273624
rect 111985 273590 111989 273624
rect 111989 273590 112019 273624
rect 112057 273590 112091 273624
rect 112129 273590 112159 273624
rect 112159 273590 112163 273624
rect 112201 273590 112227 273624
rect 112227 273590 112235 273624
rect 112273 273590 112295 273624
rect 112295 273590 112307 273624
rect 112345 273590 112363 273624
rect 112363 273590 112379 273624
rect 112417 273590 112431 273624
rect 112431 273590 112451 273624
rect 112489 273590 112499 273624
rect 112499 273590 112523 273624
rect 112561 273590 112567 273624
rect 112567 273590 112595 273624
rect 112999 273752 113027 273786
rect 113027 273752 113033 273786
rect 113071 273752 113095 273786
rect 113095 273752 113105 273786
rect 113143 273752 113163 273786
rect 113163 273752 113177 273786
rect 113215 273752 113231 273786
rect 113231 273752 113249 273786
rect 113287 273752 113299 273786
rect 113299 273752 113321 273786
rect 113359 273752 113367 273786
rect 113367 273752 113393 273786
rect 113431 273752 113435 273786
rect 113435 273752 113465 273786
rect 113503 273752 113537 273786
rect 113575 273752 113605 273786
rect 113605 273752 113609 273786
rect 113647 273752 113673 273786
rect 113673 273752 113681 273786
rect 113719 273752 113741 273786
rect 113741 273752 113753 273786
rect 113791 273752 113809 273786
rect 113809 273752 113825 273786
rect 113863 273752 113877 273786
rect 113877 273752 113897 273786
rect 113935 273752 113945 273786
rect 113945 273752 113969 273786
rect 114007 273752 114013 273786
rect 114013 273752 114041 273786
rect 112898 273691 112932 273693
rect 112898 273659 112932 273691
rect 112898 273589 112932 273621
rect 112898 273587 112932 273589
rect 114108 273691 114142 273693
rect 114108 273659 114142 273691
rect 114108 273589 114142 273621
rect 114108 273587 114142 273589
rect 112999 273494 113027 273528
rect 113027 273494 113033 273528
rect 113071 273494 113095 273528
rect 113095 273494 113105 273528
rect 113143 273494 113163 273528
rect 113163 273494 113177 273528
rect 113215 273494 113231 273528
rect 113231 273494 113249 273528
rect 113287 273494 113299 273528
rect 113299 273494 113321 273528
rect 113359 273494 113367 273528
rect 113367 273494 113393 273528
rect 113431 273494 113435 273528
rect 113435 273494 113465 273528
rect 113503 273494 113537 273528
rect 113575 273494 113605 273528
rect 113605 273494 113609 273528
rect 113647 273494 113673 273528
rect 113673 273494 113681 273528
rect 113719 273494 113741 273528
rect 113741 273494 113753 273528
rect 113791 273494 113809 273528
rect 113809 273494 113825 273528
rect 113863 273494 113877 273528
rect 113877 273494 113897 273528
rect 113935 273494 113945 273528
rect 113945 273494 113969 273528
rect 114007 273494 114013 273528
rect 114013 273494 114041 273528
rect 111553 273448 111581 273482
rect 111581 273448 111587 273482
rect 111625 273448 111649 273482
rect 111649 273448 111659 273482
rect 111697 273448 111717 273482
rect 111717 273448 111731 273482
rect 111769 273448 111785 273482
rect 111785 273448 111803 273482
rect 111841 273448 111853 273482
rect 111853 273448 111875 273482
rect 111913 273448 111921 273482
rect 111921 273448 111947 273482
rect 111985 273448 111989 273482
rect 111989 273448 112019 273482
rect 112057 273448 112091 273482
rect 112129 273448 112159 273482
rect 112159 273448 112163 273482
rect 112201 273448 112227 273482
rect 112227 273448 112235 273482
rect 112273 273448 112295 273482
rect 112295 273448 112307 273482
rect 112345 273448 112363 273482
rect 112363 273448 112379 273482
rect 112417 273448 112431 273482
rect 112431 273448 112451 273482
rect 112489 273448 112499 273482
rect 112499 273448 112523 273482
rect 112561 273448 112567 273482
rect 112567 273448 112595 273482
rect 111452 273407 111486 273409
rect 111452 273375 111486 273407
rect 111452 273305 111486 273337
rect 111452 273303 111486 273305
rect 112662 273407 112696 273409
rect 112662 273375 112696 273407
rect 112662 273305 112696 273337
rect 112662 273303 112696 273305
rect 111553 273230 111581 273264
rect 111581 273230 111587 273264
rect 111625 273230 111649 273264
rect 111649 273230 111659 273264
rect 111697 273230 111717 273264
rect 111717 273230 111731 273264
rect 111769 273230 111785 273264
rect 111785 273230 111803 273264
rect 111841 273230 111853 273264
rect 111853 273230 111875 273264
rect 111913 273230 111921 273264
rect 111921 273230 111947 273264
rect 111985 273230 111989 273264
rect 111989 273230 112019 273264
rect 112057 273230 112091 273264
rect 112129 273230 112159 273264
rect 112159 273230 112163 273264
rect 112201 273230 112227 273264
rect 112227 273230 112235 273264
rect 112273 273230 112295 273264
rect 112295 273230 112307 273264
rect 112345 273230 112363 273264
rect 112363 273230 112379 273264
rect 112417 273230 112431 273264
rect 112431 273230 112451 273264
rect 112489 273230 112499 273264
rect 112499 273230 112523 273264
rect 112561 273230 112567 273264
rect 112567 273230 112595 273264
rect 113029 273350 113057 273384
rect 113057 273350 113063 273384
rect 113101 273350 113125 273384
rect 113125 273350 113135 273384
rect 113173 273350 113193 273384
rect 113193 273350 113207 273384
rect 113245 273350 113261 273384
rect 113261 273350 113279 273384
rect 113317 273350 113329 273384
rect 113329 273350 113351 273384
rect 113389 273350 113397 273384
rect 113397 273350 113423 273384
rect 113461 273350 113465 273384
rect 113465 273350 113495 273384
rect 113533 273350 113567 273384
rect 113605 273350 113635 273384
rect 113635 273350 113639 273384
rect 113677 273350 113703 273384
rect 113703 273350 113711 273384
rect 113749 273350 113771 273384
rect 113771 273350 113783 273384
rect 113821 273350 113839 273384
rect 113839 273350 113855 273384
rect 113893 273350 113907 273384
rect 113907 273350 113927 273384
rect 113965 273350 113975 273384
rect 113975 273350 113999 273384
rect 114037 273350 114043 273384
rect 114043 273350 114071 273384
rect 112928 273281 112962 273315
rect 114138 273281 114172 273315
rect 114342 273253 114376 273287
rect 113029 273212 113057 273246
rect 113057 273212 113063 273246
rect 113101 273212 113125 273246
rect 113125 273212 113135 273246
rect 113173 273212 113193 273246
rect 113193 273212 113207 273246
rect 113245 273212 113261 273246
rect 113261 273212 113279 273246
rect 113317 273212 113329 273246
rect 113329 273212 113351 273246
rect 113389 273212 113397 273246
rect 113397 273212 113423 273246
rect 113461 273212 113465 273246
rect 113465 273212 113495 273246
rect 113533 273212 113567 273246
rect 113605 273212 113635 273246
rect 113635 273212 113639 273246
rect 113677 273212 113703 273246
rect 113703 273212 113711 273246
rect 113749 273212 113771 273246
rect 113771 273212 113783 273246
rect 113821 273212 113839 273246
rect 113839 273212 113855 273246
rect 113893 273212 113907 273246
rect 113907 273212 113927 273246
rect 113965 273212 113975 273246
rect 113975 273212 113999 273246
rect 114037 273212 114043 273246
rect 114043 273212 114071 273246
rect 114576 274092 114610 274100
rect 114576 274066 114610 274092
rect 114576 274024 114610 274028
rect 114576 273994 114610 274024
rect 114576 273922 114610 273956
rect 114576 273854 114610 273884
rect 114576 273850 114610 273854
rect 114576 273786 114610 273812
rect 114576 273778 114610 273786
rect 114904 274092 114938 274100
rect 114904 274066 114938 274092
rect 114904 274024 114938 274028
rect 114904 273994 114938 274024
rect 114904 273922 114938 273956
rect 114904 273854 114938 273884
rect 114904 273850 114938 273854
rect 114904 273786 114938 273812
rect 114904 273778 114938 273786
rect 114704 273693 114706 273727
rect 114706 273693 114738 273727
rect 114776 273693 114808 273727
rect 114808 273693 114810 273727
rect 115395 274151 115397 274185
rect 115397 274151 115429 274185
rect 115467 274151 115499 274185
rect 115499 274151 115501 274185
rect 114899 273579 114933 273613
rect 115267 274092 115301 274100
rect 115267 274066 115301 274092
rect 115267 274024 115301 274028
rect 115267 273994 115301 274024
rect 115267 273922 115301 273956
rect 115267 273854 115301 273884
rect 115267 273850 115301 273854
rect 115267 273786 115301 273812
rect 115267 273778 115301 273786
rect 115595 274092 115629 274100
rect 115595 274066 115629 274092
rect 115595 274024 115629 274028
rect 115595 273994 115629 274024
rect 115595 273922 115629 273956
rect 115595 273854 115629 273884
rect 115595 273850 115629 273854
rect 115595 273786 115629 273812
rect 115595 273778 115629 273786
rect 115395 273693 115397 273727
rect 115397 273693 115429 273727
rect 115467 273693 115499 273727
rect 115499 273693 115501 273727
rect 114704 273465 114706 273499
rect 114706 273465 114738 273499
rect 114776 273465 114808 273499
rect 114808 273465 114810 273499
rect 114576 273424 114610 273426
rect 114576 273392 114610 273424
rect 114576 273322 114610 273354
rect 114576 273320 114610 273322
rect 114904 273424 114938 273426
rect 114904 273392 114938 273424
rect 114904 273322 114938 273354
rect 114904 273320 114938 273322
rect 115271 273579 115305 273613
rect 115395 273465 115397 273499
rect 115397 273465 115429 273499
rect 115467 273465 115499 273499
rect 115499 273465 115501 273499
rect 115267 273424 115301 273426
rect 115267 273392 115301 273424
rect 115267 273322 115301 273354
rect 115267 273320 115301 273322
rect 115595 273424 115629 273426
rect 115595 273392 115629 273424
rect 115595 273322 115629 273354
rect 115595 273320 115629 273322
rect 116164 274176 116192 274210
rect 116192 274176 116198 274210
rect 116236 274176 116260 274210
rect 116260 274176 116270 274210
rect 116308 274176 116328 274210
rect 116328 274176 116342 274210
rect 116380 274176 116396 274210
rect 116396 274176 116414 274210
rect 116452 274176 116464 274210
rect 116464 274176 116486 274210
rect 116524 274176 116532 274210
rect 116532 274176 116558 274210
rect 116596 274176 116600 274210
rect 116600 274176 116630 274210
rect 116668 274176 116702 274210
rect 116740 274176 116770 274210
rect 116770 274176 116774 274210
rect 116812 274176 116838 274210
rect 116838 274176 116846 274210
rect 116884 274176 116906 274210
rect 116906 274176 116918 274210
rect 116956 274176 116974 274210
rect 116974 274176 116990 274210
rect 117028 274176 117042 274210
rect 117042 274176 117062 274210
rect 117100 274176 117110 274210
rect 117110 274176 117134 274210
rect 117172 274176 117178 274210
rect 117178 274176 117206 274210
rect 116063 274115 116097 274117
rect 116063 274083 116097 274115
rect 116063 274013 116097 274045
rect 116063 274011 116097 274013
rect 117273 274115 117307 274117
rect 117273 274083 117307 274115
rect 117273 274013 117307 274045
rect 117273 274011 117307 274013
rect 116164 273918 116192 273952
rect 116192 273918 116198 273952
rect 116236 273918 116260 273952
rect 116260 273918 116270 273952
rect 116308 273918 116328 273952
rect 116328 273918 116342 273952
rect 116380 273918 116396 273952
rect 116396 273918 116414 273952
rect 116452 273918 116464 273952
rect 116464 273918 116486 273952
rect 116524 273918 116532 273952
rect 116532 273918 116558 273952
rect 116596 273918 116600 273952
rect 116600 273918 116630 273952
rect 116668 273918 116702 273952
rect 116740 273918 116770 273952
rect 116770 273918 116774 273952
rect 116812 273918 116838 273952
rect 116838 273918 116846 273952
rect 116884 273918 116906 273952
rect 116906 273918 116918 273952
rect 116956 273918 116974 273952
rect 116974 273918 116990 273952
rect 117028 273918 117042 273952
rect 117042 273918 117062 273952
rect 117100 273918 117110 273952
rect 117110 273918 117134 273952
rect 117172 273918 117178 273952
rect 117178 273918 117206 273952
rect 117610 274168 117638 274202
rect 117638 274168 117644 274202
rect 117682 274168 117706 274202
rect 117706 274168 117716 274202
rect 117754 274168 117774 274202
rect 117774 274168 117788 274202
rect 117826 274168 117842 274202
rect 117842 274168 117860 274202
rect 117898 274168 117910 274202
rect 117910 274168 117932 274202
rect 117970 274168 117978 274202
rect 117978 274168 118004 274202
rect 118042 274168 118046 274202
rect 118046 274168 118076 274202
rect 118114 274168 118148 274202
rect 118186 274168 118216 274202
rect 118216 274168 118220 274202
rect 118258 274168 118284 274202
rect 118284 274168 118292 274202
rect 118330 274168 118352 274202
rect 118352 274168 118364 274202
rect 118402 274168 118420 274202
rect 118420 274168 118436 274202
rect 118474 274168 118488 274202
rect 118488 274168 118508 274202
rect 118546 274168 118556 274202
rect 118556 274168 118580 274202
rect 118618 274168 118624 274202
rect 118624 274168 118652 274202
rect 117509 274127 117543 274129
rect 117509 274095 117543 274127
rect 117509 274025 117543 274057
rect 117509 274023 117543 274025
rect 118719 274127 118753 274129
rect 118719 274095 118753 274127
rect 118719 274025 118753 274057
rect 118719 274023 118753 274025
rect 117610 273950 117638 273984
rect 117638 273950 117644 273984
rect 117682 273950 117706 273984
rect 117706 273950 117716 273984
rect 117754 273950 117774 273984
rect 117774 273950 117788 273984
rect 117826 273950 117842 273984
rect 117842 273950 117860 273984
rect 117898 273950 117910 273984
rect 117910 273950 117932 273984
rect 117970 273950 117978 273984
rect 117978 273950 118004 273984
rect 118042 273950 118046 273984
rect 118046 273950 118076 273984
rect 118114 273950 118148 273984
rect 118186 273950 118216 273984
rect 118216 273950 118220 273984
rect 118258 273950 118284 273984
rect 118284 273950 118292 273984
rect 118330 273950 118352 273984
rect 118352 273950 118364 273984
rect 118402 273950 118420 273984
rect 118420 273950 118436 273984
rect 118474 273950 118488 273984
rect 118488 273950 118508 273984
rect 118546 273950 118556 273984
rect 118556 273950 118580 273984
rect 118618 273950 118624 273984
rect 118624 273950 118652 273984
rect 116164 273752 116192 273786
rect 116192 273752 116198 273786
rect 116236 273752 116260 273786
rect 116260 273752 116270 273786
rect 116308 273752 116328 273786
rect 116328 273752 116342 273786
rect 116380 273752 116396 273786
rect 116396 273752 116414 273786
rect 116452 273752 116464 273786
rect 116464 273752 116486 273786
rect 116524 273752 116532 273786
rect 116532 273752 116558 273786
rect 116596 273752 116600 273786
rect 116600 273752 116630 273786
rect 116668 273752 116702 273786
rect 116740 273752 116770 273786
rect 116770 273752 116774 273786
rect 116812 273752 116838 273786
rect 116838 273752 116846 273786
rect 116884 273752 116906 273786
rect 116906 273752 116918 273786
rect 116956 273752 116974 273786
rect 116974 273752 116990 273786
rect 117028 273752 117042 273786
rect 117042 273752 117062 273786
rect 117100 273752 117110 273786
rect 117110 273752 117134 273786
rect 117172 273752 117178 273786
rect 117178 273752 117206 273786
rect 116063 273691 116097 273693
rect 116063 273659 116097 273691
rect 116063 273589 116097 273621
rect 116063 273587 116097 273589
rect 117273 273691 117307 273693
rect 117273 273659 117307 273691
rect 117273 273589 117307 273621
rect 117273 273587 117307 273589
rect 116164 273494 116192 273528
rect 116192 273494 116198 273528
rect 116236 273494 116260 273528
rect 116260 273494 116270 273528
rect 116308 273494 116328 273528
rect 116328 273494 116342 273528
rect 116380 273494 116396 273528
rect 116396 273494 116414 273528
rect 116452 273494 116464 273528
rect 116464 273494 116486 273528
rect 116524 273494 116532 273528
rect 116532 273494 116558 273528
rect 116596 273494 116600 273528
rect 116600 273494 116630 273528
rect 116668 273494 116702 273528
rect 116740 273494 116770 273528
rect 116770 273494 116774 273528
rect 116812 273494 116838 273528
rect 116838 273494 116846 273528
rect 116884 273494 116906 273528
rect 116906 273494 116918 273528
rect 116956 273494 116974 273528
rect 116974 273494 116990 273528
rect 117028 273494 117042 273528
rect 117042 273494 117062 273528
rect 117100 273494 117110 273528
rect 117110 273494 117134 273528
rect 117172 273494 117178 273528
rect 117178 273494 117206 273528
rect 117610 273808 117638 273842
rect 117638 273808 117644 273842
rect 117682 273808 117706 273842
rect 117706 273808 117716 273842
rect 117754 273808 117774 273842
rect 117774 273808 117788 273842
rect 117826 273808 117842 273842
rect 117842 273808 117860 273842
rect 117898 273808 117910 273842
rect 117910 273808 117932 273842
rect 117970 273808 117978 273842
rect 117978 273808 118004 273842
rect 118042 273808 118046 273842
rect 118046 273808 118076 273842
rect 118114 273808 118148 273842
rect 118186 273808 118216 273842
rect 118216 273808 118220 273842
rect 118258 273808 118284 273842
rect 118284 273808 118292 273842
rect 118330 273808 118352 273842
rect 118352 273808 118364 273842
rect 118402 273808 118420 273842
rect 118420 273808 118436 273842
rect 118474 273808 118488 273842
rect 118488 273808 118508 273842
rect 118546 273808 118556 273842
rect 118556 273808 118580 273842
rect 118618 273808 118624 273842
rect 118624 273808 118652 273842
rect 117509 273767 117543 273769
rect 117509 273735 117543 273767
rect 117509 273665 117543 273697
rect 117509 273663 117543 273665
rect 118719 273767 118753 273769
rect 118719 273735 118753 273767
rect 118719 273665 118753 273697
rect 118719 273663 118753 273665
rect 117610 273590 117638 273624
rect 117638 273590 117644 273624
rect 117682 273590 117706 273624
rect 117706 273590 117716 273624
rect 117754 273590 117774 273624
rect 117774 273590 117788 273624
rect 117826 273590 117842 273624
rect 117842 273590 117860 273624
rect 117898 273590 117910 273624
rect 117910 273590 117932 273624
rect 117970 273590 117978 273624
rect 117978 273590 118004 273624
rect 118042 273590 118046 273624
rect 118046 273590 118076 273624
rect 118114 273590 118148 273624
rect 118186 273590 118216 273624
rect 118216 273590 118220 273624
rect 118258 273590 118284 273624
rect 118284 273590 118292 273624
rect 118330 273590 118352 273624
rect 118352 273590 118364 273624
rect 118402 273590 118420 273624
rect 118420 273590 118436 273624
rect 118474 273590 118488 273624
rect 118488 273590 118508 273624
rect 118546 273590 118556 273624
rect 118556 273590 118580 273624
rect 118618 273590 118624 273624
rect 118624 273590 118652 273624
rect 111553 273088 111581 273122
rect 111581 273088 111587 273122
rect 111625 273088 111649 273122
rect 111649 273088 111659 273122
rect 111697 273088 111717 273122
rect 111717 273088 111731 273122
rect 111769 273088 111785 273122
rect 111785 273088 111803 273122
rect 111841 273088 111853 273122
rect 111853 273088 111875 273122
rect 111913 273088 111921 273122
rect 111921 273088 111947 273122
rect 111985 273088 111989 273122
rect 111989 273088 112019 273122
rect 112057 273088 112091 273122
rect 112129 273088 112159 273122
rect 112159 273088 112163 273122
rect 112201 273088 112227 273122
rect 112227 273088 112235 273122
rect 112273 273088 112295 273122
rect 112295 273088 112307 273122
rect 112345 273088 112363 273122
rect 112363 273088 112379 273122
rect 112417 273088 112431 273122
rect 112431 273088 112451 273122
rect 112489 273088 112499 273122
rect 112499 273088 112523 273122
rect 112561 273088 112567 273122
rect 112567 273088 112595 273122
rect 111452 273047 111486 273049
rect 111452 273015 111486 273047
rect 111452 272945 111486 272977
rect 111452 272943 111486 272945
rect 113029 273052 113057 273086
rect 113057 273052 113063 273086
rect 113101 273052 113125 273086
rect 113125 273052 113135 273086
rect 113173 273052 113193 273086
rect 113193 273052 113207 273086
rect 113245 273052 113261 273086
rect 113261 273052 113279 273086
rect 113317 273052 113329 273086
rect 113329 273052 113351 273086
rect 113389 273052 113397 273086
rect 113397 273052 113423 273086
rect 113461 273052 113465 273086
rect 113465 273052 113495 273086
rect 113533 273052 113567 273086
rect 113605 273052 113635 273086
rect 113635 273052 113639 273086
rect 113677 273052 113703 273086
rect 113703 273052 113711 273086
rect 113749 273052 113771 273086
rect 113771 273052 113783 273086
rect 113821 273052 113839 273086
rect 113839 273052 113855 273086
rect 113893 273052 113907 273086
rect 113907 273052 113927 273086
rect 113965 273052 113975 273086
rect 113975 273052 113999 273086
rect 114037 273052 114043 273086
rect 114043 273052 114071 273086
rect 112662 273047 112696 273049
rect 112662 273015 112696 273047
rect 112662 272945 112696 272977
rect 112928 272983 112962 273017
rect 114138 272983 114172 273017
rect 112662 272943 112696 272945
rect 113029 272914 113057 272948
rect 113057 272914 113063 272948
rect 113101 272914 113125 272948
rect 113125 272914 113135 272948
rect 113173 272914 113193 272948
rect 113193 272914 113207 272948
rect 113245 272914 113261 272948
rect 113261 272914 113279 272948
rect 113317 272914 113329 272948
rect 113329 272914 113351 272948
rect 113389 272914 113397 272948
rect 113397 272914 113423 272948
rect 113461 272914 113465 272948
rect 113465 272914 113495 272948
rect 113533 272914 113567 272948
rect 113605 272914 113635 272948
rect 113635 272914 113639 272948
rect 113677 272914 113703 272948
rect 113703 272914 113711 272948
rect 113749 272914 113771 272948
rect 113771 272914 113783 272948
rect 113821 272914 113839 272948
rect 113839 272914 113855 272948
rect 113893 272914 113907 272948
rect 113907 272914 113927 272948
rect 113965 272914 113975 272948
rect 113975 272914 113999 272948
rect 114037 272914 114043 272948
rect 114043 272914 114071 272948
rect 114704 273247 114706 273281
rect 114706 273247 114738 273281
rect 114776 273247 114808 273281
rect 114808 273247 114810 273281
rect 111553 272870 111581 272904
rect 111581 272870 111587 272904
rect 111625 272870 111649 272904
rect 111649 272870 111659 272904
rect 111697 272870 111717 272904
rect 111717 272870 111731 272904
rect 111769 272870 111785 272904
rect 111785 272870 111803 272904
rect 111841 272870 111853 272904
rect 111853 272870 111875 272904
rect 111913 272870 111921 272904
rect 111921 272870 111947 272904
rect 111985 272870 111989 272904
rect 111989 272870 112019 272904
rect 112057 272870 112091 272904
rect 112129 272870 112159 272904
rect 112159 272870 112163 272904
rect 112201 272870 112227 272904
rect 112227 272870 112235 272904
rect 112273 272870 112295 272904
rect 112295 272870 112307 272904
rect 112345 272870 112363 272904
rect 112363 272870 112379 272904
rect 112417 272870 112431 272904
rect 112431 272870 112451 272904
rect 112489 272870 112499 272904
rect 112499 272870 112523 272904
rect 112561 272870 112567 272904
rect 112567 272870 112595 272904
rect 114899 273156 114933 273190
rect 115395 273247 115397 273281
rect 115397 273247 115429 273281
rect 115467 273247 115499 273281
rect 115499 273247 115501 273281
rect 114704 273057 114706 273091
rect 114706 273057 114738 273091
rect 114776 273057 114808 273091
rect 114808 273057 114810 273091
rect 114576 273016 114610 273018
rect 114576 272984 114610 273016
rect 114576 272914 114610 272946
rect 114576 272912 114610 272914
rect 114904 273016 114938 273018
rect 114904 272984 114938 273016
rect 114904 272914 114938 272946
rect 114904 272912 114938 272914
rect 115271 273156 115305 273190
rect 115395 273057 115397 273091
rect 115397 273057 115429 273091
rect 115467 273057 115499 273091
rect 115499 273057 115501 273091
rect 115267 273016 115301 273018
rect 115267 272984 115301 273016
rect 115267 272914 115301 272946
rect 115267 272912 115301 272914
rect 115595 273016 115629 273018
rect 115595 272984 115629 273016
rect 115595 272914 115629 272946
rect 115595 272912 115629 272914
rect 116134 273350 116162 273384
rect 116162 273350 116168 273384
rect 116206 273350 116230 273384
rect 116230 273350 116240 273384
rect 116278 273350 116298 273384
rect 116298 273350 116312 273384
rect 116350 273350 116366 273384
rect 116366 273350 116384 273384
rect 116422 273350 116434 273384
rect 116434 273350 116456 273384
rect 116494 273350 116502 273384
rect 116502 273350 116528 273384
rect 116566 273350 116570 273384
rect 116570 273350 116600 273384
rect 116638 273350 116672 273384
rect 116710 273350 116740 273384
rect 116740 273350 116744 273384
rect 116782 273350 116808 273384
rect 116808 273350 116816 273384
rect 116854 273350 116876 273384
rect 116876 273350 116888 273384
rect 116926 273350 116944 273384
rect 116944 273350 116960 273384
rect 116998 273350 117012 273384
rect 117012 273350 117032 273384
rect 117070 273350 117080 273384
rect 117080 273350 117104 273384
rect 117142 273350 117148 273384
rect 117148 273350 117176 273384
rect 115828 273253 115862 273287
rect 116033 273281 116067 273315
rect 117243 273281 117277 273315
rect 116134 273212 116162 273246
rect 116162 273212 116168 273246
rect 116206 273212 116230 273246
rect 116230 273212 116240 273246
rect 116278 273212 116298 273246
rect 116298 273212 116312 273246
rect 116350 273212 116366 273246
rect 116366 273212 116384 273246
rect 116422 273212 116434 273246
rect 116434 273212 116456 273246
rect 116494 273212 116502 273246
rect 116502 273212 116528 273246
rect 116566 273212 116570 273246
rect 116570 273212 116600 273246
rect 116638 273212 116672 273246
rect 116710 273212 116740 273246
rect 116740 273212 116744 273246
rect 116782 273212 116808 273246
rect 116808 273212 116816 273246
rect 116854 273212 116876 273246
rect 116876 273212 116888 273246
rect 116926 273212 116944 273246
rect 116944 273212 116960 273246
rect 116998 273212 117012 273246
rect 117012 273212 117032 273246
rect 117070 273212 117080 273246
rect 117080 273212 117104 273246
rect 117142 273212 117148 273246
rect 117148 273212 117176 273246
rect 117610 273448 117638 273482
rect 117638 273448 117644 273482
rect 117682 273448 117706 273482
rect 117706 273448 117716 273482
rect 117754 273448 117774 273482
rect 117774 273448 117788 273482
rect 117826 273448 117842 273482
rect 117842 273448 117860 273482
rect 117898 273448 117910 273482
rect 117910 273448 117932 273482
rect 117970 273448 117978 273482
rect 117978 273448 118004 273482
rect 118042 273448 118046 273482
rect 118046 273448 118076 273482
rect 118114 273448 118148 273482
rect 118186 273448 118216 273482
rect 118216 273448 118220 273482
rect 118258 273448 118284 273482
rect 118284 273448 118292 273482
rect 118330 273448 118352 273482
rect 118352 273448 118364 273482
rect 118402 273448 118420 273482
rect 118420 273448 118436 273482
rect 118474 273448 118488 273482
rect 118488 273448 118508 273482
rect 118546 273448 118556 273482
rect 118556 273448 118580 273482
rect 118618 273448 118624 273482
rect 118624 273448 118652 273482
rect 117509 273407 117543 273409
rect 117509 273375 117543 273407
rect 117509 273305 117543 273337
rect 117509 273303 117543 273305
rect 118719 273407 118753 273409
rect 118719 273375 118753 273407
rect 118719 273305 118753 273337
rect 118719 273303 118753 273305
rect 117610 273230 117638 273264
rect 117638 273230 117644 273264
rect 117682 273230 117706 273264
rect 117706 273230 117716 273264
rect 117754 273230 117774 273264
rect 117774 273230 117788 273264
rect 117826 273230 117842 273264
rect 117842 273230 117860 273264
rect 117898 273230 117910 273264
rect 117910 273230 117932 273264
rect 117970 273230 117978 273264
rect 117978 273230 118004 273264
rect 118042 273230 118046 273264
rect 118046 273230 118076 273264
rect 118114 273230 118148 273264
rect 118186 273230 118216 273264
rect 118216 273230 118220 273264
rect 118258 273230 118284 273264
rect 118284 273230 118292 273264
rect 118330 273230 118352 273264
rect 118352 273230 118364 273264
rect 118402 273230 118420 273264
rect 118420 273230 118436 273264
rect 118474 273230 118488 273264
rect 118488 273230 118508 273264
rect 118546 273230 118556 273264
rect 118556 273230 118580 273264
rect 118618 273230 118624 273264
rect 118624 273230 118652 273264
rect 117610 273088 117638 273122
rect 117638 273088 117644 273122
rect 117682 273088 117706 273122
rect 117706 273088 117716 273122
rect 117754 273088 117774 273122
rect 117774 273088 117788 273122
rect 117826 273088 117842 273122
rect 117842 273088 117860 273122
rect 117898 273088 117910 273122
rect 117910 273088 117932 273122
rect 117970 273088 117978 273122
rect 117978 273088 118004 273122
rect 118042 273088 118046 273122
rect 118046 273088 118076 273122
rect 118114 273088 118148 273122
rect 118186 273088 118216 273122
rect 118216 273088 118220 273122
rect 118258 273088 118284 273122
rect 118284 273088 118292 273122
rect 118330 273088 118352 273122
rect 118352 273088 118364 273122
rect 118402 273088 118420 273122
rect 118420 273088 118436 273122
rect 118474 273088 118488 273122
rect 118488 273088 118508 273122
rect 118546 273088 118556 273122
rect 118556 273088 118580 273122
rect 118618 273088 118624 273122
rect 118624 273088 118652 273122
rect 116134 273052 116162 273086
rect 116162 273052 116168 273086
rect 116206 273052 116230 273086
rect 116230 273052 116240 273086
rect 116278 273052 116298 273086
rect 116298 273052 116312 273086
rect 116350 273052 116366 273086
rect 116366 273052 116384 273086
rect 116422 273052 116434 273086
rect 116434 273052 116456 273086
rect 116494 273052 116502 273086
rect 116502 273052 116528 273086
rect 116566 273052 116570 273086
rect 116570 273052 116600 273086
rect 116638 273052 116672 273086
rect 116710 273052 116740 273086
rect 116740 273052 116744 273086
rect 116782 273052 116808 273086
rect 116808 273052 116816 273086
rect 116854 273052 116876 273086
rect 116876 273052 116888 273086
rect 116926 273052 116944 273086
rect 116944 273052 116960 273086
rect 116998 273052 117012 273086
rect 117012 273052 117032 273086
rect 117070 273052 117080 273086
rect 117080 273052 117104 273086
rect 117142 273052 117148 273086
rect 117148 273052 117176 273086
rect 117509 273047 117543 273049
rect 116033 272983 116067 273017
rect 117243 272983 117277 273017
rect 117509 273015 117543 273047
rect 116134 272914 116162 272948
rect 116162 272914 116168 272948
rect 116206 272914 116230 272948
rect 116230 272914 116240 272948
rect 116278 272914 116298 272948
rect 116298 272914 116312 272948
rect 116350 272914 116366 272948
rect 116366 272914 116384 272948
rect 116422 272914 116434 272948
rect 116434 272914 116456 272948
rect 116494 272914 116502 272948
rect 116502 272914 116528 272948
rect 116566 272914 116570 272948
rect 116570 272914 116600 272948
rect 116638 272914 116672 272948
rect 116710 272914 116740 272948
rect 116740 272914 116744 272948
rect 116782 272914 116808 272948
rect 116808 272914 116816 272948
rect 116854 272914 116876 272948
rect 116876 272914 116888 272948
rect 116926 272914 116944 272948
rect 116944 272914 116960 272948
rect 116998 272914 117012 272948
rect 117012 272914 117032 272948
rect 117070 272914 117080 272948
rect 117080 272914 117104 272948
rect 117142 272914 117148 272948
rect 117148 272914 117176 272948
rect 117509 272945 117543 272977
rect 117509 272943 117543 272945
rect 118719 273047 118753 273049
rect 118719 273015 118753 273047
rect 118719 272945 118753 272977
rect 118719 272943 118753 272945
rect 114704 272839 114706 272873
rect 114706 272839 114738 272873
rect 114776 272839 114808 272873
rect 114808 272839 114810 272873
rect 115395 272839 115397 272873
rect 115397 272839 115429 272873
rect 115467 272839 115499 272873
rect 115499 272839 115501 272873
rect 117610 272870 117638 272904
rect 117638 272870 117644 272904
rect 117682 272870 117706 272904
rect 117706 272870 117716 272904
rect 117754 272870 117774 272904
rect 117774 272870 117788 272904
rect 117826 272870 117842 272904
rect 117842 272870 117860 272904
rect 117898 272870 117910 272904
rect 117910 272870 117932 272904
rect 117970 272870 117978 272904
rect 117978 272870 118004 272904
rect 118042 272870 118046 272904
rect 118046 272870 118076 272904
rect 118114 272870 118148 272904
rect 118186 272870 118216 272904
rect 118216 272870 118220 272904
rect 118258 272870 118284 272904
rect 118284 272870 118292 272904
rect 118330 272870 118352 272904
rect 118352 272870 118364 272904
rect 118402 272870 118420 272904
rect 118420 272870 118436 272904
rect 118474 272870 118488 272904
rect 118488 272870 118508 272904
rect 118546 272870 118556 272904
rect 118556 272870 118580 272904
rect 118618 272870 118624 272904
rect 118624 272870 118652 272904
rect 114034 272733 114068 272735
rect 114106 272733 114140 272735
rect 114178 272733 114212 272735
rect 114034 272701 114060 272733
rect 114060 272701 114068 272733
rect 114106 272701 114128 272733
rect 114128 272701 114140 272733
rect 114178 272701 114196 272733
rect 114196 272701 114212 272733
rect 115016 272444 115194 272766
rect 115992 272733 116026 272735
rect 116064 272733 116098 272735
rect 116136 272733 116170 272735
rect 115992 272701 116009 272733
rect 116009 272701 116026 272733
rect 116064 272701 116077 272733
rect 116077 272701 116098 272733
rect 116136 272701 116145 272733
rect 116145 272701 116170 272733
rect 116644 272159 116678 272193
rect 116716 272159 116750 272193
rect 116788 272159 116822 272193
rect 116860 272159 116894 272193
rect 116932 272159 116966 272193
rect 117004 272159 117038 272193
rect 117076 272159 117110 272193
rect 117148 272159 117182 272193
rect 117220 272159 117254 272193
rect 117292 272159 117326 272193
rect 117364 272159 117398 272193
rect 117436 272159 117470 272193
rect 117508 272159 117542 272193
rect 117580 272159 117614 272193
rect 117652 272159 117686 272193
rect 117724 272159 117758 272193
rect 117796 272159 117830 272193
rect 117868 272159 117902 272193
rect 117940 272159 117974 272193
rect 118012 272159 118046 272193
rect 118084 272159 118118 272193
rect 113863 271731 114041 271981
rect 115019 271950 115053 271984
rect 115091 271950 115125 271984
rect 115163 271950 115197 271984
rect 115235 271950 115269 271984
rect 115307 271950 115341 271984
rect 115379 271950 115413 271984
rect 115451 271950 115485 271984
rect 115523 271950 115557 271984
rect 113100 271567 113134 271601
rect 113172 271567 113206 271601
rect 113244 271567 113278 271601
rect 113316 271567 113350 271601
rect 113388 271567 113422 271601
rect 112605 271353 112607 271387
rect 112607 271353 112639 271387
rect 112677 271353 112709 271387
rect 112709 271353 112711 271387
rect 113005 271353 113007 271387
rect 113007 271353 113039 271387
rect 113077 271353 113109 271387
rect 113109 271353 113111 271387
rect 113405 271353 113407 271387
rect 113407 271353 113439 271387
rect 113477 271353 113509 271387
rect 113509 271353 113511 271387
rect 113805 271353 113807 271387
rect 113807 271353 113839 271387
rect 113877 271353 113909 271387
rect 113909 271353 113911 271387
rect 112532 271257 112566 271259
rect 112532 271225 112566 271257
rect 112532 271155 112566 271187
rect 112532 271153 112566 271155
rect 112750 271257 112784 271259
rect 112750 271225 112784 271257
rect 112750 271155 112784 271187
rect 112750 271153 112784 271155
rect 112932 271257 112966 271259
rect 112932 271225 112966 271257
rect 112932 271155 112966 271187
rect 112932 271153 112966 271155
rect 113150 271257 113184 271259
rect 113150 271225 113184 271257
rect 113150 271155 113184 271187
rect 113150 271153 113184 271155
rect 113332 271257 113366 271259
rect 113332 271225 113366 271257
rect 113332 271155 113366 271187
rect 113332 271153 113366 271155
rect 113550 271257 113584 271259
rect 113550 271225 113584 271257
rect 113550 271155 113584 271187
rect 113550 271153 113584 271155
rect 114664 271324 114666 271358
rect 114666 271324 114698 271358
rect 114736 271324 114768 271358
rect 114768 271324 114770 271358
rect 113732 271257 113766 271259
rect 113732 271225 113766 271257
rect 113732 271155 113766 271187
rect 113732 271153 113766 271155
rect 113950 271257 113984 271259
rect 113950 271225 113984 271257
rect 113950 271155 113984 271187
rect 113950 271153 113984 271155
rect 114591 271228 114625 271230
rect 114591 271196 114625 271228
rect 114591 271126 114625 271158
rect 114591 271124 114625 271126
rect 115064 271324 115066 271358
rect 115066 271324 115098 271358
rect 115136 271324 115168 271358
rect 115168 271324 115170 271358
rect 114809 271228 114843 271230
rect 114809 271196 114843 271228
rect 114809 271126 114843 271158
rect 114809 271124 114843 271126
rect 114991 271228 115025 271230
rect 114991 271196 115025 271228
rect 114991 271126 115025 271158
rect 114991 271124 115025 271126
rect 115209 271228 115243 271230
rect 115209 271196 115243 271228
rect 115209 271126 115243 271158
rect 115209 271124 115243 271126
rect 112605 271025 112607 271059
rect 112607 271025 112639 271059
rect 112677 271025 112709 271059
rect 112709 271025 112711 271059
rect 113005 271025 113007 271059
rect 113007 271025 113039 271059
rect 113077 271025 113109 271059
rect 113109 271025 113111 271059
rect 113405 271025 113407 271059
rect 113407 271025 113439 271059
rect 113477 271025 113509 271059
rect 113509 271025 113511 271059
rect 113805 271025 113807 271059
rect 113807 271025 113839 271059
rect 113877 271025 113909 271059
rect 113909 271025 113911 271059
rect 114664 270996 114666 271030
rect 114666 270996 114698 271030
rect 114736 270996 114768 271030
rect 114768 270996 114770 271030
rect 115064 270996 115066 271030
rect 115066 270996 115098 271030
rect 115136 270996 115168 271030
rect 115168 270996 115170 271030
rect 115908 271962 115910 271996
rect 115910 271962 115942 271996
rect 115980 271962 116012 271996
rect 116012 271962 116014 271996
rect 116308 271962 116310 271996
rect 116310 271962 116342 271996
rect 116380 271962 116412 271996
rect 116412 271962 116414 271996
rect 116708 271962 116710 271996
rect 116710 271962 116742 271996
rect 116780 271962 116812 271996
rect 116812 271962 116814 271996
rect 117108 271962 117110 271996
rect 117110 271962 117142 271996
rect 117180 271962 117212 271996
rect 117212 271962 117214 271996
rect 117508 271962 117510 271996
rect 117510 271962 117542 271996
rect 117580 271962 117612 271996
rect 117612 271962 117614 271996
rect 117908 271962 117910 271996
rect 117910 271962 117942 271996
rect 117980 271962 118012 271996
rect 118012 271962 118014 271996
rect 118308 271962 118310 271996
rect 118310 271962 118342 271996
rect 118380 271962 118412 271996
rect 118412 271962 118414 271996
rect 118708 271962 118710 271996
rect 118710 271962 118742 271996
rect 118780 271962 118812 271996
rect 118812 271962 118814 271996
rect 115835 271867 115869 271895
rect 115835 271861 115869 271867
rect 115835 271799 115869 271823
rect 115835 271789 115869 271799
rect 115835 271731 115869 271751
rect 115835 271717 115869 271731
rect 115835 271663 115869 271679
rect 115835 271645 115869 271663
rect 115835 271595 115869 271607
rect 115835 271573 115869 271595
rect 115835 271527 115869 271535
rect 115835 271501 115869 271527
rect 115835 271459 115869 271463
rect 115835 271429 115869 271459
rect 115835 271357 115869 271391
rect 115835 271289 115869 271319
rect 115835 271285 115869 271289
rect 115835 271221 115869 271247
rect 115835 271213 115869 271221
rect 115835 271153 115869 271175
rect 115835 271141 115869 271153
rect 115835 271085 115869 271103
rect 115835 271069 115869 271085
rect 115835 271017 115869 271031
rect 115835 270997 115869 271017
rect 115835 270949 115869 270959
rect 115835 270925 115869 270949
rect 115835 270881 115869 270887
rect 115835 270853 115869 270881
rect 116053 271867 116087 271895
rect 116053 271861 116087 271867
rect 116053 271799 116087 271823
rect 116053 271789 116087 271799
rect 116053 271731 116087 271751
rect 116053 271717 116087 271731
rect 116053 271663 116087 271679
rect 116053 271645 116087 271663
rect 116053 271595 116087 271607
rect 116053 271573 116087 271595
rect 116053 271527 116087 271535
rect 116053 271501 116087 271527
rect 116053 271459 116087 271463
rect 116053 271429 116087 271459
rect 116053 271357 116087 271391
rect 116053 271289 116087 271319
rect 116053 271285 116087 271289
rect 116053 271221 116087 271247
rect 116053 271213 116087 271221
rect 116053 271153 116087 271175
rect 116053 271141 116087 271153
rect 116053 271085 116087 271103
rect 116053 271069 116087 271085
rect 116053 271017 116087 271031
rect 116053 270997 116087 271017
rect 116053 270949 116087 270959
rect 116053 270925 116087 270949
rect 116053 270881 116087 270887
rect 116053 270853 116087 270881
rect 116235 271867 116269 271895
rect 116235 271861 116269 271867
rect 116235 271799 116269 271823
rect 116235 271789 116269 271799
rect 116235 271731 116269 271751
rect 116235 271717 116269 271731
rect 116235 271663 116269 271679
rect 116235 271645 116269 271663
rect 116235 271595 116269 271607
rect 116235 271573 116269 271595
rect 116235 271527 116269 271535
rect 116235 271501 116269 271527
rect 116235 271459 116269 271463
rect 116235 271429 116269 271459
rect 116235 271357 116269 271391
rect 116235 271289 116269 271319
rect 116235 271285 116269 271289
rect 116235 271221 116269 271247
rect 116235 271213 116269 271221
rect 116235 271153 116269 271175
rect 116235 271141 116269 271153
rect 116235 271085 116269 271103
rect 116235 271069 116269 271085
rect 116235 271017 116269 271031
rect 116235 270997 116269 271017
rect 116235 270949 116269 270959
rect 116235 270925 116269 270949
rect 116235 270881 116269 270887
rect 116235 270853 116269 270881
rect 116453 271867 116487 271895
rect 116453 271861 116487 271867
rect 116453 271799 116487 271823
rect 116453 271789 116487 271799
rect 116453 271731 116487 271751
rect 116453 271717 116487 271731
rect 116453 271663 116487 271679
rect 116453 271645 116487 271663
rect 116453 271595 116487 271607
rect 116453 271573 116487 271595
rect 116453 271527 116487 271535
rect 116453 271501 116487 271527
rect 116453 271459 116487 271463
rect 116453 271429 116487 271459
rect 116453 271357 116487 271391
rect 116453 271289 116487 271319
rect 116453 271285 116487 271289
rect 116453 271221 116487 271247
rect 116453 271213 116487 271221
rect 116453 271153 116487 271175
rect 116453 271141 116487 271153
rect 116453 271085 116487 271103
rect 116453 271069 116487 271085
rect 116453 271017 116487 271031
rect 116453 270997 116487 271017
rect 116453 270949 116487 270959
rect 116453 270925 116487 270949
rect 116453 270881 116487 270887
rect 116453 270853 116487 270881
rect 116635 271867 116669 271895
rect 116635 271861 116669 271867
rect 116635 271799 116669 271823
rect 116635 271789 116669 271799
rect 116635 271731 116669 271751
rect 116635 271717 116669 271731
rect 116635 271663 116669 271679
rect 116635 271645 116669 271663
rect 116635 271595 116669 271607
rect 116635 271573 116669 271595
rect 116635 271527 116669 271535
rect 116635 271501 116669 271527
rect 116635 271459 116669 271463
rect 116635 271429 116669 271459
rect 116635 271357 116669 271391
rect 116635 271289 116669 271319
rect 116635 271285 116669 271289
rect 116635 271221 116669 271247
rect 116635 271213 116669 271221
rect 116635 271153 116669 271175
rect 116635 271141 116669 271153
rect 116635 271085 116669 271103
rect 116635 271069 116669 271085
rect 116635 271017 116669 271031
rect 116635 270997 116669 271017
rect 116635 270949 116669 270959
rect 116635 270925 116669 270949
rect 116635 270881 116669 270887
rect 116635 270853 116669 270881
rect 116853 271867 116887 271895
rect 116853 271861 116887 271867
rect 116853 271799 116887 271823
rect 116853 271789 116887 271799
rect 116853 271731 116887 271751
rect 116853 271717 116887 271731
rect 116853 271663 116887 271679
rect 116853 271645 116887 271663
rect 116853 271595 116887 271607
rect 116853 271573 116887 271595
rect 116853 271527 116887 271535
rect 116853 271501 116887 271527
rect 116853 271459 116887 271463
rect 116853 271429 116887 271459
rect 116853 271357 116887 271391
rect 116853 271289 116887 271319
rect 116853 271285 116887 271289
rect 116853 271221 116887 271247
rect 116853 271213 116887 271221
rect 116853 271153 116887 271175
rect 116853 271141 116887 271153
rect 116853 271085 116887 271103
rect 116853 271069 116887 271085
rect 116853 271017 116887 271031
rect 116853 270997 116887 271017
rect 116853 270949 116887 270959
rect 116853 270925 116887 270949
rect 116853 270881 116887 270887
rect 116853 270853 116887 270881
rect 117035 271867 117069 271895
rect 117035 271861 117069 271867
rect 117035 271799 117069 271823
rect 117035 271789 117069 271799
rect 117035 271731 117069 271751
rect 117035 271717 117069 271731
rect 117035 271663 117069 271679
rect 117035 271645 117069 271663
rect 117035 271595 117069 271607
rect 117035 271573 117069 271595
rect 117035 271527 117069 271535
rect 117035 271501 117069 271527
rect 117035 271459 117069 271463
rect 117035 271429 117069 271459
rect 117035 271357 117069 271391
rect 117035 271289 117069 271319
rect 117035 271285 117069 271289
rect 117035 271221 117069 271247
rect 117035 271213 117069 271221
rect 117035 271153 117069 271175
rect 117035 271141 117069 271153
rect 117035 271085 117069 271103
rect 117035 271069 117069 271085
rect 117035 271017 117069 271031
rect 117035 270997 117069 271017
rect 117035 270949 117069 270959
rect 117035 270925 117069 270949
rect 117035 270881 117069 270887
rect 117035 270853 117069 270881
rect 117253 271867 117287 271895
rect 117253 271861 117287 271867
rect 117253 271799 117287 271823
rect 117253 271789 117287 271799
rect 117253 271731 117287 271751
rect 117253 271717 117287 271731
rect 117253 271663 117287 271679
rect 117253 271645 117287 271663
rect 117253 271595 117287 271607
rect 117253 271573 117287 271595
rect 117253 271527 117287 271535
rect 117253 271501 117287 271527
rect 117253 271459 117287 271463
rect 117253 271429 117287 271459
rect 117253 271357 117287 271391
rect 117253 271289 117287 271319
rect 117253 271285 117287 271289
rect 117253 271221 117287 271247
rect 117253 271213 117287 271221
rect 117253 271153 117287 271175
rect 117253 271141 117287 271153
rect 117253 271085 117287 271103
rect 117253 271069 117287 271085
rect 117253 271017 117287 271031
rect 117253 270997 117287 271017
rect 117253 270949 117287 270959
rect 117253 270925 117287 270949
rect 117253 270881 117287 270887
rect 117253 270853 117287 270881
rect 117435 271867 117469 271895
rect 117435 271861 117469 271867
rect 117435 271799 117469 271823
rect 117435 271789 117469 271799
rect 117435 271731 117469 271751
rect 117435 271717 117469 271731
rect 117435 271663 117469 271679
rect 117435 271645 117469 271663
rect 117435 271595 117469 271607
rect 117435 271573 117469 271595
rect 117435 271527 117469 271535
rect 117435 271501 117469 271527
rect 117435 271459 117469 271463
rect 117435 271429 117469 271459
rect 117435 271357 117469 271391
rect 117435 271289 117469 271319
rect 117435 271285 117469 271289
rect 117435 271221 117469 271247
rect 117435 271213 117469 271221
rect 117435 271153 117469 271175
rect 117435 271141 117469 271153
rect 117435 271085 117469 271103
rect 117435 271069 117469 271085
rect 117435 271017 117469 271031
rect 117435 270997 117469 271017
rect 117435 270949 117469 270959
rect 117435 270925 117469 270949
rect 117435 270881 117469 270887
rect 117435 270853 117469 270881
rect 117653 271867 117687 271895
rect 117653 271861 117687 271867
rect 117653 271799 117687 271823
rect 117653 271789 117687 271799
rect 117653 271731 117687 271751
rect 117653 271717 117687 271731
rect 117653 271663 117687 271679
rect 117653 271645 117687 271663
rect 117653 271595 117687 271607
rect 117653 271573 117687 271595
rect 117653 271527 117687 271535
rect 117653 271501 117687 271527
rect 117653 271459 117687 271463
rect 117653 271429 117687 271459
rect 117653 271357 117687 271391
rect 117653 271289 117687 271319
rect 117653 271285 117687 271289
rect 117653 271221 117687 271247
rect 117653 271213 117687 271221
rect 117653 271153 117687 271175
rect 117653 271141 117687 271153
rect 117653 271085 117687 271103
rect 117653 271069 117687 271085
rect 117653 271017 117687 271031
rect 117653 270997 117687 271017
rect 117653 270949 117687 270959
rect 117653 270925 117687 270949
rect 117653 270881 117687 270887
rect 117653 270853 117687 270881
rect 117835 271867 117869 271895
rect 117835 271861 117869 271867
rect 117835 271799 117869 271823
rect 117835 271789 117869 271799
rect 117835 271731 117869 271751
rect 117835 271717 117869 271731
rect 117835 271663 117869 271679
rect 117835 271645 117869 271663
rect 117835 271595 117869 271607
rect 117835 271573 117869 271595
rect 117835 271527 117869 271535
rect 117835 271501 117869 271527
rect 117835 271459 117869 271463
rect 117835 271429 117869 271459
rect 117835 271357 117869 271391
rect 117835 271289 117869 271319
rect 117835 271285 117869 271289
rect 117835 271221 117869 271247
rect 117835 271213 117869 271221
rect 117835 271153 117869 271175
rect 117835 271141 117869 271153
rect 117835 271085 117869 271103
rect 117835 271069 117869 271085
rect 117835 271017 117869 271031
rect 117835 270997 117869 271017
rect 117835 270949 117869 270959
rect 117835 270925 117869 270949
rect 117835 270881 117869 270887
rect 117835 270853 117869 270881
rect 118053 271867 118087 271895
rect 118053 271861 118087 271867
rect 118053 271799 118087 271823
rect 118053 271789 118087 271799
rect 118053 271731 118087 271751
rect 118053 271717 118087 271731
rect 118053 271663 118087 271679
rect 118053 271645 118087 271663
rect 118053 271595 118087 271607
rect 118053 271573 118087 271595
rect 118053 271527 118087 271535
rect 118053 271501 118087 271527
rect 118053 271459 118087 271463
rect 118053 271429 118087 271459
rect 118053 271357 118087 271391
rect 118053 271289 118087 271319
rect 118053 271285 118087 271289
rect 118053 271221 118087 271247
rect 118053 271213 118087 271221
rect 118053 271153 118087 271175
rect 118053 271141 118087 271153
rect 118053 271085 118087 271103
rect 118053 271069 118087 271085
rect 118053 271017 118087 271031
rect 118053 270997 118087 271017
rect 118053 270949 118087 270959
rect 118053 270925 118087 270949
rect 118053 270881 118087 270887
rect 118053 270853 118087 270881
rect 118235 271867 118269 271895
rect 118235 271861 118269 271867
rect 118235 271799 118269 271823
rect 118235 271789 118269 271799
rect 118235 271731 118269 271751
rect 118235 271717 118269 271731
rect 118235 271663 118269 271679
rect 118235 271645 118269 271663
rect 118235 271595 118269 271607
rect 118235 271573 118269 271595
rect 118235 271527 118269 271535
rect 118235 271501 118269 271527
rect 118235 271459 118269 271463
rect 118235 271429 118269 271459
rect 118235 271357 118269 271391
rect 118235 271289 118269 271319
rect 118235 271285 118269 271289
rect 118235 271221 118269 271247
rect 118235 271213 118269 271221
rect 118235 271153 118269 271175
rect 118235 271141 118269 271153
rect 118235 271085 118269 271103
rect 118235 271069 118269 271085
rect 118235 271017 118269 271031
rect 118235 270997 118269 271017
rect 118235 270949 118269 270959
rect 118235 270925 118269 270949
rect 118235 270881 118269 270887
rect 118235 270853 118269 270881
rect 118453 271867 118487 271895
rect 118453 271861 118487 271867
rect 118453 271799 118487 271823
rect 118453 271789 118487 271799
rect 118453 271731 118487 271751
rect 118453 271717 118487 271731
rect 118453 271663 118487 271679
rect 118453 271645 118487 271663
rect 118453 271595 118487 271607
rect 118453 271573 118487 271595
rect 118453 271527 118487 271535
rect 118453 271501 118487 271527
rect 118453 271459 118487 271463
rect 118453 271429 118487 271459
rect 118453 271357 118487 271391
rect 118453 271289 118487 271319
rect 118453 271285 118487 271289
rect 118453 271221 118487 271247
rect 118453 271213 118487 271221
rect 118453 271153 118487 271175
rect 118453 271141 118487 271153
rect 118453 271085 118487 271103
rect 118453 271069 118487 271085
rect 118453 271017 118487 271031
rect 118453 270997 118487 271017
rect 118453 270949 118487 270959
rect 118453 270925 118487 270949
rect 118453 270881 118487 270887
rect 118453 270853 118487 270881
rect 118635 271867 118669 271895
rect 118635 271861 118669 271867
rect 118635 271799 118669 271823
rect 118635 271789 118669 271799
rect 118635 271731 118669 271751
rect 118635 271717 118669 271731
rect 118635 271663 118669 271679
rect 118635 271645 118669 271663
rect 118635 271595 118669 271607
rect 118635 271573 118669 271595
rect 118635 271527 118669 271535
rect 118635 271501 118669 271527
rect 118635 271459 118669 271463
rect 118635 271429 118669 271459
rect 118635 271357 118669 271391
rect 118635 271289 118669 271319
rect 118635 271285 118669 271289
rect 118635 271221 118669 271247
rect 118635 271213 118669 271221
rect 118635 271153 118669 271175
rect 118635 271141 118669 271153
rect 118635 271085 118669 271103
rect 118635 271069 118669 271085
rect 118635 271017 118669 271031
rect 118635 270997 118669 271017
rect 118635 270949 118669 270959
rect 118635 270925 118669 270949
rect 118635 270881 118669 270887
rect 118635 270853 118669 270881
rect 118853 271867 118887 271895
rect 118853 271861 118887 271867
rect 118853 271799 118887 271823
rect 118853 271789 118887 271799
rect 118853 271731 118887 271751
rect 118853 271717 118887 271731
rect 118853 271663 118887 271679
rect 118853 271645 118887 271663
rect 118853 271595 118887 271607
rect 118853 271573 118887 271595
rect 118853 271527 118887 271535
rect 118853 271501 118887 271527
rect 118853 271459 118887 271463
rect 118853 271429 118887 271459
rect 118853 271357 118887 271391
rect 118853 271289 118887 271319
rect 118853 271285 118887 271289
rect 118853 271221 118887 271247
rect 118853 271213 118887 271221
rect 118853 271153 118887 271175
rect 118853 271141 118887 271153
rect 118853 271085 118887 271103
rect 118853 271069 118887 271085
rect 118853 271017 118887 271031
rect 118853 270997 118887 271017
rect 118853 270949 118887 270959
rect 118853 270925 118887 270949
rect 118853 270881 118887 270887
rect 118853 270853 118887 270881
rect 115908 270752 115910 270786
rect 115910 270752 115942 270786
rect 115980 270752 116012 270786
rect 116012 270752 116014 270786
rect 116308 270752 116310 270786
rect 116310 270752 116342 270786
rect 116380 270752 116412 270786
rect 116412 270752 116414 270786
rect 116708 270752 116710 270786
rect 116710 270752 116742 270786
rect 116780 270752 116812 270786
rect 116812 270752 116814 270786
rect 117108 270752 117110 270786
rect 117110 270752 117142 270786
rect 117180 270752 117212 270786
rect 117212 270752 117214 270786
rect 117508 270752 117510 270786
rect 117510 270752 117542 270786
rect 117580 270752 117612 270786
rect 117612 270752 117614 270786
rect 117908 270752 117910 270786
rect 117910 270752 117942 270786
rect 117980 270752 118012 270786
rect 118012 270752 118014 270786
rect 118308 270752 118310 270786
rect 118310 270752 118342 270786
rect 118380 270752 118412 270786
rect 118412 270752 118414 270786
rect 118708 270752 118710 270786
rect 118710 270752 118742 270786
rect 118780 270752 118812 270786
rect 118812 270752 118814 270786
rect 114096 270607 114130 270641
rect 114168 270607 114202 270641
rect 114240 270607 114274 270641
rect 114312 270607 114346 270641
rect 114384 270607 114418 270641
rect 114456 270607 114490 270641
rect 112587 270262 112589 270296
rect 112589 270262 112621 270296
rect 112659 270262 112691 270296
rect 112691 270262 112693 270296
rect 112987 270262 112989 270296
rect 112989 270262 113021 270296
rect 113059 270262 113091 270296
rect 113091 270262 113093 270296
rect 113387 270262 113389 270296
rect 113389 270262 113421 270296
rect 113459 270262 113491 270296
rect 113491 270262 113493 270296
rect 113787 270262 113789 270296
rect 113789 270262 113821 270296
rect 113859 270262 113891 270296
rect 113891 270262 113893 270296
rect 114187 270262 114189 270296
rect 114189 270262 114221 270296
rect 114259 270262 114291 270296
rect 114291 270262 114293 270296
rect 114587 270262 114589 270296
rect 114589 270262 114621 270296
rect 114659 270262 114691 270296
rect 114691 270262 114693 270296
rect 114987 270262 114989 270296
rect 114989 270262 115021 270296
rect 115059 270262 115091 270296
rect 115091 270262 115093 270296
rect 115387 270262 115389 270296
rect 115389 270262 115421 270296
rect 115459 270262 115491 270296
rect 115491 270262 115493 270296
rect 115787 270262 115789 270296
rect 115789 270262 115821 270296
rect 115859 270262 115891 270296
rect 115891 270262 115893 270296
rect 116187 270262 116189 270296
rect 116189 270262 116221 270296
rect 116259 270262 116291 270296
rect 116291 270262 116293 270296
rect 116587 270262 116589 270296
rect 116589 270262 116621 270296
rect 116659 270262 116691 270296
rect 116691 270262 116693 270296
rect 116987 270262 116989 270296
rect 116989 270262 117021 270296
rect 117059 270262 117091 270296
rect 117091 270262 117093 270296
rect 117387 270262 117389 270296
rect 117389 270262 117421 270296
rect 117459 270262 117491 270296
rect 117491 270262 117493 270296
rect 117787 270262 117789 270296
rect 117789 270262 117821 270296
rect 117859 270262 117891 270296
rect 117891 270262 117893 270296
rect 118187 270262 118189 270296
rect 118189 270262 118221 270296
rect 118259 270262 118291 270296
rect 118291 270262 118293 270296
rect 118587 270262 118589 270296
rect 118589 270262 118621 270296
rect 118659 270262 118691 270296
rect 118691 270262 118693 270296
rect 112514 270167 112548 270195
rect 112514 270161 112548 270167
rect 112514 270099 112548 270123
rect 112514 270089 112548 270099
rect 112514 270031 112548 270051
rect 112514 270017 112548 270031
rect 112514 269963 112548 269979
rect 112514 269945 112548 269963
rect 112514 269895 112548 269907
rect 112514 269873 112548 269895
rect 112514 269827 112548 269835
rect 112514 269801 112548 269827
rect 112514 269759 112548 269763
rect 112514 269729 112548 269759
rect 112514 269657 112548 269691
rect 112514 269589 112548 269619
rect 112514 269585 112548 269589
rect 112514 269521 112548 269547
rect 112514 269513 112548 269521
rect 112514 269453 112548 269475
rect 112514 269441 112548 269453
rect 112514 269385 112548 269403
rect 112514 269369 112548 269385
rect 112514 269317 112548 269331
rect 112514 269297 112548 269317
rect 112514 269249 112548 269259
rect 112514 269225 112548 269249
rect 112514 269181 112548 269187
rect 112514 269153 112548 269181
rect 112732 270167 112766 270195
rect 112732 270161 112766 270167
rect 112732 270099 112766 270123
rect 112732 270089 112766 270099
rect 112732 270031 112766 270051
rect 112732 270017 112766 270031
rect 112732 269963 112766 269979
rect 112732 269945 112766 269963
rect 112732 269895 112766 269907
rect 112732 269873 112766 269895
rect 112732 269827 112766 269835
rect 112732 269801 112766 269827
rect 112732 269759 112766 269763
rect 112732 269729 112766 269759
rect 112732 269657 112766 269691
rect 112732 269589 112766 269619
rect 112732 269585 112766 269589
rect 112732 269521 112766 269547
rect 112732 269513 112766 269521
rect 112732 269453 112766 269475
rect 112732 269441 112766 269453
rect 112732 269385 112766 269403
rect 112732 269369 112766 269385
rect 112732 269317 112766 269331
rect 112732 269297 112766 269317
rect 112732 269249 112766 269259
rect 112732 269225 112766 269249
rect 112732 269181 112766 269187
rect 112732 269153 112766 269181
rect 112914 270167 112948 270195
rect 112914 270161 112948 270167
rect 112914 270099 112948 270123
rect 112914 270089 112948 270099
rect 112914 270031 112948 270051
rect 112914 270017 112948 270031
rect 112914 269963 112948 269979
rect 112914 269945 112948 269963
rect 112914 269895 112948 269907
rect 112914 269873 112948 269895
rect 112914 269827 112948 269835
rect 112914 269801 112948 269827
rect 112914 269759 112948 269763
rect 112914 269729 112948 269759
rect 112914 269657 112948 269691
rect 112914 269589 112948 269619
rect 112914 269585 112948 269589
rect 112914 269521 112948 269547
rect 112914 269513 112948 269521
rect 112914 269453 112948 269475
rect 112914 269441 112948 269453
rect 112914 269385 112948 269403
rect 112914 269369 112948 269385
rect 112914 269317 112948 269331
rect 112914 269297 112948 269317
rect 112914 269249 112948 269259
rect 112914 269225 112948 269249
rect 112914 269181 112948 269187
rect 112914 269153 112948 269181
rect 113132 270167 113166 270195
rect 113132 270161 113166 270167
rect 113132 270099 113166 270123
rect 113132 270089 113166 270099
rect 113132 270031 113166 270051
rect 113132 270017 113166 270031
rect 113132 269963 113166 269979
rect 113132 269945 113166 269963
rect 113132 269895 113166 269907
rect 113132 269873 113166 269895
rect 113132 269827 113166 269835
rect 113132 269801 113166 269827
rect 113132 269759 113166 269763
rect 113132 269729 113166 269759
rect 113132 269657 113166 269691
rect 113132 269589 113166 269619
rect 113132 269585 113166 269589
rect 113132 269521 113166 269547
rect 113132 269513 113166 269521
rect 113132 269453 113166 269475
rect 113132 269441 113166 269453
rect 113132 269385 113166 269403
rect 113132 269369 113166 269385
rect 113132 269317 113166 269331
rect 113132 269297 113166 269317
rect 113132 269249 113166 269259
rect 113132 269225 113166 269249
rect 113132 269181 113166 269187
rect 113132 269153 113166 269181
rect 113314 270167 113348 270195
rect 113314 270161 113348 270167
rect 113314 270099 113348 270123
rect 113314 270089 113348 270099
rect 113314 270031 113348 270051
rect 113314 270017 113348 270031
rect 113314 269963 113348 269979
rect 113314 269945 113348 269963
rect 113314 269895 113348 269907
rect 113314 269873 113348 269895
rect 113314 269827 113348 269835
rect 113314 269801 113348 269827
rect 113314 269759 113348 269763
rect 113314 269729 113348 269759
rect 113314 269657 113348 269691
rect 113314 269589 113348 269619
rect 113314 269585 113348 269589
rect 113314 269521 113348 269547
rect 113314 269513 113348 269521
rect 113314 269453 113348 269475
rect 113314 269441 113348 269453
rect 113314 269385 113348 269403
rect 113314 269369 113348 269385
rect 113314 269317 113348 269331
rect 113314 269297 113348 269317
rect 113314 269249 113348 269259
rect 113314 269225 113348 269249
rect 113314 269181 113348 269187
rect 113314 269153 113348 269181
rect 113532 270167 113566 270195
rect 113532 270161 113566 270167
rect 113532 270099 113566 270123
rect 113532 270089 113566 270099
rect 113532 270031 113566 270051
rect 113532 270017 113566 270031
rect 113532 269963 113566 269979
rect 113532 269945 113566 269963
rect 113532 269895 113566 269907
rect 113532 269873 113566 269895
rect 113532 269827 113566 269835
rect 113532 269801 113566 269827
rect 113532 269759 113566 269763
rect 113532 269729 113566 269759
rect 113532 269657 113566 269691
rect 113532 269589 113566 269619
rect 113532 269585 113566 269589
rect 113532 269521 113566 269547
rect 113532 269513 113566 269521
rect 113532 269453 113566 269475
rect 113532 269441 113566 269453
rect 113532 269385 113566 269403
rect 113532 269369 113566 269385
rect 113532 269317 113566 269331
rect 113532 269297 113566 269317
rect 113532 269249 113566 269259
rect 113532 269225 113566 269249
rect 113532 269181 113566 269187
rect 113532 269153 113566 269181
rect 113714 270167 113748 270195
rect 113714 270161 113748 270167
rect 113714 270099 113748 270123
rect 113714 270089 113748 270099
rect 113714 270031 113748 270051
rect 113714 270017 113748 270031
rect 113714 269963 113748 269979
rect 113714 269945 113748 269963
rect 113714 269895 113748 269907
rect 113714 269873 113748 269895
rect 113714 269827 113748 269835
rect 113714 269801 113748 269827
rect 113714 269759 113748 269763
rect 113714 269729 113748 269759
rect 113714 269657 113748 269691
rect 113714 269589 113748 269619
rect 113714 269585 113748 269589
rect 113714 269521 113748 269547
rect 113714 269513 113748 269521
rect 113714 269453 113748 269475
rect 113714 269441 113748 269453
rect 113714 269385 113748 269403
rect 113714 269369 113748 269385
rect 113714 269317 113748 269331
rect 113714 269297 113748 269317
rect 113714 269249 113748 269259
rect 113714 269225 113748 269249
rect 113714 269181 113748 269187
rect 113714 269153 113748 269181
rect 113932 270167 113966 270195
rect 113932 270161 113966 270167
rect 113932 270099 113966 270123
rect 113932 270089 113966 270099
rect 113932 270031 113966 270051
rect 113932 270017 113966 270031
rect 113932 269963 113966 269979
rect 113932 269945 113966 269963
rect 113932 269895 113966 269907
rect 113932 269873 113966 269895
rect 113932 269827 113966 269835
rect 113932 269801 113966 269827
rect 113932 269759 113966 269763
rect 113932 269729 113966 269759
rect 113932 269657 113966 269691
rect 113932 269589 113966 269619
rect 113932 269585 113966 269589
rect 113932 269521 113966 269547
rect 113932 269513 113966 269521
rect 113932 269453 113966 269475
rect 113932 269441 113966 269453
rect 113932 269385 113966 269403
rect 113932 269369 113966 269385
rect 113932 269317 113966 269331
rect 113932 269297 113966 269317
rect 113932 269249 113966 269259
rect 113932 269225 113966 269249
rect 113932 269181 113966 269187
rect 113932 269153 113966 269181
rect 114114 270167 114148 270195
rect 114114 270161 114148 270167
rect 114114 270099 114148 270123
rect 114114 270089 114148 270099
rect 114114 270031 114148 270051
rect 114114 270017 114148 270031
rect 114114 269963 114148 269979
rect 114114 269945 114148 269963
rect 114114 269895 114148 269907
rect 114114 269873 114148 269895
rect 114114 269827 114148 269835
rect 114114 269801 114148 269827
rect 114114 269759 114148 269763
rect 114114 269729 114148 269759
rect 114114 269657 114148 269691
rect 114114 269589 114148 269619
rect 114114 269585 114148 269589
rect 114114 269521 114148 269547
rect 114114 269513 114148 269521
rect 114114 269453 114148 269475
rect 114114 269441 114148 269453
rect 114114 269385 114148 269403
rect 114114 269369 114148 269385
rect 114114 269317 114148 269331
rect 114114 269297 114148 269317
rect 114114 269249 114148 269259
rect 114114 269225 114148 269249
rect 114114 269181 114148 269187
rect 114114 269153 114148 269181
rect 114332 270167 114366 270195
rect 114332 270161 114366 270167
rect 114332 270099 114366 270123
rect 114332 270089 114366 270099
rect 114332 270031 114366 270051
rect 114332 270017 114366 270031
rect 114332 269963 114366 269979
rect 114332 269945 114366 269963
rect 114332 269895 114366 269907
rect 114332 269873 114366 269895
rect 114332 269827 114366 269835
rect 114332 269801 114366 269827
rect 114332 269759 114366 269763
rect 114332 269729 114366 269759
rect 114332 269657 114366 269691
rect 114332 269589 114366 269619
rect 114332 269585 114366 269589
rect 114332 269521 114366 269547
rect 114332 269513 114366 269521
rect 114332 269453 114366 269475
rect 114332 269441 114366 269453
rect 114332 269385 114366 269403
rect 114332 269369 114366 269385
rect 114332 269317 114366 269331
rect 114332 269297 114366 269317
rect 114332 269249 114366 269259
rect 114332 269225 114366 269249
rect 114332 269181 114366 269187
rect 114332 269153 114366 269181
rect 114514 270167 114548 270195
rect 114514 270161 114548 270167
rect 114514 270099 114548 270123
rect 114514 270089 114548 270099
rect 114514 270031 114548 270051
rect 114514 270017 114548 270031
rect 114514 269963 114548 269979
rect 114514 269945 114548 269963
rect 114514 269895 114548 269907
rect 114514 269873 114548 269895
rect 114514 269827 114548 269835
rect 114514 269801 114548 269827
rect 114514 269759 114548 269763
rect 114514 269729 114548 269759
rect 114514 269657 114548 269691
rect 114514 269589 114548 269619
rect 114514 269585 114548 269589
rect 114514 269521 114548 269547
rect 114514 269513 114548 269521
rect 114514 269453 114548 269475
rect 114514 269441 114548 269453
rect 114514 269385 114548 269403
rect 114514 269369 114548 269385
rect 114514 269317 114548 269331
rect 114514 269297 114548 269317
rect 114514 269249 114548 269259
rect 114514 269225 114548 269249
rect 114514 269181 114548 269187
rect 114514 269153 114548 269181
rect 114732 270167 114766 270195
rect 114732 270161 114766 270167
rect 114732 270099 114766 270123
rect 114732 270089 114766 270099
rect 114732 270031 114766 270051
rect 114732 270017 114766 270031
rect 114732 269963 114766 269979
rect 114732 269945 114766 269963
rect 114732 269895 114766 269907
rect 114732 269873 114766 269895
rect 114732 269827 114766 269835
rect 114732 269801 114766 269827
rect 114732 269759 114766 269763
rect 114732 269729 114766 269759
rect 114732 269657 114766 269691
rect 114732 269589 114766 269619
rect 114732 269585 114766 269589
rect 114732 269521 114766 269547
rect 114732 269513 114766 269521
rect 114732 269453 114766 269475
rect 114732 269441 114766 269453
rect 114732 269385 114766 269403
rect 114732 269369 114766 269385
rect 114732 269317 114766 269331
rect 114732 269297 114766 269317
rect 114732 269249 114766 269259
rect 114732 269225 114766 269249
rect 114732 269181 114766 269187
rect 114732 269153 114766 269181
rect 114914 270167 114948 270195
rect 114914 270161 114948 270167
rect 114914 270099 114948 270123
rect 114914 270089 114948 270099
rect 114914 270031 114948 270051
rect 114914 270017 114948 270031
rect 114914 269963 114948 269979
rect 114914 269945 114948 269963
rect 114914 269895 114948 269907
rect 114914 269873 114948 269895
rect 114914 269827 114948 269835
rect 114914 269801 114948 269827
rect 114914 269759 114948 269763
rect 114914 269729 114948 269759
rect 114914 269657 114948 269691
rect 114914 269589 114948 269619
rect 114914 269585 114948 269589
rect 114914 269521 114948 269547
rect 114914 269513 114948 269521
rect 114914 269453 114948 269475
rect 114914 269441 114948 269453
rect 114914 269385 114948 269403
rect 114914 269369 114948 269385
rect 114914 269317 114948 269331
rect 114914 269297 114948 269317
rect 114914 269249 114948 269259
rect 114914 269225 114948 269249
rect 114914 269181 114948 269187
rect 114914 269153 114948 269181
rect 115132 270167 115166 270195
rect 115132 270161 115166 270167
rect 115132 270099 115166 270123
rect 115132 270089 115166 270099
rect 115132 270031 115166 270051
rect 115132 270017 115166 270031
rect 115132 269963 115166 269979
rect 115132 269945 115166 269963
rect 115132 269895 115166 269907
rect 115132 269873 115166 269895
rect 115132 269827 115166 269835
rect 115132 269801 115166 269827
rect 115132 269759 115166 269763
rect 115132 269729 115166 269759
rect 115132 269657 115166 269691
rect 115132 269589 115166 269619
rect 115132 269585 115166 269589
rect 115132 269521 115166 269547
rect 115132 269513 115166 269521
rect 115132 269453 115166 269475
rect 115132 269441 115166 269453
rect 115132 269385 115166 269403
rect 115132 269369 115166 269385
rect 115132 269317 115166 269331
rect 115132 269297 115166 269317
rect 115132 269249 115166 269259
rect 115132 269225 115166 269249
rect 115132 269181 115166 269187
rect 115132 269153 115166 269181
rect 115314 270167 115348 270195
rect 115314 270161 115348 270167
rect 115314 270099 115348 270123
rect 115314 270089 115348 270099
rect 115314 270031 115348 270051
rect 115314 270017 115348 270031
rect 115314 269963 115348 269979
rect 115314 269945 115348 269963
rect 115314 269895 115348 269907
rect 115314 269873 115348 269895
rect 115314 269827 115348 269835
rect 115314 269801 115348 269827
rect 115314 269759 115348 269763
rect 115314 269729 115348 269759
rect 115314 269657 115348 269691
rect 115314 269589 115348 269619
rect 115314 269585 115348 269589
rect 115314 269521 115348 269547
rect 115314 269513 115348 269521
rect 115314 269453 115348 269475
rect 115314 269441 115348 269453
rect 115314 269385 115348 269403
rect 115314 269369 115348 269385
rect 115314 269317 115348 269331
rect 115314 269297 115348 269317
rect 115314 269249 115348 269259
rect 115314 269225 115348 269249
rect 115314 269181 115348 269187
rect 115314 269153 115348 269181
rect 115532 270167 115566 270195
rect 115532 270161 115566 270167
rect 115532 270099 115566 270123
rect 115532 270089 115566 270099
rect 115532 270031 115566 270051
rect 115532 270017 115566 270031
rect 115532 269963 115566 269979
rect 115532 269945 115566 269963
rect 115532 269895 115566 269907
rect 115532 269873 115566 269895
rect 115532 269827 115566 269835
rect 115532 269801 115566 269827
rect 115532 269759 115566 269763
rect 115532 269729 115566 269759
rect 115532 269657 115566 269691
rect 115532 269589 115566 269619
rect 115532 269585 115566 269589
rect 115532 269521 115566 269547
rect 115532 269513 115566 269521
rect 115532 269453 115566 269475
rect 115532 269441 115566 269453
rect 115532 269385 115566 269403
rect 115532 269369 115566 269385
rect 115532 269317 115566 269331
rect 115532 269297 115566 269317
rect 115532 269249 115566 269259
rect 115532 269225 115566 269249
rect 115532 269181 115566 269187
rect 115532 269153 115566 269181
rect 115714 270167 115748 270195
rect 115714 270161 115748 270167
rect 115714 270099 115748 270123
rect 115714 270089 115748 270099
rect 115714 270031 115748 270051
rect 115714 270017 115748 270031
rect 115714 269963 115748 269979
rect 115714 269945 115748 269963
rect 115714 269895 115748 269907
rect 115714 269873 115748 269895
rect 115714 269827 115748 269835
rect 115714 269801 115748 269827
rect 115714 269759 115748 269763
rect 115714 269729 115748 269759
rect 115714 269657 115748 269691
rect 115714 269589 115748 269619
rect 115714 269585 115748 269589
rect 115714 269521 115748 269547
rect 115714 269513 115748 269521
rect 115714 269453 115748 269475
rect 115714 269441 115748 269453
rect 115714 269385 115748 269403
rect 115714 269369 115748 269385
rect 115714 269317 115748 269331
rect 115714 269297 115748 269317
rect 115714 269249 115748 269259
rect 115714 269225 115748 269249
rect 115714 269181 115748 269187
rect 115714 269153 115748 269181
rect 115932 270167 115966 270195
rect 115932 270161 115966 270167
rect 115932 270099 115966 270123
rect 115932 270089 115966 270099
rect 115932 270031 115966 270051
rect 115932 270017 115966 270031
rect 115932 269963 115966 269979
rect 115932 269945 115966 269963
rect 115932 269895 115966 269907
rect 115932 269873 115966 269895
rect 115932 269827 115966 269835
rect 115932 269801 115966 269827
rect 115932 269759 115966 269763
rect 115932 269729 115966 269759
rect 115932 269657 115966 269691
rect 115932 269589 115966 269619
rect 115932 269585 115966 269589
rect 115932 269521 115966 269547
rect 115932 269513 115966 269521
rect 115932 269453 115966 269475
rect 115932 269441 115966 269453
rect 115932 269385 115966 269403
rect 115932 269369 115966 269385
rect 115932 269317 115966 269331
rect 115932 269297 115966 269317
rect 115932 269249 115966 269259
rect 115932 269225 115966 269249
rect 115932 269181 115966 269187
rect 115932 269153 115966 269181
rect 116114 270167 116148 270195
rect 116114 270161 116148 270167
rect 116114 270099 116148 270123
rect 116114 270089 116148 270099
rect 116114 270031 116148 270051
rect 116114 270017 116148 270031
rect 116114 269963 116148 269979
rect 116114 269945 116148 269963
rect 116114 269895 116148 269907
rect 116114 269873 116148 269895
rect 116114 269827 116148 269835
rect 116114 269801 116148 269827
rect 116114 269759 116148 269763
rect 116114 269729 116148 269759
rect 116114 269657 116148 269691
rect 116114 269589 116148 269619
rect 116114 269585 116148 269589
rect 116114 269521 116148 269547
rect 116114 269513 116148 269521
rect 116114 269453 116148 269475
rect 116114 269441 116148 269453
rect 116114 269385 116148 269403
rect 116114 269369 116148 269385
rect 116114 269317 116148 269331
rect 116114 269297 116148 269317
rect 116114 269249 116148 269259
rect 116114 269225 116148 269249
rect 116114 269181 116148 269187
rect 116114 269153 116148 269181
rect 116332 270167 116366 270195
rect 116332 270161 116366 270167
rect 116332 270099 116366 270123
rect 116332 270089 116366 270099
rect 116332 270031 116366 270051
rect 116332 270017 116366 270031
rect 116332 269963 116366 269979
rect 116332 269945 116366 269963
rect 116332 269895 116366 269907
rect 116332 269873 116366 269895
rect 116332 269827 116366 269835
rect 116332 269801 116366 269827
rect 116332 269759 116366 269763
rect 116332 269729 116366 269759
rect 116332 269657 116366 269691
rect 116332 269589 116366 269619
rect 116332 269585 116366 269589
rect 116332 269521 116366 269547
rect 116332 269513 116366 269521
rect 116332 269453 116366 269475
rect 116332 269441 116366 269453
rect 116332 269385 116366 269403
rect 116332 269369 116366 269385
rect 116332 269317 116366 269331
rect 116332 269297 116366 269317
rect 116332 269249 116366 269259
rect 116332 269225 116366 269249
rect 116332 269181 116366 269187
rect 116332 269153 116366 269181
rect 116514 270167 116548 270195
rect 116514 270161 116548 270167
rect 116514 270099 116548 270123
rect 116514 270089 116548 270099
rect 116514 270031 116548 270051
rect 116514 270017 116548 270031
rect 116514 269963 116548 269979
rect 116514 269945 116548 269963
rect 116514 269895 116548 269907
rect 116514 269873 116548 269895
rect 116514 269827 116548 269835
rect 116514 269801 116548 269827
rect 116514 269759 116548 269763
rect 116514 269729 116548 269759
rect 116514 269657 116548 269691
rect 116514 269589 116548 269619
rect 116514 269585 116548 269589
rect 116514 269521 116548 269547
rect 116514 269513 116548 269521
rect 116514 269453 116548 269475
rect 116514 269441 116548 269453
rect 116514 269385 116548 269403
rect 116514 269369 116548 269385
rect 116514 269317 116548 269331
rect 116514 269297 116548 269317
rect 116514 269249 116548 269259
rect 116514 269225 116548 269249
rect 116514 269181 116548 269187
rect 116514 269153 116548 269181
rect 116732 270167 116766 270195
rect 116732 270161 116766 270167
rect 116732 270099 116766 270123
rect 116732 270089 116766 270099
rect 116732 270031 116766 270051
rect 116732 270017 116766 270031
rect 116732 269963 116766 269979
rect 116732 269945 116766 269963
rect 116732 269895 116766 269907
rect 116732 269873 116766 269895
rect 116732 269827 116766 269835
rect 116732 269801 116766 269827
rect 116732 269759 116766 269763
rect 116732 269729 116766 269759
rect 116732 269657 116766 269691
rect 116732 269589 116766 269619
rect 116732 269585 116766 269589
rect 116732 269521 116766 269547
rect 116732 269513 116766 269521
rect 116732 269453 116766 269475
rect 116732 269441 116766 269453
rect 116732 269385 116766 269403
rect 116732 269369 116766 269385
rect 116732 269317 116766 269331
rect 116732 269297 116766 269317
rect 116732 269249 116766 269259
rect 116732 269225 116766 269249
rect 116732 269181 116766 269187
rect 116732 269153 116766 269181
rect 116914 270167 116948 270195
rect 116914 270161 116948 270167
rect 116914 270099 116948 270123
rect 116914 270089 116948 270099
rect 116914 270031 116948 270051
rect 116914 270017 116948 270031
rect 116914 269963 116948 269979
rect 116914 269945 116948 269963
rect 116914 269895 116948 269907
rect 116914 269873 116948 269895
rect 116914 269827 116948 269835
rect 116914 269801 116948 269827
rect 116914 269759 116948 269763
rect 116914 269729 116948 269759
rect 116914 269657 116948 269691
rect 116914 269589 116948 269619
rect 116914 269585 116948 269589
rect 116914 269521 116948 269547
rect 116914 269513 116948 269521
rect 116914 269453 116948 269475
rect 116914 269441 116948 269453
rect 116914 269385 116948 269403
rect 116914 269369 116948 269385
rect 116914 269317 116948 269331
rect 116914 269297 116948 269317
rect 116914 269249 116948 269259
rect 116914 269225 116948 269249
rect 116914 269181 116948 269187
rect 116914 269153 116948 269181
rect 117132 270167 117166 270195
rect 117132 270161 117166 270167
rect 117132 270099 117166 270123
rect 117132 270089 117166 270099
rect 117132 270031 117166 270051
rect 117132 270017 117166 270031
rect 117132 269963 117166 269979
rect 117132 269945 117166 269963
rect 117132 269895 117166 269907
rect 117132 269873 117166 269895
rect 117132 269827 117166 269835
rect 117132 269801 117166 269827
rect 117132 269759 117166 269763
rect 117132 269729 117166 269759
rect 117132 269657 117166 269691
rect 117132 269589 117166 269619
rect 117132 269585 117166 269589
rect 117132 269521 117166 269547
rect 117132 269513 117166 269521
rect 117132 269453 117166 269475
rect 117132 269441 117166 269453
rect 117132 269385 117166 269403
rect 117132 269369 117166 269385
rect 117132 269317 117166 269331
rect 117132 269297 117166 269317
rect 117132 269249 117166 269259
rect 117132 269225 117166 269249
rect 117132 269181 117166 269187
rect 117132 269153 117166 269181
rect 117314 270167 117348 270195
rect 117314 270161 117348 270167
rect 117314 270099 117348 270123
rect 117314 270089 117348 270099
rect 117314 270031 117348 270051
rect 117314 270017 117348 270031
rect 117314 269963 117348 269979
rect 117314 269945 117348 269963
rect 117314 269895 117348 269907
rect 117314 269873 117348 269895
rect 117314 269827 117348 269835
rect 117314 269801 117348 269827
rect 117314 269759 117348 269763
rect 117314 269729 117348 269759
rect 117314 269657 117348 269691
rect 117314 269589 117348 269619
rect 117314 269585 117348 269589
rect 117314 269521 117348 269547
rect 117314 269513 117348 269521
rect 117314 269453 117348 269475
rect 117314 269441 117348 269453
rect 117314 269385 117348 269403
rect 117314 269369 117348 269385
rect 117314 269317 117348 269331
rect 117314 269297 117348 269317
rect 117314 269249 117348 269259
rect 117314 269225 117348 269249
rect 117314 269181 117348 269187
rect 117314 269153 117348 269181
rect 117532 270167 117566 270195
rect 117532 270161 117566 270167
rect 117532 270099 117566 270123
rect 117532 270089 117566 270099
rect 117532 270031 117566 270051
rect 117532 270017 117566 270031
rect 117532 269963 117566 269979
rect 117532 269945 117566 269963
rect 117532 269895 117566 269907
rect 117532 269873 117566 269895
rect 117532 269827 117566 269835
rect 117532 269801 117566 269827
rect 117532 269759 117566 269763
rect 117532 269729 117566 269759
rect 117532 269657 117566 269691
rect 117532 269589 117566 269619
rect 117532 269585 117566 269589
rect 117532 269521 117566 269547
rect 117532 269513 117566 269521
rect 117532 269453 117566 269475
rect 117532 269441 117566 269453
rect 117532 269385 117566 269403
rect 117532 269369 117566 269385
rect 117532 269317 117566 269331
rect 117532 269297 117566 269317
rect 117532 269249 117566 269259
rect 117532 269225 117566 269249
rect 117532 269181 117566 269187
rect 117532 269153 117566 269181
rect 117714 270167 117748 270195
rect 117714 270161 117748 270167
rect 117714 270099 117748 270123
rect 117714 270089 117748 270099
rect 117714 270031 117748 270051
rect 117714 270017 117748 270031
rect 117714 269963 117748 269979
rect 117714 269945 117748 269963
rect 117714 269895 117748 269907
rect 117714 269873 117748 269895
rect 117714 269827 117748 269835
rect 117714 269801 117748 269827
rect 117714 269759 117748 269763
rect 117714 269729 117748 269759
rect 117714 269657 117748 269691
rect 117714 269589 117748 269619
rect 117714 269585 117748 269589
rect 117714 269521 117748 269547
rect 117714 269513 117748 269521
rect 117714 269453 117748 269475
rect 117714 269441 117748 269453
rect 117714 269385 117748 269403
rect 117714 269369 117748 269385
rect 117714 269317 117748 269331
rect 117714 269297 117748 269317
rect 117714 269249 117748 269259
rect 117714 269225 117748 269249
rect 117714 269181 117748 269187
rect 117714 269153 117748 269181
rect 117932 270167 117966 270195
rect 117932 270161 117966 270167
rect 117932 270099 117966 270123
rect 117932 270089 117966 270099
rect 117932 270031 117966 270051
rect 117932 270017 117966 270031
rect 117932 269963 117966 269979
rect 117932 269945 117966 269963
rect 117932 269895 117966 269907
rect 117932 269873 117966 269895
rect 117932 269827 117966 269835
rect 117932 269801 117966 269827
rect 117932 269759 117966 269763
rect 117932 269729 117966 269759
rect 117932 269657 117966 269691
rect 117932 269589 117966 269619
rect 117932 269585 117966 269589
rect 117932 269521 117966 269547
rect 117932 269513 117966 269521
rect 117932 269453 117966 269475
rect 117932 269441 117966 269453
rect 117932 269385 117966 269403
rect 117932 269369 117966 269385
rect 117932 269317 117966 269331
rect 117932 269297 117966 269317
rect 117932 269249 117966 269259
rect 117932 269225 117966 269249
rect 117932 269181 117966 269187
rect 117932 269153 117966 269181
rect 118114 270167 118148 270195
rect 118114 270161 118148 270167
rect 118114 270099 118148 270123
rect 118114 270089 118148 270099
rect 118114 270031 118148 270051
rect 118114 270017 118148 270031
rect 118114 269963 118148 269979
rect 118114 269945 118148 269963
rect 118114 269895 118148 269907
rect 118114 269873 118148 269895
rect 118114 269827 118148 269835
rect 118114 269801 118148 269827
rect 118114 269759 118148 269763
rect 118114 269729 118148 269759
rect 118114 269657 118148 269691
rect 118114 269589 118148 269619
rect 118114 269585 118148 269589
rect 118114 269521 118148 269547
rect 118114 269513 118148 269521
rect 118114 269453 118148 269475
rect 118114 269441 118148 269453
rect 118114 269385 118148 269403
rect 118114 269369 118148 269385
rect 118114 269317 118148 269331
rect 118114 269297 118148 269317
rect 118114 269249 118148 269259
rect 118114 269225 118148 269249
rect 118114 269181 118148 269187
rect 118114 269153 118148 269181
rect 118332 270167 118366 270195
rect 118332 270161 118366 270167
rect 118332 270099 118366 270123
rect 118332 270089 118366 270099
rect 118332 270031 118366 270051
rect 118332 270017 118366 270031
rect 118332 269963 118366 269979
rect 118332 269945 118366 269963
rect 118332 269895 118366 269907
rect 118332 269873 118366 269895
rect 118332 269827 118366 269835
rect 118332 269801 118366 269827
rect 118332 269759 118366 269763
rect 118332 269729 118366 269759
rect 118332 269657 118366 269691
rect 118332 269589 118366 269619
rect 118332 269585 118366 269589
rect 118332 269521 118366 269547
rect 118332 269513 118366 269521
rect 118332 269453 118366 269475
rect 118332 269441 118366 269453
rect 118332 269385 118366 269403
rect 118332 269369 118366 269385
rect 118332 269317 118366 269331
rect 118332 269297 118366 269317
rect 118332 269249 118366 269259
rect 118332 269225 118366 269249
rect 118332 269181 118366 269187
rect 118332 269153 118366 269181
rect 118514 270167 118548 270195
rect 118514 270161 118548 270167
rect 118514 270099 118548 270123
rect 118514 270089 118548 270099
rect 118514 270031 118548 270051
rect 118514 270017 118548 270031
rect 118514 269963 118548 269979
rect 118514 269945 118548 269963
rect 118514 269895 118548 269907
rect 118514 269873 118548 269895
rect 118514 269827 118548 269835
rect 118514 269801 118548 269827
rect 118514 269759 118548 269763
rect 118514 269729 118548 269759
rect 118514 269657 118548 269691
rect 118514 269589 118548 269619
rect 118514 269585 118548 269589
rect 118514 269521 118548 269547
rect 118514 269513 118548 269521
rect 118514 269453 118548 269475
rect 118514 269441 118548 269453
rect 118514 269385 118548 269403
rect 118514 269369 118548 269385
rect 118514 269317 118548 269331
rect 118514 269297 118548 269317
rect 118514 269249 118548 269259
rect 118514 269225 118548 269249
rect 118514 269181 118548 269187
rect 118514 269153 118548 269181
rect 118732 270167 118766 270195
rect 118732 270161 118766 270167
rect 118732 270099 118766 270123
rect 118732 270089 118766 270099
rect 118732 270031 118766 270051
rect 118732 270017 118766 270031
rect 118732 269963 118766 269979
rect 118732 269945 118766 269963
rect 118732 269895 118766 269907
rect 118732 269873 118766 269895
rect 118732 269827 118766 269835
rect 118732 269801 118766 269827
rect 118732 269759 118766 269763
rect 118732 269729 118766 269759
rect 118732 269657 118766 269691
rect 118732 269589 118766 269619
rect 118732 269585 118766 269589
rect 118732 269521 118766 269547
rect 118732 269513 118766 269521
rect 118732 269453 118766 269475
rect 118732 269441 118766 269453
rect 118732 269385 118766 269403
rect 118732 269369 118766 269385
rect 118732 269317 118766 269331
rect 118732 269297 118766 269317
rect 118732 269249 118766 269259
rect 118732 269225 118766 269249
rect 118732 269181 118766 269187
rect 118732 269153 118766 269181
rect 112587 269052 112589 269086
rect 112589 269052 112621 269086
rect 112659 269052 112691 269086
rect 112691 269052 112693 269086
rect 112987 269052 112989 269086
rect 112989 269052 113021 269086
rect 113059 269052 113091 269086
rect 113091 269052 113093 269086
rect 113387 269052 113389 269086
rect 113389 269052 113421 269086
rect 113459 269052 113491 269086
rect 113491 269052 113493 269086
rect 113787 269052 113789 269086
rect 113789 269052 113821 269086
rect 113859 269052 113891 269086
rect 113891 269052 113893 269086
rect 114187 269052 114189 269086
rect 114189 269052 114221 269086
rect 114259 269052 114291 269086
rect 114291 269052 114293 269086
rect 114587 269052 114589 269086
rect 114589 269052 114621 269086
rect 114659 269052 114691 269086
rect 114691 269052 114693 269086
rect 114987 269052 114989 269086
rect 114989 269052 115021 269086
rect 115059 269052 115091 269086
rect 115091 269052 115093 269086
rect 115387 269052 115389 269086
rect 115389 269052 115421 269086
rect 115459 269052 115491 269086
rect 115491 269052 115493 269086
rect 115787 269052 115789 269086
rect 115789 269052 115821 269086
rect 115859 269052 115891 269086
rect 115891 269052 115893 269086
rect 116187 269052 116189 269086
rect 116189 269052 116221 269086
rect 116259 269052 116291 269086
rect 116291 269052 116293 269086
rect 116587 269052 116589 269086
rect 116589 269052 116621 269086
rect 116659 269052 116691 269086
rect 116691 269052 116693 269086
rect 116987 269052 116989 269086
rect 116989 269052 117021 269086
rect 117059 269052 117091 269086
rect 117091 269052 117093 269086
rect 117387 269052 117389 269086
rect 117389 269052 117421 269086
rect 117459 269052 117491 269086
rect 117491 269052 117493 269086
rect 117787 269052 117789 269086
rect 117789 269052 117821 269086
rect 117859 269052 117891 269086
rect 117891 269052 117893 269086
rect 118187 269052 118189 269086
rect 118189 269052 118221 269086
rect 118259 269052 118291 269086
rect 118291 269052 118293 269086
rect 118587 269052 118589 269086
rect 118589 269052 118621 269086
rect 118659 269052 118691 269086
rect 118691 269052 118693 269086
rect 114345 268815 117475 268868
rect 114345 268762 117475 268815
rect 120468 280684 120476 280718
rect 120476 280684 120502 280718
rect 120540 280684 120544 280718
rect 120544 280684 120574 280718
rect 120612 280684 120646 280718
rect 120684 280684 120714 280718
rect 120714 280684 120718 280718
rect 120756 280684 120782 280718
rect 120782 280684 120790 280718
rect 120383 280570 120417 280604
rect 120841 280570 120875 280604
rect 121168 280684 121176 280718
rect 121176 280684 121202 280718
rect 121240 280684 121244 280718
rect 121244 280684 121274 280718
rect 121312 280684 121346 280718
rect 121384 280684 121414 280718
rect 121414 280684 121418 280718
rect 121456 280684 121482 280718
rect 121482 280684 121490 280718
rect 121083 280570 121117 280604
rect 121541 280570 121575 280604
rect 120468 280456 120476 280490
rect 120476 280456 120502 280490
rect 120540 280456 120544 280490
rect 120544 280456 120574 280490
rect 120612 280456 120646 280490
rect 120684 280456 120714 280490
rect 120714 280456 120718 280490
rect 120756 280456 120782 280490
rect 120782 280456 120790 280490
rect 121168 280456 121176 280490
rect 121176 280456 121202 280490
rect 121240 280456 121244 280490
rect 121244 280456 121274 280490
rect 121312 280456 121346 280490
rect 121384 280456 121414 280490
rect 121414 280456 121418 280490
rect 121456 280456 121482 280490
rect 121482 280456 121490 280490
rect 120468 280300 120476 280334
rect 120476 280300 120502 280334
rect 120540 280300 120544 280334
rect 120544 280300 120574 280334
rect 120612 280300 120646 280334
rect 120684 280300 120714 280334
rect 120714 280300 120718 280334
rect 120756 280300 120782 280334
rect 120782 280300 120790 280334
rect 121168 280300 121176 280334
rect 121176 280300 121202 280334
rect 121240 280300 121244 280334
rect 121244 280300 121274 280334
rect 121312 280300 121346 280334
rect 121384 280300 121414 280334
rect 121414 280300 121418 280334
rect 121456 280300 121482 280334
rect 121482 280300 121490 280334
rect 120383 280224 120417 280236
rect 120383 280202 120417 280224
rect 120383 280156 120417 280164
rect 120383 280130 120417 280156
rect 120383 280088 120417 280092
rect 120383 280058 120417 280088
rect 120383 279986 120417 280020
rect 120383 279918 120417 279948
rect 120383 279914 120417 279918
rect 120383 279850 120417 279876
rect 120383 279842 120417 279850
rect 120383 279782 120417 279804
rect 120383 279770 120417 279782
rect 120841 280224 120875 280236
rect 120841 280202 120875 280224
rect 120841 280156 120875 280164
rect 120841 280130 120875 280156
rect 120841 280088 120875 280092
rect 120841 280058 120875 280088
rect 120841 279986 120875 280020
rect 120841 279918 120875 279948
rect 120841 279914 120875 279918
rect 120841 279850 120875 279876
rect 120841 279842 120875 279850
rect 120841 279782 120875 279804
rect 120841 279770 120875 279782
rect 121083 280224 121117 280236
rect 121083 280202 121117 280224
rect 121083 280156 121117 280164
rect 121083 280130 121117 280156
rect 121083 280088 121117 280092
rect 121083 280058 121117 280088
rect 121083 279986 121117 280020
rect 121083 279918 121117 279948
rect 121083 279914 121117 279918
rect 121083 279850 121117 279876
rect 121083 279842 121117 279850
rect 121083 279782 121117 279804
rect 121083 279770 121117 279782
rect 121541 280224 121575 280236
rect 121541 280202 121575 280224
rect 121541 280156 121575 280164
rect 121541 280130 121575 280156
rect 121541 280088 121575 280092
rect 121541 280058 121575 280088
rect 121541 279986 121575 280020
rect 121541 279918 121575 279948
rect 121541 279914 121575 279918
rect 121541 279850 121575 279876
rect 121541 279842 121575 279850
rect 121541 279782 121575 279804
rect 121541 279770 121575 279782
rect 122395 280470 122403 280504
rect 122403 280470 122429 280504
rect 122467 280470 122471 280504
rect 122471 280470 122501 280504
rect 122539 280470 122573 280504
rect 122611 280470 122641 280504
rect 122641 280470 122645 280504
rect 122683 280470 122709 280504
rect 122709 280470 122717 280504
rect 123095 280470 123103 280504
rect 123103 280470 123129 280504
rect 123167 280470 123171 280504
rect 123171 280470 123201 280504
rect 123239 280470 123273 280504
rect 123311 280470 123341 280504
rect 123341 280470 123345 280504
rect 123383 280470 123409 280504
rect 123409 280470 123417 280504
rect 122310 280394 122344 280406
rect 122310 280372 122344 280394
rect 122310 280326 122344 280334
rect 122310 280300 122344 280326
rect 122310 280258 122344 280262
rect 122310 280228 122344 280258
rect 122310 280156 122344 280190
rect 122310 280088 122344 280118
rect 122310 280084 122344 280088
rect 122310 280020 122344 280046
rect 122310 280012 122344 280020
rect 122310 279952 122344 279974
rect 122310 279940 122344 279952
rect 122768 280394 122802 280406
rect 122768 280372 122802 280394
rect 122768 280326 122802 280334
rect 122768 280300 122802 280326
rect 122768 280258 122802 280262
rect 122768 280228 122802 280258
rect 122768 280156 122802 280190
rect 122768 280088 122802 280118
rect 122768 280084 122802 280088
rect 122768 280020 122802 280046
rect 122768 280012 122802 280020
rect 122768 279952 122802 279974
rect 122768 279940 122802 279952
rect 123010 280394 123044 280406
rect 123010 280372 123044 280394
rect 123010 280326 123044 280334
rect 123010 280300 123044 280326
rect 123010 280258 123044 280262
rect 123010 280228 123044 280258
rect 123010 280156 123044 280190
rect 123010 280088 123044 280118
rect 123010 280084 123044 280088
rect 123010 280020 123044 280046
rect 123010 280012 123044 280020
rect 123010 279952 123044 279974
rect 123010 279940 123044 279952
rect 123468 280394 123502 280406
rect 123468 280372 123502 280394
rect 123468 280326 123502 280334
rect 123468 280300 123502 280326
rect 123468 280258 123502 280262
rect 123468 280228 123502 280258
rect 123468 280156 123502 280190
rect 123468 280088 123502 280118
rect 123468 280084 123502 280088
rect 123468 280020 123502 280046
rect 123468 280012 123502 280020
rect 123468 279952 123502 279974
rect 123468 279940 123502 279952
rect 121859 279872 122178 279886
rect 122178 279872 122181 279886
rect 121859 279838 122181 279872
rect 122395 279842 122403 279876
rect 122403 279842 122429 279876
rect 122467 279842 122471 279876
rect 122471 279842 122501 279876
rect 122539 279842 122573 279876
rect 122611 279842 122641 279876
rect 122641 279842 122645 279876
rect 122683 279842 122709 279876
rect 122709 279842 122717 279876
rect 123095 279842 123103 279876
rect 123103 279842 123129 279876
rect 123167 279842 123171 279876
rect 123171 279842 123201 279876
rect 123239 279842 123273 279876
rect 123311 279842 123341 279876
rect 123341 279842 123345 279876
rect 123383 279842 123409 279876
rect 123409 279842 123417 279876
rect 121859 279804 122178 279838
rect 122178 279804 122181 279838
rect 121859 279770 122181 279804
rect 121859 279736 122178 279770
rect 122178 279736 122181 279770
rect 120468 279672 120476 279706
rect 120476 279672 120502 279706
rect 120540 279672 120544 279706
rect 120544 279672 120574 279706
rect 120612 279672 120646 279706
rect 120684 279672 120714 279706
rect 120714 279672 120718 279706
rect 120756 279672 120782 279706
rect 120782 279672 120790 279706
rect 121168 279672 121176 279706
rect 121176 279672 121202 279706
rect 121240 279672 121244 279706
rect 121244 279672 121274 279706
rect 121312 279672 121346 279706
rect 121384 279672 121414 279706
rect 121414 279672 121418 279706
rect 121456 279672 121482 279706
rect 121482 279672 121490 279706
rect 121859 279702 122181 279736
rect 121859 279668 122178 279702
rect 122178 279668 122181 279702
rect 122395 279686 122403 279720
rect 122403 279686 122429 279720
rect 122467 279686 122471 279720
rect 122471 279686 122501 279720
rect 122539 279686 122573 279720
rect 122611 279686 122641 279720
rect 122641 279686 122645 279720
rect 122683 279686 122709 279720
rect 122709 279686 122717 279720
rect 123095 279686 123103 279720
rect 123103 279686 123129 279720
rect 123167 279686 123171 279720
rect 123171 279686 123201 279720
rect 123239 279686 123273 279720
rect 123311 279686 123341 279720
rect 123341 279686 123345 279720
rect 123383 279686 123409 279720
rect 123409 279686 123417 279720
rect 121859 279634 122181 279668
rect 121859 279600 122178 279634
rect 122178 279600 122181 279634
rect 122310 279610 122344 279622
rect 120468 279516 120476 279550
rect 120476 279516 120502 279550
rect 120540 279516 120544 279550
rect 120544 279516 120574 279550
rect 120612 279516 120646 279550
rect 120684 279516 120714 279550
rect 120714 279516 120718 279550
rect 120756 279516 120782 279550
rect 120782 279516 120790 279550
rect 121168 279516 121176 279550
rect 121176 279516 121202 279550
rect 121240 279516 121244 279550
rect 121244 279516 121274 279550
rect 121312 279516 121346 279550
rect 121384 279516 121414 279550
rect 121414 279516 121418 279550
rect 121456 279516 121482 279550
rect 121482 279516 121490 279550
rect 121859 279566 122181 279600
rect 122310 279588 122344 279610
rect 121859 279532 122178 279566
rect 122178 279532 122181 279566
rect 122310 279542 122344 279550
rect 120383 279440 120417 279452
rect 120383 279418 120417 279440
rect 120383 279372 120417 279380
rect 120383 279346 120417 279372
rect 120383 279304 120417 279308
rect 120383 279274 120417 279304
rect 120383 279202 120417 279236
rect 120383 279134 120417 279164
rect 120383 279130 120417 279134
rect 120383 279066 120417 279092
rect 120383 279058 120417 279066
rect 120383 278998 120417 279020
rect 120383 278986 120417 278998
rect 120841 279440 120875 279452
rect 120841 279418 120875 279440
rect 120841 279372 120875 279380
rect 120841 279346 120875 279372
rect 120841 279304 120875 279308
rect 120841 279274 120875 279304
rect 120841 279202 120875 279236
rect 120841 279134 120875 279164
rect 120841 279130 120875 279134
rect 120841 279066 120875 279092
rect 120841 279058 120875 279066
rect 120841 278998 120875 279020
rect 120841 278986 120875 278998
rect 121083 279440 121117 279452
rect 121083 279418 121117 279440
rect 121083 279372 121117 279380
rect 121083 279346 121117 279372
rect 121083 279304 121117 279308
rect 121083 279274 121117 279304
rect 121083 279202 121117 279236
rect 121083 279134 121117 279164
rect 121083 279130 121117 279134
rect 121083 279066 121117 279092
rect 121083 279058 121117 279066
rect 121083 278998 121117 279020
rect 121083 278986 121117 278998
rect 121541 279440 121575 279452
rect 121541 279418 121575 279440
rect 121541 279372 121575 279380
rect 121541 279346 121575 279372
rect 121541 279304 121575 279308
rect 121541 279274 121575 279304
rect 121541 279202 121575 279236
rect 121541 279134 121575 279164
rect 121541 279130 121575 279134
rect 121541 279066 121575 279092
rect 121541 279058 121575 279066
rect 121541 278998 121575 279020
rect 121541 278986 121575 278998
rect 121859 279498 122181 279532
rect 122310 279516 122344 279542
rect 121859 279464 122178 279498
rect 122178 279464 122181 279498
rect 122310 279474 122344 279478
rect 121859 279430 122181 279464
rect 122310 279444 122344 279474
rect 121859 279396 122178 279430
rect 122178 279396 122181 279430
rect 121859 279362 122181 279396
rect 122310 279372 122344 279406
rect 121859 279328 122178 279362
rect 122178 279328 122181 279362
rect 121859 279294 122181 279328
rect 122310 279304 122344 279334
rect 122310 279300 122344 279304
rect 121859 279276 122178 279294
rect 122178 279276 122181 279294
rect 122310 279236 122344 279262
rect 122310 279228 122344 279236
rect 122310 279168 122344 279190
rect 122310 279156 122344 279168
rect 122768 279610 122802 279622
rect 122768 279588 122802 279610
rect 122768 279542 122802 279550
rect 122768 279516 122802 279542
rect 122768 279474 122802 279478
rect 122768 279444 122802 279474
rect 122768 279372 122802 279406
rect 122768 279304 122802 279334
rect 122768 279300 122802 279304
rect 122768 279236 122802 279262
rect 122768 279228 122802 279236
rect 122768 279168 122802 279190
rect 122768 279156 122802 279168
rect 123010 279610 123044 279622
rect 123010 279588 123044 279610
rect 123010 279542 123044 279550
rect 123010 279516 123044 279542
rect 123010 279474 123044 279478
rect 123010 279444 123044 279474
rect 123010 279372 123044 279406
rect 123010 279304 123044 279334
rect 123010 279300 123044 279304
rect 123010 279236 123044 279262
rect 123010 279228 123044 279236
rect 123010 279168 123044 279190
rect 123010 279156 123044 279168
rect 123468 279610 123502 279622
rect 123468 279588 123502 279610
rect 123468 279542 123502 279550
rect 123468 279516 123502 279542
rect 123468 279474 123502 279478
rect 123468 279444 123502 279474
rect 123468 279372 123502 279406
rect 123468 279304 123502 279334
rect 123468 279300 123502 279304
rect 123468 279236 123502 279262
rect 123468 279228 123502 279236
rect 123468 279168 123502 279190
rect 123468 279156 123502 279168
rect 122395 279058 122403 279092
rect 122403 279058 122429 279092
rect 122467 279058 122471 279092
rect 122471 279058 122501 279092
rect 122539 279058 122573 279092
rect 122611 279058 122641 279092
rect 122641 279058 122645 279092
rect 122683 279058 122709 279092
rect 122709 279058 122717 279092
rect 123095 279058 123103 279092
rect 123103 279058 123129 279092
rect 123167 279058 123171 279092
rect 123171 279058 123201 279092
rect 123239 279058 123273 279092
rect 123311 279058 123341 279092
rect 123341 279058 123345 279092
rect 123383 279058 123409 279092
rect 123409 279058 123417 279092
rect 120468 278888 120476 278922
rect 120476 278888 120502 278922
rect 120540 278888 120544 278922
rect 120544 278888 120574 278922
rect 120612 278888 120646 278922
rect 120684 278888 120714 278922
rect 120714 278888 120718 278922
rect 120756 278888 120782 278922
rect 120782 278888 120790 278922
rect 121168 278888 121176 278922
rect 121176 278888 121202 278922
rect 121240 278888 121244 278922
rect 121244 278888 121274 278922
rect 121312 278888 121346 278922
rect 121384 278888 121414 278922
rect 121414 278888 121418 278922
rect 121456 278888 121482 278922
rect 121482 278888 121490 278922
rect 120468 278732 120476 278766
rect 120476 278732 120502 278766
rect 120540 278732 120544 278766
rect 120544 278732 120574 278766
rect 120612 278732 120646 278766
rect 120684 278732 120714 278766
rect 120714 278732 120718 278766
rect 120756 278732 120782 278766
rect 120782 278732 120790 278766
rect 121168 278732 121176 278766
rect 121176 278732 121202 278766
rect 121240 278732 121244 278766
rect 121244 278732 121274 278766
rect 121312 278732 121346 278766
rect 121384 278732 121414 278766
rect 121414 278732 121418 278766
rect 121456 278732 121482 278766
rect 121482 278732 121490 278766
rect 120383 278656 120417 278668
rect 120383 278634 120417 278656
rect 120383 278588 120417 278596
rect 120383 278562 120417 278588
rect 120383 278520 120417 278524
rect 120383 278490 120417 278520
rect 120383 278418 120417 278452
rect 120383 278350 120417 278380
rect 120383 278346 120417 278350
rect 120383 278282 120417 278308
rect 120383 278274 120417 278282
rect 120383 278214 120417 278236
rect 120383 278202 120417 278214
rect 120841 278656 120875 278668
rect 120841 278634 120875 278656
rect 120841 278588 120875 278596
rect 120841 278562 120875 278588
rect 120841 278520 120875 278524
rect 120841 278490 120875 278520
rect 120841 278418 120875 278452
rect 120841 278350 120875 278380
rect 120841 278346 120875 278350
rect 120841 278282 120875 278308
rect 120841 278274 120875 278282
rect 120841 278214 120875 278236
rect 120841 278202 120875 278214
rect 121083 278656 121117 278668
rect 121083 278634 121117 278656
rect 121083 278588 121117 278596
rect 121083 278562 121117 278588
rect 121083 278520 121117 278524
rect 121083 278490 121117 278520
rect 121083 278418 121117 278452
rect 121083 278350 121117 278380
rect 121083 278346 121117 278350
rect 121083 278282 121117 278308
rect 121083 278274 121117 278282
rect 121083 278214 121117 278236
rect 121083 278202 121117 278214
rect 121541 278656 121575 278668
rect 121541 278634 121575 278656
rect 121541 278588 121575 278596
rect 121541 278562 121575 278588
rect 121541 278520 121575 278524
rect 121541 278490 121575 278520
rect 121541 278418 121575 278452
rect 121541 278350 121575 278380
rect 121541 278346 121575 278350
rect 121541 278282 121575 278308
rect 121541 278274 121575 278282
rect 121541 278214 121575 278236
rect 121541 278202 121575 278214
rect 120468 278104 120476 278138
rect 120476 278104 120502 278138
rect 120540 278104 120544 278138
rect 120544 278104 120574 278138
rect 120612 278104 120646 278138
rect 120684 278104 120714 278138
rect 120714 278104 120718 278138
rect 120756 278104 120782 278138
rect 120782 278104 120790 278138
rect 121168 278104 121176 278138
rect 121176 278104 121202 278138
rect 121240 278104 121244 278138
rect 121244 278104 121274 278138
rect 121312 278104 121346 278138
rect 121384 278104 121414 278138
rect 121414 278104 121418 278138
rect 121456 278104 121482 278138
rect 121482 278104 121490 278138
rect 120468 277948 120476 277982
rect 120476 277948 120502 277982
rect 120540 277948 120544 277982
rect 120544 277948 120574 277982
rect 120612 277948 120646 277982
rect 120684 277948 120714 277982
rect 120714 277948 120718 277982
rect 120756 277948 120782 277982
rect 120782 277948 120790 277982
rect 121168 277948 121176 277982
rect 121176 277948 121202 277982
rect 121240 277948 121244 277982
rect 121244 277948 121274 277982
rect 121312 277948 121346 277982
rect 121384 277948 121414 277982
rect 121414 277948 121418 277982
rect 121456 277948 121482 277982
rect 121482 277948 121490 277982
rect 120383 277872 120417 277884
rect 120383 277850 120417 277872
rect 120383 277804 120417 277812
rect 120383 277778 120417 277804
rect 120383 277736 120417 277740
rect 120383 277706 120417 277736
rect 120383 277634 120417 277668
rect 120383 277566 120417 277596
rect 120383 277562 120417 277566
rect 120383 277498 120417 277524
rect 120383 277490 120417 277498
rect 120383 277430 120417 277452
rect 120383 277418 120417 277430
rect 120841 277872 120875 277884
rect 120841 277850 120875 277872
rect 120841 277804 120875 277812
rect 120841 277778 120875 277804
rect 120841 277736 120875 277740
rect 120841 277706 120875 277736
rect 120841 277634 120875 277668
rect 120841 277566 120875 277596
rect 120841 277562 120875 277566
rect 120841 277498 120875 277524
rect 120841 277490 120875 277498
rect 120841 277430 120875 277452
rect 120841 277418 120875 277430
rect 121083 277872 121117 277884
rect 121083 277850 121117 277872
rect 121083 277804 121117 277812
rect 121083 277778 121117 277804
rect 121083 277736 121117 277740
rect 121083 277706 121117 277736
rect 121083 277634 121117 277668
rect 121083 277566 121117 277596
rect 121083 277562 121117 277566
rect 121083 277498 121117 277524
rect 121083 277490 121117 277498
rect 121083 277430 121117 277452
rect 121083 277418 121117 277430
rect 121541 277872 121575 277884
rect 121541 277850 121575 277872
rect 121541 277804 121575 277812
rect 121541 277778 121575 277804
rect 121541 277736 121575 277740
rect 121541 277706 121575 277736
rect 121541 277634 121575 277668
rect 121541 277566 121575 277596
rect 121541 277562 121575 277566
rect 121541 277498 121575 277524
rect 121541 277490 121575 277498
rect 121541 277430 121575 277452
rect 121541 277418 121575 277430
rect 120468 277320 120476 277354
rect 120476 277320 120502 277354
rect 120540 277320 120544 277354
rect 120544 277320 120574 277354
rect 120612 277320 120646 277354
rect 120684 277320 120714 277354
rect 120714 277320 120718 277354
rect 120756 277320 120782 277354
rect 120782 277320 120790 277354
rect 121168 277320 121176 277354
rect 121176 277320 121202 277354
rect 121240 277320 121244 277354
rect 121244 277320 121274 277354
rect 121312 277320 121346 277354
rect 121384 277320 121414 277354
rect 121414 277320 121418 277354
rect 121456 277320 121482 277354
rect 121482 277320 121490 277354
rect 120468 277164 120476 277198
rect 120476 277164 120502 277198
rect 120540 277164 120544 277198
rect 120544 277164 120574 277198
rect 120612 277164 120646 277198
rect 120684 277164 120714 277198
rect 120714 277164 120718 277198
rect 120756 277164 120782 277198
rect 120782 277164 120790 277198
rect 121168 277164 121176 277198
rect 121176 277164 121202 277198
rect 121240 277164 121244 277198
rect 121244 277164 121274 277198
rect 121312 277164 121346 277198
rect 121384 277164 121414 277198
rect 121414 277164 121418 277198
rect 121456 277164 121482 277198
rect 121482 277164 121490 277198
rect 120383 277088 120417 277100
rect 120383 277066 120417 277088
rect 120383 277020 120417 277028
rect 120383 276994 120417 277020
rect 120383 276952 120417 276956
rect 120383 276922 120417 276952
rect 120383 276850 120417 276884
rect 120383 276782 120417 276812
rect 120383 276778 120417 276782
rect 120383 276714 120417 276740
rect 120383 276706 120417 276714
rect 120383 276646 120417 276668
rect 120383 276634 120417 276646
rect 120841 277088 120875 277100
rect 120841 277066 120875 277088
rect 120841 277020 120875 277028
rect 120841 276994 120875 277020
rect 120841 276952 120875 276956
rect 120841 276922 120875 276952
rect 120841 276850 120875 276884
rect 120841 276782 120875 276812
rect 120841 276778 120875 276782
rect 120841 276714 120875 276740
rect 120841 276706 120875 276714
rect 120841 276646 120875 276668
rect 120841 276634 120875 276646
rect 121083 277088 121117 277100
rect 121083 277066 121117 277088
rect 121083 277020 121117 277028
rect 121083 276994 121117 277020
rect 121083 276952 121117 276956
rect 121083 276922 121117 276952
rect 121083 276850 121117 276884
rect 121083 276782 121117 276812
rect 121083 276778 121117 276782
rect 121083 276714 121117 276740
rect 121083 276706 121117 276714
rect 121083 276646 121117 276668
rect 121083 276634 121117 276646
rect 121541 277088 121575 277100
rect 121541 277066 121575 277088
rect 121541 277020 121575 277028
rect 121541 276994 121575 277020
rect 121541 276952 121575 276956
rect 121541 276922 121575 276952
rect 121541 276850 121575 276884
rect 121541 276782 121575 276812
rect 121541 276778 121575 276782
rect 121541 276714 121575 276740
rect 121541 276706 121575 276714
rect 121541 276646 121575 276668
rect 121541 276634 121575 276646
rect 120468 276536 120476 276570
rect 120476 276536 120502 276570
rect 120540 276536 120544 276570
rect 120544 276536 120574 276570
rect 120612 276536 120646 276570
rect 120684 276536 120714 276570
rect 120714 276536 120718 276570
rect 120756 276536 120782 276570
rect 120782 276536 120790 276570
rect 121168 276536 121176 276570
rect 121176 276536 121202 276570
rect 121240 276536 121244 276570
rect 121244 276536 121274 276570
rect 121312 276536 121346 276570
rect 121384 276536 121414 276570
rect 121414 276536 121418 276570
rect 121456 276536 121482 276570
rect 121482 276536 121490 276570
rect 120468 276380 120476 276414
rect 120476 276380 120502 276414
rect 120540 276380 120544 276414
rect 120544 276380 120574 276414
rect 120612 276380 120646 276414
rect 120684 276380 120714 276414
rect 120714 276380 120718 276414
rect 120756 276380 120782 276414
rect 120782 276380 120790 276414
rect 121168 276380 121176 276414
rect 121176 276380 121202 276414
rect 121240 276380 121244 276414
rect 121244 276380 121274 276414
rect 121312 276380 121346 276414
rect 121384 276380 121414 276414
rect 121414 276380 121418 276414
rect 121456 276380 121482 276414
rect 121482 276380 121490 276414
rect 120383 276304 120417 276316
rect 120383 276282 120417 276304
rect 120383 276236 120417 276244
rect 120383 276210 120417 276236
rect 120383 276168 120417 276172
rect 120383 276138 120417 276168
rect 120383 276066 120417 276100
rect 120383 275998 120417 276028
rect 120383 275994 120417 275998
rect 120383 275930 120417 275956
rect 120383 275922 120417 275930
rect 120383 275862 120417 275884
rect 120383 275850 120417 275862
rect 120841 276304 120875 276316
rect 120841 276282 120875 276304
rect 120841 276236 120875 276244
rect 120841 276210 120875 276236
rect 120841 276168 120875 276172
rect 120841 276138 120875 276168
rect 121083 276304 121117 276316
rect 121083 276282 121117 276304
rect 121083 276236 121117 276244
rect 121083 276210 121117 276236
rect 121083 276168 121117 276172
rect 121083 276138 121117 276168
rect 120841 276066 120875 276100
rect 120969 276069 121003 276103
rect 121083 276066 121117 276100
rect 120841 275998 120875 276028
rect 120841 275994 120875 275998
rect 120841 275930 120875 275956
rect 120841 275922 120875 275930
rect 120841 275862 120875 275884
rect 120841 275850 120875 275862
rect 121083 275998 121117 276028
rect 121083 275994 121117 275998
rect 121083 275930 121117 275956
rect 121083 275922 121117 275930
rect 121083 275862 121117 275884
rect 121083 275850 121117 275862
rect 121541 276304 121575 276316
rect 121541 276282 121575 276304
rect 121541 276236 121575 276244
rect 121541 276210 121575 276236
rect 121541 276168 121575 276172
rect 121541 276138 121575 276168
rect 121541 276066 121575 276100
rect 121541 275998 121575 276028
rect 121541 275994 121575 275998
rect 121541 275930 121575 275956
rect 121541 275922 121575 275930
rect 121541 275862 121575 275884
rect 121541 275850 121575 275862
rect 120468 275752 120476 275786
rect 120476 275752 120502 275786
rect 120540 275752 120544 275786
rect 120544 275752 120574 275786
rect 120612 275752 120646 275786
rect 120684 275752 120714 275786
rect 120714 275752 120718 275786
rect 120756 275752 120782 275786
rect 120782 275752 120790 275786
rect 121168 275752 121176 275786
rect 121176 275752 121202 275786
rect 121240 275752 121244 275786
rect 121244 275752 121274 275786
rect 121312 275752 121346 275786
rect 121384 275752 121414 275786
rect 121414 275752 121418 275786
rect 121456 275752 121482 275786
rect 121482 275752 121490 275786
rect 120468 275596 120476 275630
rect 120476 275596 120502 275630
rect 120540 275596 120544 275630
rect 120544 275596 120574 275630
rect 120612 275596 120646 275630
rect 120684 275596 120714 275630
rect 120714 275596 120718 275630
rect 120756 275596 120782 275630
rect 120782 275596 120790 275630
rect 121168 275596 121176 275630
rect 121176 275596 121202 275630
rect 121240 275596 121244 275630
rect 121244 275596 121274 275630
rect 121312 275596 121346 275630
rect 121384 275596 121414 275630
rect 121414 275596 121418 275630
rect 121456 275596 121482 275630
rect 121482 275596 121490 275630
rect 120383 275520 120417 275532
rect 120383 275498 120417 275520
rect 120383 275452 120417 275460
rect 120383 275426 120417 275452
rect 120383 275384 120417 275388
rect 120383 275354 120417 275384
rect 120383 275282 120417 275316
rect 120383 275214 120417 275244
rect 120383 275210 120417 275214
rect 120383 275146 120417 275172
rect 120383 275138 120417 275146
rect 120383 275078 120417 275100
rect 120383 275066 120417 275078
rect 120841 275520 120875 275532
rect 120841 275498 120875 275520
rect 120841 275452 120875 275460
rect 120841 275426 120875 275452
rect 120841 275384 120875 275388
rect 120841 275354 120875 275384
rect 121083 275520 121117 275532
rect 121083 275498 121117 275520
rect 121083 275452 121117 275460
rect 121083 275426 121117 275452
rect 121083 275384 121117 275388
rect 121083 275354 121117 275384
rect 120841 275282 120875 275316
rect 121083 275282 121117 275316
rect 120841 275214 120875 275244
rect 120841 275210 120875 275214
rect 120841 275146 120875 275172
rect 120841 275138 120875 275146
rect 120841 275078 120875 275100
rect 120841 275066 120875 275078
rect 120468 274968 120476 275002
rect 120476 274968 120502 275002
rect 120540 274968 120544 275002
rect 120544 274968 120574 275002
rect 120612 274968 120646 275002
rect 120684 274968 120714 275002
rect 120714 274968 120718 275002
rect 120756 274968 120782 275002
rect 120782 274968 120790 275002
rect 120468 274812 120476 274846
rect 120476 274812 120502 274846
rect 120540 274812 120544 274846
rect 120544 274812 120574 274846
rect 120612 274812 120646 274846
rect 120684 274812 120714 274846
rect 120714 274812 120718 274846
rect 120756 274812 120782 274846
rect 120782 274812 120790 274846
rect 120383 274736 120417 274748
rect 120383 274714 120417 274736
rect 120383 274668 120417 274676
rect 120383 274642 120417 274668
rect 120383 274600 120417 274604
rect 120383 274570 120417 274600
rect 120383 274498 120417 274532
rect 120383 274430 120417 274460
rect 120383 274426 120417 274430
rect 120383 274362 120417 274388
rect 120383 274354 120417 274362
rect 120383 274294 120417 274316
rect 120383 274282 120417 274294
rect 120841 274736 120875 274748
rect 120841 274714 120875 274736
rect 120841 274668 120875 274676
rect 120841 274642 120875 274668
rect 120841 274600 120875 274604
rect 120841 274570 120875 274600
rect 121083 275214 121117 275244
rect 121083 275210 121117 275214
rect 121083 275146 121117 275172
rect 121083 275138 121117 275146
rect 121083 275078 121117 275100
rect 121083 275066 121117 275078
rect 121541 275520 121575 275532
rect 121541 275498 121575 275520
rect 121541 275452 121575 275460
rect 121541 275426 121575 275452
rect 121541 275384 121575 275388
rect 121541 275354 121575 275384
rect 121541 275282 121575 275316
rect 121541 275214 121575 275244
rect 121541 275210 121575 275214
rect 121541 275146 121575 275172
rect 121541 275138 121575 275146
rect 121541 275078 121575 275100
rect 121541 275066 121575 275078
rect 122439 278313 122461 278347
rect 122461 278313 122473 278347
rect 122511 278313 122529 278347
rect 122529 278313 122545 278347
rect 122583 278313 122597 278347
rect 122597 278313 122617 278347
rect 122655 278313 122665 278347
rect 122665 278313 122689 278347
rect 122727 278313 122733 278347
rect 122733 278313 122761 278347
rect 122799 278313 122801 278347
rect 122801 278313 122833 278347
rect 122871 278313 122903 278347
rect 122903 278313 122905 278347
rect 122943 278313 122971 278347
rect 122971 278313 122977 278347
rect 123015 278313 123039 278347
rect 123039 278313 123049 278347
rect 123087 278313 123107 278347
rect 123107 278313 123121 278347
rect 123159 278313 123175 278347
rect 123175 278313 123193 278347
rect 123231 278313 123243 278347
rect 123243 278313 123265 278347
rect 122368 278216 122402 278226
rect 122368 278192 122402 278216
rect 122368 278148 122402 278154
rect 122368 278120 122402 278148
rect 122368 278080 122402 278082
rect 122368 278048 122402 278080
rect 122368 277978 122402 278010
rect 122368 277976 122402 277978
rect 122368 277910 122402 277938
rect 122368 277904 122402 277910
rect 122368 277842 122402 277866
rect 122368 277832 122402 277842
rect 123302 278216 123336 278226
rect 123302 278192 123336 278216
rect 123302 278148 123336 278154
rect 123302 278120 123336 278148
rect 123302 278080 123336 278082
rect 123302 278048 123336 278080
rect 123302 277978 123336 278010
rect 123302 277976 123336 277978
rect 123302 277910 123336 277938
rect 123302 277904 123336 277910
rect 123302 277842 123336 277866
rect 123302 277832 123336 277842
rect 122439 277711 122461 277745
rect 122461 277711 122473 277745
rect 122511 277711 122529 277745
rect 122529 277711 122545 277745
rect 122583 277711 122597 277745
rect 122597 277711 122617 277745
rect 122655 277711 122665 277745
rect 122665 277711 122689 277745
rect 122727 277711 122733 277745
rect 122733 277711 122761 277745
rect 122799 277711 122801 277745
rect 122801 277711 122833 277745
rect 122871 277711 122903 277745
rect 122903 277711 122905 277745
rect 122943 277711 122971 277745
rect 122971 277711 122977 277745
rect 123015 277711 123039 277745
rect 123039 277711 123049 277745
rect 123087 277711 123107 277745
rect 123107 277711 123121 277745
rect 123159 277711 123175 277745
rect 123175 277711 123193 277745
rect 123231 277711 123243 277745
rect 123243 277711 123265 277745
rect 122439 277547 122459 277581
rect 122459 277547 122473 277581
rect 122511 277547 122527 277581
rect 122527 277547 122545 277581
rect 122583 277547 122595 277581
rect 122595 277547 122617 277581
rect 122655 277547 122663 277581
rect 122663 277547 122689 277581
rect 122727 277547 122731 277581
rect 122731 277547 122761 277581
rect 122799 277547 122833 277581
rect 122871 277547 122901 277581
rect 122901 277547 122905 277581
rect 122943 277547 122969 277581
rect 122969 277547 122977 277581
rect 123015 277547 123037 277581
rect 123037 277547 123049 277581
rect 123087 277547 123105 277581
rect 123105 277547 123121 277581
rect 123159 277547 123173 277581
rect 123173 277547 123193 277581
rect 122370 277433 122404 277467
rect 123228 277433 123262 277467
rect 122439 277319 122459 277353
rect 122459 277319 122473 277353
rect 122511 277319 122527 277353
rect 122527 277319 122545 277353
rect 122583 277319 122595 277353
rect 122595 277319 122617 277353
rect 122655 277319 122663 277353
rect 122663 277319 122689 277353
rect 122727 277319 122731 277353
rect 122731 277319 122761 277353
rect 122799 277319 122833 277353
rect 122871 277319 122901 277353
rect 122901 277319 122905 277353
rect 122943 277319 122969 277353
rect 122969 277319 122977 277353
rect 123015 277319 123037 277353
rect 123037 277319 123049 277353
rect 123087 277319 123105 277353
rect 123105 277319 123121 277353
rect 123159 277319 123173 277353
rect 123173 277319 123193 277353
rect 123700 278127 123712 278161
rect 123712 278127 123734 278161
rect 123772 278127 123780 278161
rect 123780 278127 123806 278161
rect 123844 278127 123848 278161
rect 123848 278127 123878 278161
rect 123916 278127 123950 278161
rect 123988 278127 124018 278161
rect 124018 278127 124022 278161
rect 124060 278127 124086 278161
rect 124086 278127 124094 278161
rect 124132 278127 124154 278161
rect 124154 278127 124166 278161
rect 123610 278026 123644 278042
rect 123610 278008 123644 278026
rect 123610 277958 123644 277970
rect 123610 277936 123644 277958
rect 123610 277890 123644 277898
rect 123610 277864 123644 277890
rect 123610 277822 123644 277826
rect 123610 277792 123644 277822
rect 123610 277720 123644 277754
rect 123610 277652 123644 277682
rect 123610 277648 123644 277652
rect 123610 277584 123644 277610
rect 123610 277576 123644 277584
rect 123610 277516 123644 277538
rect 123610 277504 123644 277516
rect 123610 277448 123644 277466
rect 123610 277432 123644 277448
rect 124222 278026 124256 278042
rect 124222 278008 124256 278026
rect 124222 277958 124256 277970
rect 124222 277936 124256 277958
rect 124222 277890 124256 277898
rect 124222 277864 124256 277890
rect 124222 277822 124256 277826
rect 124222 277792 124256 277822
rect 124222 277720 124256 277754
rect 124222 277652 124256 277682
rect 124222 277648 124256 277652
rect 124222 277584 124256 277610
rect 124222 277576 124256 277584
rect 124222 277516 124256 277538
rect 124222 277504 124256 277516
rect 124222 277448 124256 277466
rect 124222 277432 124256 277448
rect 123700 277313 123712 277347
rect 123712 277313 123734 277347
rect 123772 277313 123780 277347
rect 123780 277313 123806 277347
rect 123844 277313 123848 277347
rect 123848 277313 123878 277347
rect 123916 277313 123950 277347
rect 123988 277313 124018 277347
rect 124018 277313 124022 277347
rect 124060 277313 124086 277347
rect 124086 277313 124094 277347
rect 124132 277313 124154 277347
rect 124154 277313 124166 277347
rect 123771 276904 123877 277010
rect 122470 276715 122472 276749
rect 122472 276715 122504 276749
rect 122542 276715 122574 276749
rect 122574 276715 122576 276749
rect 122614 276715 122642 276749
rect 122642 276715 122648 276749
rect 122686 276715 122710 276749
rect 122710 276715 122720 276749
rect 122758 276715 122778 276749
rect 122778 276715 122792 276749
rect 122830 276715 122846 276749
rect 122846 276715 122864 276749
rect 122902 276715 122914 276749
rect 122914 276715 122936 276749
rect 122974 276715 122982 276749
rect 122982 276715 123008 276749
rect 123046 276715 123050 276749
rect 123050 276715 123080 276749
rect 123118 276715 123152 276749
rect 123190 276715 123220 276749
rect 123220 276715 123224 276749
rect 123262 276715 123288 276749
rect 123288 276715 123296 276749
rect 123334 276715 123356 276749
rect 123356 276715 123368 276749
rect 123406 276715 123424 276749
rect 123424 276715 123440 276749
rect 123478 276715 123492 276749
rect 123492 276715 123512 276749
rect 123550 276715 123560 276749
rect 123560 276715 123584 276749
rect 123622 276715 123628 276749
rect 123628 276715 123656 276749
rect 123694 276715 123696 276749
rect 123696 276715 123728 276749
rect 123766 276715 123798 276749
rect 123798 276715 123800 276749
rect 122392 276631 122426 276633
rect 122392 276599 122426 276631
rect 122392 276529 122426 276561
rect 122392 276527 122426 276529
rect 123844 276631 123878 276633
rect 123844 276599 123878 276631
rect 123844 276529 123878 276561
rect 123844 276527 123878 276529
rect 122470 276411 122472 276445
rect 122472 276411 122504 276445
rect 122542 276411 122574 276445
rect 122574 276411 122576 276445
rect 122614 276411 122642 276445
rect 122642 276411 122648 276445
rect 122686 276411 122710 276445
rect 122710 276411 122720 276445
rect 122758 276411 122778 276445
rect 122778 276411 122792 276445
rect 122830 276411 122846 276445
rect 122846 276411 122864 276445
rect 122902 276411 122914 276445
rect 122914 276411 122936 276445
rect 122974 276411 122982 276445
rect 122982 276411 123008 276445
rect 123046 276411 123050 276445
rect 123050 276411 123080 276445
rect 123118 276411 123152 276445
rect 123190 276411 123220 276445
rect 123220 276411 123224 276445
rect 123262 276411 123288 276445
rect 123288 276411 123296 276445
rect 123334 276411 123356 276445
rect 123356 276411 123368 276445
rect 123406 276411 123424 276445
rect 123424 276411 123440 276445
rect 123478 276411 123492 276445
rect 123492 276411 123512 276445
rect 123550 276411 123560 276445
rect 123560 276411 123584 276445
rect 123622 276411 123628 276445
rect 123628 276411 123656 276445
rect 123694 276411 123696 276445
rect 123696 276411 123728 276445
rect 123766 276411 123798 276445
rect 123798 276411 123800 276445
rect 122137 276078 122171 276112
rect 122209 276078 122243 276112
rect 122281 276078 122315 276112
rect 122353 276078 122387 276112
rect 124490 276015 124524 276049
rect 122505 275823 122513 275857
rect 122513 275823 122539 275857
rect 122577 275823 122581 275857
rect 122581 275823 122611 275857
rect 122649 275823 122683 275857
rect 122721 275823 122751 275857
rect 122751 275823 122755 275857
rect 122793 275823 122819 275857
rect 122819 275823 122827 275857
rect 123141 275823 123149 275857
rect 123149 275823 123175 275857
rect 123213 275823 123217 275857
rect 123217 275823 123247 275857
rect 123285 275823 123319 275857
rect 123357 275823 123387 275857
rect 123387 275823 123391 275857
rect 123429 275823 123455 275857
rect 123455 275823 123463 275857
rect 123777 275823 123785 275857
rect 123785 275823 123811 275857
rect 123849 275823 123853 275857
rect 123853 275823 123883 275857
rect 123921 275823 123955 275857
rect 123993 275823 124023 275857
rect 124023 275823 124027 275857
rect 124065 275823 124091 275857
rect 124091 275823 124099 275857
rect 124413 275823 124421 275857
rect 124421 275823 124447 275857
rect 124485 275823 124489 275857
rect 124489 275823 124519 275857
rect 124557 275823 124591 275857
rect 124629 275823 124659 275857
rect 124659 275823 124663 275857
rect 124701 275823 124727 275857
rect 124727 275823 124735 275857
rect 122385 275744 122419 275778
rect 122913 275744 122947 275778
rect 123021 275744 123055 275778
rect 123549 275744 123583 275778
rect 123657 275744 123691 275778
rect 124185 275744 124219 275778
rect 124293 275744 124327 275778
rect 124821 275744 124855 275778
rect 122505 275665 122513 275699
rect 122513 275665 122539 275699
rect 122577 275665 122581 275699
rect 122581 275665 122611 275699
rect 122649 275665 122683 275699
rect 122721 275665 122751 275699
rect 122751 275665 122755 275699
rect 122793 275665 122819 275699
rect 122819 275665 122827 275699
rect 123141 275665 123149 275699
rect 123149 275665 123175 275699
rect 123213 275665 123217 275699
rect 123217 275665 123247 275699
rect 123285 275665 123319 275699
rect 123357 275665 123387 275699
rect 123387 275665 123391 275699
rect 123429 275665 123455 275699
rect 123455 275665 123463 275699
rect 123777 275665 123785 275699
rect 123785 275665 123811 275699
rect 123849 275665 123853 275699
rect 123853 275665 123883 275699
rect 123921 275665 123955 275699
rect 123993 275665 124023 275699
rect 124023 275665 124027 275699
rect 124065 275665 124091 275699
rect 124091 275665 124099 275699
rect 124413 275665 124421 275699
rect 124421 275665 124447 275699
rect 124485 275665 124489 275699
rect 124489 275665 124519 275699
rect 124557 275665 124591 275699
rect 124629 275665 124659 275699
rect 124659 275665 124663 275699
rect 124701 275665 124727 275699
rect 124727 275665 124735 275699
rect 123246 275190 123424 275368
rect 121168 274968 121176 275002
rect 121176 274968 121202 275002
rect 121240 274968 121244 275002
rect 121244 274968 121274 275002
rect 121312 274968 121346 275002
rect 121384 274968 121414 275002
rect 121414 274968 121418 275002
rect 121456 274968 121482 275002
rect 121482 274968 121490 275002
rect 121168 274812 121176 274846
rect 121176 274812 121202 274846
rect 121240 274812 121244 274846
rect 121244 274812 121274 274846
rect 121312 274812 121346 274846
rect 121384 274812 121414 274846
rect 121414 274812 121418 274846
rect 121456 274812 121482 274846
rect 121482 274812 121490 274846
rect 121083 274736 121117 274748
rect 121083 274714 121117 274736
rect 121083 274668 121117 274676
rect 121083 274642 121117 274668
rect 121083 274600 121117 274604
rect 121083 274570 121117 274600
rect 120841 274498 120875 274532
rect 121083 274498 121117 274532
rect 120841 274430 120875 274460
rect 120841 274426 120875 274430
rect 120841 274362 120875 274388
rect 120841 274354 120875 274362
rect 120841 274294 120875 274316
rect 120841 274282 120875 274294
rect 121083 274430 121117 274460
rect 121083 274426 121117 274430
rect 121083 274362 121117 274388
rect 121083 274354 121117 274362
rect 121083 274294 121117 274316
rect 121083 274282 121117 274294
rect 121541 274736 121575 274748
rect 121541 274714 121575 274736
rect 121541 274668 121575 274676
rect 121541 274642 121575 274668
rect 121541 274600 121575 274604
rect 121541 274570 121575 274600
rect 121541 274498 121575 274532
rect 121541 274430 121575 274460
rect 121541 274426 121575 274430
rect 121541 274362 121575 274388
rect 121541 274354 121575 274362
rect 121541 274294 121575 274316
rect 121541 274282 121575 274294
rect 123003 274900 123027 274934
rect 123027 274900 123037 274934
rect 123075 274900 123095 274934
rect 123095 274900 123109 274934
rect 123147 274900 123163 274934
rect 123163 274900 123181 274934
rect 123219 274900 123231 274934
rect 123231 274900 123253 274934
rect 123291 274900 123299 274934
rect 123299 274900 123325 274934
rect 123363 274900 123367 274934
rect 123367 274900 123397 274934
rect 123435 274900 123469 274934
rect 123507 274900 123537 274934
rect 123537 274900 123541 274934
rect 123579 274900 123605 274934
rect 123605 274900 123613 274934
rect 123651 274900 123673 274934
rect 123673 274900 123685 274934
rect 123723 274900 123741 274934
rect 123741 274900 123757 274934
rect 123795 274900 123809 274934
rect 123809 274900 123829 274934
rect 123867 274900 123877 274934
rect 123877 274900 123901 274934
rect 122906 274813 122940 274815
rect 122906 274781 122940 274813
rect 122906 274711 122940 274743
rect 122906 274709 122940 274711
rect 123964 274813 123998 274815
rect 123964 274781 123998 274813
rect 123964 274711 123998 274743
rect 123964 274709 123998 274711
rect 123003 274590 123027 274624
rect 123027 274590 123037 274624
rect 123075 274590 123095 274624
rect 123095 274590 123109 274624
rect 123147 274590 123163 274624
rect 123163 274590 123181 274624
rect 123219 274590 123231 274624
rect 123231 274590 123253 274624
rect 123291 274590 123299 274624
rect 123299 274590 123325 274624
rect 123363 274590 123367 274624
rect 123367 274590 123397 274624
rect 123435 274590 123469 274624
rect 123507 274590 123537 274624
rect 123537 274590 123541 274624
rect 123579 274590 123605 274624
rect 123605 274590 123613 274624
rect 123651 274590 123673 274624
rect 123673 274590 123685 274624
rect 123723 274590 123741 274624
rect 123741 274590 123757 274624
rect 123795 274590 123809 274624
rect 123809 274590 123829 274624
rect 123867 274590 123877 274624
rect 123877 274590 123901 274624
rect 122324 274316 122326 274350
rect 122326 274316 122358 274350
rect 122396 274316 122428 274350
rect 122428 274316 122430 274350
rect 122740 274316 122742 274350
rect 122742 274316 122774 274350
rect 122812 274316 122844 274350
rect 122844 274316 122846 274350
rect 123534 274409 123568 274443
rect 123606 274409 123640 274443
rect 123156 274316 123158 274350
rect 123158 274316 123190 274350
rect 123228 274316 123260 274350
rect 123260 274316 123262 274350
rect 123572 274316 123574 274350
rect 123574 274316 123606 274350
rect 123644 274316 123676 274350
rect 123676 274316 123678 274350
rect 123988 274316 123990 274350
rect 123990 274316 124022 274350
rect 124060 274316 124092 274350
rect 124092 274316 124094 274350
rect 120468 274184 120476 274218
rect 120476 274184 120502 274218
rect 120540 274184 120544 274218
rect 120544 274184 120574 274218
rect 120612 274184 120646 274218
rect 120684 274184 120714 274218
rect 120714 274184 120718 274218
rect 120756 274184 120782 274218
rect 120782 274184 120790 274218
rect 121168 274184 121176 274218
rect 121176 274184 121202 274218
rect 121240 274184 121244 274218
rect 121244 274184 121274 274218
rect 121312 274184 121346 274218
rect 121384 274184 121414 274218
rect 121414 274184 121418 274218
rect 121456 274184 121482 274218
rect 121482 274184 121490 274218
rect 120468 274028 120476 274062
rect 120476 274028 120502 274062
rect 120540 274028 120544 274062
rect 120544 274028 120574 274062
rect 120612 274028 120646 274062
rect 120684 274028 120714 274062
rect 120714 274028 120718 274062
rect 120756 274028 120782 274062
rect 120782 274028 120790 274062
rect 121168 274028 121176 274062
rect 121176 274028 121202 274062
rect 121240 274028 121244 274062
rect 121244 274028 121274 274062
rect 121312 274028 121346 274062
rect 121384 274028 121414 274062
rect 121414 274028 121418 274062
rect 121456 274028 121482 274062
rect 121482 274028 121490 274062
rect 120383 273952 120417 273964
rect 120383 273930 120417 273952
rect 120383 273884 120417 273892
rect 120383 273858 120417 273884
rect 120383 273816 120417 273820
rect 120383 273786 120417 273816
rect 120383 273714 120417 273748
rect 120383 273646 120417 273676
rect 120383 273642 120417 273646
rect 120383 273578 120417 273604
rect 120383 273570 120417 273578
rect 120383 273510 120417 273532
rect 120383 273498 120417 273510
rect 120841 273952 120875 273964
rect 120841 273930 120875 273952
rect 120841 273884 120875 273892
rect 120841 273858 120875 273884
rect 120841 273816 120875 273820
rect 120841 273786 120875 273816
rect 121083 273952 121117 273964
rect 121083 273930 121117 273952
rect 121083 273884 121117 273892
rect 121083 273858 121117 273884
rect 121083 273816 121117 273820
rect 121083 273786 121117 273816
rect 120841 273714 120875 273748
rect 120972 273707 121006 273741
rect 121083 273714 121117 273748
rect 120841 273646 120875 273676
rect 120841 273642 120875 273646
rect 120841 273578 120875 273604
rect 120841 273570 120875 273578
rect 120841 273510 120875 273532
rect 120841 273498 120875 273510
rect 121083 273646 121117 273676
rect 121083 273642 121117 273646
rect 121083 273578 121117 273604
rect 121083 273570 121117 273578
rect 121083 273510 121117 273532
rect 121083 273498 121117 273510
rect 121541 273952 121575 273964
rect 121541 273930 121575 273952
rect 121541 273884 121575 273892
rect 121541 273858 121575 273884
rect 121541 273816 121575 273820
rect 121541 273786 121575 273816
rect 121541 273714 121575 273748
rect 121541 273646 121575 273676
rect 121541 273642 121575 273646
rect 121541 273578 121575 273604
rect 121541 273570 121575 273578
rect 121541 273510 121575 273532
rect 121541 273498 121575 273510
rect 122231 274249 122265 274261
rect 122231 274227 122265 274249
rect 122231 274181 122265 274189
rect 122231 274155 122265 274181
rect 122231 274113 122265 274117
rect 122231 274083 122265 274113
rect 122231 274011 122265 274045
rect 122231 273943 122265 273973
rect 122231 273939 122265 273943
rect 122231 273875 122265 273901
rect 122231 273867 122265 273875
rect 122231 273807 122265 273829
rect 122231 273795 122265 273807
rect 122489 274249 122523 274261
rect 122489 274227 122523 274249
rect 122489 274181 122523 274189
rect 122489 274155 122523 274181
rect 122489 274113 122523 274117
rect 122489 274083 122523 274113
rect 122489 274011 122523 274045
rect 122489 273943 122523 273973
rect 122489 273939 122523 273943
rect 122489 273875 122523 273901
rect 122489 273867 122523 273875
rect 122489 273807 122523 273829
rect 122489 273795 122523 273807
rect 122647 274249 122681 274261
rect 122647 274227 122681 274249
rect 122647 274181 122681 274189
rect 122647 274155 122681 274181
rect 122647 274113 122681 274117
rect 122647 274083 122681 274113
rect 122647 274011 122681 274045
rect 122647 273943 122681 273973
rect 122647 273939 122681 273943
rect 122647 273875 122681 273901
rect 122647 273867 122681 273875
rect 122647 273807 122681 273829
rect 122647 273795 122681 273807
rect 122905 274249 122939 274261
rect 122905 274227 122939 274249
rect 122905 274181 122939 274189
rect 122905 274155 122939 274181
rect 122905 274113 122939 274117
rect 122905 274083 122939 274113
rect 122905 274011 122939 274045
rect 122905 273943 122939 273973
rect 122905 273939 122939 273943
rect 122905 273875 122939 273901
rect 122905 273867 122939 273875
rect 122905 273807 122939 273829
rect 122905 273795 122939 273807
rect 123063 274249 123097 274261
rect 123063 274227 123097 274249
rect 123063 274181 123097 274189
rect 123063 274155 123097 274181
rect 123063 274113 123097 274117
rect 123063 274083 123097 274113
rect 123063 274011 123097 274045
rect 123063 273943 123097 273973
rect 123063 273939 123097 273943
rect 123063 273875 123097 273901
rect 123063 273867 123097 273875
rect 123063 273807 123097 273829
rect 123063 273795 123097 273807
rect 123321 274249 123355 274261
rect 123321 274227 123355 274249
rect 123321 274181 123355 274189
rect 123321 274155 123355 274181
rect 123321 274113 123355 274117
rect 123321 274083 123355 274113
rect 123321 274011 123355 274045
rect 123321 273943 123355 273973
rect 123321 273939 123355 273943
rect 123321 273875 123355 273901
rect 123321 273867 123355 273875
rect 123321 273807 123355 273829
rect 123321 273795 123355 273807
rect 123479 274249 123513 274261
rect 123479 274227 123513 274249
rect 123479 274181 123513 274189
rect 123479 274155 123513 274181
rect 123479 274113 123513 274117
rect 123479 274083 123513 274113
rect 123479 274011 123513 274045
rect 123479 273943 123513 273973
rect 123479 273939 123513 273943
rect 123479 273875 123513 273901
rect 123479 273867 123513 273875
rect 123479 273807 123513 273829
rect 123479 273795 123513 273807
rect 123737 274249 123771 274261
rect 123737 274227 123771 274249
rect 123737 274181 123771 274189
rect 123737 274155 123771 274181
rect 123737 274113 123771 274117
rect 123737 274083 123771 274113
rect 123737 274011 123771 274045
rect 123737 273943 123771 273973
rect 123737 273939 123771 273943
rect 123737 273875 123771 273901
rect 123737 273867 123771 273875
rect 123737 273807 123771 273829
rect 123737 273795 123771 273807
rect 123895 274249 123929 274261
rect 123895 274227 123929 274249
rect 123895 274181 123929 274189
rect 123895 274155 123929 274181
rect 123895 274113 123929 274117
rect 123895 274083 123929 274113
rect 123895 274011 123929 274045
rect 123895 273943 123929 273973
rect 123895 273939 123929 273943
rect 123895 273875 123929 273901
rect 123895 273867 123929 273875
rect 123895 273807 123929 273829
rect 123895 273795 123929 273807
rect 124153 274249 124187 274261
rect 124153 274227 124187 274249
rect 124153 274181 124187 274189
rect 124153 274155 124187 274181
rect 124153 274113 124187 274117
rect 124153 274083 124187 274113
rect 124153 274011 124187 274045
rect 124153 273943 124187 273973
rect 124153 273939 124187 273943
rect 124153 273875 124187 273901
rect 124153 273867 124187 273875
rect 124153 273807 124187 273829
rect 124153 273795 124187 273807
rect 124404 274316 124406 274350
rect 124406 274316 124438 274350
rect 124476 274316 124508 274350
rect 124508 274316 124510 274350
rect 124311 274249 124345 274261
rect 124311 274227 124345 274249
rect 124311 274181 124345 274189
rect 124311 274155 124345 274181
rect 124311 274113 124345 274117
rect 124311 274083 124345 274113
rect 124311 274011 124345 274045
rect 124311 273943 124345 273973
rect 124311 273939 124345 273943
rect 124311 273875 124345 273901
rect 124311 273867 124345 273875
rect 124311 273807 124345 273829
rect 124311 273795 124345 273807
rect 124569 274249 124603 274261
rect 124569 274227 124603 274249
rect 124569 274181 124603 274189
rect 124569 274155 124603 274181
rect 124569 274113 124603 274117
rect 124569 274083 124603 274113
rect 124569 274011 124603 274045
rect 124569 273943 124603 273973
rect 124569 273939 124603 273943
rect 124569 273875 124603 273901
rect 124569 273867 124603 273875
rect 124569 273807 124603 273829
rect 124569 273795 124603 273807
rect 122324 273706 122326 273740
rect 122326 273706 122358 273740
rect 122396 273706 122428 273740
rect 122428 273706 122430 273740
rect 122740 273706 122742 273740
rect 122742 273706 122774 273740
rect 122812 273706 122844 273740
rect 122844 273706 122846 273740
rect 123156 273706 123158 273740
rect 123158 273706 123190 273740
rect 123228 273706 123260 273740
rect 123260 273706 123262 273740
rect 123572 273706 123574 273740
rect 123574 273706 123606 273740
rect 123644 273706 123676 273740
rect 123676 273706 123678 273740
rect 123988 273706 123990 273740
rect 123990 273706 124022 273740
rect 124060 273706 124092 273740
rect 124092 273706 124094 273740
rect 124404 273706 124406 273740
rect 124406 273706 124438 273740
rect 124476 273706 124508 273740
rect 124508 273706 124510 273740
rect 120468 273400 120476 273434
rect 120476 273400 120502 273434
rect 120540 273400 120544 273434
rect 120544 273400 120574 273434
rect 120612 273400 120646 273434
rect 120684 273400 120714 273434
rect 120714 273400 120718 273434
rect 120756 273400 120782 273434
rect 120782 273400 120790 273434
rect 121168 273400 121176 273434
rect 121176 273400 121202 273434
rect 121240 273400 121244 273434
rect 121244 273400 121274 273434
rect 121312 273400 121346 273434
rect 121384 273400 121414 273434
rect 121414 273400 121418 273434
rect 121456 273400 121482 273434
rect 121482 273400 121490 273434
rect 120468 273244 120476 273278
rect 120476 273244 120502 273278
rect 120540 273244 120544 273278
rect 120544 273244 120574 273278
rect 120612 273244 120646 273278
rect 120684 273244 120714 273278
rect 120714 273244 120718 273278
rect 120756 273244 120782 273278
rect 120782 273244 120790 273278
rect 121168 273244 121176 273278
rect 121176 273244 121202 273278
rect 121240 273244 121244 273278
rect 121244 273244 121274 273278
rect 121312 273244 121346 273278
rect 121384 273244 121414 273278
rect 121414 273244 121418 273278
rect 121456 273244 121482 273278
rect 121482 273244 121490 273278
rect 120383 273168 120417 273180
rect 120383 273146 120417 273168
rect 120383 273100 120417 273108
rect 120383 273074 120417 273100
rect 120383 273032 120417 273036
rect 120383 273002 120417 273032
rect 120383 272930 120417 272964
rect 120383 272862 120417 272892
rect 120383 272858 120417 272862
rect 120383 272794 120417 272820
rect 120383 272786 120417 272794
rect 120383 272726 120417 272748
rect 120383 272714 120417 272726
rect 120841 273168 120875 273180
rect 120841 273146 120875 273168
rect 120841 273100 120875 273108
rect 120841 273074 120875 273100
rect 120841 273032 120875 273036
rect 120841 273002 120875 273032
rect 120841 272930 120875 272964
rect 120841 272862 120875 272892
rect 120841 272858 120875 272862
rect 120841 272794 120875 272820
rect 120841 272786 120875 272794
rect 120841 272726 120875 272748
rect 120841 272714 120875 272726
rect 121083 273168 121117 273180
rect 121083 273146 121117 273168
rect 121083 273100 121117 273108
rect 121083 273074 121117 273100
rect 121083 273032 121117 273036
rect 121083 273002 121117 273032
rect 121083 272930 121117 272964
rect 121083 272862 121117 272892
rect 121083 272858 121117 272862
rect 121083 272794 121117 272820
rect 121083 272786 121117 272794
rect 121083 272726 121117 272748
rect 121083 272714 121117 272726
rect 121541 273168 121575 273180
rect 121541 273146 121575 273168
rect 121541 273100 121575 273108
rect 121541 273074 121575 273100
rect 121541 273032 121575 273036
rect 121541 273002 121575 273032
rect 121541 272930 121575 272964
rect 121541 272862 121575 272892
rect 121541 272858 121575 272862
rect 121541 272794 121575 272820
rect 121541 272786 121575 272794
rect 121541 272726 121575 272748
rect 121541 272714 121575 272726
rect 120468 272616 120476 272650
rect 120476 272616 120502 272650
rect 120540 272616 120544 272650
rect 120544 272616 120574 272650
rect 120612 272616 120646 272650
rect 120684 272616 120714 272650
rect 120714 272616 120718 272650
rect 120756 272616 120782 272650
rect 120782 272616 120790 272650
rect 121168 272616 121176 272650
rect 121176 272616 121202 272650
rect 121240 272616 121244 272650
rect 121244 272616 121274 272650
rect 121312 272616 121346 272650
rect 121384 272616 121414 272650
rect 121414 272616 121418 272650
rect 121456 272616 121482 272650
rect 121482 272616 121490 272650
rect 122164 272860 122172 272894
rect 122172 272860 122198 272894
rect 122236 272860 122240 272894
rect 122240 272860 122270 272894
rect 122308 272860 122342 272894
rect 122380 272860 122410 272894
rect 122410 272860 122414 272894
rect 122452 272860 122478 272894
rect 122478 272860 122486 272894
rect 122079 272746 122113 272780
rect 122537 272746 122571 272780
rect 122164 272632 122172 272666
rect 122172 272632 122198 272666
rect 122236 272632 122240 272666
rect 122240 272632 122270 272666
rect 122308 272632 122342 272666
rect 122380 272632 122410 272666
rect 122410 272632 122414 272666
rect 122452 272632 122478 272666
rect 122478 272632 122486 272666
rect 122864 272860 122872 272894
rect 122872 272860 122898 272894
rect 122936 272860 122940 272894
rect 122940 272860 122970 272894
rect 123008 272860 123042 272894
rect 123080 272860 123110 272894
rect 123110 272860 123114 272894
rect 123152 272860 123178 272894
rect 123178 272860 123186 272894
rect 122779 272746 122813 272780
rect 123237 272746 123271 272780
rect 122864 272632 122872 272666
rect 122872 272632 122898 272666
rect 122936 272632 122940 272666
rect 122940 272632 122970 272666
rect 123008 272632 123042 272666
rect 123080 272632 123110 272666
rect 123110 272632 123114 272666
rect 123152 272632 123178 272666
rect 123178 272632 123186 272666
rect 123382 272591 123416 272625
rect 123382 272519 123416 272553
rect 120468 272460 120476 272494
rect 120476 272460 120502 272494
rect 120540 272460 120544 272494
rect 120544 272460 120574 272494
rect 120612 272460 120646 272494
rect 120684 272460 120714 272494
rect 120714 272460 120718 272494
rect 120756 272460 120782 272494
rect 120782 272460 120790 272494
rect 121168 272460 121176 272494
rect 121176 272460 121202 272494
rect 121240 272460 121244 272494
rect 121244 272460 121274 272494
rect 121312 272460 121346 272494
rect 121384 272460 121414 272494
rect 121414 272460 121418 272494
rect 121456 272460 121482 272494
rect 121482 272460 121490 272494
rect 122164 272476 122172 272510
rect 122172 272476 122198 272510
rect 122236 272476 122240 272510
rect 122240 272476 122270 272510
rect 122308 272476 122342 272510
rect 122380 272476 122410 272510
rect 122410 272476 122414 272510
rect 122452 272476 122478 272510
rect 122478 272476 122486 272510
rect 122864 272476 122872 272510
rect 122872 272476 122898 272510
rect 122936 272476 122940 272510
rect 122940 272476 122970 272510
rect 123008 272476 123042 272510
rect 123080 272476 123110 272510
rect 123110 272476 123114 272510
rect 123152 272476 123178 272510
rect 123178 272476 123186 272510
rect 120383 272384 120417 272396
rect 120383 272362 120417 272384
rect 120383 272316 120417 272324
rect 120383 272290 120417 272316
rect 120383 272248 120417 272252
rect 120383 272218 120417 272248
rect 120383 272146 120417 272180
rect 120383 272078 120417 272108
rect 120383 272074 120417 272078
rect 120383 272010 120417 272036
rect 120383 272002 120417 272010
rect 120383 271942 120417 271964
rect 120383 271930 120417 271942
rect 120841 272384 120875 272396
rect 120841 272362 120875 272384
rect 120841 272316 120875 272324
rect 120841 272290 120875 272316
rect 120841 272248 120875 272252
rect 120841 272218 120875 272248
rect 120841 272146 120875 272180
rect 120841 272078 120875 272108
rect 120841 272074 120875 272078
rect 120841 272010 120875 272036
rect 120841 272002 120875 272010
rect 120841 271942 120875 271964
rect 120841 271930 120875 271942
rect 121083 272384 121117 272396
rect 121083 272362 121117 272384
rect 121083 272316 121117 272324
rect 121083 272290 121117 272316
rect 121083 272248 121117 272252
rect 121083 272218 121117 272248
rect 121083 272146 121117 272180
rect 121083 272078 121117 272108
rect 121083 272074 121117 272078
rect 121083 272010 121117 272036
rect 121083 272002 121117 272010
rect 121083 271942 121117 271964
rect 121083 271930 121117 271942
rect 121541 272384 121575 272396
rect 121541 272362 121575 272384
rect 121541 272316 121575 272324
rect 121541 272290 121575 272316
rect 121541 272248 121575 272252
rect 121541 272218 121575 272248
rect 121541 272146 121575 272180
rect 121541 272078 121575 272108
rect 121541 272074 121575 272078
rect 121541 272010 121575 272036
rect 121541 272002 121575 272010
rect 121541 271942 121575 271964
rect 121541 271930 121575 271942
rect 123382 272447 123416 272481
rect 122079 272400 122113 272412
rect 122079 272378 122113 272400
rect 122079 272332 122113 272340
rect 122079 272306 122113 272332
rect 122079 272264 122113 272268
rect 122079 272234 122113 272264
rect 122079 272162 122113 272196
rect 122079 272094 122113 272124
rect 122079 272090 122113 272094
rect 122079 272026 122113 272052
rect 122079 272018 122113 272026
rect 122079 271958 122113 271980
rect 122079 271946 122113 271958
rect 122537 272400 122571 272412
rect 122537 272378 122571 272400
rect 122537 272332 122571 272340
rect 122537 272306 122571 272332
rect 122537 272264 122571 272268
rect 122537 272234 122571 272264
rect 122779 272400 122813 272412
rect 122779 272378 122813 272400
rect 122779 272332 122813 272340
rect 122779 272306 122813 272332
rect 122779 272264 122813 272268
rect 122779 272234 122813 272264
rect 122537 272162 122571 272196
rect 122665 272165 122699 272199
rect 122779 272162 122813 272196
rect 122537 272094 122571 272124
rect 122537 272090 122571 272094
rect 122537 272026 122571 272052
rect 122537 272018 122571 272026
rect 122537 271958 122571 271980
rect 122537 271946 122571 271958
rect 122779 272094 122813 272124
rect 122779 272090 122813 272094
rect 122779 272026 122813 272052
rect 122779 272018 122813 272026
rect 122779 271958 122813 271980
rect 122779 271946 122813 271958
rect 123237 272400 123271 272412
rect 123237 272378 123271 272400
rect 123237 272332 123271 272340
rect 123237 272306 123271 272332
rect 123237 272264 123271 272268
rect 123237 272234 123271 272264
rect 123237 272162 123271 272196
rect 123237 272094 123271 272124
rect 123237 272090 123271 272094
rect 123237 272026 123271 272052
rect 123237 272018 123271 272026
rect 123237 271958 123271 271980
rect 123237 271946 123271 271958
rect 120468 271832 120476 271866
rect 120476 271832 120502 271866
rect 120540 271832 120544 271866
rect 120544 271832 120574 271866
rect 120612 271832 120646 271866
rect 120684 271832 120714 271866
rect 120714 271832 120718 271866
rect 120756 271832 120782 271866
rect 120782 271832 120790 271866
rect 121168 271832 121176 271866
rect 121176 271832 121202 271866
rect 121240 271832 121244 271866
rect 121244 271832 121274 271866
rect 121312 271832 121346 271866
rect 121384 271832 121414 271866
rect 121414 271832 121418 271866
rect 121456 271832 121482 271866
rect 121482 271832 121490 271866
rect 122164 271848 122172 271882
rect 122172 271848 122198 271882
rect 122236 271848 122240 271882
rect 122240 271848 122270 271882
rect 122308 271848 122342 271882
rect 122380 271848 122410 271882
rect 122410 271848 122414 271882
rect 122452 271848 122478 271882
rect 122478 271848 122486 271882
rect 122864 271848 122872 271882
rect 122872 271848 122898 271882
rect 122936 271848 122940 271882
rect 122940 271848 122970 271882
rect 123008 271848 123042 271882
rect 123080 271848 123110 271882
rect 123110 271848 123114 271882
rect 123152 271848 123178 271882
rect 123178 271848 123186 271882
rect 120468 271676 120476 271710
rect 120476 271676 120502 271710
rect 120540 271676 120544 271710
rect 120544 271676 120574 271710
rect 120612 271676 120646 271710
rect 120684 271676 120714 271710
rect 120714 271676 120718 271710
rect 120756 271676 120782 271710
rect 120782 271676 120790 271710
rect 121168 271676 121176 271710
rect 121176 271676 121202 271710
rect 121240 271676 121244 271710
rect 121244 271676 121274 271710
rect 121312 271676 121346 271710
rect 121384 271676 121414 271710
rect 121414 271676 121418 271710
rect 121456 271676 121482 271710
rect 121482 271676 121490 271710
rect 122164 271692 122172 271726
rect 122172 271692 122198 271726
rect 122236 271692 122240 271726
rect 122240 271692 122270 271726
rect 122308 271692 122342 271726
rect 122380 271692 122410 271726
rect 122410 271692 122414 271726
rect 122452 271692 122478 271726
rect 122478 271692 122486 271726
rect 122864 271692 122872 271726
rect 122872 271692 122898 271726
rect 122936 271692 122940 271726
rect 122940 271692 122970 271726
rect 123008 271692 123042 271726
rect 123080 271692 123110 271726
rect 123110 271692 123114 271726
rect 123152 271692 123178 271726
rect 123178 271692 123186 271726
rect 120383 271600 120417 271612
rect 120383 271578 120417 271600
rect 120383 271532 120417 271540
rect 120383 271506 120417 271532
rect 120383 271464 120417 271468
rect 120383 271434 120417 271464
rect 120383 271362 120417 271396
rect 120383 271294 120417 271324
rect 120383 271290 120417 271294
rect 120383 271226 120417 271252
rect 120383 271218 120417 271226
rect 120383 271158 120417 271180
rect 120383 271146 120417 271158
rect 120841 271600 120875 271612
rect 120841 271578 120875 271600
rect 120841 271532 120875 271540
rect 120841 271506 120875 271532
rect 120841 271464 120875 271468
rect 120841 271434 120875 271464
rect 120841 271362 120875 271396
rect 120841 271294 120875 271324
rect 120841 271290 120875 271294
rect 120841 271226 120875 271252
rect 120841 271218 120875 271226
rect 120841 271158 120875 271180
rect 120841 271146 120875 271158
rect 121083 271600 121117 271612
rect 121083 271578 121117 271600
rect 121083 271532 121117 271540
rect 121083 271506 121117 271532
rect 121083 271464 121117 271468
rect 121083 271434 121117 271464
rect 121083 271362 121117 271396
rect 121083 271294 121117 271324
rect 121083 271290 121117 271294
rect 121083 271226 121117 271252
rect 121083 271218 121117 271226
rect 121083 271158 121117 271180
rect 121083 271146 121117 271158
rect 121541 271600 121575 271612
rect 121541 271578 121575 271600
rect 121541 271532 121575 271540
rect 121541 271506 121575 271532
rect 121541 271464 121575 271468
rect 121541 271434 121575 271464
rect 121541 271362 121575 271396
rect 121541 271294 121575 271324
rect 121541 271290 121575 271294
rect 121541 271226 121575 271252
rect 121541 271218 121575 271226
rect 121541 271158 121575 271180
rect 121541 271146 121575 271158
rect 122079 271616 122113 271628
rect 122079 271594 122113 271616
rect 122079 271548 122113 271556
rect 122079 271522 122113 271548
rect 122079 271480 122113 271484
rect 122079 271450 122113 271480
rect 122079 271378 122113 271412
rect 122079 271310 122113 271340
rect 122079 271306 122113 271310
rect 122079 271242 122113 271268
rect 122079 271234 122113 271242
rect 122079 271174 122113 271196
rect 122079 271162 122113 271174
rect 122537 271616 122571 271628
rect 122537 271594 122571 271616
rect 122537 271548 122571 271556
rect 122537 271522 122571 271548
rect 122537 271480 122571 271484
rect 122537 271450 122571 271480
rect 122779 271616 122813 271628
rect 122779 271594 122813 271616
rect 122779 271548 122813 271556
rect 122779 271522 122813 271548
rect 122779 271480 122813 271484
rect 122779 271450 122813 271480
rect 122537 271378 122571 271412
rect 122779 271378 122813 271412
rect 122537 271310 122571 271340
rect 122537 271306 122571 271310
rect 122537 271242 122571 271268
rect 122537 271234 122571 271242
rect 122537 271174 122571 271196
rect 122537 271162 122571 271174
rect 120468 271048 120476 271082
rect 120476 271048 120502 271082
rect 120540 271048 120544 271082
rect 120544 271048 120574 271082
rect 120612 271048 120646 271082
rect 120684 271048 120714 271082
rect 120714 271048 120718 271082
rect 120756 271048 120782 271082
rect 120782 271048 120790 271082
rect 121168 271048 121176 271082
rect 121176 271048 121202 271082
rect 121240 271048 121244 271082
rect 121244 271048 121274 271082
rect 121312 271048 121346 271082
rect 121384 271048 121414 271082
rect 121414 271048 121418 271082
rect 121456 271048 121482 271082
rect 121482 271048 121490 271082
rect 122164 271064 122172 271098
rect 122172 271064 122198 271098
rect 122236 271064 122240 271098
rect 122240 271064 122270 271098
rect 122308 271064 122342 271098
rect 122380 271064 122410 271098
rect 122410 271064 122414 271098
rect 122452 271064 122478 271098
rect 122478 271064 122486 271098
rect 120468 270892 120476 270926
rect 120476 270892 120502 270926
rect 120540 270892 120544 270926
rect 120544 270892 120574 270926
rect 120612 270892 120646 270926
rect 120684 270892 120714 270926
rect 120714 270892 120718 270926
rect 120756 270892 120782 270926
rect 120782 270892 120790 270926
rect 121168 270892 121176 270926
rect 121176 270892 121202 270926
rect 121240 270892 121244 270926
rect 121244 270892 121274 270926
rect 121312 270892 121346 270926
rect 121384 270892 121414 270926
rect 121414 270892 121418 270926
rect 121456 270892 121482 270926
rect 121482 270892 121490 270926
rect 122164 270908 122172 270942
rect 122172 270908 122198 270942
rect 122236 270908 122240 270942
rect 122240 270908 122270 270942
rect 122308 270908 122342 270942
rect 122380 270908 122410 270942
rect 122410 270908 122414 270942
rect 122452 270908 122478 270942
rect 122478 270908 122486 270942
rect 120383 270816 120417 270828
rect 120383 270794 120417 270816
rect 120383 270748 120417 270756
rect 120383 270722 120417 270748
rect 120383 270680 120417 270684
rect 120383 270650 120417 270680
rect 120383 270578 120417 270612
rect 120383 270510 120417 270540
rect 120383 270506 120417 270510
rect 120383 270442 120417 270468
rect 120383 270434 120417 270442
rect 120383 270374 120417 270396
rect 120383 270362 120417 270374
rect 120841 270816 120875 270828
rect 120841 270794 120875 270816
rect 120841 270748 120875 270756
rect 120841 270722 120875 270748
rect 120841 270680 120875 270684
rect 120841 270650 120875 270680
rect 120841 270578 120875 270612
rect 120841 270510 120875 270540
rect 120841 270506 120875 270510
rect 120841 270442 120875 270468
rect 120841 270434 120875 270442
rect 120841 270374 120875 270396
rect 120841 270362 120875 270374
rect 121083 270816 121117 270828
rect 121083 270794 121117 270816
rect 121083 270748 121117 270756
rect 121083 270722 121117 270748
rect 121083 270680 121117 270684
rect 121083 270650 121117 270680
rect 121083 270578 121117 270612
rect 121083 270510 121117 270540
rect 121083 270506 121117 270510
rect 121083 270442 121117 270468
rect 121083 270434 121117 270442
rect 121083 270374 121117 270396
rect 121083 270362 121117 270374
rect 121541 270816 121575 270828
rect 121541 270794 121575 270816
rect 121541 270748 121575 270756
rect 121541 270722 121575 270748
rect 121541 270680 121575 270684
rect 121541 270650 121575 270680
rect 121541 270578 121575 270612
rect 121541 270510 121575 270540
rect 121541 270506 121575 270510
rect 121541 270442 121575 270468
rect 121541 270434 121575 270442
rect 121541 270374 121575 270396
rect 121541 270362 121575 270374
rect 122079 270832 122113 270844
rect 122079 270810 122113 270832
rect 122079 270764 122113 270772
rect 122079 270738 122113 270764
rect 122079 270696 122113 270700
rect 122079 270666 122113 270696
rect 122079 270594 122113 270628
rect 122079 270526 122113 270556
rect 122079 270522 122113 270526
rect 122079 270458 122113 270484
rect 122079 270450 122113 270458
rect 122079 270390 122113 270412
rect 122079 270378 122113 270390
rect 122537 270832 122571 270844
rect 122537 270810 122571 270832
rect 122537 270764 122571 270772
rect 122537 270738 122571 270764
rect 122537 270696 122571 270700
rect 122537 270666 122571 270696
rect 122779 271310 122813 271340
rect 122779 271306 122813 271310
rect 122779 271242 122813 271268
rect 122779 271234 122813 271242
rect 122779 271174 122813 271196
rect 122779 271162 122813 271174
rect 123237 271616 123271 271628
rect 123237 271594 123271 271616
rect 123237 271548 123271 271556
rect 123237 271522 123271 271548
rect 123237 271480 123271 271484
rect 123237 271450 123271 271480
rect 123237 271378 123271 271412
rect 123237 271310 123271 271340
rect 123237 271306 123271 271310
rect 123237 271242 123271 271268
rect 123237 271234 123271 271242
rect 123237 271174 123271 271196
rect 123237 271162 123271 271174
rect 122864 271064 122872 271098
rect 122872 271064 122898 271098
rect 122936 271064 122940 271098
rect 122940 271064 122970 271098
rect 123008 271064 123042 271098
rect 123080 271064 123110 271098
rect 123110 271064 123114 271098
rect 123152 271064 123178 271098
rect 123178 271064 123186 271098
rect 122864 270908 122872 270942
rect 122872 270908 122898 270942
rect 122936 270908 122940 270942
rect 122940 270908 122970 270942
rect 123008 270908 123042 270942
rect 123080 270908 123110 270942
rect 123110 270908 123114 270942
rect 123152 270908 123178 270942
rect 123178 270908 123186 270942
rect 122779 270832 122813 270844
rect 122779 270810 122813 270832
rect 122779 270764 122813 270772
rect 122779 270738 122813 270764
rect 122779 270696 122813 270700
rect 122779 270666 122813 270696
rect 122537 270594 122571 270628
rect 122779 270594 122813 270628
rect 122537 270526 122571 270556
rect 122537 270522 122571 270526
rect 122537 270458 122571 270484
rect 122537 270450 122571 270458
rect 122537 270390 122571 270412
rect 122537 270378 122571 270390
rect 122779 270526 122813 270556
rect 122779 270522 122813 270526
rect 122779 270458 122813 270484
rect 122779 270450 122813 270458
rect 122779 270390 122813 270412
rect 122779 270378 122813 270390
rect 123237 270832 123271 270844
rect 123237 270810 123271 270832
rect 123237 270764 123271 270772
rect 123237 270738 123271 270764
rect 123237 270696 123271 270700
rect 123237 270666 123271 270696
rect 123237 270594 123271 270628
rect 123237 270526 123271 270556
rect 123237 270522 123271 270526
rect 123237 270458 123271 270484
rect 123237 270450 123271 270458
rect 123237 270390 123271 270412
rect 123237 270378 123271 270390
rect 120468 270264 120476 270298
rect 120476 270264 120502 270298
rect 120540 270264 120544 270298
rect 120544 270264 120574 270298
rect 120612 270264 120646 270298
rect 120684 270264 120714 270298
rect 120714 270264 120718 270298
rect 120756 270264 120782 270298
rect 120782 270264 120790 270298
rect 121168 270264 121176 270298
rect 121176 270264 121202 270298
rect 121240 270264 121244 270298
rect 121244 270264 121274 270298
rect 121312 270264 121346 270298
rect 121384 270264 121414 270298
rect 121414 270264 121418 270298
rect 121456 270264 121482 270298
rect 121482 270264 121490 270298
rect 122164 270280 122172 270314
rect 122172 270280 122198 270314
rect 122236 270280 122240 270314
rect 122240 270280 122270 270314
rect 122308 270280 122342 270314
rect 122380 270280 122410 270314
rect 122410 270280 122414 270314
rect 122452 270280 122478 270314
rect 122478 270280 122486 270314
rect 122864 270280 122872 270314
rect 122872 270280 122898 270314
rect 122936 270280 122940 270314
rect 122940 270280 122970 270314
rect 123008 270280 123042 270314
rect 123080 270280 123110 270314
rect 123110 270280 123114 270314
rect 123152 270280 123178 270314
rect 123178 270280 123186 270314
rect 120468 270108 120476 270142
rect 120476 270108 120502 270142
rect 120540 270108 120544 270142
rect 120544 270108 120574 270142
rect 120612 270108 120646 270142
rect 120684 270108 120714 270142
rect 120714 270108 120718 270142
rect 120756 270108 120782 270142
rect 120782 270108 120790 270142
rect 121168 270108 121176 270142
rect 121176 270108 121202 270142
rect 121240 270108 121244 270142
rect 121244 270108 121274 270142
rect 121312 270108 121346 270142
rect 121384 270108 121414 270142
rect 121414 270108 121418 270142
rect 121456 270108 121482 270142
rect 121482 270108 121490 270142
rect 122164 270124 122172 270158
rect 122172 270124 122198 270158
rect 122236 270124 122240 270158
rect 122240 270124 122270 270158
rect 122308 270124 122342 270158
rect 122380 270124 122410 270158
rect 122410 270124 122414 270158
rect 122452 270124 122478 270158
rect 122478 270124 122486 270158
rect 122864 270124 122872 270158
rect 122872 270124 122898 270158
rect 122936 270124 122940 270158
rect 122940 270124 122970 270158
rect 123008 270124 123042 270158
rect 123080 270124 123110 270158
rect 123110 270124 123114 270158
rect 123152 270124 123178 270158
rect 123178 270124 123186 270158
rect 120383 270032 120417 270044
rect 120383 270010 120417 270032
rect 120383 269964 120417 269972
rect 120383 269938 120417 269964
rect 120383 269896 120417 269900
rect 120383 269866 120417 269896
rect 120383 269794 120417 269828
rect 120383 269726 120417 269756
rect 120383 269722 120417 269726
rect 120383 269658 120417 269684
rect 120383 269650 120417 269658
rect 120383 269590 120417 269612
rect 120383 269578 120417 269590
rect 120841 270032 120875 270044
rect 120841 270010 120875 270032
rect 120841 269964 120875 269972
rect 120841 269938 120875 269964
rect 120841 269896 120875 269900
rect 120841 269866 120875 269896
rect 120841 269794 120875 269828
rect 120841 269726 120875 269756
rect 120841 269722 120875 269726
rect 120841 269658 120875 269684
rect 120841 269650 120875 269658
rect 120841 269590 120875 269612
rect 120841 269578 120875 269590
rect 121083 270032 121117 270044
rect 121083 270010 121117 270032
rect 121083 269964 121117 269972
rect 121083 269938 121117 269964
rect 121083 269896 121117 269900
rect 121083 269866 121117 269896
rect 121083 269794 121117 269828
rect 121083 269726 121117 269756
rect 121083 269722 121117 269726
rect 121083 269658 121117 269684
rect 121083 269650 121117 269658
rect 121083 269590 121117 269612
rect 121083 269578 121117 269590
rect 121541 270032 121575 270044
rect 121541 270010 121575 270032
rect 121541 269964 121575 269972
rect 121541 269938 121575 269964
rect 121541 269896 121575 269900
rect 121541 269866 121575 269896
rect 121541 269794 121575 269828
rect 121541 269726 121575 269756
rect 121541 269722 121575 269726
rect 121541 269658 121575 269684
rect 121541 269650 121575 269658
rect 121541 269590 121575 269612
rect 121541 269578 121575 269590
rect 122079 270048 122113 270060
rect 122079 270026 122113 270048
rect 122079 269980 122113 269988
rect 122079 269954 122113 269980
rect 122079 269912 122113 269916
rect 122079 269882 122113 269912
rect 122079 269810 122113 269844
rect 122079 269742 122113 269772
rect 122079 269738 122113 269742
rect 122079 269674 122113 269700
rect 122079 269666 122113 269674
rect 122079 269606 122113 269628
rect 122079 269594 122113 269606
rect 122537 270048 122571 270060
rect 122537 270026 122571 270048
rect 122537 269980 122571 269988
rect 122537 269954 122571 269980
rect 122537 269912 122571 269916
rect 122537 269882 122571 269912
rect 122779 270048 122813 270060
rect 122779 270026 122813 270048
rect 122779 269980 122813 269988
rect 122779 269954 122813 269980
rect 122779 269912 122813 269916
rect 122779 269882 122813 269912
rect 122537 269810 122571 269844
rect 122668 269803 122702 269837
rect 122779 269810 122813 269844
rect 122537 269742 122571 269772
rect 122537 269738 122571 269742
rect 122537 269674 122571 269700
rect 122537 269666 122571 269674
rect 122537 269606 122571 269628
rect 122537 269594 122571 269606
rect 122779 269742 122813 269772
rect 122779 269738 122813 269742
rect 122779 269674 122813 269700
rect 122779 269666 122813 269674
rect 122779 269606 122813 269628
rect 122779 269594 122813 269606
rect 123237 270048 123271 270060
rect 123237 270026 123271 270048
rect 123237 269980 123271 269988
rect 123237 269954 123271 269980
rect 123237 269912 123271 269916
rect 123237 269882 123271 269912
rect 123237 269810 123271 269844
rect 123237 269742 123271 269772
rect 123237 269738 123271 269742
rect 123237 269674 123271 269700
rect 123237 269666 123271 269674
rect 123237 269606 123271 269628
rect 123237 269594 123271 269606
rect 120468 269480 120476 269514
rect 120476 269480 120502 269514
rect 120540 269480 120544 269514
rect 120544 269480 120574 269514
rect 120612 269480 120646 269514
rect 120684 269480 120714 269514
rect 120714 269480 120718 269514
rect 120756 269480 120782 269514
rect 120782 269480 120790 269514
rect 121168 269480 121176 269514
rect 121176 269480 121202 269514
rect 121240 269480 121244 269514
rect 121244 269480 121274 269514
rect 121312 269480 121346 269514
rect 121384 269480 121414 269514
rect 121414 269480 121418 269514
rect 121456 269480 121482 269514
rect 121482 269480 121490 269514
rect 122164 269496 122172 269530
rect 122172 269496 122198 269530
rect 122236 269496 122240 269530
rect 122240 269496 122270 269530
rect 122308 269496 122342 269530
rect 122380 269496 122410 269530
rect 122410 269496 122414 269530
rect 122452 269496 122478 269530
rect 122478 269496 122486 269530
rect 122864 269496 122872 269530
rect 122872 269496 122898 269530
rect 122936 269496 122940 269530
rect 122940 269496 122970 269530
rect 123008 269496 123042 269530
rect 123080 269496 123110 269530
rect 123110 269496 123114 269530
rect 123152 269496 123178 269530
rect 123178 269496 123186 269530
rect 120468 269324 120476 269358
rect 120476 269324 120502 269358
rect 120540 269324 120544 269358
rect 120544 269324 120574 269358
rect 120612 269324 120646 269358
rect 120684 269324 120714 269358
rect 120714 269324 120718 269358
rect 120756 269324 120782 269358
rect 120782 269324 120790 269358
rect 121168 269324 121176 269358
rect 121176 269324 121202 269358
rect 121240 269324 121244 269358
rect 121244 269324 121274 269358
rect 121312 269324 121346 269358
rect 121384 269324 121414 269358
rect 121414 269324 121418 269358
rect 121456 269324 121482 269358
rect 121482 269324 121490 269358
rect 120383 269210 120417 269244
rect 120841 269210 120875 269244
rect 120468 269096 120476 269130
rect 120476 269096 120502 269130
rect 120540 269096 120544 269130
rect 120544 269096 120574 269130
rect 120612 269096 120646 269130
rect 120684 269096 120714 269130
rect 120714 269096 120718 269130
rect 120756 269096 120782 269130
rect 120782 269096 120790 269130
rect 121083 269210 121117 269244
rect 121541 269210 121575 269244
rect 121168 269096 121176 269130
rect 121176 269096 121202 269130
rect 121240 269096 121244 269130
rect 121244 269096 121274 269130
rect 121312 269096 121346 269130
rect 121384 269096 121414 269130
rect 121414 269096 121418 269130
rect 121456 269096 121482 269130
rect 121482 269096 121490 269130
rect 122164 269340 122172 269374
rect 122172 269340 122198 269374
rect 122236 269340 122240 269374
rect 122240 269340 122270 269374
rect 122308 269340 122342 269374
rect 122380 269340 122410 269374
rect 122410 269340 122414 269374
rect 122452 269340 122478 269374
rect 122478 269340 122486 269374
rect 122079 269226 122113 269260
rect 122537 269226 122571 269260
rect 122164 269112 122172 269146
rect 122172 269112 122198 269146
rect 122236 269112 122240 269146
rect 122240 269112 122270 269146
rect 122308 269112 122342 269146
rect 122380 269112 122410 269146
rect 122410 269112 122414 269146
rect 122452 269112 122478 269146
rect 122478 269112 122486 269146
rect 122864 269340 122872 269374
rect 122872 269340 122898 269374
rect 122936 269340 122940 269374
rect 122940 269340 122970 269374
rect 123008 269340 123042 269374
rect 123080 269340 123110 269374
rect 123110 269340 123114 269374
rect 123152 269340 123178 269374
rect 123178 269340 123186 269374
rect 122779 269226 122813 269260
rect 123237 269226 123271 269260
rect 122864 269112 122872 269146
rect 122872 269112 122898 269146
rect 122936 269112 122940 269146
rect 122940 269112 122970 269146
rect 123008 269112 123042 269146
rect 123080 269112 123110 269146
rect 123110 269112 123114 269146
rect 123152 269112 123178 269146
rect 123178 269112 123186 269146
rect 124209 272532 124221 272566
rect 124221 272532 124243 272566
rect 124281 272532 124289 272566
rect 124289 272532 124315 272566
rect 124353 272532 124357 272566
rect 124357 272532 124387 272566
rect 124425 272532 124459 272566
rect 124497 272532 124527 272566
rect 124527 272532 124531 272566
rect 124569 272532 124595 272566
rect 124595 272532 124603 272566
rect 124641 272532 124663 272566
rect 124663 272532 124675 272566
rect 124120 272471 124154 272473
rect 124120 272439 124154 272471
rect 124120 272369 124154 272401
rect 124120 272367 124154 272369
rect 124730 272471 124764 272473
rect 124730 272439 124764 272471
rect 124730 272369 124764 272401
rect 124730 272367 124764 272369
rect 124209 272274 124221 272308
rect 124221 272274 124243 272308
rect 124281 272274 124289 272308
rect 124289 272274 124315 272308
rect 124353 272274 124357 272308
rect 124357 272274 124387 272308
rect 124425 272274 124459 272308
rect 124497 272274 124527 272308
rect 124527 272274 124531 272308
rect 124569 272274 124595 272308
rect 124595 272274 124603 272308
rect 124641 272274 124663 272308
rect 124663 272274 124675 272308
rect 124209 272116 124221 272150
rect 124221 272116 124243 272150
rect 124281 272116 124289 272150
rect 124289 272116 124315 272150
rect 124353 272116 124357 272150
rect 124357 272116 124387 272150
rect 124425 272116 124459 272150
rect 124497 272116 124527 272150
rect 124527 272116 124531 272150
rect 124569 272116 124595 272150
rect 124595 272116 124603 272150
rect 124641 272116 124663 272150
rect 124663 272116 124675 272150
rect 124120 272055 124154 272057
rect 124120 272023 124154 272055
rect 124120 271953 124154 271985
rect 124120 271951 124154 271953
rect 124730 272055 124764 272057
rect 124730 272023 124764 272055
rect 124730 271953 124764 271985
rect 124730 271951 124764 271953
rect 124209 271858 124221 271892
rect 124221 271858 124243 271892
rect 124281 271858 124289 271892
rect 124289 271858 124315 271892
rect 124353 271858 124357 271892
rect 124357 271858 124387 271892
rect 124425 271858 124459 271892
rect 124497 271858 124527 271892
rect 124527 271858 124531 271892
rect 124569 271858 124595 271892
rect 124595 271858 124603 271892
rect 124641 271858 124663 271892
rect 124663 271858 124675 271892
rect 124209 271700 124221 271734
rect 124221 271700 124243 271734
rect 124281 271700 124289 271734
rect 124289 271700 124315 271734
rect 124353 271700 124357 271734
rect 124357 271700 124387 271734
rect 124425 271700 124459 271734
rect 124497 271700 124527 271734
rect 124527 271700 124531 271734
rect 124569 271700 124595 271734
rect 124595 271700 124603 271734
rect 124641 271700 124663 271734
rect 124663 271700 124675 271734
rect 124120 271639 124154 271641
rect 124120 271607 124154 271639
rect 124120 271537 124154 271569
rect 124120 271535 124154 271537
rect 124730 271639 124764 271641
rect 124730 271607 124764 271639
rect 124730 271537 124764 271569
rect 124730 271535 124764 271537
rect 124209 271442 124221 271476
rect 124221 271442 124243 271476
rect 124281 271442 124289 271476
rect 124289 271442 124315 271476
rect 124353 271442 124357 271476
rect 124357 271442 124387 271476
rect 124425 271442 124459 271476
rect 124497 271442 124527 271476
rect 124527 271442 124531 271476
rect 124569 271442 124595 271476
rect 124595 271442 124603 271476
rect 124641 271442 124663 271476
rect 124663 271442 124675 271476
rect 124209 271284 124221 271318
rect 124221 271284 124243 271318
rect 124281 271284 124289 271318
rect 124289 271284 124315 271318
rect 124353 271284 124357 271318
rect 124357 271284 124387 271318
rect 124425 271284 124459 271318
rect 124497 271284 124527 271318
rect 124527 271284 124531 271318
rect 124569 271284 124595 271318
rect 124595 271284 124603 271318
rect 124641 271284 124663 271318
rect 124663 271284 124675 271318
rect 124120 271223 124154 271225
rect 124120 271191 124154 271223
rect 124120 271121 124154 271153
rect 124120 271119 124154 271121
rect 124730 271223 124764 271225
rect 124730 271191 124764 271223
rect 124730 271121 124764 271153
rect 124730 271119 124764 271121
rect 124209 271026 124221 271060
rect 124221 271026 124243 271060
rect 124281 271026 124289 271060
rect 124289 271026 124315 271060
rect 124353 271026 124357 271060
rect 124357 271026 124387 271060
rect 124425 271026 124459 271060
rect 124497 271026 124527 271060
rect 124527 271026 124531 271060
rect 124569 271026 124595 271060
rect 124595 271026 124603 271060
rect 124641 271026 124663 271060
rect 124663 271026 124675 271060
rect 124209 270868 124221 270902
rect 124221 270868 124243 270902
rect 124281 270868 124289 270902
rect 124289 270868 124315 270902
rect 124353 270868 124357 270902
rect 124357 270868 124387 270902
rect 124425 270868 124459 270902
rect 124497 270868 124527 270902
rect 124527 270868 124531 270902
rect 124569 270868 124595 270902
rect 124595 270868 124603 270902
rect 124641 270868 124663 270902
rect 124663 270868 124675 270902
rect 124120 270807 124154 270809
rect 124120 270775 124154 270807
rect 124120 270705 124154 270737
rect 124120 270703 124154 270705
rect 124730 270807 124764 270809
rect 124730 270775 124764 270807
rect 124730 270705 124764 270737
rect 124730 270703 124764 270705
rect 124209 270610 124221 270644
rect 124221 270610 124243 270644
rect 124281 270610 124289 270644
rect 124289 270610 124315 270644
rect 124353 270610 124357 270644
rect 124357 270610 124387 270644
rect 124425 270610 124459 270644
rect 124497 270610 124527 270644
rect 124527 270610 124531 270644
rect 124569 270610 124595 270644
rect 124595 270610 124603 270644
rect 124641 270610 124663 270644
rect 124663 270610 124675 270644
rect 124209 270452 124221 270486
rect 124221 270452 124243 270486
rect 124281 270452 124289 270486
rect 124289 270452 124315 270486
rect 124353 270452 124357 270486
rect 124357 270452 124387 270486
rect 124425 270452 124459 270486
rect 124497 270452 124527 270486
rect 124527 270452 124531 270486
rect 124569 270452 124595 270486
rect 124595 270452 124603 270486
rect 124641 270452 124663 270486
rect 124663 270452 124675 270486
rect 124120 270391 124154 270393
rect 124120 270359 124154 270391
rect 124120 270289 124154 270321
rect 124120 270287 124154 270289
rect 124730 270391 124764 270393
rect 124730 270359 124764 270391
rect 124730 270289 124764 270321
rect 124730 270287 124764 270289
rect 124209 270194 124221 270228
rect 124221 270194 124243 270228
rect 124281 270194 124289 270228
rect 124289 270194 124315 270228
rect 124353 270194 124357 270228
rect 124357 270194 124387 270228
rect 124425 270194 124459 270228
rect 124497 270194 124527 270228
rect 124527 270194 124531 270228
rect 124569 270194 124595 270228
rect 124595 270194 124603 270228
rect 124641 270194 124663 270228
rect 124663 270194 124675 270228
rect 124209 270036 124221 270070
rect 124221 270036 124243 270070
rect 124281 270036 124289 270070
rect 124289 270036 124315 270070
rect 124353 270036 124357 270070
rect 124357 270036 124387 270070
rect 124425 270036 124459 270070
rect 124497 270036 124527 270070
rect 124527 270036 124531 270070
rect 124569 270036 124595 270070
rect 124595 270036 124603 270070
rect 124641 270036 124663 270070
rect 124663 270036 124675 270070
rect 124120 269975 124154 269977
rect 124120 269943 124154 269975
rect 124120 269873 124154 269905
rect 124120 269871 124154 269873
rect 124730 269975 124764 269977
rect 124730 269943 124764 269975
rect 124730 269873 124764 269905
rect 124730 269871 124764 269873
rect 124209 269778 124221 269812
rect 124221 269778 124243 269812
rect 124281 269778 124289 269812
rect 124289 269778 124315 269812
rect 124353 269778 124357 269812
rect 124357 269778 124387 269812
rect 124425 269778 124459 269812
rect 124497 269778 124527 269812
rect 124527 269778 124531 269812
rect 124569 269778 124595 269812
rect 124595 269778 124603 269812
rect 124641 269778 124663 269812
rect 124663 269778 124675 269812
rect 124209 269620 124221 269654
rect 124221 269620 124243 269654
rect 124281 269620 124289 269654
rect 124289 269620 124315 269654
rect 124353 269620 124357 269654
rect 124357 269620 124387 269654
rect 124425 269620 124459 269654
rect 124497 269620 124527 269654
rect 124527 269620 124531 269654
rect 124569 269620 124595 269654
rect 124595 269620 124603 269654
rect 124641 269620 124663 269654
rect 124663 269620 124675 269654
rect 124120 269559 124154 269561
rect 124120 269527 124154 269559
rect 124120 269457 124154 269489
rect 124120 269455 124154 269457
rect 124730 269559 124764 269561
rect 124730 269527 124764 269559
rect 124730 269457 124764 269489
rect 124730 269455 124764 269457
rect 124209 269362 124221 269396
rect 124221 269362 124243 269396
rect 124281 269362 124289 269396
rect 124289 269362 124315 269396
rect 124353 269362 124357 269396
rect 124357 269362 124387 269396
rect 124425 269362 124459 269396
rect 124497 269362 124527 269396
rect 124527 269362 124531 269396
rect 124569 269362 124595 269396
rect 124595 269362 124603 269396
rect 124641 269362 124663 269396
rect 124663 269362 124675 269396
rect 125825 268349 128019 275151
<< metal1 >>
rect 105796 283650 113672 283895
rect 105796 282446 106167 283650
rect 113387 282909 113672 283650
rect 113387 282446 125337 282909
rect 105796 282251 125337 282446
rect 102098 281628 103259 281810
rect 102098 280872 102272 281628
rect 103092 281274 103259 281628
rect 103092 281095 108300 281274
rect 103092 280872 103259 281095
rect 108146 281064 108300 281095
rect 108146 280949 108295 281064
rect 102098 280720 103259 280872
rect 106361 280885 106485 280891
rect 106361 280851 106406 280885
rect 106440 280851 106485 280885
rect 106361 280845 106485 280851
rect 106761 280885 109685 280949
rect 106761 280851 106806 280885
rect 106840 280879 107206 280885
rect 106840 280851 106885 280879
rect 106761 280845 106885 280851
rect 107161 280851 107206 280879
rect 107240 280879 107606 280885
rect 107240 280851 107285 280879
rect 107161 280845 107285 280851
rect 107561 280851 107606 280879
rect 107640 280879 108006 280885
rect 107640 280851 107685 280879
rect 107561 280845 107685 280851
rect 107961 280851 108006 280879
rect 108040 280879 108406 280885
rect 108040 280851 108085 280879
rect 107961 280845 108085 280851
rect 108196 280813 108255 280879
rect 108361 280851 108406 280879
rect 108440 280879 108806 280885
rect 108440 280851 108485 280879
rect 108361 280845 108485 280851
rect 108761 280851 108806 280879
rect 108840 280879 109206 280885
rect 108840 280851 108885 280879
rect 108761 280845 108885 280851
rect 109161 280851 109206 280879
rect 109240 280879 109606 280885
rect 109240 280851 109285 280879
rect 109161 280845 109285 280851
rect 109561 280851 109606 280879
rect 109640 280851 109685 280885
rect 109561 280845 109685 280851
rect 109961 280885 110085 280891
rect 109961 280851 110006 280885
rect 110040 280851 110085 280885
rect 109961 280845 110085 280851
rect 106305 280788 106351 280813
rect 106305 280754 106311 280788
rect 106345 280754 106351 280788
rect 106305 280716 106351 280754
rect 106305 280682 106311 280716
rect 106345 280682 106351 280716
rect 106305 280644 106351 280682
rect 106305 280610 106311 280644
rect 106345 280610 106351 280644
rect 106305 280572 106351 280610
rect 106305 280538 106311 280572
rect 106345 280538 106351 280572
rect 106305 280500 106351 280538
rect 106305 280466 106311 280500
rect 106345 280466 106351 280500
rect 106305 280428 106351 280466
rect 106305 280394 106311 280428
rect 106345 280394 106351 280428
rect 106305 280356 106351 280394
rect 106305 280322 106311 280356
rect 106345 280322 106351 280356
rect 106305 280284 106351 280322
rect 106305 280250 106311 280284
rect 106345 280250 106351 280284
rect 106305 280212 106351 280250
rect 106305 280178 106311 280212
rect 106345 280178 106351 280212
rect 106305 280140 106351 280178
rect 106305 280106 106311 280140
rect 106345 280106 106351 280140
rect 106305 280068 106351 280106
rect 106305 280034 106311 280068
rect 106345 280034 106351 280068
rect 106305 279996 106351 280034
rect 106305 279962 106311 279996
rect 106345 279962 106351 279996
rect 106305 279924 106351 279962
rect 106305 279890 106311 279924
rect 106345 279890 106351 279924
rect 106305 279852 106351 279890
rect 106305 279818 106311 279852
rect 106345 279818 106351 279852
rect 106305 279793 106351 279818
rect 106495 280788 106541 280813
rect 106495 280754 106501 280788
rect 106535 280754 106541 280788
rect 106495 280716 106541 280754
rect 106495 280682 106501 280716
rect 106535 280682 106541 280716
rect 106495 280644 106541 280682
rect 106495 280610 106501 280644
rect 106535 280610 106541 280644
rect 106495 280572 106541 280610
rect 106495 280538 106501 280572
rect 106535 280538 106541 280572
rect 106495 280500 106541 280538
rect 106495 280466 106501 280500
rect 106535 280466 106541 280500
rect 106495 280428 106541 280466
rect 106495 280394 106501 280428
rect 106535 280394 106541 280428
rect 106495 280356 106541 280394
rect 106495 280322 106501 280356
rect 106535 280322 106541 280356
rect 106495 280284 106541 280322
rect 106495 280250 106501 280284
rect 106535 280250 106541 280284
rect 106495 280212 106541 280250
rect 106495 280178 106501 280212
rect 106535 280178 106541 280212
rect 106495 280140 106541 280178
rect 106495 280106 106501 280140
rect 106535 280106 106541 280140
rect 106495 280068 106541 280106
rect 106495 280034 106501 280068
rect 106535 280034 106541 280068
rect 106495 279996 106541 280034
rect 106495 279962 106501 279996
rect 106535 279962 106541 279996
rect 106495 279924 106541 279962
rect 106495 279890 106501 279924
rect 106535 279890 106541 279924
rect 106495 279852 106541 279890
rect 106495 279818 106501 279852
rect 106535 279818 106541 279852
rect 106495 279793 106541 279818
rect 106705 280788 106751 280813
rect 106705 280754 106711 280788
rect 106745 280754 106751 280788
rect 106705 280716 106751 280754
rect 106705 280682 106711 280716
rect 106745 280682 106751 280716
rect 106705 280644 106751 280682
rect 106705 280610 106711 280644
rect 106745 280610 106751 280644
rect 106705 280572 106751 280610
rect 106705 280538 106711 280572
rect 106745 280538 106751 280572
rect 106705 280500 106751 280538
rect 106705 280466 106711 280500
rect 106745 280466 106751 280500
rect 106705 280428 106751 280466
rect 106705 280394 106711 280428
rect 106745 280394 106751 280428
rect 106705 280356 106751 280394
rect 106705 280322 106711 280356
rect 106745 280322 106751 280356
rect 106705 280284 106751 280322
rect 106705 280250 106711 280284
rect 106745 280250 106751 280284
rect 106705 280212 106751 280250
rect 106705 280178 106711 280212
rect 106745 280178 106751 280212
rect 106705 280140 106751 280178
rect 106705 280106 106711 280140
rect 106745 280106 106751 280140
rect 106705 280068 106751 280106
rect 106705 280034 106711 280068
rect 106745 280034 106751 280068
rect 106705 279996 106751 280034
rect 106705 279962 106711 279996
rect 106745 279962 106751 279996
rect 106705 279924 106751 279962
rect 106705 279890 106711 279924
rect 106745 279890 106751 279924
rect 106705 279852 106751 279890
rect 106705 279818 106711 279852
rect 106745 279818 106751 279852
rect 106705 279793 106751 279818
rect 106895 280788 106996 280813
rect 106895 280754 106901 280788
rect 106935 280754 106996 280788
rect 106895 280716 106996 280754
rect 106895 280682 106901 280716
rect 106935 280682 106996 280716
rect 106895 280644 106996 280682
rect 106895 280610 106901 280644
rect 106935 280610 106996 280644
rect 106895 280572 106996 280610
rect 106895 280538 106901 280572
rect 106935 280538 106996 280572
rect 106895 280500 106996 280538
rect 106895 280466 106901 280500
rect 106935 280466 106996 280500
rect 106895 280428 106996 280466
rect 106895 280394 106901 280428
rect 106935 280394 106996 280428
rect 106895 280356 106996 280394
rect 106895 280322 106901 280356
rect 106935 280322 106996 280356
rect 106895 280284 106996 280322
rect 106895 280250 106901 280284
rect 106935 280250 106996 280284
rect 106895 280212 106996 280250
rect 106895 280178 106901 280212
rect 106935 280178 106996 280212
rect 106895 280140 106996 280178
rect 106895 280106 106901 280140
rect 106935 280106 106996 280140
rect 106895 280068 106996 280106
rect 106895 280034 106901 280068
rect 106935 280034 106996 280068
rect 106895 279996 106996 280034
rect 106895 279962 106901 279996
rect 106935 279962 106996 279996
rect 106895 279924 106996 279962
rect 106895 279890 106901 279924
rect 106935 279890 106996 279924
rect 106895 279852 106996 279890
rect 106895 279818 106901 279852
rect 106935 279818 106996 279852
rect 106895 279793 106996 279818
rect 107105 280788 107151 280813
rect 107105 280754 107111 280788
rect 107145 280754 107151 280788
rect 107105 280716 107151 280754
rect 107105 280682 107111 280716
rect 107145 280682 107151 280716
rect 107105 280644 107151 280682
rect 107105 280610 107111 280644
rect 107145 280610 107151 280644
rect 107105 280572 107151 280610
rect 107105 280538 107111 280572
rect 107145 280538 107151 280572
rect 107105 280500 107151 280538
rect 107105 280466 107111 280500
rect 107145 280466 107151 280500
rect 107105 280428 107151 280466
rect 107105 280394 107111 280428
rect 107145 280394 107151 280428
rect 107105 280356 107151 280394
rect 107105 280322 107111 280356
rect 107145 280322 107151 280356
rect 107105 280284 107151 280322
rect 107105 280250 107111 280284
rect 107145 280250 107151 280284
rect 107105 280212 107151 280250
rect 107105 280178 107111 280212
rect 107145 280178 107151 280212
rect 107105 280140 107151 280178
rect 107105 280106 107111 280140
rect 107145 280106 107151 280140
rect 107105 280068 107151 280106
rect 107105 280034 107111 280068
rect 107145 280034 107151 280068
rect 107105 279996 107151 280034
rect 107105 279962 107111 279996
rect 107145 279962 107151 279996
rect 107105 279924 107151 279962
rect 107105 279890 107111 279924
rect 107145 279890 107151 279924
rect 107105 279852 107151 279890
rect 107105 279818 107111 279852
rect 107145 279818 107151 279852
rect 107105 279793 107151 279818
rect 107295 280788 107396 280813
rect 107295 280754 107301 280788
rect 107335 280754 107396 280788
rect 107295 280716 107396 280754
rect 107295 280682 107301 280716
rect 107335 280682 107396 280716
rect 107295 280644 107396 280682
rect 107295 280610 107301 280644
rect 107335 280610 107396 280644
rect 107295 280572 107396 280610
rect 107295 280538 107301 280572
rect 107335 280538 107396 280572
rect 107295 280500 107396 280538
rect 107295 280466 107301 280500
rect 107335 280466 107396 280500
rect 107295 280428 107396 280466
rect 107295 280394 107301 280428
rect 107335 280394 107396 280428
rect 107295 280356 107396 280394
rect 107295 280322 107301 280356
rect 107335 280322 107396 280356
rect 107295 280284 107396 280322
rect 107295 280250 107301 280284
rect 107335 280250 107396 280284
rect 107295 280212 107396 280250
rect 107295 280178 107301 280212
rect 107335 280178 107396 280212
rect 107295 280140 107396 280178
rect 107295 280106 107301 280140
rect 107335 280106 107396 280140
rect 107295 280068 107396 280106
rect 107295 280034 107301 280068
rect 107335 280034 107396 280068
rect 107295 279996 107396 280034
rect 107295 279962 107301 279996
rect 107335 279962 107396 279996
rect 107295 279924 107396 279962
rect 107295 279890 107301 279924
rect 107335 279890 107396 279924
rect 107295 279852 107396 279890
rect 107295 279818 107301 279852
rect 107335 279818 107396 279852
rect 107295 279793 107396 279818
rect 107505 280788 107551 280813
rect 107505 280754 107511 280788
rect 107545 280754 107551 280788
rect 107505 280716 107551 280754
rect 107505 280682 107511 280716
rect 107545 280682 107551 280716
rect 107505 280644 107551 280682
rect 107505 280610 107511 280644
rect 107545 280610 107551 280644
rect 107505 280572 107551 280610
rect 107505 280538 107511 280572
rect 107545 280538 107551 280572
rect 107505 280500 107551 280538
rect 107505 280466 107511 280500
rect 107545 280466 107551 280500
rect 107505 280428 107551 280466
rect 107505 280394 107511 280428
rect 107545 280394 107551 280428
rect 107505 280356 107551 280394
rect 107505 280322 107511 280356
rect 107545 280322 107551 280356
rect 107505 280284 107551 280322
rect 107505 280250 107511 280284
rect 107545 280250 107551 280284
rect 107505 280212 107551 280250
rect 107505 280178 107511 280212
rect 107545 280178 107551 280212
rect 107505 280140 107551 280178
rect 107505 280106 107511 280140
rect 107545 280106 107551 280140
rect 107505 280068 107551 280106
rect 107505 280034 107511 280068
rect 107545 280034 107551 280068
rect 107505 279996 107551 280034
rect 107505 279962 107511 279996
rect 107545 279962 107551 279996
rect 107505 279924 107551 279962
rect 107505 279890 107511 279924
rect 107545 279890 107551 279924
rect 107505 279852 107551 279890
rect 107505 279818 107511 279852
rect 107545 279818 107551 279852
rect 107505 279793 107551 279818
rect 107695 280788 107796 280813
rect 107695 280754 107701 280788
rect 107735 280754 107796 280788
rect 107695 280716 107796 280754
rect 107695 280682 107701 280716
rect 107735 280682 107796 280716
rect 107695 280644 107796 280682
rect 107695 280610 107701 280644
rect 107735 280610 107796 280644
rect 107695 280572 107796 280610
rect 107695 280538 107701 280572
rect 107735 280538 107796 280572
rect 107695 280500 107796 280538
rect 107695 280466 107701 280500
rect 107735 280466 107796 280500
rect 107695 280428 107796 280466
rect 107695 280394 107701 280428
rect 107735 280394 107796 280428
rect 107695 280356 107796 280394
rect 107695 280322 107701 280356
rect 107735 280322 107796 280356
rect 107695 280284 107796 280322
rect 107695 280250 107701 280284
rect 107735 280250 107796 280284
rect 107695 280212 107796 280250
rect 107695 280178 107701 280212
rect 107735 280178 107796 280212
rect 107695 280140 107796 280178
rect 107695 280106 107701 280140
rect 107735 280106 107796 280140
rect 107695 280068 107796 280106
rect 107695 280034 107701 280068
rect 107735 280034 107796 280068
rect 107695 279996 107796 280034
rect 107695 279962 107701 279996
rect 107735 279962 107796 279996
rect 107695 279924 107796 279962
rect 107695 279890 107701 279924
rect 107735 279890 107796 279924
rect 107695 279852 107796 279890
rect 107695 279818 107701 279852
rect 107735 279818 107796 279852
rect 107695 279793 107796 279818
rect 107905 280788 107951 280813
rect 107905 280754 107911 280788
rect 107945 280754 107951 280788
rect 107905 280716 107951 280754
rect 107905 280682 107911 280716
rect 107945 280682 107951 280716
rect 107905 280644 107951 280682
rect 107905 280610 107911 280644
rect 107945 280610 107951 280644
rect 107905 280572 107951 280610
rect 107905 280538 107911 280572
rect 107945 280538 107951 280572
rect 107905 280500 107951 280538
rect 107905 280466 107911 280500
rect 107945 280466 107951 280500
rect 107905 280428 107951 280466
rect 107905 280394 107911 280428
rect 107945 280394 107951 280428
rect 107905 280356 107951 280394
rect 107905 280322 107911 280356
rect 107945 280322 107951 280356
rect 107905 280284 107951 280322
rect 107905 280250 107911 280284
rect 107945 280250 107951 280284
rect 107905 280212 107951 280250
rect 107905 280178 107911 280212
rect 107945 280178 107951 280212
rect 107905 280140 107951 280178
rect 107905 280106 107911 280140
rect 107945 280106 107951 280140
rect 107905 280068 107951 280106
rect 107905 280034 107911 280068
rect 107945 280034 107951 280068
rect 107905 279996 107951 280034
rect 107905 279962 107911 279996
rect 107945 279962 107951 279996
rect 107905 279924 107951 279962
rect 107905 279890 107911 279924
rect 107945 279890 107951 279924
rect 107905 279852 107951 279890
rect 107905 279818 107911 279852
rect 107945 279818 107951 279852
rect 107905 279793 107951 279818
rect 108095 280788 108351 280813
rect 108095 280754 108101 280788
rect 108135 280754 108311 280788
rect 108345 280754 108351 280788
rect 108095 280716 108351 280754
rect 108095 280682 108101 280716
rect 108135 280682 108311 280716
rect 108345 280682 108351 280716
rect 108095 280644 108351 280682
rect 108095 280610 108101 280644
rect 108135 280610 108311 280644
rect 108345 280610 108351 280644
rect 108095 280572 108351 280610
rect 108095 280538 108101 280572
rect 108135 280538 108311 280572
rect 108345 280538 108351 280572
rect 108095 280500 108351 280538
rect 108095 280466 108101 280500
rect 108135 280466 108311 280500
rect 108345 280466 108351 280500
rect 108095 280428 108351 280466
rect 108095 280394 108101 280428
rect 108135 280394 108311 280428
rect 108345 280394 108351 280428
rect 108095 280356 108351 280394
rect 108095 280322 108101 280356
rect 108135 280322 108311 280356
rect 108345 280322 108351 280356
rect 108095 280284 108351 280322
rect 108095 280250 108101 280284
rect 108135 280250 108311 280284
rect 108345 280250 108351 280284
rect 108095 280212 108351 280250
rect 108095 280178 108101 280212
rect 108135 280178 108311 280212
rect 108345 280178 108351 280212
rect 108095 280140 108351 280178
rect 108095 280106 108101 280140
rect 108135 280106 108311 280140
rect 108345 280106 108351 280140
rect 108095 280068 108351 280106
rect 108095 280034 108101 280068
rect 108135 280034 108311 280068
rect 108345 280034 108351 280068
rect 108095 279996 108351 280034
rect 108095 279962 108101 279996
rect 108135 279962 108311 279996
rect 108345 279962 108351 279996
rect 108095 279924 108351 279962
rect 108095 279890 108101 279924
rect 108135 279890 108311 279924
rect 108345 279890 108351 279924
rect 108095 279852 108351 279890
rect 108095 279818 108101 279852
rect 108135 279818 108311 279852
rect 108345 279818 108351 279852
rect 108095 279793 108351 279818
rect 108495 280788 108541 280813
rect 108495 280754 108501 280788
rect 108535 280754 108541 280788
rect 108495 280716 108541 280754
rect 108495 280682 108501 280716
rect 108535 280682 108541 280716
rect 108495 280644 108541 280682
rect 108495 280610 108501 280644
rect 108535 280610 108541 280644
rect 108495 280572 108541 280610
rect 108495 280538 108501 280572
rect 108535 280538 108541 280572
rect 108495 280500 108541 280538
rect 108495 280466 108501 280500
rect 108535 280466 108541 280500
rect 108495 280428 108541 280466
rect 108495 280394 108501 280428
rect 108535 280394 108541 280428
rect 108495 280356 108541 280394
rect 108495 280322 108501 280356
rect 108535 280322 108541 280356
rect 108495 280284 108541 280322
rect 108495 280250 108501 280284
rect 108535 280250 108541 280284
rect 108495 280212 108541 280250
rect 108495 280178 108501 280212
rect 108535 280178 108541 280212
rect 108495 280140 108541 280178
rect 108495 280106 108501 280140
rect 108535 280106 108541 280140
rect 108495 280068 108541 280106
rect 108495 280034 108501 280068
rect 108535 280034 108541 280068
rect 108495 279996 108541 280034
rect 108495 279962 108501 279996
rect 108535 279962 108541 279996
rect 108495 279924 108541 279962
rect 108495 279890 108501 279924
rect 108535 279890 108541 279924
rect 108495 279852 108541 279890
rect 108495 279818 108501 279852
rect 108535 279818 108541 279852
rect 108495 279793 108541 279818
rect 108650 280788 108751 280813
rect 108650 280754 108711 280788
rect 108745 280754 108751 280788
rect 108650 280716 108751 280754
rect 108650 280682 108711 280716
rect 108745 280682 108751 280716
rect 108650 280644 108751 280682
rect 108650 280610 108711 280644
rect 108745 280610 108751 280644
rect 108650 280572 108751 280610
rect 108650 280538 108711 280572
rect 108745 280538 108751 280572
rect 108650 280500 108751 280538
rect 108650 280466 108711 280500
rect 108745 280466 108751 280500
rect 108650 280428 108751 280466
rect 108650 280394 108711 280428
rect 108745 280394 108751 280428
rect 108650 280356 108751 280394
rect 108650 280322 108711 280356
rect 108745 280322 108751 280356
rect 108650 280284 108751 280322
rect 108650 280250 108711 280284
rect 108745 280250 108751 280284
rect 108650 280212 108751 280250
rect 108650 280178 108711 280212
rect 108745 280178 108751 280212
rect 108650 280140 108751 280178
rect 108650 280106 108711 280140
rect 108745 280106 108751 280140
rect 108650 280068 108751 280106
rect 108650 280034 108711 280068
rect 108745 280034 108751 280068
rect 108650 279996 108751 280034
rect 108650 279962 108711 279996
rect 108745 279962 108751 279996
rect 108650 279924 108751 279962
rect 108650 279890 108711 279924
rect 108745 279890 108751 279924
rect 108650 279852 108751 279890
rect 108650 279818 108711 279852
rect 108745 279818 108751 279852
rect 108650 279793 108751 279818
rect 108895 280788 108941 280813
rect 108895 280754 108901 280788
rect 108935 280754 108941 280788
rect 108895 280716 108941 280754
rect 108895 280682 108901 280716
rect 108935 280682 108941 280716
rect 108895 280644 108941 280682
rect 108895 280610 108901 280644
rect 108935 280610 108941 280644
rect 108895 280572 108941 280610
rect 108895 280538 108901 280572
rect 108935 280538 108941 280572
rect 108895 280500 108941 280538
rect 108895 280466 108901 280500
rect 108935 280466 108941 280500
rect 108895 280428 108941 280466
rect 108895 280394 108901 280428
rect 108935 280394 108941 280428
rect 108895 280356 108941 280394
rect 108895 280322 108901 280356
rect 108935 280322 108941 280356
rect 108895 280284 108941 280322
rect 108895 280250 108901 280284
rect 108935 280250 108941 280284
rect 108895 280212 108941 280250
rect 108895 280178 108901 280212
rect 108935 280178 108941 280212
rect 108895 280140 108941 280178
rect 108895 280106 108901 280140
rect 108935 280106 108941 280140
rect 108895 280068 108941 280106
rect 108895 280034 108901 280068
rect 108935 280034 108941 280068
rect 108895 279996 108941 280034
rect 108895 279962 108901 279996
rect 108935 279962 108941 279996
rect 108895 279924 108941 279962
rect 108895 279890 108901 279924
rect 108935 279890 108941 279924
rect 108895 279852 108941 279890
rect 108895 279818 108901 279852
rect 108935 279818 108941 279852
rect 108895 279793 108941 279818
rect 109050 280788 109151 280813
rect 109050 280754 109111 280788
rect 109145 280754 109151 280788
rect 109050 280716 109151 280754
rect 109050 280682 109111 280716
rect 109145 280682 109151 280716
rect 109050 280644 109151 280682
rect 109050 280610 109111 280644
rect 109145 280610 109151 280644
rect 109050 280572 109151 280610
rect 109050 280538 109111 280572
rect 109145 280538 109151 280572
rect 109050 280500 109151 280538
rect 109050 280466 109111 280500
rect 109145 280466 109151 280500
rect 109050 280428 109151 280466
rect 109050 280394 109111 280428
rect 109145 280394 109151 280428
rect 109050 280356 109151 280394
rect 109050 280322 109111 280356
rect 109145 280322 109151 280356
rect 109050 280284 109151 280322
rect 109050 280250 109111 280284
rect 109145 280250 109151 280284
rect 109050 280212 109151 280250
rect 109050 280178 109111 280212
rect 109145 280178 109151 280212
rect 109050 280140 109151 280178
rect 109050 280106 109111 280140
rect 109145 280106 109151 280140
rect 109050 280068 109151 280106
rect 109050 280034 109111 280068
rect 109145 280034 109151 280068
rect 109050 279996 109151 280034
rect 109050 279962 109111 279996
rect 109145 279962 109151 279996
rect 109050 279924 109151 279962
rect 109050 279890 109111 279924
rect 109145 279890 109151 279924
rect 109050 279852 109151 279890
rect 109050 279818 109111 279852
rect 109145 279818 109151 279852
rect 109050 279793 109151 279818
rect 109295 280788 109341 280813
rect 109295 280754 109301 280788
rect 109335 280754 109341 280788
rect 109295 280716 109341 280754
rect 109295 280682 109301 280716
rect 109335 280682 109341 280716
rect 109295 280644 109341 280682
rect 109295 280610 109301 280644
rect 109335 280610 109341 280644
rect 109295 280572 109341 280610
rect 109295 280538 109301 280572
rect 109335 280538 109341 280572
rect 109295 280500 109341 280538
rect 109295 280466 109301 280500
rect 109335 280466 109341 280500
rect 109295 280428 109341 280466
rect 109295 280394 109301 280428
rect 109335 280394 109341 280428
rect 109295 280356 109341 280394
rect 109295 280322 109301 280356
rect 109335 280322 109341 280356
rect 109295 280284 109341 280322
rect 109295 280250 109301 280284
rect 109335 280250 109341 280284
rect 109295 280212 109341 280250
rect 109295 280178 109301 280212
rect 109335 280178 109341 280212
rect 109295 280140 109341 280178
rect 109295 280106 109301 280140
rect 109335 280106 109341 280140
rect 109295 280068 109341 280106
rect 109295 280034 109301 280068
rect 109335 280034 109341 280068
rect 109295 279996 109341 280034
rect 109295 279962 109301 279996
rect 109335 279962 109341 279996
rect 109295 279924 109341 279962
rect 109295 279890 109301 279924
rect 109335 279890 109341 279924
rect 109295 279852 109341 279890
rect 109295 279818 109301 279852
rect 109335 279818 109341 279852
rect 109295 279793 109341 279818
rect 109450 280788 109551 280813
rect 109450 280754 109511 280788
rect 109545 280754 109551 280788
rect 109450 280716 109551 280754
rect 109450 280682 109511 280716
rect 109545 280682 109551 280716
rect 109450 280644 109551 280682
rect 109450 280610 109511 280644
rect 109545 280610 109551 280644
rect 109450 280572 109551 280610
rect 109450 280538 109511 280572
rect 109545 280538 109551 280572
rect 109450 280500 109551 280538
rect 109450 280466 109511 280500
rect 109545 280466 109551 280500
rect 109450 280428 109551 280466
rect 109450 280394 109511 280428
rect 109545 280394 109551 280428
rect 109450 280356 109551 280394
rect 109450 280322 109511 280356
rect 109545 280322 109551 280356
rect 109450 280284 109551 280322
rect 109450 280250 109511 280284
rect 109545 280250 109551 280284
rect 109450 280212 109551 280250
rect 109450 280178 109511 280212
rect 109545 280178 109551 280212
rect 109450 280140 109551 280178
rect 109450 280106 109511 280140
rect 109545 280106 109551 280140
rect 109450 280068 109551 280106
rect 109450 280034 109511 280068
rect 109545 280034 109551 280068
rect 109450 279996 109551 280034
rect 109450 279962 109511 279996
rect 109545 279962 109551 279996
rect 109450 279924 109551 279962
rect 109450 279890 109511 279924
rect 109545 279890 109551 279924
rect 109450 279852 109551 279890
rect 109450 279818 109511 279852
rect 109545 279818 109551 279852
rect 109450 279793 109551 279818
rect 109695 280788 109741 280813
rect 109695 280754 109701 280788
rect 109735 280754 109741 280788
rect 109695 280716 109741 280754
rect 109695 280682 109701 280716
rect 109735 280682 109741 280716
rect 109695 280644 109741 280682
rect 109695 280610 109701 280644
rect 109735 280610 109741 280644
rect 109695 280572 109741 280610
rect 109695 280538 109701 280572
rect 109735 280538 109741 280572
rect 109695 280500 109741 280538
rect 109695 280466 109701 280500
rect 109735 280466 109741 280500
rect 109695 280428 109741 280466
rect 109695 280394 109701 280428
rect 109735 280394 109741 280428
rect 109695 280356 109741 280394
rect 109695 280322 109701 280356
rect 109735 280322 109741 280356
rect 109695 280284 109741 280322
rect 109695 280250 109701 280284
rect 109735 280250 109741 280284
rect 109695 280212 109741 280250
rect 109695 280178 109701 280212
rect 109735 280178 109741 280212
rect 109695 280140 109741 280178
rect 109695 280106 109701 280140
rect 109735 280106 109741 280140
rect 109695 280068 109741 280106
rect 109695 280034 109701 280068
rect 109735 280034 109741 280068
rect 109695 279996 109741 280034
rect 109695 279962 109701 279996
rect 109735 279962 109741 279996
rect 109695 279924 109741 279962
rect 109695 279890 109701 279924
rect 109735 279890 109741 279924
rect 109695 279852 109741 279890
rect 109695 279818 109701 279852
rect 109735 279818 109741 279852
rect 109695 279793 109741 279818
rect 109905 280788 109951 280813
rect 109905 280754 109911 280788
rect 109945 280754 109951 280788
rect 109905 280716 109951 280754
rect 109905 280682 109911 280716
rect 109945 280682 109951 280716
rect 109905 280644 109951 280682
rect 109905 280610 109911 280644
rect 109945 280610 109951 280644
rect 109905 280572 109951 280610
rect 109905 280538 109911 280572
rect 109945 280538 109951 280572
rect 109905 280500 109951 280538
rect 109905 280466 109911 280500
rect 109945 280466 109951 280500
rect 109905 280428 109951 280466
rect 109905 280394 109911 280428
rect 109945 280394 109951 280428
rect 109905 280356 109951 280394
rect 109905 280322 109911 280356
rect 109945 280322 109951 280356
rect 109905 280284 109951 280322
rect 109905 280250 109911 280284
rect 109945 280250 109951 280284
rect 109905 280212 109951 280250
rect 109905 280178 109911 280212
rect 109945 280178 109951 280212
rect 109905 280140 109951 280178
rect 109905 280106 109911 280140
rect 109945 280106 109951 280140
rect 109905 280068 109951 280106
rect 109905 280034 109911 280068
rect 109945 280034 109951 280068
rect 109905 279996 109951 280034
rect 109905 279962 109911 279996
rect 109945 279962 109951 279996
rect 109905 279924 109951 279962
rect 109905 279890 109911 279924
rect 109945 279890 109951 279924
rect 109905 279852 109951 279890
rect 109905 279818 109911 279852
rect 109945 279818 109951 279852
rect 109905 279793 109951 279818
rect 110095 280788 110141 280813
rect 110095 280754 110101 280788
rect 110135 280754 110141 280788
rect 110095 280716 110141 280754
rect 110095 280682 110101 280716
rect 110135 280682 110141 280716
rect 110095 280644 110141 280682
rect 110095 280610 110101 280644
rect 110135 280610 110141 280644
rect 110095 280572 110141 280610
rect 110095 280538 110101 280572
rect 110135 280538 110141 280572
rect 110095 280500 110141 280538
rect 110095 280466 110101 280500
rect 110135 280466 110141 280500
rect 110095 280428 110141 280466
rect 110095 280394 110101 280428
rect 110135 280394 110141 280428
rect 110095 280356 110141 280394
rect 110095 280322 110101 280356
rect 110135 280322 110141 280356
rect 110095 280284 110141 280322
rect 110095 280250 110101 280284
rect 110135 280250 110141 280284
rect 110095 280212 110141 280250
rect 110095 280178 110101 280212
rect 110135 280178 110141 280212
rect 110095 280140 110141 280178
rect 110095 280106 110101 280140
rect 110135 280106 110141 280140
rect 110095 280068 110141 280106
rect 110095 280034 110101 280068
rect 110135 280034 110141 280068
rect 110095 279996 110141 280034
rect 110095 279962 110101 279996
rect 110135 279962 110141 279996
rect 110095 279924 110141 279962
rect 110095 279890 110101 279924
rect 110135 279890 110141 279924
rect 110095 279852 110141 279890
rect 110095 279818 110101 279852
rect 110135 279818 110141 279852
rect 110095 279793 110141 279818
rect 106361 279755 106485 279761
rect 106361 279721 106406 279755
rect 106440 279721 106485 279755
rect 106361 279715 106485 279721
rect 106761 279755 106885 279761
rect 106761 279721 106806 279755
rect 106840 279721 106885 279755
rect 106761 279715 106885 279721
rect 106941 279401 106996 279793
rect 107161 279755 107285 279761
rect 107161 279721 107206 279755
rect 107240 279721 107285 279755
rect 107161 279715 107285 279721
rect 107341 279642 107396 279793
rect 107561 279755 107685 279761
rect 107561 279721 107606 279755
rect 107640 279721 107685 279755
rect 107561 279715 107685 279721
rect 107741 279642 107796 279793
rect 107961 279755 108085 279761
rect 107961 279721 108006 279755
rect 108040 279721 108085 279755
rect 107961 279715 108085 279721
rect 108361 279755 108485 279761
rect 108361 279721 108406 279755
rect 108440 279721 108485 279755
rect 108361 279715 108485 279721
rect 107341 279581 107796 279642
rect 107341 279529 107449 279581
rect 107501 279529 107513 279581
rect 107565 279529 107577 279581
rect 107629 279529 107641 279581
rect 107693 279529 107796 279581
rect 107341 279519 107796 279529
rect 108650 279641 108705 279793
rect 108761 279755 108885 279761
rect 108761 279721 108806 279755
rect 108840 279721 108885 279755
rect 108761 279715 108885 279721
rect 109050 279641 109105 279793
rect 109161 279755 109285 279761
rect 109161 279721 109206 279755
rect 109240 279721 109285 279755
rect 109161 279715 109285 279721
rect 108650 279581 109105 279641
rect 108650 279529 108759 279581
rect 108811 279529 108823 279581
rect 108875 279529 108887 279581
rect 108939 279529 108951 279581
rect 109003 279529 109105 279581
rect 108650 279519 109105 279529
rect 107341 279471 109105 279519
rect 109450 279401 109505 279793
rect 109561 279755 109685 279761
rect 109561 279721 109606 279755
rect 109640 279721 109685 279755
rect 109561 279715 109685 279721
rect 109961 279755 110085 279761
rect 109961 279721 110006 279755
rect 110040 279721 110085 279755
rect 109961 279715 110085 279721
rect 106941 279348 109505 279401
rect 107340 279231 107584 279258
rect 107340 279130 107409 279231
rect 106148 279115 107409 279130
rect 107525 279115 107584 279231
rect 106148 279065 107584 279115
rect 106148 279063 107582 279065
rect 106148 278530 106235 279063
rect 106368 279057 107582 279063
rect 106368 279023 106382 279057
rect 106416 279023 106454 279057
rect 106488 279023 106526 279057
rect 106560 279023 106598 279057
rect 106632 279023 106670 279057
rect 106704 279023 106742 279057
rect 106776 279023 106814 279057
rect 106848 279023 106886 279057
rect 106920 279023 106958 279057
rect 106992 279023 107030 279057
rect 107064 279023 107102 279057
rect 107136 279023 107174 279057
rect 107208 279023 107246 279057
rect 107280 279023 107318 279057
rect 107352 279023 107390 279057
rect 107424 279023 107462 279057
rect 107496 279023 107534 279057
rect 107568 279023 107582 279057
rect 106368 279017 107582 279023
rect 106281 278973 106327 279007
rect 106281 278939 106287 278973
rect 106321 278939 106327 278973
rect 106281 278901 106327 278939
rect 106281 278867 106287 278901
rect 106321 278867 106327 278901
rect 106281 278829 106327 278867
rect 106281 278795 106287 278829
rect 106321 278795 106327 278829
rect 106281 278761 106327 278795
rect 107623 278973 107669 279007
rect 107623 278939 107629 278973
rect 107663 278939 107669 278973
rect 107623 278901 107669 278939
rect 107623 278867 107629 278901
rect 107663 278867 107669 278901
rect 107623 278829 107669 278867
rect 107623 278795 107629 278829
rect 107663 278795 107669 278829
rect 107623 278761 107669 278795
rect 106368 278745 107582 278751
rect 106368 278711 106382 278745
rect 106416 278711 106454 278745
rect 106488 278711 106526 278745
rect 106560 278711 106598 278745
rect 106632 278711 106670 278745
rect 106704 278711 106742 278745
rect 106776 278711 106814 278745
rect 106848 278711 106886 278745
rect 106920 278711 106958 278745
rect 106992 278711 107030 278745
rect 107064 278711 107102 278745
rect 107136 278711 107174 278745
rect 107208 278711 107246 278745
rect 107280 278711 107318 278745
rect 107352 278711 107390 278745
rect 107424 278711 107462 278745
rect 107496 278711 107534 278745
rect 107568 278711 107582 278745
rect 106368 278705 107582 278711
rect 106368 278638 107796 278705
rect 106148 278463 107582 278530
rect 106368 278457 107582 278463
rect 106368 278423 106382 278457
rect 106416 278423 106454 278457
rect 106488 278423 106526 278457
rect 106560 278423 106598 278457
rect 106632 278423 106670 278457
rect 106704 278423 106742 278457
rect 106776 278423 106814 278457
rect 106848 278423 106886 278457
rect 106920 278423 106958 278457
rect 106992 278423 107030 278457
rect 107064 278423 107102 278457
rect 107136 278423 107174 278457
rect 107208 278423 107246 278457
rect 107280 278423 107318 278457
rect 107352 278423 107390 278457
rect 107424 278423 107462 278457
rect 107496 278423 107534 278457
rect 107568 278423 107582 278457
rect 106368 278417 107582 278423
rect 104099 278379 106210 278382
rect 106281 278379 106327 278407
rect 104099 278373 106327 278379
rect 104099 278339 106287 278373
rect 106321 278339 106327 278373
rect 104099 278301 106327 278339
rect 104099 278267 106287 278301
rect 106321 278267 106327 278301
rect 104099 278229 106327 278267
rect 104099 278195 106287 278229
rect 106321 278195 106327 278229
rect 104099 278179 106327 278195
rect 104099 278177 106210 278179
rect 102098 276457 103259 276621
rect 102098 275701 102266 276457
rect 103086 276209 103259 276457
rect 104099 276209 104304 278177
rect 106281 278161 106327 278179
rect 107623 278373 107669 278407
rect 107623 278339 107629 278373
rect 107663 278339 107669 278373
rect 107623 278301 107669 278339
rect 107623 278267 107629 278301
rect 107663 278267 107669 278301
rect 107623 278229 107669 278267
rect 107623 278195 107629 278229
rect 107663 278195 107669 278229
rect 107623 278161 107669 278195
rect 106368 278145 107582 278151
rect 106368 278111 106382 278145
rect 106416 278111 106454 278145
rect 106488 278111 106526 278145
rect 106560 278111 106598 278145
rect 106632 278111 106670 278145
rect 106704 278111 106742 278145
rect 106776 278111 106814 278145
rect 106848 278111 106886 278145
rect 106920 278111 106958 278145
rect 106992 278111 107030 278145
rect 107064 278111 107102 278145
rect 107136 278111 107174 278145
rect 107208 278111 107246 278145
rect 107280 278111 107318 278145
rect 107352 278111 107390 278145
rect 107424 278111 107462 278145
rect 107496 278111 107534 278145
rect 107568 278111 107582 278145
rect 106368 278105 107582 278111
rect 107709 278105 107796 278638
rect 106368 278053 107796 278105
rect 106368 278038 106966 278053
rect 103086 276004 104304 276209
rect 104854 277825 106544 277826
rect 104854 277627 106760 277825
rect 106902 277803 106966 278038
rect 107072 278038 107796 278053
rect 107072 277803 107130 278038
rect 106902 277799 107130 277803
rect 106902 277724 107553 277799
rect 106957 277722 107553 277724
rect 106957 277627 107033 277722
rect 104854 277478 107033 277627
rect 107469 277478 107553 277722
rect 104854 277407 107553 277478
rect 104854 277397 106760 277407
rect 106957 277403 107553 277407
rect 103086 275701 103259 276004
rect 102098 275531 103259 275701
rect 102557 274145 104316 274146
rect 104854 274145 105283 277397
rect 106959 277216 107081 277403
rect 106491 277210 107525 277216
rect 106491 277176 106523 277210
rect 106557 277176 106595 277210
rect 106629 277176 106667 277210
rect 106701 277176 106739 277210
rect 106773 277176 106811 277210
rect 106845 277176 106883 277210
rect 106917 277176 106955 277210
rect 106989 277176 107027 277210
rect 107061 277176 107099 277210
rect 107133 277176 107171 277210
rect 107205 277176 107243 277210
rect 107277 277176 107315 277210
rect 107349 277176 107387 277210
rect 107421 277176 107459 277210
rect 107493 277176 107525 277210
rect 106491 277170 107525 277176
rect 106404 277144 106450 277160
rect 106404 277110 106410 277144
rect 106444 277110 106450 277144
rect 106404 276855 106450 277110
rect 107566 277158 107612 277160
rect 107566 277144 107889 277158
rect 107566 277110 107572 277144
rect 107606 277110 107889 277144
rect 107566 277105 107889 277110
rect 107566 277102 107795 277105
rect 107566 277094 107612 277102
rect 106491 277078 107525 277084
rect 106491 277044 106523 277078
rect 106557 277044 106595 277078
rect 106629 277044 106667 277078
rect 106701 277044 106739 277078
rect 106773 277044 106811 277078
rect 106845 277044 106883 277078
rect 106917 277044 106955 277078
rect 106989 277044 107027 277078
rect 107061 277044 107099 277078
rect 107133 277044 107171 277078
rect 107205 277044 107243 277078
rect 107277 277044 107315 277078
rect 107349 277044 107387 277078
rect 107421 277044 107459 277078
rect 107493 277044 107525 277078
rect 106491 277038 107525 277044
rect 107754 277053 107795 277102
rect 107847 277053 107889 277105
rect 107754 277041 107889 277053
rect 107754 276989 107795 277041
rect 107847 276989 107889 277041
rect 107754 276977 107889 276989
rect 107754 276925 107795 276977
rect 107847 276925 107889 276977
rect 107754 276913 107889 276925
rect 107754 276861 107795 276913
rect 107847 276861 107889 276913
rect 107754 276855 107889 276861
rect 106404 276808 107889 276855
rect 106294 276272 106623 276403
rect 106294 275337 106409 276272
rect 106100 274870 106409 275337
rect 106515 274870 106623 276272
rect 107947 276126 108079 276165
rect 107947 276074 107987 276126
rect 108039 276074 108079 276126
rect 107947 276062 108079 276074
rect 107947 276010 107987 276062
rect 108039 276010 108079 276062
rect 107947 275882 108079 276010
rect 109196 275969 109291 279348
rect 109517 279089 110059 279151
rect 109517 277895 109569 279089
rect 109781 279083 110059 279089
rect 109781 279049 109795 279083
rect 109829 279049 109867 279083
rect 109901 279049 109939 279083
rect 109973 279049 110011 279083
rect 110045 279049 110059 279083
rect 109781 279043 110059 279049
rect 109725 278977 109771 279011
rect 109725 278943 109731 278977
rect 109765 278943 109771 278977
rect 109725 278905 109771 278943
rect 109725 278903 109731 278905
rect 109659 278871 109731 278903
rect 109765 278871 109771 278905
rect 109659 278850 109771 278871
rect 109659 278798 109692 278850
rect 109744 278833 109771 278850
rect 109765 278799 109771 278833
rect 109744 278798 109771 278799
rect 109659 278786 109771 278798
rect 109659 278734 109692 278786
rect 109744 278761 109771 278786
rect 109659 278727 109731 278734
rect 109765 278727 109771 278761
rect 109659 278722 109771 278727
rect 109659 278670 109692 278722
rect 109744 278689 109771 278722
rect 109659 278658 109731 278670
rect 109659 278606 109692 278658
rect 109765 278655 109771 278689
rect 109744 278617 109771 278655
rect 109659 278594 109731 278606
rect 109659 278542 109692 278594
rect 109765 278583 109771 278617
rect 109744 278545 109771 278583
rect 109659 278530 109731 278542
rect 109659 278478 109692 278530
rect 109765 278511 109771 278545
rect 109744 278478 109771 278511
rect 109659 278473 109771 278478
rect 109659 278466 109731 278473
rect 109659 278414 109692 278466
rect 109765 278439 109771 278473
rect 109744 278414 109771 278439
rect 109659 278402 109771 278414
rect 109659 278350 109692 278402
rect 109744 278401 109771 278402
rect 109765 278367 109771 278401
rect 109744 278350 109771 278367
rect 109659 278338 109771 278350
rect 109659 278286 109692 278338
rect 109744 278329 109771 278338
rect 109765 278295 109771 278329
rect 109744 278286 109771 278295
rect 109659 278274 109771 278286
rect 109659 278222 109692 278274
rect 109744 278257 109771 278274
rect 109765 278223 109771 278257
rect 109744 278222 109771 278223
rect 109659 278210 109771 278222
rect 109659 278158 109692 278210
rect 109744 278185 109771 278210
rect 109659 278151 109731 278158
rect 109765 278151 109771 278185
rect 109659 278146 109771 278151
rect 109659 278094 109692 278146
rect 109744 278113 109771 278146
rect 109659 278082 109731 278094
rect 109659 278030 109692 278082
rect 109765 278079 109771 278113
rect 109744 278041 109771 278079
rect 109659 278007 109731 278030
rect 109765 278007 109771 278041
rect 109659 277973 109771 278007
rect 110069 278977 110165 279011
rect 110069 278943 110075 278977
rect 110109 278943 110165 278977
rect 110069 278905 110165 278943
rect 110069 278871 110075 278905
rect 110109 278871 110165 278905
rect 110069 278833 110165 278871
rect 110069 278799 110075 278833
rect 110109 278799 110165 278833
rect 110069 278761 110165 278799
rect 110069 278727 110075 278761
rect 110109 278727 110165 278761
rect 110069 278689 110165 278727
rect 110069 278655 110075 278689
rect 110109 278655 110165 278689
rect 110069 278617 110165 278655
rect 110069 278583 110075 278617
rect 110109 278583 110165 278617
rect 110069 278545 110165 278583
rect 110069 278511 110075 278545
rect 110109 278511 110165 278545
rect 110069 278473 110165 278511
rect 110069 278439 110075 278473
rect 110109 278439 110165 278473
rect 110069 278401 110165 278439
rect 110069 278367 110075 278401
rect 110109 278367 110165 278401
rect 110069 278329 110165 278367
rect 110069 278295 110075 278329
rect 110109 278295 110165 278329
rect 110069 278257 110165 278295
rect 110069 278223 110075 278257
rect 110109 278223 110165 278257
rect 110069 278185 110165 278223
rect 110069 278151 110075 278185
rect 110109 278151 110165 278185
rect 110069 278113 110165 278151
rect 110069 278079 110075 278113
rect 110109 278079 110165 278113
rect 110069 278060 110165 278079
rect 110069 278041 110256 278060
rect 110069 278007 110075 278041
rect 110109 278007 110256 278041
rect 110069 277973 110256 278007
rect 109781 277935 110059 277941
rect 109781 277901 109795 277935
rect 109829 277901 109867 277935
rect 109901 277901 109939 277935
rect 109973 277901 110011 277935
rect 110045 277901 110059 277935
rect 109781 277895 110059 277901
rect 109517 277833 110059 277895
rect 109517 277341 109569 277833
rect 109781 277827 110059 277833
rect 109781 277793 109795 277827
rect 109829 277793 109867 277827
rect 109901 277793 109939 277827
rect 109973 277793 110011 277827
rect 110045 277793 110059 277827
rect 109781 277787 110059 277793
rect 110115 277755 110256 277973
rect 109413 277275 109569 277341
rect 109413 277223 109466 277275
rect 109518 277223 109569 277275
rect 109413 277211 109569 277223
rect 109413 277159 109466 277211
rect 109518 277159 109569 277211
rect 109413 277147 109569 277159
rect 109413 277095 109466 277147
rect 109518 277095 109569 277147
rect 109413 277083 109569 277095
rect 109413 277031 109466 277083
rect 109518 277031 109569 277083
rect 109413 277019 109569 277031
rect 109413 276967 109466 277019
rect 109518 276967 109569 277019
rect 109413 276955 109569 276967
rect 109413 276903 109466 276955
rect 109518 276903 109569 276955
rect 109413 276891 109569 276903
rect 109413 276839 109466 276891
rect 109518 276839 109569 276891
rect 109413 276827 109569 276839
rect 109413 276775 109466 276827
rect 109518 276775 109569 276827
rect 109659 277721 109771 277755
rect 109659 277696 109731 277721
rect 109659 277644 109687 277696
rect 109765 277687 109771 277721
rect 109739 277649 109771 277687
rect 109659 277632 109731 277644
rect 109659 277580 109687 277632
rect 109765 277615 109771 277649
rect 109739 277580 109771 277615
rect 109659 277577 109771 277580
rect 109659 277568 109731 277577
rect 109659 277516 109687 277568
rect 109765 277543 109771 277577
rect 109739 277516 109771 277543
rect 109659 277505 109771 277516
rect 109659 277504 109731 277505
rect 109659 277452 109687 277504
rect 109765 277471 109771 277505
rect 109739 277452 109771 277471
rect 109659 277440 109771 277452
rect 109659 277388 109687 277440
rect 109739 277433 109771 277440
rect 109765 277399 109771 277433
rect 109739 277388 109771 277399
rect 109659 277376 109771 277388
rect 109659 277324 109687 277376
rect 109739 277361 109771 277376
rect 109765 277327 109771 277361
rect 109739 277324 109771 277327
rect 109659 277312 109771 277324
rect 109659 277260 109687 277312
rect 109739 277289 109771 277312
rect 109659 277255 109731 277260
rect 109765 277255 109771 277289
rect 109659 277248 109771 277255
rect 109659 277196 109687 277248
rect 109739 277217 109771 277248
rect 109659 277184 109731 277196
rect 109659 277132 109687 277184
rect 109765 277183 109771 277217
rect 109739 277145 109771 277183
rect 109659 277120 109731 277132
rect 109659 277068 109687 277120
rect 109765 277111 109771 277145
rect 109739 277073 109771 277111
rect 109659 277056 109731 277068
rect 109659 277004 109687 277056
rect 109765 277039 109771 277073
rect 109739 277004 109771 277039
rect 109659 277001 109771 277004
rect 109659 276992 109731 277001
rect 109659 276940 109687 276992
rect 109765 276967 109771 277001
rect 109739 276940 109771 276967
rect 109659 276929 109771 276940
rect 109659 276928 109731 276929
rect 109659 276876 109687 276928
rect 109765 276895 109771 276929
rect 109739 276876 109771 276895
rect 109659 276857 109771 276876
rect 109659 276825 109731 276857
rect 109413 276763 109569 276775
rect 109413 276711 109466 276763
rect 109518 276711 109569 276763
rect 109725 276823 109731 276825
rect 109765 276823 109771 276857
rect 109725 276785 109771 276823
rect 109725 276751 109731 276785
rect 109765 276751 109771 276785
rect 109725 276717 109771 276751
rect 110069 277721 110256 277755
rect 110069 277687 110075 277721
rect 110109 277687 110256 277721
rect 110069 277649 110256 277687
rect 110069 277615 110075 277649
rect 110109 277615 110256 277649
rect 110069 277577 110256 277615
rect 110069 277543 110075 277577
rect 110109 277543 110256 277577
rect 110069 277505 110256 277543
rect 110069 277471 110075 277505
rect 110109 277471 110256 277505
rect 110069 277433 110256 277471
rect 110069 277399 110075 277433
rect 110109 277399 110256 277433
rect 110069 277361 110256 277399
rect 110069 277327 110075 277361
rect 110109 277327 110256 277361
rect 110069 277289 110256 277327
rect 110069 277255 110075 277289
rect 110109 277255 110256 277289
rect 110069 277217 110256 277255
rect 110069 277183 110075 277217
rect 110109 277183 110256 277217
rect 110069 277145 110256 277183
rect 110069 277111 110075 277145
rect 110109 277111 110256 277145
rect 110069 277073 110256 277111
rect 110069 277039 110075 277073
rect 110109 277039 110256 277073
rect 110069 277001 110256 277039
rect 110069 276967 110075 277001
rect 110109 276967 110256 277001
rect 110069 276929 110256 276967
rect 110069 276895 110075 276929
rect 110109 276895 110256 276929
rect 110069 276857 110256 276895
rect 110069 276823 110075 276857
rect 110109 276823 110256 276857
rect 110069 276785 110256 276823
rect 110069 276751 110075 276785
rect 110109 276751 110256 276785
rect 110069 276717 110256 276751
rect 109413 276699 109569 276711
rect 109413 276647 109466 276699
rect 109518 276647 109569 276699
rect 109413 276639 109569 276647
rect 109781 276679 110059 276685
rect 109781 276645 109795 276679
rect 109829 276645 109867 276679
rect 109901 276645 109939 276679
rect 109973 276645 110011 276679
rect 110045 276645 110059 276679
rect 109781 276639 110059 276645
rect 109413 276577 110059 276639
rect 110149 276420 110256 276717
rect 109824 276347 110271 276420
rect 109824 276167 109927 276347
rect 110171 276167 110271 276347
rect 109824 276093 110271 276167
rect 109193 275930 109712 275969
rect 107507 275832 109067 275882
rect 109193 275878 109263 275930
rect 109315 275878 109327 275930
rect 109379 275878 109391 275930
rect 109443 275878 109455 275930
rect 109507 275878 109519 275930
rect 109571 275878 109583 275930
rect 109635 275878 109712 275930
rect 109193 275836 109712 275878
rect 107507 275765 107567 275832
rect 109007 275765 109067 275832
rect 106951 275759 107129 275765
rect 106951 275725 106987 275759
rect 107021 275725 107059 275759
rect 107093 275725 107129 275759
rect 106951 275719 107129 275725
rect 107451 275759 107629 275765
rect 107451 275725 107487 275759
rect 107521 275725 107559 275759
rect 107593 275725 107629 275759
rect 107451 275719 107629 275725
rect 107951 275759 108629 275765
rect 107951 275725 107987 275759
rect 108021 275725 108059 275759
rect 108093 275725 108487 275759
rect 108521 275725 108559 275759
rect 108593 275725 108629 275759
rect 107951 275719 108629 275725
rect 108951 275759 109129 275765
rect 108951 275725 108987 275759
rect 109021 275725 109059 275759
rect 109093 275725 109129 275759
rect 108951 275719 109129 275725
rect 109451 275759 109629 275765
rect 109451 275725 109487 275759
rect 109521 275725 109559 275759
rect 109593 275725 109629 275759
rect 109451 275719 109629 275725
rect 108129 275709 108451 275719
rect 106864 275665 106910 275709
rect 106864 275631 106870 275665
rect 106904 275631 106910 275665
rect 106864 275593 106910 275631
rect 106864 275559 106870 275593
rect 106904 275559 106910 275593
rect 106864 275521 106910 275559
rect 106864 275487 106870 275521
rect 106904 275487 106910 275521
rect 106864 275449 106910 275487
rect 106864 275415 106870 275449
rect 106904 275415 106910 275449
rect 106864 275377 106910 275415
rect 106864 275343 106870 275377
rect 106904 275343 106910 275377
rect 106864 275305 106910 275343
rect 106864 275271 106870 275305
rect 106904 275271 106910 275305
rect 106864 275233 106910 275271
rect 106864 275199 106870 275233
rect 106904 275199 106910 275233
rect 106864 275161 106910 275199
rect 106864 275127 106870 275161
rect 106904 275127 106910 275161
rect 106864 275089 106910 275127
rect 106864 275055 106870 275089
rect 106904 275055 106910 275089
rect 106864 275017 106910 275055
rect 106864 274983 106870 275017
rect 106904 274983 106910 275017
rect 106864 274939 106910 274983
rect 107170 275665 107216 275709
rect 107170 275631 107176 275665
rect 107210 275631 107216 275665
rect 107170 275593 107216 275631
rect 107170 275559 107176 275593
rect 107210 275559 107216 275593
rect 107170 275521 107216 275559
rect 107170 275487 107176 275521
rect 107210 275487 107216 275521
rect 107170 275449 107216 275487
rect 107170 275415 107176 275449
rect 107210 275415 107216 275449
rect 107170 275377 107216 275415
rect 107170 275343 107176 275377
rect 107210 275343 107216 275377
rect 107170 275305 107216 275343
rect 107170 275271 107176 275305
rect 107210 275271 107216 275305
rect 107170 275233 107216 275271
rect 107170 275199 107176 275233
rect 107210 275199 107216 275233
rect 107170 275161 107216 275199
rect 107170 275127 107176 275161
rect 107210 275127 107216 275161
rect 107170 275089 107216 275127
rect 107170 275055 107176 275089
rect 107210 275055 107216 275089
rect 107170 275017 107216 275055
rect 107170 274983 107176 275017
rect 107210 274983 107216 275017
rect 107170 274939 107216 274983
rect 107364 275665 107410 275709
rect 107364 275631 107370 275665
rect 107404 275631 107410 275665
rect 107364 275593 107410 275631
rect 107364 275559 107370 275593
rect 107404 275559 107410 275593
rect 107364 275521 107410 275559
rect 107364 275487 107370 275521
rect 107404 275487 107410 275521
rect 107364 275449 107410 275487
rect 107364 275415 107370 275449
rect 107404 275415 107410 275449
rect 107364 275377 107410 275415
rect 107364 275343 107370 275377
rect 107404 275343 107410 275377
rect 107364 275305 107410 275343
rect 107364 275271 107370 275305
rect 107404 275271 107410 275305
rect 107364 275233 107410 275271
rect 107364 275199 107370 275233
rect 107404 275199 107410 275233
rect 107364 275161 107410 275199
rect 107364 275127 107370 275161
rect 107404 275127 107410 275161
rect 107364 275089 107410 275127
rect 107364 275055 107370 275089
rect 107404 275055 107410 275089
rect 107364 275017 107410 275055
rect 107364 274983 107370 275017
rect 107404 274983 107410 275017
rect 107364 274939 107410 274983
rect 107670 275665 107716 275709
rect 107670 275631 107676 275665
rect 107710 275631 107716 275665
rect 107670 275593 107716 275631
rect 107670 275559 107676 275593
rect 107710 275559 107716 275593
rect 107670 275521 107716 275559
rect 107670 275487 107676 275521
rect 107710 275487 107716 275521
rect 107670 275449 107716 275487
rect 107670 275415 107676 275449
rect 107710 275415 107716 275449
rect 107670 275393 107716 275415
rect 107864 275665 107910 275709
rect 107864 275631 107870 275665
rect 107904 275631 107910 275665
rect 107864 275593 107910 275631
rect 107864 275559 107870 275593
rect 107904 275559 107910 275593
rect 107864 275521 107910 275559
rect 107864 275487 107870 275521
rect 107904 275487 107910 275521
rect 107864 275449 107910 275487
rect 107864 275415 107870 275449
rect 107904 275415 107910 275449
rect 107864 275393 107910 275415
rect 107670 275377 107910 275393
rect 107670 275343 107676 275377
rect 107710 275343 107870 275377
rect 107904 275343 107910 275377
rect 107670 275305 107910 275343
rect 107670 275271 107676 275305
rect 107710 275271 107870 275305
rect 107904 275271 107910 275305
rect 107670 275259 107910 275271
rect 107670 275233 107716 275259
rect 107670 275199 107676 275233
rect 107710 275199 107716 275233
rect 107670 275161 107716 275199
rect 107670 275127 107676 275161
rect 107710 275127 107716 275161
rect 107670 275089 107716 275127
rect 107670 275055 107676 275089
rect 107710 275055 107716 275089
rect 107670 275017 107716 275055
rect 107670 274983 107676 275017
rect 107710 274983 107716 275017
rect 107670 274939 107716 274983
rect 107864 275233 107910 275259
rect 107864 275199 107870 275233
rect 107904 275199 107910 275233
rect 107864 275161 107910 275199
rect 107864 275127 107870 275161
rect 107904 275127 107910 275161
rect 107864 275089 107910 275127
rect 107864 275055 107870 275089
rect 107904 275055 107910 275089
rect 107864 275017 107910 275055
rect 107864 274983 107870 275017
rect 107904 274983 107910 275017
rect 107864 274939 107910 274983
rect 108170 275665 108232 275709
rect 108170 275631 108176 275665
rect 108210 275631 108232 275665
rect 108170 275593 108232 275631
rect 108348 275665 108410 275709
rect 108348 275631 108370 275665
rect 108404 275631 108410 275665
rect 108348 275593 108410 275631
rect 108170 275559 108176 275593
rect 108210 275559 108370 275593
rect 108404 275559 108410 275593
rect 108170 275522 108410 275559
rect 108170 275521 108216 275522
rect 108170 275487 108176 275521
rect 108210 275487 108216 275521
rect 108170 275449 108216 275487
rect 108170 275415 108176 275449
rect 108210 275415 108216 275449
rect 108170 275393 108216 275415
rect 108364 275521 108410 275522
rect 108364 275487 108370 275521
rect 108404 275487 108410 275521
rect 108364 275449 108410 275487
rect 108364 275415 108370 275449
rect 108404 275415 108410 275449
rect 108364 275393 108410 275415
rect 108170 275377 108410 275393
rect 108170 275343 108176 275377
rect 108210 275343 108370 275377
rect 108404 275343 108410 275377
rect 108170 275305 108410 275343
rect 108170 275271 108176 275305
rect 108210 275271 108370 275305
rect 108404 275271 108410 275305
rect 108170 275259 108410 275271
rect 108170 275233 108216 275259
rect 108170 275199 108176 275233
rect 108210 275199 108216 275233
rect 108170 275161 108216 275199
rect 108170 275127 108176 275161
rect 108210 275127 108216 275161
rect 108170 275089 108216 275127
rect 108170 275055 108176 275089
rect 108210 275055 108216 275089
rect 108170 275017 108216 275055
rect 108170 274983 108176 275017
rect 108210 274983 108216 275017
rect 108170 274939 108216 274983
rect 108364 275233 108410 275259
rect 108364 275199 108370 275233
rect 108404 275199 108410 275233
rect 108364 275161 108410 275199
rect 108364 275127 108370 275161
rect 108404 275127 108410 275161
rect 108364 275089 108410 275127
rect 108364 275055 108370 275089
rect 108404 275055 108410 275089
rect 108364 275017 108410 275055
rect 108364 274983 108370 275017
rect 108404 274983 108410 275017
rect 108364 274939 108410 274983
rect 108670 275665 108716 275709
rect 108670 275631 108676 275665
rect 108710 275631 108716 275665
rect 108670 275593 108716 275631
rect 108670 275559 108676 275593
rect 108710 275559 108716 275593
rect 108670 275521 108716 275559
rect 108670 275487 108676 275521
rect 108710 275487 108716 275521
rect 108670 275449 108716 275487
rect 108670 275415 108676 275449
rect 108710 275415 108716 275449
rect 108670 275393 108716 275415
rect 108864 275665 108910 275709
rect 108864 275631 108870 275665
rect 108904 275631 108910 275665
rect 108864 275593 108910 275631
rect 108864 275559 108870 275593
rect 108904 275559 108910 275593
rect 108864 275521 108910 275559
rect 108864 275487 108870 275521
rect 108904 275487 108910 275521
rect 108864 275449 108910 275487
rect 108864 275415 108870 275449
rect 108904 275415 108910 275449
rect 108864 275393 108910 275415
rect 108670 275377 108910 275393
rect 108670 275343 108676 275377
rect 108710 275343 108870 275377
rect 108904 275343 108910 275377
rect 108670 275305 108910 275343
rect 108670 275271 108676 275305
rect 108710 275271 108870 275305
rect 108904 275271 108910 275305
rect 108670 275259 108910 275271
rect 108670 275233 108716 275259
rect 108670 275199 108676 275233
rect 108710 275199 108716 275233
rect 108670 275161 108716 275199
rect 108670 275127 108676 275161
rect 108710 275127 108716 275161
rect 108670 275089 108716 275127
rect 108670 275055 108676 275089
rect 108710 275055 108716 275089
rect 108670 275017 108716 275055
rect 108670 274983 108676 275017
rect 108710 274983 108716 275017
rect 108670 274939 108716 274983
rect 108864 275233 108910 275259
rect 108864 275199 108870 275233
rect 108904 275199 108910 275233
rect 108864 275161 108910 275199
rect 108864 275127 108870 275161
rect 108904 275127 108910 275161
rect 108864 275089 108910 275127
rect 108864 275055 108870 275089
rect 108904 275055 108910 275089
rect 108864 275017 108910 275055
rect 108864 274983 108870 275017
rect 108904 274983 108910 275017
rect 108864 274939 108910 274983
rect 109170 275665 109216 275709
rect 109170 275631 109176 275665
rect 109210 275631 109216 275665
rect 109170 275593 109216 275631
rect 109170 275559 109176 275593
rect 109210 275559 109216 275593
rect 109170 275521 109216 275559
rect 109170 275487 109176 275521
rect 109210 275487 109216 275521
rect 109170 275449 109216 275487
rect 109170 275415 109176 275449
rect 109210 275415 109216 275449
rect 109170 275377 109216 275415
rect 109170 275343 109176 275377
rect 109210 275343 109216 275377
rect 109170 275305 109216 275343
rect 109170 275271 109176 275305
rect 109210 275271 109216 275305
rect 109170 275233 109216 275271
rect 109170 275199 109176 275233
rect 109210 275199 109216 275233
rect 109170 275161 109216 275199
rect 109170 275127 109176 275161
rect 109210 275127 109216 275161
rect 109170 275089 109216 275127
rect 109170 275055 109176 275089
rect 109210 275055 109216 275089
rect 109170 275017 109216 275055
rect 109170 274983 109176 275017
rect 109210 274983 109216 275017
rect 109170 274939 109216 274983
rect 109364 275665 109410 275709
rect 109364 275631 109370 275665
rect 109404 275631 109410 275665
rect 109364 275593 109410 275631
rect 109364 275559 109370 275593
rect 109404 275559 109410 275593
rect 109364 275521 109410 275559
rect 109364 275487 109370 275521
rect 109404 275487 109410 275521
rect 109364 275449 109410 275487
rect 109364 275415 109370 275449
rect 109404 275415 109410 275449
rect 109364 275377 109410 275415
rect 109364 275343 109370 275377
rect 109404 275343 109410 275377
rect 109364 275305 109410 275343
rect 109364 275271 109370 275305
rect 109404 275271 109410 275305
rect 109364 275233 109410 275271
rect 109364 275199 109370 275233
rect 109404 275199 109410 275233
rect 109364 275161 109410 275199
rect 109364 275127 109370 275161
rect 109404 275127 109410 275161
rect 109364 275089 109410 275127
rect 109364 275055 109370 275089
rect 109404 275055 109410 275089
rect 109364 275017 109410 275055
rect 109364 274983 109370 275017
rect 109404 274983 109410 275017
rect 109364 274939 109410 274983
rect 109670 275665 109716 275709
rect 109670 275631 109676 275665
rect 109710 275631 109716 275665
rect 109670 275593 109716 275631
rect 109670 275559 109676 275593
rect 109710 275559 109716 275593
rect 109670 275521 109716 275559
rect 109670 275487 109676 275521
rect 109710 275487 109716 275521
rect 109670 275449 109716 275487
rect 109670 275415 109676 275449
rect 109710 275415 109716 275449
rect 109670 275377 109716 275415
rect 109670 275343 109676 275377
rect 109710 275343 109716 275377
rect 109670 275305 109716 275343
rect 109670 275271 109676 275305
rect 109710 275271 109716 275305
rect 109670 275233 109716 275271
rect 109670 275199 109676 275233
rect 109710 275199 109716 275233
rect 109670 275161 109716 275199
rect 109670 275127 109676 275161
rect 109710 275127 109716 275161
rect 109670 275089 109716 275127
rect 109670 275055 109676 275089
rect 109710 275055 109716 275089
rect 109670 275017 109716 275055
rect 109670 274983 109676 275017
rect 109710 274983 109716 275017
rect 109670 274939 109716 274983
rect 106951 274923 107129 274929
rect 106951 274889 106987 274923
rect 107021 274889 107059 274923
rect 107093 274889 107129 274923
rect 106951 274883 107129 274889
rect 107451 274923 107629 274929
rect 107451 274889 107487 274923
rect 107521 274889 107559 274923
rect 107593 274889 107629 274923
rect 107451 274883 107629 274889
rect 107951 274923 108129 274929
rect 107951 274889 107987 274923
rect 108021 274889 108059 274923
rect 108093 274889 108129 274923
rect 107951 274883 108129 274889
rect 108451 274923 108629 274929
rect 108451 274889 108487 274923
rect 108521 274889 108559 274923
rect 108593 274889 108629 274923
rect 108451 274883 108629 274889
rect 108951 274923 109129 274929
rect 108951 274889 108987 274923
rect 109021 274889 109059 274923
rect 109093 274889 109129 274923
rect 108951 274883 109129 274889
rect 109451 274923 109629 274929
rect 109451 274889 109487 274923
rect 109521 274889 109559 274923
rect 109593 274889 109629 274923
rect 109451 274883 109629 274889
rect 106100 274731 106623 274870
rect 106100 274505 106622 274731
rect 110521 274509 111012 282251
rect 119259 281225 119845 282251
rect 119257 281140 119845 281225
rect 112970 280874 114070 280880
rect 111524 280866 112624 280872
rect 111524 280832 111553 280866
rect 111587 280832 111625 280866
rect 111659 280832 111697 280866
rect 111731 280832 111769 280866
rect 111803 280832 111841 280866
rect 111875 280832 111913 280866
rect 111947 280832 111985 280866
rect 112019 280832 112057 280866
rect 112091 280832 112129 280866
rect 112163 280832 112201 280866
rect 112235 280832 112273 280866
rect 112307 280832 112345 280866
rect 112379 280832 112417 280866
rect 112451 280832 112489 280866
rect 112523 280832 112561 280866
rect 112595 280832 112624 280866
rect 112970 280840 112999 280874
rect 113033 280840 113071 280874
rect 113105 280840 113143 280874
rect 113177 280840 113215 280874
rect 113249 280840 113287 280874
rect 113321 280840 113359 280874
rect 113393 280840 113431 280874
rect 113465 280840 113503 280874
rect 113537 280840 113575 280874
rect 113609 280840 113647 280874
rect 113681 280840 113719 280874
rect 113753 280840 113791 280874
rect 113825 280840 113863 280874
rect 113897 280840 113935 280874
rect 113969 280840 114007 280874
rect 114041 280840 114070 280874
rect 116135 280874 117235 280880
rect 112970 280834 114070 280840
rect 114657 280849 114857 280855
rect 111524 280826 112624 280832
rect 111404 280793 111492 280816
rect 111404 280759 111452 280793
rect 111486 280759 111492 280793
rect 111404 280721 111492 280759
rect 111404 280687 111452 280721
rect 111486 280687 111492 280721
rect 111404 280664 111492 280687
rect 112656 280793 112744 280816
rect 112656 280759 112662 280793
rect 112696 280759 112744 280793
rect 112656 280748 112744 280759
rect 112850 280781 112938 280824
rect 112850 280748 112898 280781
rect 112656 280747 112898 280748
rect 112932 280747 112938 280781
rect 112656 280721 112938 280747
rect 112656 280687 112662 280721
rect 112696 280709 112938 280721
rect 112696 280687 112898 280709
rect 112656 280686 112898 280687
rect 112656 280664 112744 280686
rect 111404 280456 111446 280664
rect 111524 280648 112624 280654
rect 111524 280614 111553 280648
rect 111587 280614 111625 280648
rect 111659 280614 111697 280648
rect 111731 280614 111769 280648
rect 111803 280614 111841 280648
rect 111875 280614 111913 280648
rect 111947 280614 111985 280648
rect 112019 280614 112057 280648
rect 112091 280614 112129 280648
rect 112163 280614 112201 280648
rect 112235 280614 112273 280648
rect 112307 280614 112345 280648
rect 112379 280614 112417 280648
rect 112451 280614 112489 280648
rect 112523 280614 112561 280648
rect 112595 280614 112624 280648
rect 111524 280608 112624 280614
rect 112702 280632 112744 280664
rect 112850 280675 112898 280686
rect 112932 280675 112938 280709
rect 112850 280632 112938 280675
rect 114102 280781 114190 280824
rect 114657 280815 114704 280849
rect 114738 280815 114776 280849
rect 114810 280815 114857 280849
rect 114657 280809 114857 280815
rect 115348 280849 115548 280855
rect 115348 280815 115395 280849
rect 115429 280815 115467 280849
rect 115501 280815 115548 280849
rect 116135 280840 116164 280874
rect 116198 280840 116236 280874
rect 116270 280840 116308 280874
rect 116342 280840 116380 280874
rect 116414 280840 116452 280874
rect 116486 280840 116524 280874
rect 116558 280840 116596 280874
rect 116630 280840 116668 280874
rect 116702 280840 116740 280874
rect 116774 280840 116812 280874
rect 116846 280840 116884 280874
rect 116918 280840 116956 280874
rect 116990 280840 117028 280874
rect 117062 280840 117100 280874
rect 117134 280840 117172 280874
rect 117206 280840 117235 280874
rect 116135 280834 117235 280840
rect 117581 280866 118681 280872
rect 117581 280832 117610 280866
rect 117644 280832 117682 280866
rect 117716 280832 117754 280866
rect 117788 280832 117826 280866
rect 117860 280832 117898 280866
rect 117932 280832 117970 280866
rect 118004 280832 118042 280866
rect 118076 280832 118114 280866
rect 118148 280832 118186 280866
rect 118220 280832 118258 280866
rect 118292 280832 118330 280866
rect 118364 280832 118402 280866
rect 118436 280832 118474 280866
rect 118508 280832 118546 280866
rect 118580 280832 118618 280866
rect 118652 280832 118681 280866
rect 117581 280826 118681 280832
rect 115348 280809 115548 280815
rect 114102 280747 114108 280781
rect 114142 280758 114190 280781
rect 114570 280764 114616 280799
rect 114570 280758 114576 280764
rect 114142 280747 114576 280758
rect 114102 280730 114576 280747
rect 114610 280730 114616 280764
rect 114102 280709 114616 280730
rect 114102 280675 114108 280709
rect 114142 280692 114616 280709
rect 114142 280675 114576 280692
rect 114102 280658 114576 280675
rect 114610 280658 114616 280692
rect 114102 280632 114616 280658
rect 111524 280506 112624 280512
rect 111524 280472 111553 280506
rect 111587 280472 111625 280506
rect 111659 280472 111697 280506
rect 111731 280472 111769 280506
rect 111803 280472 111841 280506
rect 111875 280472 111913 280506
rect 111947 280472 111985 280506
rect 112019 280472 112057 280506
rect 112091 280472 112129 280506
rect 112163 280472 112201 280506
rect 112235 280472 112273 280506
rect 112307 280472 112345 280506
rect 112379 280472 112417 280506
rect 112451 280472 112489 280506
rect 112523 280472 112561 280506
rect 112595 280472 112624 280506
rect 111524 280466 112624 280472
rect 112702 280456 112746 280632
rect 111404 280433 111492 280456
rect 111404 280399 111452 280433
rect 111486 280399 111492 280433
rect 111404 280361 111492 280399
rect 111404 280327 111452 280361
rect 111486 280327 111492 280361
rect 111404 280304 111492 280327
rect 112656 280433 112746 280456
rect 112656 280399 112662 280433
rect 112696 280412 112746 280433
rect 112850 280532 112892 280632
rect 114148 280625 114616 280632
rect 112970 280616 114070 280622
rect 112970 280582 112999 280616
rect 113033 280582 113071 280616
rect 113105 280582 113143 280616
rect 113177 280582 113215 280616
rect 113249 280582 113287 280616
rect 113321 280582 113359 280616
rect 113393 280582 113431 280616
rect 113465 280582 113503 280616
rect 113537 280582 113575 280616
rect 113609 280582 113647 280616
rect 113681 280582 113719 280616
rect 113753 280582 113791 280616
rect 113825 280582 113863 280616
rect 113897 280582 113935 280616
rect 113969 280582 114007 280616
rect 114041 280582 114070 280616
rect 112970 280576 114070 280582
rect 114148 280532 114190 280625
rect 112850 280494 114190 280532
rect 112696 280399 112744 280412
rect 112656 280364 112744 280399
rect 112850 280400 112892 280494
rect 112970 280450 114070 280456
rect 112970 280416 112999 280450
rect 113033 280416 113071 280450
rect 113105 280416 113143 280450
rect 113177 280416 113215 280450
rect 113249 280416 113287 280450
rect 113321 280416 113359 280450
rect 113393 280416 113431 280450
rect 113465 280416 113503 280450
rect 113537 280416 113575 280450
rect 113609 280416 113647 280450
rect 113681 280416 113719 280450
rect 113753 280416 113791 280450
rect 113825 280416 113863 280450
rect 113897 280416 113935 280450
rect 113969 280416 114007 280450
rect 114041 280416 114070 280450
rect 112970 280410 114070 280416
rect 114148 280400 114190 280494
rect 114570 280620 114616 280625
rect 114570 280586 114576 280620
rect 114610 280586 114616 280620
rect 114570 280548 114616 280586
rect 114570 280514 114576 280548
rect 114610 280514 114616 280548
rect 114570 280476 114616 280514
rect 114570 280442 114576 280476
rect 114610 280442 114616 280476
rect 114570 280407 114616 280442
rect 114898 280764 114944 280799
rect 114898 280730 114904 280764
rect 114938 280730 114944 280764
rect 114898 280692 114944 280730
rect 114898 280658 114904 280692
rect 114938 280658 114944 280692
rect 114898 280620 114944 280658
rect 114898 280586 114904 280620
rect 114938 280586 114944 280620
rect 114898 280548 114944 280586
rect 114898 280514 114904 280548
rect 114938 280514 114944 280548
rect 114898 280476 114944 280514
rect 114898 280442 114904 280476
rect 114938 280442 114944 280476
rect 114898 280407 114944 280442
rect 115261 280764 115307 280799
rect 115261 280730 115267 280764
rect 115301 280730 115307 280764
rect 115261 280692 115307 280730
rect 115261 280658 115267 280692
rect 115301 280658 115307 280692
rect 115261 280620 115307 280658
rect 115261 280586 115267 280620
rect 115301 280586 115307 280620
rect 115261 280548 115307 280586
rect 115261 280514 115267 280548
rect 115301 280514 115307 280548
rect 115261 280476 115307 280514
rect 115261 280442 115267 280476
rect 115301 280442 115307 280476
rect 115261 280407 115307 280442
rect 115589 280764 115635 280799
rect 115589 280730 115595 280764
rect 115629 280758 115635 280764
rect 116015 280781 116103 280824
rect 116015 280758 116063 280781
rect 115629 280747 116063 280758
rect 116097 280747 116103 280781
rect 115629 280730 116103 280747
rect 115589 280709 116103 280730
rect 115589 280692 116063 280709
rect 115589 280658 115595 280692
rect 115629 280675 116063 280692
rect 116097 280675 116103 280709
rect 115629 280658 116103 280675
rect 115589 280632 116103 280658
rect 117267 280781 117355 280824
rect 117267 280747 117273 280781
rect 117307 280748 117355 280781
rect 117461 280793 117549 280816
rect 117461 280759 117509 280793
rect 117543 280759 117549 280793
rect 117461 280748 117549 280759
rect 117307 280747 117549 280748
rect 117267 280721 117549 280747
rect 117267 280709 117509 280721
rect 117267 280675 117273 280709
rect 117307 280687 117509 280709
rect 117543 280687 117549 280721
rect 117307 280686 117549 280687
rect 117307 280675 117355 280686
rect 117267 280632 117355 280675
rect 117461 280664 117549 280686
rect 118713 280793 118801 280816
rect 118713 280759 118719 280793
rect 118753 280759 118801 280793
rect 118713 280721 118801 280759
rect 118713 280687 118719 280721
rect 118753 280687 118801 280721
rect 118713 280664 118801 280687
rect 117461 280632 117503 280664
rect 115589 280625 116057 280632
rect 115589 280620 115635 280625
rect 115589 280586 115595 280620
rect 115629 280586 115635 280620
rect 115589 280548 115635 280586
rect 115589 280514 115595 280548
rect 115629 280514 115635 280548
rect 115589 280476 115635 280514
rect 115589 280442 115595 280476
rect 115629 280442 115635 280476
rect 115589 280407 115635 280442
rect 116015 280532 116057 280625
rect 116135 280616 117235 280622
rect 116135 280582 116164 280616
rect 116198 280582 116236 280616
rect 116270 280582 116308 280616
rect 116342 280582 116380 280616
rect 116414 280582 116452 280616
rect 116486 280582 116524 280616
rect 116558 280582 116596 280616
rect 116630 280582 116668 280616
rect 116702 280582 116740 280616
rect 116774 280582 116812 280616
rect 116846 280582 116884 280616
rect 116918 280582 116956 280616
rect 116990 280582 117028 280616
rect 117062 280582 117100 280616
rect 117134 280582 117172 280616
rect 117206 280582 117235 280616
rect 116135 280576 117235 280582
rect 117313 280532 117355 280632
rect 116015 280494 117355 280532
rect 112850 280364 112938 280400
rect 112656 280361 112938 280364
rect 112656 280327 112662 280361
rect 112696 280357 112938 280361
rect 112696 280327 112898 280357
rect 112656 280323 112898 280327
rect 112932 280323 112938 280357
rect 112656 280304 112938 280323
rect 111404 280096 111446 280304
rect 112702 280302 112938 280304
rect 111524 280288 112624 280294
rect 111524 280254 111553 280288
rect 111587 280254 111625 280288
rect 111659 280254 111697 280288
rect 111731 280254 111769 280288
rect 111803 280254 111841 280288
rect 111875 280254 111913 280288
rect 111947 280254 111985 280288
rect 112019 280254 112057 280288
rect 112091 280254 112129 280288
rect 112163 280254 112201 280288
rect 112235 280254 112273 280288
rect 112307 280254 112345 280288
rect 112379 280254 112417 280288
rect 112451 280254 112489 280288
rect 112523 280254 112561 280288
rect 112595 280254 112624 280288
rect 111524 280248 112624 280254
rect 111524 280146 112624 280152
rect 111524 280112 111553 280146
rect 111587 280112 111625 280146
rect 111659 280112 111697 280146
rect 111731 280112 111769 280146
rect 111803 280112 111841 280146
rect 111875 280112 111913 280146
rect 111947 280112 111985 280146
rect 112019 280112 112057 280146
rect 112091 280112 112129 280146
rect 112163 280112 112201 280146
rect 112235 280112 112273 280146
rect 112307 280112 112345 280146
rect 112379 280112 112417 280146
rect 112451 280112 112489 280146
rect 112523 280112 112561 280146
rect 112595 280112 112624 280146
rect 111524 280106 112624 280112
rect 112702 280096 112744 280302
rect 112850 280285 112938 280302
rect 112850 280251 112898 280285
rect 112932 280251 112938 280285
rect 112850 280208 112938 280251
rect 114102 280357 114190 280400
rect 116015 280400 116057 280494
rect 116135 280450 117235 280456
rect 116135 280416 116164 280450
rect 116198 280416 116236 280450
rect 116270 280416 116308 280450
rect 116342 280416 116380 280450
rect 116414 280416 116452 280450
rect 116486 280416 116524 280450
rect 116558 280416 116596 280450
rect 116630 280416 116668 280450
rect 116702 280416 116740 280450
rect 116774 280416 116812 280450
rect 116846 280416 116884 280450
rect 116918 280416 116956 280450
rect 116990 280416 117028 280450
rect 117062 280416 117100 280450
rect 117134 280416 117172 280450
rect 117206 280416 117235 280450
rect 116135 280410 117235 280416
rect 117313 280400 117355 280494
rect 117459 280456 117503 280632
rect 117581 280648 118681 280654
rect 117581 280614 117610 280648
rect 117644 280614 117682 280648
rect 117716 280614 117754 280648
rect 117788 280614 117826 280648
rect 117860 280614 117898 280648
rect 117932 280614 117970 280648
rect 118004 280614 118042 280648
rect 118076 280614 118114 280648
rect 118148 280614 118186 280648
rect 118220 280614 118258 280648
rect 118292 280614 118330 280648
rect 118364 280614 118402 280648
rect 118436 280614 118474 280648
rect 118508 280614 118546 280648
rect 118580 280614 118618 280648
rect 118652 280614 118681 280648
rect 117581 280608 118681 280614
rect 117581 280506 118681 280512
rect 117581 280472 117610 280506
rect 117644 280472 117682 280506
rect 117716 280472 117754 280506
rect 117788 280472 117826 280506
rect 117860 280472 117898 280506
rect 117932 280472 117970 280506
rect 118004 280472 118042 280506
rect 118076 280472 118114 280506
rect 118148 280472 118186 280506
rect 118220 280472 118258 280506
rect 118292 280472 118330 280506
rect 118364 280472 118402 280506
rect 118436 280472 118474 280506
rect 118508 280472 118546 280506
rect 118580 280472 118618 280506
rect 118652 280472 118681 280506
rect 117581 280466 118681 280472
rect 118759 280456 118801 280664
rect 117459 280433 117549 280456
rect 117459 280412 117509 280433
rect 114102 280323 114108 280357
rect 114142 280323 114190 280357
rect 114657 280391 114857 280397
rect 114657 280357 114704 280391
rect 114738 280357 114776 280391
rect 114810 280357 114857 280391
rect 114657 280351 114857 280357
rect 115348 280391 115548 280397
rect 115348 280357 115395 280391
rect 115429 280357 115467 280391
rect 115501 280357 115548 280391
rect 115348 280351 115548 280357
rect 116015 280357 116103 280400
rect 114102 280285 114190 280323
rect 114102 280251 114108 280285
rect 114142 280251 114190 280285
rect 114720 280283 114790 280351
rect 114102 280208 114190 280251
rect 114308 280199 114790 280283
rect 114865 280286 114970 280311
rect 114865 280234 114890 280286
rect 114942 280234 114970 280286
rect 114865 280204 114970 280234
rect 115235 280286 115340 280311
rect 115235 280234 115262 280286
rect 115314 280234 115340 280286
rect 115235 280204 115340 280234
rect 115415 280283 115485 280351
rect 116015 280323 116063 280357
rect 116097 280323 116103 280357
rect 116015 280285 116103 280323
rect 112970 280192 114070 280198
rect 112970 280158 112999 280192
rect 113033 280158 113071 280192
rect 113105 280158 113143 280192
rect 113177 280158 113215 280192
rect 113249 280158 113287 280192
rect 113321 280158 113359 280192
rect 113393 280158 113431 280192
rect 113465 280158 113503 280192
rect 113537 280158 113575 280192
rect 113609 280158 113647 280192
rect 113681 280158 113719 280192
rect 113753 280158 113791 280192
rect 113825 280158 113863 280192
rect 113897 280158 113935 280192
rect 113969 280158 114007 280192
rect 114041 280158 114070 280192
rect 112970 280152 114070 280158
rect 111404 280073 111492 280096
rect 111404 280039 111452 280073
rect 111486 280039 111492 280073
rect 111404 280001 111492 280039
rect 111404 279967 111452 280001
rect 111486 279967 111492 280001
rect 111404 279944 111492 279967
rect 112656 280073 112744 280096
rect 114308 280084 114343 280199
rect 114720 280169 114790 280199
rect 115415 280199 115897 280283
rect 116015 280251 116063 280285
rect 116097 280251 116103 280285
rect 116015 280208 116103 280251
rect 117267 280364 117355 280400
rect 117461 280399 117509 280412
rect 117543 280399 117549 280433
rect 117461 280364 117549 280399
rect 117267 280361 117549 280364
rect 117267 280357 117509 280361
rect 117267 280323 117273 280357
rect 117307 280327 117509 280357
rect 117543 280327 117549 280361
rect 117307 280323 117549 280327
rect 117267 280304 117549 280323
rect 118713 280433 118801 280456
rect 118713 280399 118719 280433
rect 118753 280399 118801 280433
rect 118713 280361 118801 280399
rect 118713 280327 118719 280361
rect 118753 280327 118801 280361
rect 118713 280304 118801 280327
rect 117267 280302 117503 280304
rect 117267 280285 117355 280302
rect 117267 280251 117273 280285
rect 117307 280251 117355 280285
rect 117267 280208 117355 280251
rect 115415 280169 115485 280199
rect 114657 280163 114857 280169
rect 114657 280129 114704 280163
rect 114738 280129 114776 280163
rect 114810 280129 114857 280163
rect 114657 280123 114857 280129
rect 115348 280163 115548 280169
rect 115348 280129 115395 280163
rect 115429 280129 115467 280163
rect 115501 280129 115548 280163
rect 115348 280123 115548 280129
rect 112656 280039 112662 280073
rect 112696 280039 112744 280073
rect 113843 280054 114343 280084
rect 112656 280001 112744 280039
rect 113000 280048 114343 280054
rect 113000 280014 113029 280048
rect 113063 280014 113101 280048
rect 113135 280014 113173 280048
rect 113207 280014 113245 280048
rect 113279 280014 113317 280048
rect 113351 280014 113389 280048
rect 113423 280014 113461 280048
rect 113495 280014 113533 280048
rect 113567 280014 113605 280048
rect 113639 280014 113677 280048
rect 113711 280014 113749 280048
rect 113783 280014 113821 280048
rect 113855 280014 113893 280048
rect 113927 280014 113965 280048
rect 113999 280014 114037 280048
rect 114071 280043 114343 280048
rect 114570 280090 114616 280113
rect 114570 280056 114576 280090
rect 114610 280056 114616 280090
rect 114071 280014 114100 280043
rect 113000 280008 114100 280014
rect 114570 280018 114616 280056
rect 112656 279967 112662 280001
rect 112696 279967 112744 280001
rect 112656 279944 112744 279967
rect 111404 279736 111446 279944
rect 111524 279928 112624 279934
rect 111524 279894 111553 279928
rect 111587 279894 111625 279928
rect 111659 279894 111697 279928
rect 111731 279894 111769 279928
rect 111803 279894 111841 279928
rect 111875 279894 111913 279928
rect 111947 279894 111985 279928
rect 112019 279894 112057 279928
rect 112091 279894 112129 279928
rect 112163 279894 112201 279928
rect 112235 279894 112273 279928
rect 112307 279894 112345 279928
rect 112379 279894 112417 279928
rect 112451 279894 112489 279928
rect 112523 279894 112561 279928
rect 112595 279894 112624 279928
rect 111524 279888 112624 279894
rect 111524 279786 112624 279792
rect 111524 279752 111553 279786
rect 111587 279752 111625 279786
rect 111659 279752 111697 279786
rect 111731 279752 111769 279786
rect 111803 279752 111841 279786
rect 111875 279752 111913 279786
rect 111947 279752 111985 279786
rect 112019 279752 112057 279786
rect 112091 279752 112129 279786
rect 112163 279752 112201 279786
rect 112235 279752 112273 279786
rect 112307 279752 112345 279786
rect 112379 279752 112417 279786
rect 112451 279752 112489 279786
rect 112523 279752 112561 279786
rect 112595 279752 112624 279786
rect 111524 279746 112624 279752
rect 112702 279736 112744 279944
rect 111404 279713 111492 279736
rect 111404 279679 111452 279713
rect 111486 279679 111492 279713
rect 111404 279641 111492 279679
rect 111404 279607 111452 279641
rect 111486 279607 111492 279641
rect 111404 279584 111492 279607
rect 112656 279713 112744 279736
rect 112656 279679 112662 279713
rect 112696 279679 112744 279713
rect 112656 279641 112744 279679
rect 112656 279607 112662 279641
rect 112696 279607 112744 279641
rect 112656 279584 112744 279607
rect 112874 279979 112968 279998
rect 112874 279945 112928 279979
rect 112962 279945 112968 279979
rect 112874 279926 112968 279945
rect 114132 279979 114226 279998
rect 114132 279945 114138 279979
rect 114172 279945 114226 279979
rect 114132 279926 114226 279945
rect 112874 279834 112922 279926
rect 113000 279910 114100 279916
rect 113000 279876 113029 279910
rect 113063 279876 113101 279910
rect 113135 279876 113173 279910
rect 113207 279876 113245 279910
rect 113279 279876 113317 279910
rect 113351 279876 113389 279910
rect 113423 279876 113461 279910
rect 113495 279876 113533 279910
rect 113567 279876 113605 279910
rect 113639 279876 113677 279910
rect 113711 279876 113749 279910
rect 113783 279876 113821 279910
rect 113855 279876 113893 279910
rect 113927 279876 113965 279910
rect 113999 279876 114037 279910
rect 114071 279876 114100 279910
rect 113000 279870 114100 279876
rect 114178 279834 114226 279926
rect 112874 279790 114226 279834
rect 114324 279951 114396 279992
rect 114570 279984 114576 280018
rect 114610 279984 114616 280018
rect 114570 279961 114616 279984
rect 114898 280090 114944 280113
rect 114898 280056 114904 280090
rect 114938 280056 114944 280090
rect 114898 280018 114944 280056
rect 114898 279984 114904 280018
rect 114938 279984 114944 280018
rect 114898 279961 114944 279984
rect 115261 280090 115307 280113
rect 115261 280056 115267 280090
rect 115301 280056 115307 280090
rect 115261 280018 115307 280056
rect 115261 279984 115267 280018
rect 115301 279984 115307 280018
rect 115261 279961 115307 279984
rect 115589 280090 115635 280113
rect 115589 280056 115595 280090
rect 115629 280056 115635 280090
rect 115589 280018 115635 280056
rect 115862 280084 115897 280199
rect 116135 280192 117235 280198
rect 116135 280158 116164 280192
rect 116198 280158 116236 280192
rect 116270 280158 116308 280192
rect 116342 280158 116380 280192
rect 116414 280158 116452 280192
rect 116486 280158 116524 280192
rect 116558 280158 116596 280192
rect 116630 280158 116668 280192
rect 116702 280158 116740 280192
rect 116774 280158 116812 280192
rect 116846 280158 116884 280192
rect 116918 280158 116956 280192
rect 116990 280158 117028 280192
rect 117062 280158 117100 280192
rect 117134 280158 117172 280192
rect 117206 280158 117235 280192
rect 116135 280152 117235 280158
rect 117461 280096 117503 280302
rect 117581 280288 118681 280294
rect 117581 280254 117610 280288
rect 117644 280254 117682 280288
rect 117716 280254 117754 280288
rect 117788 280254 117826 280288
rect 117860 280254 117898 280288
rect 117932 280254 117970 280288
rect 118004 280254 118042 280288
rect 118076 280254 118114 280288
rect 118148 280254 118186 280288
rect 118220 280254 118258 280288
rect 118292 280254 118330 280288
rect 118364 280254 118402 280288
rect 118436 280254 118474 280288
rect 118508 280254 118546 280288
rect 118580 280254 118618 280288
rect 118652 280254 118681 280288
rect 117581 280248 118681 280254
rect 117581 280146 118681 280152
rect 117581 280112 117610 280146
rect 117644 280112 117682 280146
rect 117716 280112 117754 280146
rect 117788 280112 117826 280146
rect 117860 280112 117898 280146
rect 117932 280112 117970 280146
rect 118004 280112 118042 280146
rect 118076 280112 118114 280146
rect 118148 280112 118186 280146
rect 118220 280112 118258 280146
rect 118292 280112 118330 280146
rect 118364 280112 118402 280146
rect 118436 280112 118474 280146
rect 118508 280112 118546 280146
rect 118580 280112 118618 280146
rect 118652 280112 118681 280146
rect 117581 280106 118681 280112
rect 118759 280096 118801 280304
rect 115862 280054 116362 280084
rect 117461 280073 117549 280096
rect 115862 280048 117205 280054
rect 115862 280043 116134 280048
rect 115589 279984 115595 280018
rect 115629 279984 115635 280018
rect 116105 280014 116134 280043
rect 116168 280014 116206 280048
rect 116240 280014 116278 280048
rect 116312 280014 116350 280048
rect 116384 280014 116422 280048
rect 116456 280014 116494 280048
rect 116528 280014 116566 280048
rect 116600 280014 116638 280048
rect 116672 280014 116710 280048
rect 116744 280014 116782 280048
rect 116816 280014 116854 280048
rect 116888 280014 116926 280048
rect 116960 280014 116998 280048
rect 117032 280014 117070 280048
rect 117104 280014 117142 280048
rect 117176 280014 117205 280048
rect 116105 280008 117205 280014
rect 117461 280039 117509 280073
rect 117543 280039 117549 280073
rect 117461 280001 117549 280039
rect 115589 279961 115635 279984
rect 115809 279951 115881 279992
rect 114324 279917 114342 279951
rect 114376 279917 114396 279951
rect 114324 279861 114396 279917
rect 114657 279945 114857 279951
rect 114657 279911 114704 279945
rect 114738 279911 114776 279945
rect 114810 279911 114857 279945
rect 114657 279905 114857 279911
rect 115348 279945 115548 279951
rect 115348 279911 115395 279945
rect 115429 279911 115467 279945
rect 115501 279911 115548 279945
rect 115348 279905 115548 279911
rect 115809 279917 115828 279951
rect 115862 279917 115881 279951
rect 114843 279861 115030 279876
rect 114324 279816 114781 279861
rect 112874 279700 112922 279790
rect 113000 279750 114100 279756
rect 113000 279716 113029 279750
rect 113063 279716 113101 279750
rect 113135 279716 113173 279750
rect 113207 279716 113245 279750
rect 113279 279716 113317 279750
rect 113351 279716 113389 279750
rect 113423 279716 113461 279750
rect 113495 279716 113533 279750
rect 113567 279716 113605 279750
rect 113639 279716 113677 279750
rect 113711 279716 113749 279750
rect 113783 279716 113821 279750
rect 113855 279716 113893 279750
rect 113927 279716 113965 279750
rect 113999 279716 114037 279750
rect 114071 279716 114100 279750
rect 113000 279710 114100 279716
rect 114178 279700 114226 279790
rect 114737 279761 114781 279816
rect 114843 279809 114891 279861
rect 114943 279809 115030 279861
rect 114843 279791 115030 279809
rect 115175 279861 115362 279876
rect 115809 279861 115881 279917
rect 115175 279809 115262 279861
rect 115314 279809 115362 279861
rect 115175 279791 115362 279809
rect 115424 279816 115881 279861
rect 115979 279979 116073 279998
rect 115979 279945 116033 279979
rect 116067 279945 116073 279979
rect 115979 279926 116073 279945
rect 117237 279979 117331 279998
rect 117237 279945 117243 279979
rect 117277 279945 117331 279979
rect 117237 279926 117331 279945
rect 115979 279834 116027 279926
rect 116105 279910 117205 279916
rect 116105 279876 116134 279910
rect 116168 279876 116206 279910
rect 116240 279876 116278 279910
rect 116312 279876 116350 279910
rect 116384 279876 116422 279910
rect 116456 279876 116494 279910
rect 116528 279876 116566 279910
rect 116600 279876 116638 279910
rect 116672 279876 116710 279910
rect 116744 279876 116782 279910
rect 116816 279876 116854 279910
rect 116888 279876 116926 279910
rect 116960 279876 116998 279910
rect 117032 279876 117070 279910
rect 117104 279876 117142 279910
rect 117176 279876 117205 279910
rect 116105 279870 117205 279876
rect 117283 279834 117331 279926
rect 115424 279761 115468 279816
rect 115979 279790 117331 279834
rect 114657 279755 114857 279761
rect 114657 279721 114704 279755
rect 114738 279721 114776 279755
rect 114810 279721 114857 279755
rect 114657 279715 114857 279721
rect 115348 279755 115548 279761
rect 115348 279721 115395 279755
rect 115429 279721 115467 279755
rect 115501 279721 115548 279755
rect 115348 279715 115548 279721
rect 112874 279681 112968 279700
rect 112874 279647 112928 279681
rect 112962 279647 112968 279681
rect 112874 279628 112968 279647
rect 114132 279681 114226 279700
rect 114132 279647 114138 279681
rect 114172 279647 114226 279681
rect 114132 279628 114226 279647
rect 114570 279682 114616 279705
rect 114570 279648 114576 279682
rect 114610 279648 114616 279682
rect 111524 279568 112624 279574
rect 111524 279534 111553 279568
rect 111587 279534 111625 279568
rect 111659 279534 111697 279568
rect 111731 279534 111769 279568
rect 111803 279534 111841 279568
rect 111875 279534 111913 279568
rect 111947 279534 111985 279568
rect 112019 279534 112057 279568
rect 112091 279534 112129 279568
rect 112163 279534 112201 279568
rect 112235 279534 112273 279568
rect 112307 279534 112345 279568
rect 112379 279534 112417 279568
rect 112451 279534 112489 279568
rect 112523 279534 112561 279568
rect 112595 279534 112624 279568
rect 111524 279530 112624 279534
rect 112874 279534 112922 279628
rect 114327 279623 114395 279624
rect 114570 279623 114616 279648
rect 113000 279612 114100 279618
rect 113000 279578 113029 279612
rect 113063 279578 113101 279612
rect 113135 279578 113173 279612
rect 113207 279578 113245 279612
rect 113279 279578 113317 279612
rect 113351 279578 113389 279612
rect 113423 279578 113461 279612
rect 113495 279578 113533 279612
rect 113567 279578 113605 279612
rect 113639 279578 113677 279612
rect 113711 279578 113749 279612
rect 113783 279578 113821 279612
rect 113855 279578 113893 279612
rect 113927 279578 113965 279612
rect 113999 279578 114037 279612
rect 114071 279578 114100 279612
rect 113000 279572 114100 279578
rect 114327 279610 114616 279623
rect 114327 279576 114576 279610
rect 114610 279576 114616 279610
rect 114327 279563 114616 279576
rect 114327 279534 114395 279563
rect 114570 279553 114616 279563
rect 114898 279682 114944 279705
rect 114898 279648 114904 279682
rect 114938 279648 114944 279682
rect 114898 279610 114944 279648
rect 114898 279576 114904 279610
rect 114938 279576 114944 279610
rect 114898 279553 114944 279576
rect 115261 279682 115307 279705
rect 115261 279648 115267 279682
rect 115301 279648 115307 279682
rect 115261 279610 115307 279648
rect 115261 279576 115267 279610
rect 115301 279576 115307 279610
rect 115261 279553 115307 279576
rect 115589 279682 115635 279705
rect 115589 279648 115595 279682
rect 115629 279648 115635 279682
rect 115589 279623 115635 279648
rect 115979 279700 116027 279790
rect 116105 279750 117205 279756
rect 116105 279716 116134 279750
rect 116168 279716 116206 279750
rect 116240 279716 116278 279750
rect 116312 279716 116350 279750
rect 116384 279716 116422 279750
rect 116456 279716 116494 279750
rect 116528 279716 116566 279750
rect 116600 279716 116638 279750
rect 116672 279716 116710 279750
rect 116744 279716 116782 279750
rect 116816 279716 116854 279750
rect 116888 279716 116926 279750
rect 116960 279716 116998 279750
rect 117032 279716 117070 279750
rect 117104 279716 117142 279750
rect 117176 279716 117205 279750
rect 116105 279710 117205 279716
rect 117283 279700 117331 279790
rect 115979 279681 116073 279700
rect 115979 279647 116033 279681
rect 116067 279647 116073 279681
rect 115979 279628 116073 279647
rect 117237 279681 117331 279700
rect 117237 279647 117243 279681
rect 117277 279647 117331 279681
rect 117237 279628 117331 279647
rect 115810 279623 115878 279624
rect 115589 279610 115878 279623
rect 115589 279576 115595 279610
rect 115629 279576 115878 279610
rect 115589 279563 115878 279576
rect 116105 279612 117205 279618
rect 116105 279578 116134 279612
rect 116168 279578 116206 279612
rect 116240 279578 116278 279612
rect 116312 279578 116350 279612
rect 116384 279578 116422 279612
rect 116456 279578 116494 279612
rect 116528 279578 116566 279612
rect 116600 279578 116638 279612
rect 116672 279578 116710 279612
rect 116744 279578 116782 279612
rect 116816 279578 116854 279612
rect 116888 279578 116926 279612
rect 116960 279578 116998 279612
rect 117032 279578 117070 279612
rect 117104 279578 117142 279612
rect 117176 279578 117205 279612
rect 116105 279572 117205 279578
rect 115589 279553 115635 279563
rect 112874 279530 114395 279534
rect 111524 279528 114395 279530
rect 112044 279494 114395 279528
rect 114657 279537 114857 279543
rect 114657 279503 114704 279537
rect 114738 279503 114776 279537
rect 114810 279503 114857 279537
rect 114657 279497 114857 279503
rect 115348 279537 115548 279543
rect 115348 279503 115395 279537
rect 115429 279503 115467 279537
rect 115501 279503 115548 279537
rect 115348 279497 115548 279503
rect 115810 279534 115878 279563
rect 117283 279534 117331 279628
rect 117461 279967 117509 280001
rect 117543 279967 117549 280001
rect 117461 279944 117549 279967
rect 118713 280073 118801 280096
rect 118713 280039 118719 280073
rect 118753 280039 118801 280073
rect 118713 280001 118801 280039
rect 118713 279967 118719 280001
rect 118753 279967 118801 280001
rect 118713 279944 118801 279967
rect 117461 279736 117503 279944
rect 117581 279928 118681 279934
rect 117581 279894 117610 279928
rect 117644 279894 117682 279928
rect 117716 279894 117754 279928
rect 117788 279894 117826 279928
rect 117860 279894 117898 279928
rect 117932 279894 117970 279928
rect 118004 279894 118042 279928
rect 118076 279894 118114 279928
rect 118148 279894 118186 279928
rect 118220 279894 118258 279928
rect 118292 279894 118330 279928
rect 118364 279894 118402 279928
rect 118436 279894 118474 279928
rect 118508 279894 118546 279928
rect 118580 279894 118618 279928
rect 118652 279894 118681 279928
rect 117581 279888 118681 279894
rect 117581 279786 118681 279792
rect 117581 279752 117610 279786
rect 117644 279752 117682 279786
rect 117716 279752 117754 279786
rect 117788 279752 117826 279786
rect 117860 279752 117898 279786
rect 117932 279752 117970 279786
rect 118004 279752 118042 279786
rect 118076 279752 118114 279786
rect 118148 279752 118186 279786
rect 118220 279752 118258 279786
rect 118292 279752 118330 279786
rect 118364 279752 118402 279786
rect 118436 279752 118474 279786
rect 118508 279752 118546 279786
rect 118580 279752 118618 279786
rect 118652 279752 118681 279786
rect 117581 279746 118681 279752
rect 118759 279736 118801 279944
rect 117461 279713 117549 279736
rect 117461 279679 117509 279713
rect 117543 279679 117549 279713
rect 117461 279641 117549 279679
rect 117461 279607 117509 279641
rect 117543 279607 117549 279641
rect 117461 279584 117549 279607
rect 118713 279713 118801 279736
rect 118713 279679 118719 279713
rect 118753 279679 118801 279713
rect 118713 279641 118801 279679
rect 118713 279607 118719 279641
rect 118753 279607 118801 279641
rect 118713 279584 118801 279607
rect 115810 279530 117331 279534
rect 117581 279568 118681 279574
rect 117581 279534 117610 279568
rect 117644 279534 117682 279568
rect 117716 279534 117754 279568
rect 117788 279534 117826 279568
rect 117860 279534 117898 279568
rect 117932 279534 117970 279568
rect 118004 279534 118042 279568
rect 118076 279534 118114 279568
rect 118148 279534 118186 279568
rect 118220 279534 118258 279568
rect 118292 279534 118330 279568
rect 118364 279534 118402 279568
rect 118436 279534 118474 279568
rect 118508 279534 118546 279568
rect 118580 279534 118618 279568
rect 118652 279534 118681 279568
rect 117581 279530 118681 279534
rect 115810 279528 118681 279530
rect 112719 279452 112924 279494
rect 113982 279420 114266 279430
rect 114724 279420 114783 279497
rect 113982 279399 114783 279420
rect 113982 279365 114034 279399
rect 114068 279365 114106 279399
rect 114140 279365 114178 279399
rect 114212 279365 114783 279399
rect 113982 279331 114783 279365
rect 115422 279420 115481 279497
rect 115810 279494 118161 279528
rect 117281 279452 117486 279494
rect 115939 279420 116223 279430
rect 115422 279399 116223 279420
rect 115422 279365 115992 279399
rect 116026 279365 116064 279399
rect 116098 279365 116136 279399
rect 116170 279365 116223 279399
rect 115422 279331 116223 279365
rect 113982 279330 114266 279331
rect 115939 279330 116223 279331
rect 112970 279208 114070 279214
rect 111524 279200 112624 279206
rect 111524 279166 111553 279200
rect 111587 279166 111625 279200
rect 111659 279166 111697 279200
rect 111731 279166 111769 279200
rect 111803 279166 111841 279200
rect 111875 279166 111913 279200
rect 111947 279166 111985 279200
rect 112019 279166 112057 279200
rect 112091 279166 112129 279200
rect 112163 279166 112201 279200
rect 112235 279166 112273 279200
rect 112307 279166 112345 279200
rect 112379 279166 112417 279200
rect 112451 279166 112489 279200
rect 112523 279166 112561 279200
rect 112595 279166 112624 279200
rect 112970 279174 112999 279208
rect 113033 279174 113071 279208
rect 113105 279174 113143 279208
rect 113177 279174 113215 279208
rect 113249 279174 113287 279208
rect 113321 279174 113359 279208
rect 113393 279174 113431 279208
rect 113465 279174 113503 279208
rect 113537 279174 113575 279208
rect 113609 279174 113647 279208
rect 113681 279174 113719 279208
rect 113753 279174 113791 279208
rect 113825 279174 113863 279208
rect 113897 279174 113935 279208
rect 113969 279174 114007 279208
rect 114041 279174 114070 279208
rect 116135 279208 117235 279214
rect 112970 279168 114070 279174
rect 114657 279183 114857 279189
rect 111524 279160 112624 279166
rect 111404 279127 111492 279150
rect 111404 279093 111452 279127
rect 111486 279093 111492 279127
rect 111404 279055 111492 279093
rect 111404 279021 111452 279055
rect 111486 279021 111492 279055
rect 111404 278998 111492 279021
rect 112656 279127 112744 279150
rect 112656 279093 112662 279127
rect 112696 279093 112744 279127
rect 112656 279082 112744 279093
rect 112850 279115 112938 279158
rect 112850 279082 112898 279115
rect 112656 279081 112898 279082
rect 112932 279081 112938 279115
rect 112656 279055 112938 279081
rect 112656 279021 112662 279055
rect 112696 279043 112938 279055
rect 112696 279021 112898 279043
rect 112656 279020 112898 279021
rect 112656 278998 112744 279020
rect 111404 278790 111446 278998
rect 111524 278982 112624 278988
rect 111524 278948 111553 278982
rect 111587 278948 111625 278982
rect 111659 278948 111697 278982
rect 111731 278948 111769 278982
rect 111803 278948 111841 278982
rect 111875 278948 111913 278982
rect 111947 278948 111985 278982
rect 112019 278948 112057 278982
rect 112091 278948 112129 278982
rect 112163 278948 112201 278982
rect 112235 278948 112273 278982
rect 112307 278948 112345 278982
rect 112379 278948 112417 278982
rect 112451 278948 112489 278982
rect 112523 278948 112561 278982
rect 112595 278948 112624 278982
rect 111524 278942 112624 278948
rect 112702 278966 112744 278998
rect 112850 279009 112898 279020
rect 112932 279009 112938 279043
rect 112850 278966 112938 279009
rect 114102 279115 114190 279158
rect 114657 279149 114704 279183
rect 114738 279149 114776 279183
rect 114810 279149 114857 279183
rect 114657 279143 114857 279149
rect 115348 279183 115548 279189
rect 115348 279149 115395 279183
rect 115429 279149 115467 279183
rect 115501 279149 115548 279183
rect 116135 279174 116164 279208
rect 116198 279174 116236 279208
rect 116270 279174 116308 279208
rect 116342 279174 116380 279208
rect 116414 279174 116452 279208
rect 116486 279174 116524 279208
rect 116558 279174 116596 279208
rect 116630 279174 116668 279208
rect 116702 279174 116740 279208
rect 116774 279174 116812 279208
rect 116846 279174 116884 279208
rect 116918 279174 116956 279208
rect 116990 279174 117028 279208
rect 117062 279174 117100 279208
rect 117134 279174 117172 279208
rect 117206 279174 117235 279208
rect 116135 279168 117235 279174
rect 117581 279200 118681 279206
rect 117581 279166 117610 279200
rect 117644 279166 117682 279200
rect 117716 279166 117754 279200
rect 117788 279166 117826 279200
rect 117860 279166 117898 279200
rect 117932 279166 117970 279200
rect 118004 279166 118042 279200
rect 118076 279166 118114 279200
rect 118148 279166 118186 279200
rect 118220 279166 118258 279200
rect 118292 279166 118330 279200
rect 118364 279166 118402 279200
rect 118436 279166 118474 279200
rect 118508 279166 118546 279200
rect 118580 279166 118618 279200
rect 118652 279166 118681 279200
rect 117581 279160 118681 279166
rect 115348 279143 115548 279149
rect 114102 279081 114108 279115
rect 114142 279092 114190 279115
rect 114570 279098 114616 279133
rect 114570 279092 114576 279098
rect 114142 279081 114576 279092
rect 114102 279064 114576 279081
rect 114610 279064 114616 279098
rect 114102 279043 114616 279064
rect 114102 279009 114108 279043
rect 114142 279026 114616 279043
rect 114142 279009 114576 279026
rect 114102 278992 114576 279009
rect 114610 278992 114616 279026
rect 114102 278966 114616 278992
rect 111524 278840 112624 278846
rect 111524 278806 111553 278840
rect 111587 278806 111625 278840
rect 111659 278806 111697 278840
rect 111731 278806 111769 278840
rect 111803 278806 111841 278840
rect 111875 278806 111913 278840
rect 111947 278806 111985 278840
rect 112019 278806 112057 278840
rect 112091 278806 112129 278840
rect 112163 278806 112201 278840
rect 112235 278806 112273 278840
rect 112307 278806 112345 278840
rect 112379 278806 112417 278840
rect 112451 278806 112489 278840
rect 112523 278806 112561 278840
rect 112595 278806 112624 278840
rect 111524 278800 112624 278806
rect 112702 278790 112746 278966
rect 111404 278767 111492 278790
rect 111404 278733 111452 278767
rect 111486 278733 111492 278767
rect 111404 278695 111492 278733
rect 111404 278661 111452 278695
rect 111486 278661 111492 278695
rect 111404 278638 111492 278661
rect 112656 278767 112746 278790
rect 112656 278733 112662 278767
rect 112696 278746 112746 278767
rect 112850 278866 112892 278966
rect 114148 278959 114616 278966
rect 112970 278950 114070 278956
rect 112970 278916 112999 278950
rect 113033 278916 113071 278950
rect 113105 278916 113143 278950
rect 113177 278916 113215 278950
rect 113249 278916 113287 278950
rect 113321 278916 113359 278950
rect 113393 278916 113431 278950
rect 113465 278916 113503 278950
rect 113537 278916 113575 278950
rect 113609 278916 113647 278950
rect 113681 278916 113719 278950
rect 113753 278916 113791 278950
rect 113825 278916 113863 278950
rect 113897 278916 113935 278950
rect 113969 278916 114007 278950
rect 114041 278916 114070 278950
rect 112970 278910 114070 278916
rect 114148 278866 114190 278959
rect 112850 278828 114190 278866
rect 112696 278733 112744 278746
rect 112656 278698 112744 278733
rect 112850 278734 112892 278828
rect 112970 278784 114070 278790
rect 112970 278750 112999 278784
rect 113033 278750 113071 278784
rect 113105 278750 113143 278784
rect 113177 278750 113215 278784
rect 113249 278750 113287 278784
rect 113321 278750 113359 278784
rect 113393 278750 113431 278784
rect 113465 278750 113503 278784
rect 113537 278750 113575 278784
rect 113609 278750 113647 278784
rect 113681 278750 113719 278784
rect 113753 278750 113791 278784
rect 113825 278750 113863 278784
rect 113897 278750 113935 278784
rect 113969 278750 114007 278784
rect 114041 278750 114070 278784
rect 112970 278744 114070 278750
rect 114148 278734 114190 278828
rect 114570 278954 114616 278959
rect 114570 278920 114576 278954
rect 114610 278920 114616 278954
rect 114570 278882 114616 278920
rect 114570 278848 114576 278882
rect 114610 278848 114616 278882
rect 114570 278810 114616 278848
rect 114570 278776 114576 278810
rect 114610 278776 114616 278810
rect 114570 278741 114616 278776
rect 114898 279098 114944 279133
rect 114898 279064 114904 279098
rect 114938 279064 114944 279098
rect 114898 279026 114944 279064
rect 114898 278992 114904 279026
rect 114938 278992 114944 279026
rect 114898 278954 114944 278992
rect 114898 278920 114904 278954
rect 114938 278920 114944 278954
rect 114898 278882 114944 278920
rect 114898 278848 114904 278882
rect 114938 278848 114944 278882
rect 114898 278810 114944 278848
rect 114898 278776 114904 278810
rect 114938 278776 114944 278810
rect 114898 278741 114944 278776
rect 115261 279098 115307 279133
rect 115261 279064 115267 279098
rect 115301 279064 115307 279098
rect 115261 279026 115307 279064
rect 115261 278992 115267 279026
rect 115301 278992 115307 279026
rect 115261 278954 115307 278992
rect 115261 278920 115267 278954
rect 115301 278920 115307 278954
rect 115261 278882 115307 278920
rect 115261 278848 115267 278882
rect 115301 278848 115307 278882
rect 115261 278810 115307 278848
rect 115261 278776 115267 278810
rect 115301 278776 115307 278810
rect 115261 278741 115307 278776
rect 115589 279098 115635 279133
rect 115589 279064 115595 279098
rect 115629 279092 115635 279098
rect 116015 279115 116103 279158
rect 116015 279092 116063 279115
rect 115629 279081 116063 279092
rect 116097 279081 116103 279115
rect 115629 279064 116103 279081
rect 115589 279043 116103 279064
rect 115589 279026 116063 279043
rect 115589 278992 115595 279026
rect 115629 279009 116063 279026
rect 116097 279009 116103 279043
rect 115629 278992 116103 279009
rect 115589 278966 116103 278992
rect 117267 279115 117355 279158
rect 117267 279081 117273 279115
rect 117307 279082 117355 279115
rect 117461 279127 117549 279150
rect 117461 279093 117509 279127
rect 117543 279093 117549 279127
rect 117461 279082 117549 279093
rect 117307 279081 117549 279082
rect 117267 279055 117549 279081
rect 117267 279043 117509 279055
rect 117267 279009 117273 279043
rect 117307 279021 117509 279043
rect 117543 279021 117549 279055
rect 117307 279020 117549 279021
rect 117307 279009 117355 279020
rect 117267 278966 117355 279009
rect 117461 278998 117549 279020
rect 118713 279127 118801 279150
rect 118713 279093 118719 279127
rect 118753 279093 118801 279127
rect 118713 279055 118801 279093
rect 118713 279021 118719 279055
rect 118753 279021 118801 279055
rect 118713 278998 118801 279021
rect 117461 278966 117503 278998
rect 115589 278959 116057 278966
rect 115589 278954 115635 278959
rect 115589 278920 115595 278954
rect 115629 278920 115635 278954
rect 115589 278882 115635 278920
rect 115589 278848 115595 278882
rect 115629 278848 115635 278882
rect 115589 278810 115635 278848
rect 115589 278776 115595 278810
rect 115629 278776 115635 278810
rect 115589 278741 115635 278776
rect 116015 278866 116057 278959
rect 116135 278950 117235 278956
rect 116135 278916 116164 278950
rect 116198 278916 116236 278950
rect 116270 278916 116308 278950
rect 116342 278916 116380 278950
rect 116414 278916 116452 278950
rect 116486 278916 116524 278950
rect 116558 278916 116596 278950
rect 116630 278916 116668 278950
rect 116702 278916 116740 278950
rect 116774 278916 116812 278950
rect 116846 278916 116884 278950
rect 116918 278916 116956 278950
rect 116990 278916 117028 278950
rect 117062 278916 117100 278950
rect 117134 278916 117172 278950
rect 117206 278916 117235 278950
rect 116135 278910 117235 278916
rect 117313 278866 117355 278966
rect 116015 278828 117355 278866
rect 112850 278698 112938 278734
rect 112656 278695 112938 278698
rect 112656 278661 112662 278695
rect 112696 278691 112938 278695
rect 112696 278661 112898 278691
rect 112656 278657 112898 278661
rect 112932 278657 112938 278691
rect 112656 278638 112938 278657
rect 111404 278430 111446 278638
rect 112702 278636 112938 278638
rect 111524 278622 112624 278628
rect 111524 278588 111553 278622
rect 111587 278588 111625 278622
rect 111659 278588 111697 278622
rect 111731 278588 111769 278622
rect 111803 278588 111841 278622
rect 111875 278588 111913 278622
rect 111947 278588 111985 278622
rect 112019 278588 112057 278622
rect 112091 278588 112129 278622
rect 112163 278588 112201 278622
rect 112235 278588 112273 278622
rect 112307 278588 112345 278622
rect 112379 278588 112417 278622
rect 112451 278588 112489 278622
rect 112523 278588 112561 278622
rect 112595 278588 112624 278622
rect 111524 278582 112624 278588
rect 111524 278480 112624 278486
rect 111524 278446 111553 278480
rect 111587 278446 111625 278480
rect 111659 278446 111697 278480
rect 111731 278446 111769 278480
rect 111803 278446 111841 278480
rect 111875 278446 111913 278480
rect 111947 278446 111985 278480
rect 112019 278446 112057 278480
rect 112091 278446 112129 278480
rect 112163 278446 112201 278480
rect 112235 278446 112273 278480
rect 112307 278446 112345 278480
rect 112379 278446 112417 278480
rect 112451 278446 112489 278480
rect 112523 278446 112561 278480
rect 112595 278446 112624 278480
rect 111524 278440 112624 278446
rect 112702 278430 112744 278636
rect 112850 278619 112938 278636
rect 112850 278585 112898 278619
rect 112932 278585 112938 278619
rect 112850 278542 112938 278585
rect 114102 278691 114190 278734
rect 116015 278734 116057 278828
rect 116135 278784 117235 278790
rect 116135 278750 116164 278784
rect 116198 278750 116236 278784
rect 116270 278750 116308 278784
rect 116342 278750 116380 278784
rect 116414 278750 116452 278784
rect 116486 278750 116524 278784
rect 116558 278750 116596 278784
rect 116630 278750 116668 278784
rect 116702 278750 116740 278784
rect 116774 278750 116812 278784
rect 116846 278750 116884 278784
rect 116918 278750 116956 278784
rect 116990 278750 117028 278784
rect 117062 278750 117100 278784
rect 117134 278750 117172 278784
rect 117206 278750 117235 278784
rect 116135 278744 117235 278750
rect 117313 278734 117355 278828
rect 117459 278790 117503 278966
rect 117581 278982 118681 278988
rect 117581 278948 117610 278982
rect 117644 278948 117682 278982
rect 117716 278948 117754 278982
rect 117788 278948 117826 278982
rect 117860 278948 117898 278982
rect 117932 278948 117970 278982
rect 118004 278948 118042 278982
rect 118076 278948 118114 278982
rect 118148 278948 118186 278982
rect 118220 278948 118258 278982
rect 118292 278948 118330 278982
rect 118364 278948 118402 278982
rect 118436 278948 118474 278982
rect 118508 278948 118546 278982
rect 118580 278948 118618 278982
rect 118652 278948 118681 278982
rect 117581 278942 118681 278948
rect 117581 278840 118681 278846
rect 117581 278806 117610 278840
rect 117644 278806 117682 278840
rect 117716 278806 117754 278840
rect 117788 278806 117826 278840
rect 117860 278806 117898 278840
rect 117932 278806 117970 278840
rect 118004 278806 118042 278840
rect 118076 278806 118114 278840
rect 118148 278806 118186 278840
rect 118220 278806 118258 278840
rect 118292 278806 118330 278840
rect 118364 278806 118402 278840
rect 118436 278806 118474 278840
rect 118508 278806 118546 278840
rect 118580 278806 118618 278840
rect 118652 278806 118681 278840
rect 117581 278800 118681 278806
rect 118759 278790 118801 278998
rect 117459 278767 117549 278790
rect 117459 278746 117509 278767
rect 114102 278657 114108 278691
rect 114142 278657 114190 278691
rect 114657 278725 114857 278731
rect 114657 278691 114704 278725
rect 114738 278691 114776 278725
rect 114810 278691 114857 278725
rect 114657 278685 114857 278691
rect 115348 278725 115548 278731
rect 115348 278691 115395 278725
rect 115429 278691 115467 278725
rect 115501 278691 115548 278725
rect 115348 278685 115548 278691
rect 116015 278691 116103 278734
rect 114102 278619 114190 278657
rect 114102 278585 114108 278619
rect 114142 278585 114190 278619
rect 114720 278617 114790 278685
rect 114102 278542 114190 278585
rect 114308 278533 114790 278617
rect 114865 278620 114970 278645
rect 114865 278568 114890 278620
rect 114942 278568 114970 278620
rect 114865 278538 114970 278568
rect 115235 278620 115340 278645
rect 115235 278568 115262 278620
rect 115314 278568 115340 278620
rect 115235 278538 115340 278568
rect 115415 278617 115485 278685
rect 116015 278657 116063 278691
rect 116097 278657 116103 278691
rect 116015 278619 116103 278657
rect 112970 278526 114070 278532
rect 112970 278492 112999 278526
rect 113033 278492 113071 278526
rect 113105 278492 113143 278526
rect 113177 278492 113215 278526
rect 113249 278492 113287 278526
rect 113321 278492 113359 278526
rect 113393 278492 113431 278526
rect 113465 278492 113503 278526
rect 113537 278492 113575 278526
rect 113609 278492 113647 278526
rect 113681 278492 113719 278526
rect 113753 278492 113791 278526
rect 113825 278492 113863 278526
rect 113897 278492 113935 278526
rect 113969 278492 114007 278526
rect 114041 278492 114070 278526
rect 112970 278486 114070 278492
rect 111404 278407 111492 278430
rect 111404 278373 111452 278407
rect 111486 278373 111492 278407
rect 111404 278335 111492 278373
rect 111404 278301 111452 278335
rect 111486 278301 111492 278335
rect 111404 278278 111492 278301
rect 112656 278407 112744 278430
rect 114308 278418 114343 278533
rect 114720 278503 114790 278533
rect 115415 278533 115897 278617
rect 116015 278585 116063 278619
rect 116097 278585 116103 278619
rect 116015 278542 116103 278585
rect 117267 278698 117355 278734
rect 117461 278733 117509 278746
rect 117543 278733 117549 278767
rect 117461 278698 117549 278733
rect 117267 278695 117549 278698
rect 117267 278691 117509 278695
rect 117267 278657 117273 278691
rect 117307 278661 117509 278691
rect 117543 278661 117549 278695
rect 117307 278657 117549 278661
rect 117267 278638 117549 278657
rect 118713 278767 118801 278790
rect 118713 278733 118719 278767
rect 118753 278733 118801 278767
rect 118713 278695 118801 278733
rect 118713 278661 118719 278695
rect 118753 278661 118801 278695
rect 118713 278638 118801 278661
rect 117267 278636 117503 278638
rect 117267 278619 117355 278636
rect 117267 278585 117273 278619
rect 117307 278585 117355 278619
rect 117267 278542 117355 278585
rect 115415 278503 115485 278533
rect 114657 278497 114857 278503
rect 114657 278463 114704 278497
rect 114738 278463 114776 278497
rect 114810 278463 114857 278497
rect 114657 278457 114857 278463
rect 115348 278497 115548 278503
rect 115348 278463 115395 278497
rect 115429 278463 115467 278497
rect 115501 278463 115548 278497
rect 115348 278457 115548 278463
rect 112656 278373 112662 278407
rect 112696 278373 112744 278407
rect 113843 278388 114343 278418
rect 112656 278335 112744 278373
rect 113000 278382 114343 278388
rect 113000 278348 113029 278382
rect 113063 278348 113101 278382
rect 113135 278348 113173 278382
rect 113207 278348 113245 278382
rect 113279 278348 113317 278382
rect 113351 278348 113389 278382
rect 113423 278348 113461 278382
rect 113495 278348 113533 278382
rect 113567 278348 113605 278382
rect 113639 278348 113677 278382
rect 113711 278348 113749 278382
rect 113783 278348 113821 278382
rect 113855 278348 113893 278382
rect 113927 278348 113965 278382
rect 113999 278348 114037 278382
rect 114071 278377 114343 278382
rect 114570 278424 114616 278447
rect 114570 278390 114576 278424
rect 114610 278390 114616 278424
rect 114071 278348 114100 278377
rect 113000 278342 114100 278348
rect 114570 278352 114616 278390
rect 112656 278301 112662 278335
rect 112696 278301 112744 278335
rect 112656 278278 112744 278301
rect 111404 278070 111446 278278
rect 111524 278262 112624 278268
rect 111524 278228 111553 278262
rect 111587 278228 111625 278262
rect 111659 278228 111697 278262
rect 111731 278228 111769 278262
rect 111803 278228 111841 278262
rect 111875 278228 111913 278262
rect 111947 278228 111985 278262
rect 112019 278228 112057 278262
rect 112091 278228 112129 278262
rect 112163 278228 112201 278262
rect 112235 278228 112273 278262
rect 112307 278228 112345 278262
rect 112379 278228 112417 278262
rect 112451 278228 112489 278262
rect 112523 278228 112561 278262
rect 112595 278228 112624 278262
rect 111524 278222 112624 278228
rect 111524 278120 112624 278126
rect 111524 278086 111553 278120
rect 111587 278086 111625 278120
rect 111659 278086 111697 278120
rect 111731 278086 111769 278120
rect 111803 278086 111841 278120
rect 111875 278086 111913 278120
rect 111947 278086 111985 278120
rect 112019 278086 112057 278120
rect 112091 278086 112129 278120
rect 112163 278086 112201 278120
rect 112235 278086 112273 278120
rect 112307 278086 112345 278120
rect 112379 278086 112417 278120
rect 112451 278086 112489 278120
rect 112523 278086 112561 278120
rect 112595 278086 112624 278120
rect 111524 278080 112624 278086
rect 112702 278070 112744 278278
rect 111404 278047 111492 278070
rect 111404 278013 111452 278047
rect 111486 278013 111492 278047
rect 111404 277975 111492 278013
rect 111404 277941 111452 277975
rect 111486 277941 111492 277975
rect 111404 277918 111492 277941
rect 112656 278047 112744 278070
rect 112656 278013 112662 278047
rect 112696 278013 112744 278047
rect 112656 277975 112744 278013
rect 112656 277941 112662 277975
rect 112696 277941 112744 277975
rect 112656 277918 112744 277941
rect 112874 278313 112968 278332
rect 112874 278279 112928 278313
rect 112962 278279 112968 278313
rect 112874 278260 112968 278279
rect 114132 278313 114226 278332
rect 114132 278279 114138 278313
rect 114172 278279 114226 278313
rect 114132 278260 114226 278279
rect 112874 278168 112922 278260
rect 113000 278244 114100 278250
rect 113000 278210 113029 278244
rect 113063 278210 113101 278244
rect 113135 278210 113173 278244
rect 113207 278210 113245 278244
rect 113279 278210 113317 278244
rect 113351 278210 113389 278244
rect 113423 278210 113461 278244
rect 113495 278210 113533 278244
rect 113567 278210 113605 278244
rect 113639 278210 113677 278244
rect 113711 278210 113749 278244
rect 113783 278210 113821 278244
rect 113855 278210 113893 278244
rect 113927 278210 113965 278244
rect 113999 278210 114037 278244
rect 114071 278210 114100 278244
rect 113000 278204 114100 278210
rect 114178 278168 114226 278260
rect 112874 278124 114226 278168
rect 114324 278285 114396 278326
rect 114570 278318 114576 278352
rect 114610 278318 114616 278352
rect 114570 278295 114616 278318
rect 114898 278424 114944 278447
rect 114898 278390 114904 278424
rect 114938 278390 114944 278424
rect 114898 278352 114944 278390
rect 114898 278318 114904 278352
rect 114938 278318 114944 278352
rect 114898 278295 114944 278318
rect 115261 278424 115307 278447
rect 115261 278390 115267 278424
rect 115301 278390 115307 278424
rect 115261 278352 115307 278390
rect 115261 278318 115267 278352
rect 115301 278318 115307 278352
rect 115261 278295 115307 278318
rect 115589 278424 115635 278447
rect 115589 278390 115595 278424
rect 115629 278390 115635 278424
rect 115589 278352 115635 278390
rect 115862 278418 115897 278533
rect 116135 278526 117235 278532
rect 116135 278492 116164 278526
rect 116198 278492 116236 278526
rect 116270 278492 116308 278526
rect 116342 278492 116380 278526
rect 116414 278492 116452 278526
rect 116486 278492 116524 278526
rect 116558 278492 116596 278526
rect 116630 278492 116668 278526
rect 116702 278492 116740 278526
rect 116774 278492 116812 278526
rect 116846 278492 116884 278526
rect 116918 278492 116956 278526
rect 116990 278492 117028 278526
rect 117062 278492 117100 278526
rect 117134 278492 117172 278526
rect 117206 278492 117235 278526
rect 116135 278486 117235 278492
rect 117461 278430 117503 278636
rect 117581 278622 118681 278628
rect 117581 278588 117610 278622
rect 117644 278588 117682 278622
rect 117716 278588 117754 278622
rect 117788 278588 117826 278622
rect 117860 278588 117898 278622
rect 117932 278588 117970 278622
rect 118004 278588 118042 278622
rect 118076 278588 118114 278622
rect 118148 278588 118186 278622
rect 118220 278588 118258 278622
rect 118292 278588 118330 278622
rect 118364 278588 118402 278622
rect 118436 278588 118474 278622
rect 118508 278588 118546 278622
rect 118580 278588 118618 278622
rect 118652 278588 118681 278622
rect 117581 278582 118681 278588
rect 117581 278480 118681 278486
rect 117581 278446 117610 278480
rect 117644 278446 117682 278480
rect 117716 278446 117754 278480
rect 117788 278446 117826 278480
rect 117860 278446 117898 278480
rect 117932 278446 117970 278480
rect 118004 278446 118042 278480
rect 118076 278446 118114 278480
rect 118148 278446 118186 278480
rect 118220 278446 118258 278480
rect 118292 278446 118330 278480
rect 118364 278446 118402 278480
rect 118436 278446 118474 278480
rect 118508 278446 118546 278480
rect 118580 278446 118618 278480
rect 118652 278446 118681 278480
rect 117581 278440 118681 278446
rect 118759 278430 118801 278638
rect 119257 278720 119363 281140
rect 119735 278720 119845 281140
rect 124495 280818 124958 280846
rect 123506 280816 124958 280818
rect 123444 280811 124958 280816
rect 121846 280767 124958 280811
rect 120433 280718 120825 280724
rect 120433 280684 120468 280718
rect 120502 280684 120540 280718
rect 120574 280684 120612 280718
rect 120646 280684 120684 280718
rect 120718 280684 120756 280718
rect 120790 280684 120825 280718
rect 120433 280678 120825 280684
rect 121133 280718 121525 280724
rect 121133 280684 121168 280718
rect 121202 280684 121240 280718
rect 121274 280684 121312 280718
rect 121346 280684 121384 280718
rect 121418 280684 121456 280718
rect 121490 280684 121525 280718
rect 121133 280678 121525 280684
rect 121846 280696 124573 280767
rect 120377 280604 120423 280637
rect 120377 280570 120383 280604
rect 120417 280570 120423 280604
rect 120377 280537 120423 280570
rect 120835 280604 120881 280637
rect 120835 280570 120841 280604
rect 120875 280570 120881 280604
rect 120835 280537 120881 280570
rect 121077 280604 121123 280637
rect 121077 280570 121083 280604
rect 121117 280570 121123 280604
rect 121077 280537 121123 280570
rect 121535 280604 121581 280637
rect 121535 280570 121541 280604
rect 121575 280570 121581 280604
rect 121535 280537 121581 280570
rect 120433 280490 120825 280496
rect 120433 280456 120468 280490
rect 120502 280456 120540 280490
rect 120574 280456 120612 280490
rect 120646 280456 120684 280490
rect 120718 280456 120756 280490
rect 120790 280456 120825 280490
rect 120433 280450 120825 280456
rect 121133 280490 121525 280496
rect 121133 280456 121168 280490
rect 121202 280456 121240 280490
rect 121274 280456 121312 280490
rect 121346 280456 121384 280490
rect 121418 280456 121456 280490
rect 121490 280456 121525 280490
rect 121133 280450 121525 280456
rect 121846 280383 121915 280696
rect 123444 280632 124573 280696
rect 123444 280510 123545 280632
rect 124495 280587 124573 280632
rect 124881 280587 124958 280767
rect 122360 280504 122752 280510
rect 122360 280470 122395 280504
rect 122429 280470 122467 280504
rect 122501 280470 122539 280504
rect 122573 280470 122611 280504
rect 122645 280470 122683 280504
rect 122717 280470 122752 280504
rect 122360 280464 122752 280470
rect 123060 280504 123551 280510
rect 123060 280470 123095 280504
rect 123129 280470 123167 280504
rect 123201 280470 123239 280504
rect 123273 280470 123311 280504
rect 123345 280470 123383 280504
rect 123417 280470 123551 280504
rect 124495 280498 124958 280587
rect 123060 280464 123551 280470
rect 123452 280423 123551 280464
rect 121134 280340 121915 280383
rect 120433 280334 120825 280340
rect 120433 280300 120468 280334
rect 120502 280300 120540 280334
rect 120574 280300 120612 280334
rect 120646 280300 120684 280334
rect 120718 280300 120756 280334
rect 120790 280300 120825 280334
rect 120433 280294 120825 280300
rect 121133 280339 121915 280340
rect 122304 280406 122350 280423
rect 122304 280372 122310 280406
rect 122344 280372 122350 280406
rect 121133 280334 121525 280339
rect 121133 280300 121168 280334
rect 121202 280300 121240 280334
rect 121274 280300 121312 280334
rect 121346 280300 121384 280334
rect 121418 280300 121456 280334
rect 121490 280300 121525 280334
rect 121133 280294 121525 280300
rect 122304 280334 122350 280372
rect 122304 280300 122310 280334
rect 122344 280300 122350 280334
rect 122304 280262 122350 280300
rect 120377 280236 120423 280253
rect 120377 280202 120383 280236
rect 120417 280202 120423 280236
rect 120377 280164 120423 280202
rect 120377 280130 120383 280164
rect 120417 280130 120423 280164
rect 120377 280092 120423 280130
rect 120377 280058 120383 280092
rect 120417 280058 120423 280092
rect 120377 280020 120423 280058
rect 120377 279986 120383 280020
rect 120417 279986 120423 280020
rect 120377 279948 120423 279986
rect 120377 279914 120383 279948
rect 120417 279914 120423 279948
rect 120377 279876 120423 279914
rect 120377 279842 120383 279876
rect 120417 279842 120423 279876
rect 120377 279804 120423 279842
rect 120377 279770 120383 279804
rect 120417 279770 120423 279804
rect 120377 279753 120423 279770
rect 120835 280236 120881 280253
rect 120835 280202 120841 280236
rect 120875 280202 120881 280236
rect 120835 280164 120881 280202
rect 120835 280130 120841 280164
rect 120875 280130 120881 280164
rect 120835 280092 120881 280130
rect 120835 280058 120841 280092
rect 120875 280064 120881 280092
rect 121077 280236 121123 280253
rect 121077 280202 121083 280236
rect 121117 280202 121123 280236
rect 121077 280164 121123 280202
rect 121077 280130 121083 280164
rect 121117 280130 121123 280164
rect 121077 280092 121123 280130
rect 121077 280064 121083 280092
rect 120875 280058 121083 280064
rect 121117 280058 121123 280092
rect 120835 280020 121123 280058
rect 120835 279986 120841 280020
rect 120875 279986 121083 280020
rect 121117 279986 121123 280020
rect 120835 279948 121123 279986
rect 120835 279914 120841 279948
rect 120875 279937 121083 279948
rect 120875 279914 120881 279937
rect 120835 279876 120881 279914
rect 120835 279842 120841 279876
rect 120875 279842 120881 279876
rect 120835 279804 120881 279842
rect 120835 279770 120841 279804
rect 120875 279770 120881 279804
rect 120835 279753 120881 279770
rect 120433 279706 120825 279712
rect 120433 279672 120468 279706
rect 120502 279672 120540 279706
rect 120574 279672 120612 279706
rect 120646 279672 120684 279706
rect 120718 279672 120756 279706
rect 120790 279672 120825 279706
rect 120433 279636 120825 279672
rect 120433 279584 120529 279636
rect 120581 279584 120593 279636
rect 120645 279584 120657 279636
rect 120709 279584 120825 279636
rect 120433 279550 120825 279584
rect 120433 279516 120468 279550
rect 120502 279516 120540 279550
rect 120574 279516 120612 279550
rect 120646 279516 120684 279550
rect 120718 279516 120756 279550
rect 120790 279516 120825 279550
rect 120433 279510 120825 279516
rect 120377 279452 120423 279469
rect 120377 279418 120383 279452
rect 120417 279418 120423 279452
rect 120377 279380 120423 279418
rect 120377 279346 120383 279380
rect 120417 279346 120423 279380
rect 120377 279308 120423 279346
rect 120377 279274 120383 279308
rect 120417 279274 120423 279308
rect 120377 279236 120423 279274
rect 120377 279202 120383 279236
rect 120417 279202 120423 279236
rect 120377 279164 120423 279202
rect 120377 279130 120383 279164
rect 120417 279130 120423 279164
rect 120377 279092 120423 279130
rect 120377 279058 120383 279092
rect 120417 279058 120423 279092
rect 120377 279020 120423 279058
rect 120377 278986 120383 279020
rect 120417 278986 120423 279020
rect 120377 278969 120423 278986
rect 120835 279452 120881 279469
rect 120835 279418 120841 279452
rect 120875 279418 120881 279452
rect 120835 279380 120881 279418
rect 120835 279346 120841 279380
rect 120875 279346 120881 279380
rect 120835 279308 120881 279346
rect 120835 279274 120841 279308
rect 120875 279280 120881 279308
rect 120953 279280 121018 279937
rect 121077 279914 121083 279937
rect 121117 279914 121123 279948
rect 121077 279876 121123 279914
rect 121077 279842 121083 279876
rect 121117 279842 121123 279876
rect 121077 279804 121123 279842
rect 121077 279770 121083 279804
rect 121117 279770 121123 279804
rect 121077 279753 121123 279770
rect 121535 280236 121624 280253
rect 121535 280202 121541 280236
rect 121575 280202 121624 280236
rect 121535 280164 121624 280202
rect 121535 280130 121541 280164
rect 121575 280130 121624 280164
rect 121535 280092 121624 280130
rect 121535 280058 121541 280092
rect 121575 280058 121624 280092
rect 121535 280020 121624 280058
rect 121535 279986 121541 280020
rect 121575 279986 121624 280020
rect 121535 279948 121624 279986
rect 121535 279914 121541 279948
rect 121575 279914 121624 279948
rect 122304 280228 122310 280262
rect 122344 280228 122350 280262
rect 122304 280190 122350 280228
rect 122304 280156 122310 280190
rect 122344 280156 122350 280190
rect 122304 280118 122350 280156
rect 122304 280084 122310 280118
rect 122344 280084 122350 280118
rect 122304 280046 122350 280084
rect 122304 280012 122310 280046
rect 122344 280012 122350 280046
rect 122304 279974 122350 280012
rect 122304 279940 122310 279974
rect 122344 279940 122350 279974
rect 121535 279876 121624 279914
rect 121535 279842 121541 279876
rect 121575 279842 121624 279876
rect 121535 279804 121624 279842
rect 121535 279770 121541 279804
rect 121575 279770 121624 279804
rect 121535 279753 121624 279770
rect 121133 279706 121525 279712
rect 121133 279672 121168 279706
rect 121202 279672 121240 279706
rect 121274 279672 121312 279706
rect 121346 279672 121384 279706
rect 121418 279672 121456 279706
rect 121490 279672 121525 279706
rect 121133 279550 121525 279672
rect 121133 279516 121168 279550
rect 121202 279516 121240 279550
rect 121274 279516 121312 279550
rect 121346 279516 121384 279550
rect 121418 279516 121456 279550
rect 121490 279516 121525 279550
rect 121133 279510 121525 279516
rect 121581 279469 121624 279753
rect 121797 279886 122235 279937
rect 122304 279923 122350 279940
rect 122762 280406 123050 280423
rect 122762 280372 122768 280406
rect 122802 280372 123010 280406
rect 123044 280372 123050 280406
rect 122762 280334 123050 280372
rect 122762 280300 122768 280334
rect 122802 280300 123010 280334
rect 123044 280300 123050 280334
rect 122762 280262 123050 280300
rect 122762 280228 122768 280262
rect 122802 280228 123010 280262
rect 123044 280228 123050 280262
rect 122762 280190 123050 280228
rect 122762 280156 122768 280190
rect 122802 280156 123010 280190
rect 123044 280156 123050 280190
rect 122762 280118 123050 280156
rect 122762 280084 122768 280118
rect 122802 280084 123010 280118
rect 123044 280084 123050 280118
rect 122762 280046 123050 280084
rect 122762 280012 122768 280046
rect 122802 280012 123010 280046
rect 123044 280012 123050 280046
rect 122762 279974 123050 280012
rect 122762 279940 122768 279974
rect 122802 279940 123010 279974
rect 123044 279940 123050 279974
rect 122762 279923 123050 279940
rect 123462 280406 123551 280423
rect 123462 280372 123468 280406
rect 123502 280372 123551 280406
rect 123462 280334 123551 280372
rect 123462 280300 123468 280334
rect 123502 280300 123551 280334
rect 123462 280262 123551 280300
rect 123462 280228 123468 280262
rect 123502 280228 123551 280262
rect 123462 280190 123551 280228
rect 123462 280156 123468 280190
rect 123502 280156 123551 280190
rect 123462 280118 123551 280156
rect 123462 280084 123468 280118
rect 123502 280084 123551 280118
rect 123462 280046 123551 280084
rect 123462 280012 123468 280046
rect 123502 280012 123551 280046
rect 123462 279974 123551 280012
rect 123462 279940 123468 279974
rect 123502 279940 123551 279974
rect 123462 279923 123551 279940
rect 121077 279452 121123 279469
rect 121077 279418 121083 279452
rect 121117 279418 121123 279452
rect 121077 279380 121123 279418
rect 121077 279346 121083 279380
rect 121117 279346 121123 279380
rect 121077 279308 121123 279346
rect 121077 279280 121083 279308
rect 120875 279274 121083 279280
rect 121117 279274 121123 279308
rect 120835 279236 121123 279274
rect 120835 279202 120841 279236
rect 120875 279202 121083 279236
rect 121117 279202 121123 279236
rect 120835 279164 121123 279202
rect 120835 279130 120841 279164
rect 120875 279153 121083 279164
rect 120875 279130 120881 279153
rect 120835 279092 120881 279130
rect 120835 279058 120841 279092
rect 120875 279058 120881 279092
rect 120835 279020 120881 279058
rect 120835 278986 120841 279020
rect 120875 278986 120881 279020
rect 120835 278969 120881 278986
rect 120433 278922 120825 278928
rect 120433 278888 120468 278922
rect 120502 278888 120540 278922
rect 120574 278888 120612 278922
rect 120646 278888 120684 278922
rect 120718 278888 120756 278922
rect 120790 278888 120825 278922
rect 120433 278766 120825 278888
rect 120433 278732 120468 278766
rect 120502 278732 120540 278766
rect 120574 278732 120612 278766
rect 120646 278732 120684 278766
rect 120718 278732 120756 278766
rect 120790 278732 120825 278766
rect 120433 278726 120825 278732
rect 119257 278619 119845 278720
rect 120377 278668 120423 278685
rect 120377 278634 120383 278668
rect 120417 278634 120423 278668
rect 115862 278388 116362 278418
rect 117461 278407 117549 278430
rect 115862 278382 117205 278388
rect 115862 278377 116134 278382
rect 115589 278318 115595 278352
rect 115629 278318 115635 278352
rect 116105 278348 116134 278377
rect 116168 278348 116206 278382
rect 116240 278348 116278 278382
rect 116312 278348 116350 278382
rect 116384 278348 116422 278382
rect 116456 278348 116494 278382
rect 116528 278348 116566 278382
rect 116600 278348 116638 278382
rect 116672 278348 116710 278382
rect 116744 278348 116782 278382
rect 116816 278348 116854 278382
rect 116888 278348 116926 278382
rect 116960 278348 116998 278382
rect 117032 278348 117070 278382
rect 117104 278348 117142 278382
rect 117176 278348 117205 278382
rect 116105 278342 117205 278348
rect 117461 278373 117509 278407
rect 117543 278373 117549 278407
rect 117461 278335 117549 278373
rect 115589 278295 115635 278318
rect 115809 278285 115881 278326
rect 114324 278251 114342 278285
rect 114376 278251 114396 278285
rect 114324 278195 114396 278251
rect 114657 278279 114857 278285
rect 114657 278245 114704 278279
rect 114738 278245 114776 278279
rect 114810 278245 114857 278279
rect 114657 278239 114857 278245
rect 115348 278279 115548 278285
rect 115348 278245 115395 278279
rect 115429 278245 115467 278279
rect 115501 278245 115548 278279
rect 115348 278239 115548 278245
rect 115809 278251 115828 278285
rect 115862 278251 115881 278285
rect 114843 278195 115030 278210
rect 114324 278150 114781 278195
rect 112874 278034 112922 278124
rect 113000 278084 114100 278090
rect 113000 278050 113029 278084
rect 113063 278050 113101 278084
rect 113135 278050 113173 278084
rect 113207 278050 113245 278084
rect 113279 278050 113317 278084
rect 113351 278050 113389 278084
rect 113423 278050 113461 278084
rect 113495 278050 113533 278084
rect 113567 278050 113605 278084
rect 113639 278050 113677 278084
rect 113711 278050 113749 278084
rect 113783 278050 113821 278084
rect 113855 278050 113893 278084
rect 113927 278050 113965 278084
rect 113999 278050 114037 278084
rect 114071 278050 114100 278084
rect 113000 278044 114100 278050
rect 114178 278034 114226 278124
rect 114737 278095 114781 278150
rect 114843 278143 114891 278195
rect 114943 278143 115030 278195
rect 114843 278125 115030 278143
rect 115175 278195 115362 278210
rect 115809 278195 115881 278251
rect 115175 278143 115262 278195
rect 115314 278143 115362 278195
rect 115175 278125 115362 278143
rect 115424 278150 115881 278195
rect 115979 278313 116073 278332
rect 115979 278279 116033 278313
rect 116067 278279 116073 278313
rect 115979 278260 116073 278279
rect 117237 278313 117331 278332
rect 117237 278279 117243 278313
rect 117277 278279 117331 278313
rect 117237 278260 117331 278279
rect 115979 278168 116027 278260
rect 116105 278244 117205 278250
rect 116105 278210 116134 278244
rect 116168 278210 116206 278244
rect 116240 278210 116278 278244
rect 116312 278210 116350 278244
rect 116384 278210 116422 278244
rect 116456 278210 116494 278244
rect 116528 278210 116566 278244
rect 116600 278210 116638 278244
rect 116672 278210 116710 278244
rect 116744 278210 116782 278244
rect 116816 278210 116854 278244
rect 116888 278210 116926 278244
rect 116960 278210 116998 278244
rect 117032 278210 117070 278244
rect 117104 278210 117142 278244
rect 117176 278210 117205 278244
rect 116105 278204 117205 278210
rect 117283 278168 117331 278260
rect 115424 278095 115468 278150
rect 115979 278124 117331 278168
rect 114657 278089 114857 278095
rect 114657 278055 114704 278089
rect 114738 278055 114776 278089
rect 114810 278055 114857 278089
rect 114657 278049 114857 278055
rect 115348 278089 115548 278095
rect 115348 278055 115395 278089
rect 115429 278055 115467 278089
rect 115501 278055 115548 278089
rect 115348 278049 115548 278055
rect 112874 278015 112968 278034
rect 112874 277981 112928 278015
rect 112962 277981 112968 278015
rect 112874 277962 112968 277981
rect 114132 278015 114226 278034
rect 114132 277981 114138 278015
rect 114172 277981 114226 278015
rect 114132 277962 114226 277981
rect 114570 278016 114616 278039
rect 114570 277982 114576 278016
rect 114610 277982 114616 278016
rect 111524 277902 112624 277908
rect 111524 277868 111553 277902
rect 111587 277868 111625 277902
rect 111659 277868 111697 277902
rect 111731 277868 111769 277902
rect 111803 277868 111841 277902
rect 111875 277868 111913 277902
rect 111947 277868 111985 277902
rect 112019 277868 112057 277902
rect 112091 277868 112129 277902
rect 112163 277868 112201 277902
rect 112235 277868 112273 277902
rect 112307 277868 112345 277902
rect 112379 277868 112417 277902
rect 112451 277868 112489 277902
rect 112523 277868 112561 277902
rect 112595 277868 112624 277902
rect 111524 277864 112624 277868
rect 112874 277868 112922 277962
rect 114327 277957 114395 277958
rect 114570 277957 114616 277982
rect 113000 277946 114100 277952
rect 113000 277912 113029 277946
rect 113063 277912 113101 277946
rect 113135 277912 113173 277946
rect 113207 277912 113245 277946
rect 113279 277912 113317 277946
rect 113351 277912 113389 277946
rect 113423 277912 113461 277946
rect 113495 277912 113533 277946
rect 113567 277912 113605 277946
rect 113639 277912 113677 277946
rect 113711 277912 113749 277946
rect 113783 277912 113821 277946
rect 113855 277912 113893 277946
rect 113927 277912 113965 277946
rect 113999 277912 114037 277946
rect 114071 277912 114100 277946
rect 113000 277906 114100 277912
rect 114327 277944 114616 277957
rect 114327 277910 114576 277944
rect 114610 277910 114616 277944
rect 114327 277897 114616 277910
rect 114327 277868 114395 277897
rect 114570 277887 114616 277897
rect 114898 278016 114944 278039
rect 114898 277982 114904 278016
rect 114938 277982 114944 278016
rect 114898 277944 114944 277982
rect 114898 277910 114904 277944
rect 114938 277910 114944 277944
rect 114898 277887 114944 277910
rect 115261 278016 115307 278039
rect 115261 277982 115267 278016
rect 115301 277982 115307 278016
rect 115261 277944 115307 277982
rect 115261 277910 115267 277944
rect 115301 277910 115307 277944
rect 115261 277887 115307 277910
rect 115589 278016 115635 278039
rect 115589 277982 115595 278016
rect 115629 277982 115635 278016
rect 115589 277957 115635 277982
rect 115979 278034 116027 278124
rect 116105 278084 117205 278090
rect 116105 278050 116134 278084
rect 116168 278050 116206 278084
rect 116240 278050 116278 278084
rect 116312 278050 116350 278084
rect 116384 278050 116422 278084
rect 116456 278050 116494 278084
rect 116528 278050 116566 278084
rect 116600 278050 116638 278084
rect 116672 278050 116710 278084
rect 116744 278050 116782 278084
rect 116816 278050 116854 278084
rect 116888 278050 116926 278084
rect 116960 278050 116998 278084
rect 117032 278050 117070 278084
rect 117104 278050 117142 278084
rect 117176 278050 117205 278084
rect 116105 278044 117205 278050
rect 117283 278034 117331 278124
rect 115979 278015 116073 278034
rect 115979 277981 116033 278015
rect 116067 277981 116073 278015
rect 115979 277962 116073 277981
rect 117237 278015 117331 278034
rect 117237 277981 117243 278015
rect 117277 277981 117331 278015
rect 117237 277962 117331 277981
rect 115810 277957 115878 277958
rect 115589 277944 115878 277957
rect 115589 277910 115595 277944
rect 115629 277910 115878 277944
rect 115589 277897 115878 277910
rect 116105 277946 117205 277952
rect 116105 277912 116134 277946
rect 116168 277912 116206 277946
rect 116240 277912 116278 277946
rect 116312 277912 116350 277946
rect 116384 277912 116422 277946
rect 116456 277912 116494 277946
rect 116528 277912 116566 277946
rect 116600 277912 116638 277946
rect 116672 277912 116710 277946
rect 116744 277912 116782 277946
rect 116816 277912 116854 277946
rect 116888 277912 116926 277946
rect 116960 277912 116998 277946
rect 117032 277912 117070 277946
rect 117104 277912 117142 277946
rect 117176 277912 117205 277946
rect 116105 277906 117205 277912
rect 115589 277887 115635 277897
rect 112874 277864 114395 277868
rect 111524 277862 114395 277864
rect 112044 277828 114395 277862
rect 114657 277871 114857 277877
rect 114657 277837 114704 277871
rect 114738 277837 114776 277871
rect 114810 277837 114857 277871
rect 114657 277831 114857 277837
rect 115348 277871 115548 277877
rect 115348 277837 115395 277871
rect 115429 277837 115467 277871
rect 115501 277837 115548 277871
rect 115348 277831 115548 277837
rect 115810 277868 115878 277897
rect 117283 277868 117331 277962
rect 117461 278301 117509 278335
rect 117543 278301 117549 278335
rect 117461 278278 117549 278301
rect 118713 278407 118801 278430
rect 118713 278373 118719 278407
rect 118753 278373 118801 278407
rect 118713 278335 118801 278373
rect 118713 278301 118719 278335
rect 118753 278301 118801 278335
rect 118713 278278 118801 278301
rect 117461 278070 117503 278278
rect 117581 278262 118681 278268
rect 117581 278228 117610 278262
rect 117644 278228 117682 278262
rect 117716 278228 117754 278262
rect 117788 278228 117826 278262
rect 117860 278228 117898 278262
rect 117932 278228 117970 278262
rect 118004 278228 118042 278262
rect 118076 278228 118114 278262
rect 118148 278228 118186 278262
rect 118220 278228 118258 278262
rect 118292 278228 118330 278262
rect 118364 278228 118402 278262
rect 118436 278228 118474 278262
rect 118508 278228 118546 278262
rect 118580 278228 118618 278262
rect 118652 278228 118681 278262
rect 117581 278222 118681 278228
rect 117581 278120 118681 278126
rect 117581 278086 117610 278120
rect 117644 278086 117682 278120
rect 117716 278086 117754 278120
rect 117788 278086 117826 278120
rect 117860 278086 117898 278120
rect 117932 278086 117970 278120
rect 118004 278086 118042 278120
rect 118076 278086 118114 278120
rect 118148 278086 118186 278120
rect 118220 278086 118258 278120
rect 118292 278086 118330 278120
rect 118364 278086 118402 278120
rect 118436 278086 118474 278120
rect 118508 278086 118546 278120
rect 118580 278086 118618 278120
rect 118652 278086 118681 278120
rect 117581 278080 118681 278086
rect 118759 278070 118801 278278
rect 120377 278596 120423 278634
rect 120377 278562 120383 278596
rect 120417 278562 120423 278596
rect 120377 278524 120423 278562
rect 120377 278490 120383 278524
rect 120417 278490 120423 278524
rect 120377 278452 120423 278490
rect 120377 278418 120383 278452
rect 120417 278418 120423 278452
rect 120377 278380 120423 278418
rect 120377 278346 120383 278380
rect 120417 278346 120423 278380
rect 120377 278308 120423 278346
rect 120377 278274 120383 278308
rect 120417 278274 120423 278308
rect 120377 278236 120423 278274
rect 120377 278202 120383 278236
rect 120417 278202 120423 278236
rect 120377 278185 120423 278202
rect 120835 278668 120881 278685
rect 120835 278634 120841 278668
rect 120875 278634 120881 278668
rect 120835 278596 120881 278634
rect 120835 278562 120841 278596
rect 120875 278562 120881 278596
rect 120835 278524 120881 278562
rect 120835 278490 120841 278524
rect 120875 278496 120881 278524
rect 120953 278496 121018 279153
rect 121077 279130 121083 279153
rect 121117 279130 121123 279164
rect 121077 279092 121123 279130
rect 121077 279058 121083 279092
rect 121117 279058 121123 279092
rect 121077 279020 121123 279058
rect 121077 278986 121083 279020
rect 121117 278986 121123 279020
rect 121077 278969 121123 278986
rect 121535 279452 121677 279469
rect 121535 279418 121541 279452
rect 121575 279418 121677 279452
rect 121535 279394 121677 279418
rect 121535 279380 121605 279394
rect 121535 279346 121541 279380
rect 121575 279346 121605 279380
rect 121535 279342 121605 279346
rect 121657 279342 121677 279394
rect 121535 279330 121677 279342
rect 121535 279308 121605 279330
rect 121535 279274 121541 279308
rect 121575 279278 121605 279308
rect 121657 279278 121677 279330
rect 121575 279274 121677 279278
rect 121535 279266 121677 279274
rect 121535 279236 121605 279266
rect 121535 279202 121541 279236
rect 121575 279214 121605 279236
rect 121657 279214 121677 279266
rect 121797 279276 121859 279886
rect 122181 279276 122235 279886
rect 122360 279876 122752 279882
rect 122360 279842 122395 279876
rect 122429 279842 122467 279876
rect 122501 279842 122539 279876
rect 122573 279842 122611 279876
rect 122645 279842 122683 279876
rect 122717 279842 122752 279876
rect 122360 279836 122752 279842
rect 122808 279836 122951 279923
rect 123452 279882 123551 279923
rect 122360 279726 122951 279836
rect 122360 279720 122752 279726
rect 122360 279686 122395 279720
rect 122429 279686 122467 279720
rect 122501 279686 122539 279720
rect 122573 279686 122611 279720
rect 122645 279686 122683 279720
rect 122717 279686 122752 279720
rect 122360 279680 122752 279686
rect 122808 279639 122951 279726
rect 123060 279876 123551 279882
rect 123060 279842 123095 279876
rect 123129 279842 123167 279876
rect 123201 279842 123239 279876
rect 123273 279842 123311 279876
rect 123345 279842 123383 279876
rect 123417 279842 123551 279876
rect 123060 279720 123551 279842
rect 123060 279686 123095 279720
rect 123129 279686 123167 279720
rect 123201 279686 123239 279720
rect 123273 279686 123311 279720
rect 123345 279686 123383 279720
rect 123417 279686 123551 279720
rect 123060 279680 123551 279686
rect 123452 279639 123551 279680
rect 121797 279225 122235 279276
rect 122304 279622 122350 279639
rect 122304 279588 122310 279622
rect 122344 279588 122350 279622
rect 122304 279550 122350 279588
rect 122304 279516 122310 279550
rect 122344 279516 122350 279550
rect 122304 279478 122350 279516
rect 122304 279444 122310 279478
rect 122344 279444 122350 279478
rect 122304 279406 122350 279444
rect 122304 279372 122310 279406
rect 122344 279372 122350 279406
rect 122304 279334 122350 279372
rect 122304 279300 122310 279334
rect 122344 279300 122350 279334
rect 122304 279262 122350 279300
rect 122304 279228 122310 279262
rect 122344 279228 122350 279262
rect 121575 279202 121677 279214
rect 121535 279164 121605 279202
rect 121535 279130 121541 279164
rect 121575 279150 121605 279164
rect 121657 279150 121677 279202
rect 121575 279138 121677 279150
rect 122304 279190 122350 279228
rect 122304 279156 122310 279190
rect 122344 279156 122350 279190
rect 122304 279139 122350 279156
rect 122762 279622 123050 279639
rect 122762 279588 122768 279622
rect 122802 279588 123010 279622
rect 123044 279588 123050 279622
rect 122762 279550 123050 279588
rect 122762 279516 122768 279550
rect 122802 279516 123010 279550
rect 123044 279516 123050 279550
rect 122762 279478 123050 279516
rect 122762 279444 122768 279478
rect 122802 279444 123010 279478
rect 123044 279444 123050 279478
rect 122762 279406 123050 279444
rect 122762 279372 122768 279406
rect 122802 279372 123010 279406
rect 123044 279372 123050 279406
rect 122762 279334 123050 279372
rect 122762 279300 122768 279334
rect 122802 279300 123010 279334
rect 123044 279300 123050 279334
rect 122762 279262 123050 279300
rect 122762 279228 122768 279262
rect 122802 279228 123010 279262
rect 123044 279228 123050 279262
rect 122762 279190 123050 279228
rect 122762 279156 122768 279190
rect 122802 279156 123010 279190
rect 123044 279156 123050 279190
rect 122762 279139 123050 279156
rect 123462 279622 123551 279639
rect 123462 279588 123468 279622
rect 123502 279588 123551 279622
rect 123462 279550 123551 279588
rect 123462 279516 123468 279550
rect 123502 279516 123551 279550
rect 123462 279478 123551 279516
rect 123462 279444 123468 279478
rect 123502 279444 123551 279478
rect 123462 279406 123551 279444
rect 123462 279372 123468 279406
rect 123502 279372 123551 279406
rect 123462 279334 123551 279372
rect 123462 279300 123468 279334
rect 123502 279300 123551 279334
rect 123462 279262 123551 279300
rect 123462 279228 123468 279262
rect 123502 279228 123551 279262
rect 123462 279190 123551 279228
rect 123462 279156 123468 279190
rect 123502 279156 123551 279190
rect 123462 279139 123551 279156
rect 121575 279130 121605 279138
rect 121535 279092 121605 279130
rect 121535 279058 121541 279092
rect 121575 279086 121605 279092
rect 121657 279086 121677 279138
rect 123452 279098 123551 279139
rect 121575 279074 121677 279086
rect 121575 279058 121605 279074
rect 121535 279022 121605 279058
rect 121657 279022 121677 279074
rect 122360 279092 122752 279098
rect 122360 279058 122395 279092
rect 122429 279058 122467 279092
rect 122501 279058 122539 279092
rect 122573 279058 122611 279092
rect 122645 279058 122683 279092
rect 122717 279058 122752 279092
rect 122360 279052 122752 279058
rect 123060 279092 123551 279098
rect 123060 279058 123095 279092
rect 123129 279058 123167 279092
rect 123201 279058 123239 279092
rect 123273 279058 123311 279092
rect 123345 279058 123383 279092
rect 123417 279058 123551 279092
rect 123060 279052 123551 279058
rect 121535 279020 121677 279022
rect 121535 278986 121541 279020
rect 121575 279010 121677 279020
rect 121575 278986 121605 279010
rect 121535 278969 121605 278986
rect 121581 278958 121605 278969
rect 121657 278958 121677 279010
rect 121581 278946 121677 278958
rect 121133 278922 121525 278928
rect 121133 278888 121168 278922
rect 121202 278888 121240 278922
rect 121274 278888 121312 278922
rect 121346 278888 121384 278922
rect 121418 278888 121456 278922
rect 121490 278888 121525 278922
rect 121133 278766 121525 278888
rect 121133 278732 121168 278766
rect 121202 278732 121240 278766
rect 121274 278732 121312 278766
rect 121346 278732 121384 278766
rect 121418 278732 121456 278766
rect 121490 278732 121525 278766
rect 121133 278726 121525 278732
rect 121581 278894 121605 278946
rect 121657 278894 121677 278946
rect 121581 278882 121677 278894
rect 121581 278830 121605 278882
rect 121657 278830 121677 278882
rect 121581 278818 121677 278830
rect 121581 278766 121605 278818
rect 121657 278766 121677 278818
rect 121581 278754 121677 278766
rect 121581 278702 121605 278754
rect 121657 278702 121677 278754
rect 121581 278690 121677 278702
rect 121581 278685 121605 278690
rect 121077 278668 121123 278685
rect 121077 278634 121083 278668
rect 121117 278634 121123 278668
rect 121077 278596 121123 278634
rect 121077 278562 121083 278596
rect 121117 278562 121123 278596
rect 121077 278524 121123 278562
rect 121077 278496 121083 278524
rect 120875 278490 121083 278496
rect 121117 278490 121123 278524
rect 120835 278452 121123 278490
rect 120835 278418 120841 278452
rect 120875 278418 121083 278452
rect 121117 278418 121123 278452
rect 120835 278380 121123 278418
rect 120835 278346 120841 278380
rect 120875 278369 121083 278380
rect 120875 278346 120881 278369
rect 120835 278308 120881 278346
rect 120835 278274 120841 278308
rect 120875 278274 120881 278308
rect 120835 278236 120881 278274
rect 120835 278202 120841 278236
rect 120875 278202 120881 278236
rect 120835 278185 120881 278202
rect 117461 278047 117549 278070
rect 117461 278013 117509 278047
rect 117543 278013 117549 278047
rect 117461 277975 117549 278013
rect 117461 277941 117509 277975
rect 117543 277941 117549 277975
rect 117461 277918 117549 277941
rect 118713 278047 118801 278070
rect 118713 278013 118719 278047
rect 118753 278013 118801 278047
rect 118713 277975 118801 278013
rect 118713 277941 118719 277975
rect 118753 277941 118801 277975
rect 120433 278138 120825 278144
rect 120433 278104 120468 278138
rect 120502 278104 120540 278138
rect 120574 278104 120612 278138
rect 120646 278104 120684 278138
rect 120718 278104 120756 278138
rect 120790 278104 120825 278138
rect 120433 277982 120825 278104
rect 120433 277948 120468 277982
rect 120502 277948 120540 277982
rect 120574 277948 120612 277982
rect 120646 277948 120684 277982
rect 120718 277948 120756 277982
rect 120790 277948 120825 277982
rect 120433 277942 120825 277948
rect 118713 277918 118801 277941
rect 115810 277864 117331 277868
rect 117581 277902 118681 277908
rect 117581 277868 117610 277902
rect 117644 277868 117682 277902
rect 117716 277868 117754 277902
rect 117788 277868 117826 277902
rect 117860 277868 117898 277902
rect 117932 277868 117970 277902
rect 118004 277868 118042 277902
rect 118076 277868 118114 277902
rect 118148 277868 118186 277902
rect 118220 277868 118258 277902
rect 118292 277868 118330 277902
rect 118364 277868 118402 277902
rect 118436 277868 118474 277902
rect 118508 277868 118546 277902
rect 118580 277868 118618 277902
rect 118652 277868 118681 277902
rect 117581 277864 118681 277868
rect 115810 277862 118681 277864
rect 120377 277884 120423 277901
rect 112719 277786 112924 277828
rect 113982 277754 114266 277764
rect 114724 277754 114783 277831
rect 113982 277733 114783 277754
rect 113982 277699 114034 277733
rect 114068 277699 114106 277733
rect 114140 277699 114178 277733
rect 114212 277699 114783 277733
rect 113982 277665 114783 277699
rect 115422 277754 115481 277831
rect 115810 277828 118161 277862
rect 120377 277850 120383 277884
rect 120417 277850 120423 277884
rect 117281 277786 117486 277828
rect 120377 277812 120423 277850
rect 120377 277778 120383 277812
rect 120417 277778 120423 277812
rect 115939 277754 116223 277764
rect 115422 277733 116223 277754
rect 115422 277699 115992 277733
rect 116026 277699 116064 277733
rect 116098 277699 116136 277733
rect 116170 277699 116223 277733
rect 115422 277665 116223 277699
rect 113982 277664 114266 277665
rect 115939 277664 116223 277665
rect 120377 277740 120423 277778
rect 120377 277706 120383 277740
rect 120417 277706 120423 277740
rect 120377 277668 120423 277706
rect 120377 277634 120383 277668
rect 120417 277634 120423 277668
rect 120377 277596 120423 277634
rect 120377 277562 120383 277596
rect 120417 277562 120423 277596
rect 112970 277542 114070 277548
rect 111524 277534 112624 277540
rect 111524 277500 111553 277534
rect 111587 277500 111625 277534
rect 111659 277500 111697 277534
rect 111731 277500 111769 277534
rect 111803 277500 111841 277534
rect 111875 277500 111913 277534
rect 111947 277500 111985 277534
rect 112019 277500 112057 277534
rect 112091 277500 112129 277534
rect 112163 277500 112201 277534
rect 112235 277500 112273 277534
rect 112307 277500 112345 277534
rect 112379 277500 112417 277534
rect 112451 277500 112489 277534
rect 112523 277500 112561 277534
rect 112595 277500 112624 277534
rect 112970 277508 112999 277542
rect 113033 277508 113071 277542
rect 113105 277508 113143 277542
rect 113177 277508 113215 277542
rect 113249 277508 113287 277542
rect 113321 277508 113359 277542
rect 113393 277508 113431 277542
rect 113465 277508 113503 277542
rect 113537 277508 113575 277542
rect 113609 277508 113647 277542
rect 113681 277508 113719 277542
rect 113753 277508 113791 277542
rect 113825 277508 113863 277542
rect 113897 277508 113935 277542
rect 113969 277508 114007 277542
rect 114041 277508 114070 277542
rect 116135 277542 117235 277548
rect 112970 277502 114070 277508
rect 114657 277517 114857 277523
rect 111524 277494 112624 277500
rect 111404 277461 111492 277484
rect 111404 277427 111452 277461
rect 111486 277427 111492 277461
rect 111404 277389 111492 277427
rect 111404 277355 111452 277389
rect 111486 277355 111492 277389
rect 111404 277332 111492 277355
rect 112656 277461 112744 277484
rect 112656 277427 112662 277461
rect 112696 277427 112744 277461
rect 112656 277416 112744 277427
rect 112850 277449 112938 277492
rect 112850 277416 112898 277449
rect 112656 277415 112898 277416
rect 112932 277415 112938 277449
rect 112656 277389 112938 277415
rect 112656 277355 112662 277389
rect 112696 277377 112938 277389
rect 112696 277355 112898 277377
rect 112656 277354 112898 277355
rect 112656 277332 112744 277354
rect 111404 277124 111446 277332
rect 111524 277316 112624 277322
rect 111524 277282 111553 277316
rect 111587 277282 111625 277316
rect 111659 277282 111697 277316
rect 111731 277282 111769 277316
rect 111803 277282 111841 277316
rect 111875 277282 111913 277316
rect 111947 277282 111985 277316
rect 112019 277282 112057 277316
rect 112091 277282 112129 277316
rect 112163 277282 112201 277316
rect 112235 277282 112273 277316
rect 112307 277282 112345 277316
rect 112379 277282 112417 277316
rect 112451 277282 112489 277316
rect 112523 277282 112561 277316
rect 112595 277282 112624 277316
rect 111524 277276 112624 277282
rect 112702 277300 112744 277332
rect 112850 277343 112898 277354
rect 112932 277343 112938 277377
rect 112850 277300 112938 277343
rect 114102 277449 114190 277492
rect 114657 277483 114704 277517
rect 114738 277483 114776 277517
rect 114810 277483 114857 277517
rect 114657 277477 114857 277483
rect 115348 277517 115548 277523
rect 115348 277483 115395 277517
rect 115429 277483 115467 277517
rect 115501 277483 115548 277517
rect 116135 277508 116164 277542
rect 116198 277508 116236 277542
rect 116270 277508 116308 277542
rect 116342 277508 116380 277542
rect 116414 277508 116452 277542
rect 116486 277508 116524 277542
rect 116558 277508 116596 277542
rect 116630 277508 116668 277542
rect 116702 277508 116740 277542
rect 116774 277508 116812 277542
rect 116846 277508 116884 277542
rect 116918 277508 116956 277542
rect 116990 277508 117028 277542
rect 117062 277508 117100 277542
rect 117134 277508 117172 277542
rect 117206 277508 117235 277542
rect 116135 277502 117235 277508
rect 117581 277534 118681 277540
rect 117581 277500 117610 277534
rect 117644 277500 117682 277534
rect 117716 277500 117754 277534
rect 117788 277500 117826 277534
rect 117860 277500 117898 277534
rect 117932 277500 117970 277534
rect 118004 277500 118042 277534
rect 118076 277500 118114 277534
rect 118148 277500 118186 277534
rect 118220 277500 118258 277534
rect 118292 277500 118330 277534
rect 118364 277500 118402 277534
rect 118436 277500 118474 277534
rect 118508 277500 118546 277534
rect 118580 277500 118618 277534
rect 118652 277500 118681 277534
rect 117581 277494 118681 277500
rect 120377 277524 120423 277562
rect 115348 277477 115548 277483
rect 114102 277415 114108 277449
rect 114142 277426 114190 277449
rect 114570 277432 114616 277467
rect 114570 277426 114576 277432
rect 114142 277415 114576 277426
rect 114102 277398 114576 277415
rect 114610 277398 114616 277432
rect 114102 277377 114616 277398
rect 114102 277343 114108 277377
rect 114142 277360 114616 277377
rect 114142 277343 114576 277360
rect 114102 277326 114576 277343
rect 114610 277326 114616 277360
rect 114102 277300 114616 277326
rect 111524 277174 112624 277180
rect 111524 277140 111553 277174
rect 111587 277140 111625 277174
rect 111659 277140 111697 277174
rect 111731 277140 111769 277174
rect 111803 277140 111841 277174
rect 111875 277140 111913 277174
rect 111947 277140 111985 277174
rect 112019 277140 112057 277174
rect 112091 277140 112129 277174
rect 112163 277140 112201 277174
rect 112235 277140 112273 277174
rect 112307 277140 112345 277174
rect 112379 277140 112417 277174
rect 112451 277140 112489 277174
rect 112523 277140 112561 277174
rect 112595 277140 112624 277174
rect 111524 277134 112624 277140
rect 112702 277124 112746 277300
rect 111404 277101 111492 277124
rect 111404 277067 111452 277101
rect 111486 277067 111492 277101
rect 111404 277029 111492 277067
rect 111404 276995 111452 277029
rect 111486 276995 111492 277029
rect 111404 276972 111492 276995
rect 112656 277101 112746 277124
rect 112656 277067 112662 277101
rect 112696 277080 112746 277101
rect 112850 277200 112892 277300
rect 114148 277293 114616 277300
rect 112970 277284 114070 277290
rect 112970 277250 112999 277284
rect 113033 277250 113071 277284
rect 113105 277250 113143 277284
rect 113177 277250 113215 277284
rect 113249 277250 113287 277284
rect 113321 277250 113359 277284
rect 113393 277250 113431 277284
rect 113465 277250 113503 277284
rect 113537 277250 113575 277284
rect 113609 277250 113647 277284
rect 113681 277250 113719 277284
rect 113753 277250 113791 277284
rect 113825 277250 113863 277284
rect 113897 277250 113935 277284
rect 113969 277250 114007 277284
rect 114041 277250 114070 277284
rect 112970 277244 114070 277250
rect 114148 277200 114190 277293
rect 112850 277162 114190 277200
rect 112696 277067 112744 277080
rect 112656 277032 112744 277067
rect 112850 277068 112892 277162
rect 112970 277118 114070 277124
rect 112970 277084 112999 277118
rect 113033 277084 113071 277118
rect 113105 277084 113143 277118
rect 113177 277084 113215 277118
rect 113249 277084 113287 277118
rect 113321 277084 113359 277118
rect 113393 277084 113431 277118
rect 113465 277084 113503 277118
rect 113537 277084 113575 277118
rect 113609 277084 113647 277118
rect 113681 277084 113719 277118
rect 113753 277084 113791 277118
rect 113825 277084 113863 277118
rect 113897 277084 113935 277118
rect 113969 277084 114007 277118
rect 114041 277084 114070 277118
rect 112970 277078 114070 277084
rect 114148 277068 114190 277162
rect 114570 277288 114616 277293
rect 114570 277254 114576 277288
rect 114610 277254 114616 277288
rect 114570 277216 114616 277254
rect 114570 277182 114576 277216
rect 114610 277182 114616 277216
rect 114570 277144 114616 277182
rect 114570 277110 114576 277144
rect 114610 277110 114616 277144
rect 114570 277075 114616 277110
rect 114898 277432 114944 277467
rect 114898 277398 114904 277432
rect 114938 277398 114944 277432
rect 114898 277360 114944 277398
rect 114898 277326 114904 277360
rect 114938 277326 114944 277360
rect 114898 277288 114944 277326
rect 114898 277254 114904 277288
rect 114938 277254 114944 277288
rect 114898 277216 114944 277254
rect 114898 277182 114904 277216
rect 114938 277182 114944 277216
rect 114898 277144 114944 277182
rect 114898 277110 114904 277144
rect 114938 277110 114944 277144
rect 114898 277075 114944 277110
rect 115261 277432 115307 277467
rect 115261 277398 115267 277432
rect 115301 277398 115307 277432
rect 115261 277360 115307 277398
rect 115261 277326 115267 277360
rect 115301 277326 115307 277360
rect 115261 277288 115307 277326
rect 115261 277254 115267 277288
rect 115301 277254 115307 277288
rect 115261 277216 115307 277254
rect 115261 277182 115267 277216
rect 115301 277182 115307 277216
rect 115261 277144 115307 277182
rect 115261 277110 115267 277144
rect 115301 277110 115307 277144
rect 115261 277075 115307 277110
rect 115589 277432 115635 277467
rect 115589 277398 115595 277432
rect 115629 277426 115635 277432
rect 116015 277449 116103 277492
rect 116015 277426 116063 277449
rect 115629 277415 116063 277426
rect 116097 277415 116103 277449
rect 115629 277398 116103 277415
rect 115589 277377 116103 277398
rect 115589 277360 116063 277377
rect 115589 277326 115595 277360
rect 115629 277343 116063 277360
rect 116097 277343 116103 277377
rect 115629 277326 116103 277343
rect 115589 277300 116103 277326
rect 117267 277449 117355 277492
rect 120377 277490 120383 277524
rect 120417 277490 120423 277524
rect 117267 277415 117273 277449
rect 117307 277416 117355 277449
rect 117461 277461 117549 277484
rect 117461 277427 117509 277461
rect 117543 277427 117549 277461
rect 117461 277416 117549 277427
rect 117307 277415 117549 277416
rect 117267 277389 117549 277415
rect 117267 277377 117509 277389
rect 117267 277343 117273 277377
rect 117307 277355 117509 277377
rect 117543 277355 117549 277389
rect 117307 277354 117549 277355
rect 117307 277343 117355 277354
rect 117267 277300 117355 277343
rect 117461 277332 117549 277354
rect 118713 277461 118801 277484
rect 118713 277427 118719 277461
rect 118753 277427 118801 277461
rect 118713 277389 118801 277427
rect 120377 277452 120423 277490
rect 120377 277418 120383 277452
rect 120417 277418 120423 277452
rect 120377 277401 120423 277418
rect 120835 277884 120881 277901
rect 120835 277850 120841 277884
rect 120875 277850 120881 277884
rect 120835 277812 120881 277850
rect 120835 277778 120841 277812
rect 120875 277778 120881 277812
rect 120835 277740 120881 277778
rect 120835 277706 120841 277740
rect 120875 277712 120881 277740
rect 120953 277712 121018 278369
rect 121077 278346 121083 278369
rect 121117 278346 121123 278380
rect 121077 278308 121123 278346
rect 121077 278274 121083 278308
rect 121117 278274 121123 278308
rect 121077 278236 121123 278274
rect 121077 278202 121083 278236
rect 121117 278202 121123 278236
rect 121077 278185 121123 278202
rect 121535 278668 121605 278685
rect 121535 278634 121541 278668
rect 121575 278638 121605 278668
rect 121657 278638 121677 278690
rect 121575 278634 121677 278638
rect 121535 278626 121677 278634
rect 121535 278596 121605 278626
rect 121535 278562 121541 278596
rect 121575 278574 121605 278596
rect 121657 278574 121677 278626
rect 121575 278562 121677 278574
rect 121535 278524 121605 278562
rect 121535 278490 121541 278524
rect 121575 278510 121605 278524
rect 121657 278510 121677 278562
rect 121575 278498 121677 278510
rect 121575 278490 121605 278498
rect 121535 278452 121605 278490
rect 121535 278418 121541 278452
rect 121575 278446 121605 278452
rect 121657 278446 121677 278498
rect 121575 278434 121677 278446
rect 121575 278418 121605 278434
rect 121535 278382 121605 278418
rect 121657 278382 121677 278434
rect 121535 278380 121677 278382
rect 121535 278346 121541 278380
rect 121575 278370 121677 278380
rect 121575 278346 121605 278370
rect 121535 278318 121605 278346
rect 121657 278318 121677 278370
rect 122462 278353 123477 278384
rect 121535 278308 121677 278318
rect 121535 278274 121541 278308
rect 121575 278306 121677 278308
rect 122418 278347 123477 278353
rect 122418 278313 122439 278347
rect 122473 278313 122511 278347
rect 122545 278313 122583 278347
rect 122617 278313 122655 278347
rect 122689 278313 122727 278347
rect 122761 278313 122799 278347
rect 122833 278313 122871 278347
rect 122905 278313 122943 278347
rect 122977 278313 123015 278347
rect 123049 278313 123087 278347
rect 123121 278313 123159 278347
rect 123193 278313 123231 278347
rect 123265 278342 123477 278347
rect 123265 278313 123286 278342
rect 122418 278307 123286 278313
rect 121575 278274 121605 278306
rect 121535 278254 121605 278274
rect 121657 278254 121677 278306
rect 121535 278242 121677 278254
rect 121535 278236 121605 278242
rect 121535 278202 121541 278236
rect 121575 278202 121605 278236
rect 121535 278190 121605 278202
rect 121657 278190 121677 278242
rect 121535 278185 121677 278190
rect 121581 278178 121677 278185
rect 121133 278138 121525 278144
rect 121133 278104 121168 278138
rect 121202 278104 121240 278138
rect 121274 278104 121312 278138
rect 121346 278104 121384 278138
rect 121418 278104 121456 278138
rect 121490 278104 121525 278138
rect 121133 277982 121525 278104
rect 121133 277948 121168 277982
rect 121202 277948 121240 277982
rect 121274 277948 121312 277982
rect 121346 277948 121384 277982
rect 121418 277948 121456 277982
rect 121490 277948 121525 277982
rect 121133 277942 121525 277948
rect 121581 278126 121605 278178
rect 121657 278126 121677 278178
rect 121581 278114 121677 278126
rect 121581 278062 121605 278114
rect 121657 278062 121677 278114
rect 121581 278050 121677 278062
rect 121581 277998 121605 278050
rect 121657 277998 121677 278050
rect 121581 277986 121677 277998
rect 121581 277934 121605 277986
rect 121657 277934 121677 277986
rect 121581 277922 121677 277934
rect 121581 277901 121605 277922
rect 121077 277884 121123 277901
rect 121077 277850 121083 277884
rect 121117 277850 121123 277884
rect 121077 277812 121123 277850
rect 121077 277778 121083 277812
rect 121117 277778 121123 277812
rect 121077 277740 121123 277778
rect 121077 277712 121083 277740
rect 120875 277706 121083 277712
rect 121117 277706 121123 277740
rect 120835 277668 121123 277706
rect 120835 277634 120841 277668
rect 120875 277634 121083 277668
rect 121117 277634 121123 277668
rect 120835 277596 121123 277634
rect 120835 277562 120841 277596
rect 120875 277585 121083 277596
rect 120875 277562 120881 277585
rect 120835 277524 120881 277562
rect 120835 277490 120841 277524
rect 120875 277490 120881 277524
rect 120835 277452 120881 277490
rect 120835 277418 120841 277452
rect 120875 277418 120881 277452
rect 120835 277401 120881 277418
rect 118713 277355 118719 277389
rect 118753 277355 118801 277389
rect 118713 277332 118801 277355
rect 117461 277300 117503 277332
rect 115589 277293 116057 277300
rect 115589 277288 115635 277293
rect 115589 277254 115595 277288
rect 115629 277254 115635 277288
rect 115589 277216 115635 277254
rect 115589 277182 115595 277216
rect 115629 277182 115635 277216
rect 115589 277144 115635 277182
rect 115589 277110 115595 277144
rect 115629 277110 115635 277144
rect 115589 277075 115635 277110
rect 116015 277200 116057 277293
rect 116135 277284 117235 277290
rect 116135 277250 116164 277284
rect 116198 277250 116236 277284
rect 116270 277250 116308 277284
rect 116342 277250 116380 277284
rect 116414 277250 116452 277284
rect 116486 277250 116524 277284
rect 116558 277250 116596 277284
rect 116630 277250 116668 277284
rect 116702 277250 116740 277284
rect 116774 277250 116812 277284
rect 116846 277250 116884 277284
rect 116918 277250 116956 277284
rect 116990 277250 117028 277284
rect 117062 277250 117100 277284
rect 117134 277250 117172 277284
rect 117206 277250 117235 277284
rect 116135 277244 117235 277250
rect 117313 277200 117355 277300
rect 116015 277162 117355 277200
rect 112850 277032 112938 277068
rect 112656 277029 112938 277032
rect 112656 276995 112662 277029
rect 112696 277025 112938 277029
rect 112696 276995 112898 277025
rect 112656 276991 112898 276995
rect 112932 276991 112938 277025
rect 112656 276972 112938 276991
rect 111404 276764 111446 276972
rect 112702 276970 112938 276972
rect 111524 276956 112624 276962
rect 111524 276922 111553 276956
rect 111587 276922 111625 276956
rect 111659 276922 111697 276956
rect 111731 276922 111769 276956
rect 111803 276922 111841 276956
rect 111875 276922 111913 276956
rect 111947 276922 111985 276956
rect 112019 276922 112057 276956
rect 112091 276922 112129 276956
rect 112163 276922 112201 276956
rect 112235 276922 112273 276956
rect 112307 276922 112345 276956
rect 112379 276922 112417 276956
rect 112451 276922 112489 276956
rect 112523 276922 112561 276956
rect 112595 276922 112624 276956
rect 111524 276916 112624 276922
rect 111524 276814 112624 276820
rect 111524 276780 111553 276814
rect 111587 276780 111625 276814
rect 111659 276780 111697 276814
rect 111731 276780 111769 276814
rect 111803 276780 111841 276814
rect 111875 276780 111913 276814
rect 111947 276780 111985 276814
rect 112019 276780 112057 276814
rect 112091 276780 112129 276814
rect 112163 276780 112201 276814
rect 112235 276780 112273 276814
rect 112307 276780 112345 276814
rect 112379 276780 112417 276814
rect 112451 276780 112489 276814
rect 112523 276780 112561 276814
rect 112595 276780 112624 276814
rect 111524 276774 112624 276780
rect 112702 276764 112744 276970
rect 112850 276953 112938 276970
rect 112850 276919 112898 276953
rect 112932 276919 112938 276953
rect 112850 276876 112938 276919
rect 114102 277025 114190 277068
rect 116015 277068 116057 277162
rect 116135 277118 117235 277124
rect 116135 277084 116164 277118
rect 116198 277084 116236 277118
rect 116270 277084 116308 277118
rect 116342 277084 116380 277118
rect 116414 277084 116452 277118
rect 116486 277084 116524 277118
rect 116558 277084 116596 277118
rect 116630 277084 116668 277118
rect 116702 277084 116740 277118
rect 116774 277084 116812 277118
rect 116846 277084 116884 277118
rect 116918 277084 116956 277118
rect 116990 277084 117028 277118
rect 117062 277084 117100 277118
rect 117134 277084 117172 277118
rect 117206 277084 117235 277118
rect 116135 277078 117235 277084
rect 117313 277068 117355 277162
rect 117459 277124 117503 277300
rect 117581 277316 118681 277322
rect 117581 277282 117610 277316
rect 117644 277282 117682 277316
rect 117716 277282 117754 277316
rect 117788 277282 117826 277316
rect 117860 277282 117898 277316
rect 117932 277282 117970 277316
rect 118004 277282 118042 277316
rect 118076 277282 118114 277316
rect 118148 277282 118186 277316
rect 118220 277282 118258 277316
rect 118292 277282 118330 277316
rect 118364 277282 118402 277316
rect 118436 277282 118474 277316
rect 118508 277282 118546 277316
rect 118580 277282 118618 277316
rect 118652 277282 118681 277316
rect 117581 277276 118681 277282
rect 117581 277174 118681 277180
rect 117581 277140 117610 277174
rect 117644 277140 117682 277174
rect 117716 277140 117754 277174
rect 117788 277140 117826 277174
rect 117860 277140 117898 277174
rect 117932 277140 117970 277174
rect 118004 277140 118042 277174
rect 118076 277140 118114 277174
rect 118148 277140 118186 277174
rect 118220 277140 118258 277174
rect 118292 277140 118330 277174
rect 118364 277140 118402 277174
rect 118436 277140 118474 277174
rect 118508 277140 118546 277174
rect 118580 277140 118618 277174
rect 118652 277140 118681 277174
rect 117581 277134 118681 277140
rect 118759 277124 118801 277332
rect 120433 277354 120825 277360
rect 120433 277320 120468 277354
rect 120502 277320 120540 277354
rect 120574 277320 120612 277354
rect 120646 277320 120684 277354
rect 120718 277320 120756 277354
rect 120790 277320 120825 277354
rect 120433 277198 120825 277320
rect 120433 277164 120468 277198
rect 120502 277164 120540 277198
rect 120574 277164 120612 277198
rect 120646 277164 120684 277198
rect 120718 277164 120756 277198
rect 120790 277164 120825 277198
rect 120433 277158 120825 277164
rect 117459 277101 117549 277124
rect 117459 277080 117509 277101
rect 114102 276991 114108 277025
rect 114142 276991 114190 277025
rect 114657 277059 114857 277065
rect 114657 277025 114704 277059
rect 114738 277025 114776 277059
rect 114810 277025 114857 277059
rect 114657 277019 114857 277025
rect 115348 277059 115548 277065
rect 115348 277025 115395 277059
rect 115429 277025 115467 277059
rect 115501 277025 115548 277059
rect 115348 277019 115548 277025
rect 116015 277025 116103 277068
rect 114102 276953 114190 276991
rect 114102 276919 114108 276953
rect 114142 276919 114190 276953
rect 114720 276951 114790 277019
rect 114102 276876 114190 276919
rect 114308 276867 114790 276951
rect 114865 276954 114970 276979
rect 114865 276902 114890 276954
rect 114942 276902 114970 276954
rect 114865 276872 114970 276902
rect 115235 276954 115340 276979
rect 115235 276902 115262 276954
rect 115314 276902 115340 276954
rect 115235 276872 115340 276902
rect 115415 276951 115485 277019
rect 116015 276991 116063 277025
rect 116097 276991 116103 277025
rect 116015 276953 116103 276991
rect 112970 276860 114070 276866
rect 112970 276826 112999 276860
rect 113033 276826 113071 276860
rect 113105 276826 113143 276860
rect 113177 276826 113215 276860
rect 113249 276826 113287 276860
rect 113321 276826 113359 276860
rect 113393 276826 113431 276860
rect 113465 276826 113503 276860
rect 113537 276826 113575 276860
rect 113609 276826 113647 276860
rect 113681 276826 113719 276860
rect 113753 276826 113791 276860
rect 113825 276826 113863 276860
rect 113897 276826 113935 276860
rect 113969 276826 114007 276860
rect 114041 276826 114070 276860
rect 112970 276820 114070 276826
rect 111404 276741 111492 276764
rect 111404 276707 111452 276741
rect 111486 276707 111492 276741
rect 111404 276669 111492 276707
rect 111404 276635 111452 276669
rect 111486 276635 111492 276669
rect 111404 276612 111492 276635
rect 112656 276741 112744 276764
rect 114308 276752 114343 276867
rect 114720 276837 114790 276867
rect 115415 276867 115897 276951
rect 116015 276919 116063 276953
rect 116097 276919 116103 276953
rect 116015 276876 116103 276919
rect 117267 277032 117355 277068
rect 117461 277067 117509 277080
rect 117543 277067 117549 277101
rect 117461 277032 117549 277067
rect 117267 277029 117549 277032
rect 117267 277025 117509 277029
rect 117267 276991 117273 277025
rect 117307 276995 117509 277025
rect 117543 276995 117549 277029
rect 117307 276991 117549 276995
rect 117267 276972 117549 276991
rect 118713 277101 118801 277124
rect 118713 277067 118719 277101
rect 118753 277067 118801 277101
rect 118713 277029 118801 277067
rect 118713 276995 118719 277029
rect 118753 276995 118801 277029
rect 118713 276972 118801 276995
rect 117267 276970 117503 276972
rect 117267 276953 117355 276970
rect 117267 276919 117273 276953
rect 117307 276919 117355 276953
rect 117267 276876 117355 276919
rect 115415 276837 115485 276867
rect 114657 276831 114857 276837
rect 114657 276797 114704 276831
rect 114738 276797 114776 276831
rect 114810 276797 114857 276831
rect 114657 276791 114857 276797
rect 115348 276831 115548 276837
rect 115348 276797 115395 276831
rect 115429 276797 115467 276831
rect 115501 276797 115548 276831
rect 115348 276791 115548 276797
rect 112656 276707 112662 276741
rect 112696 276707 112744 276741
rect 113843 276722 114343 276752
rect 112656 276669 112744 276707
rect 113000 276716 114343 276722
rect 113000 276682 113029 276716
rect 113063 276682 113101 276716
rect 113135 276682 113173 276716
rect 113207 276682 113245 276716
rect 113279 276682 113317 276716
rect 113351 276682 113389 276716
rect 113423 276682 113461 276716
rect 113495 276682 113533 276716
rect 113567 276682 113605 276716
rect 113639 276682 113677 276716
rect 113711 276682 113749 276716
rect 113783 276682 113821 276716
rect 113855 276682 113893 276716
rect 113927 276682 113965 276716
rect 113999 276682 114037 276716
rect 114071 276711 114343 276716
rect 114570 276758 114616 276781
rect 114570 276724 114576 276758
rect 114610 276724 114616 276758
rect 114071 276682 114100 276711
rect 113000 276676 114100 276682
rect 114570 276686 114616 276724
rect 112656 276635 112662 276669
rect 112696 276635 112744 276669
rect 112656 276612 112744 276635
rect 111404 276404 111446 276612
rect 111524 276596 112624 276602
rect 111524 276562 111553 276596
rect 111587 276562 111625 276596
rect 111659 276562 111697 276596
rect 111731 276562 111769 276596
rect 111803 276562 111841 276596
rect 111875 276562 111913 276596
rect 111947 276562 111985 276596
rect 112019 276562 112057 276596
rect 112091 276562 112129 276596
rect 112163 276562 112201 276596
rect 112235 276562 112273 276596
rect 112307 276562 112345 276596
rect 112379 276562 112417 276596
rect 112451 276562 112489 276596
rect 112523 276562 112561 276596
rect 112595 276562 112624 276596
rect 111524 276556 112624 276562
rect 111524 276454 112624 276460
rect 111524 276420 111553 276454
rect 111587 276420 111625 276454
rect 111659 276420 111697 276454
rect 111731 276420 111769 276454
rect 111803 276420 111841 276454
rect 111875 276420 111913 276454
rect 111947 276420 111985 276454
rect 112019 276420 112057 276454
rect 112091 276420 112129 276454
rect 112163 276420 112201 276454
rect 112235 276420 112273 276454
rect 112307 276420 112345 276454
rect 112379 276420 112417 276454
rect 112451 276420 112489 276454
rect 112523 276420 112561 276454
rect 112595 276420 112624 276454
rect 111524 276414 112624 276420
rect 112702 276404 112744 276612
rect 111404 276381 111492 276404
rect 111404 276347 111452 276381
rect 111486 276347 111492 276381
rect 111404 276309 111492 276347
rect 111404 276275 111452 276309
rect 111486 276275 111492 276309
rect 111404 276252 111492 276275
rect 112656 276381 112744 276404
rect 112656 276347 112662 276381
rect 112696 276347 112744 276381
rect 112656 276309 112744 276347
rect 112656 276275 112662 276309
rect 112696 276275 112744 276309
rect 112656 276252 112744 276275
rect 112874 276647 112968 276666
rect 112874 276613 112928 276647
rect 112962 276613 112968 276647
rect 112874 276594 112968 276613
rect 114132 276647 114226 276666
rect 114132 276613 114138 276647
rect 114172 276613 114226 276647
rect 114132 276594 114226 276613
rect 112874 276502 112922 276594
rect 113000 276578 114100 276584
rect 113000 276544 113029 276578
rect 113063 276544 113101 276578
rect 113135 276544 113173 276578
rect 113207 276544 113245 276578
rect 113279 276544 113317 276578
rect 113351 276544 113389 276578
rect 113423 276544 113461 276578
rect 113495 276544 113533 276578
rect 113567 276544 113605 276578
rect 113639 276544 113677 276578
rect 113711 276544 113749 276578
rect 113783 276544 113821 276578
rect 113855 276544 113893 276578
rect 113927 276544 113965 276578
rect 113999 276544 114037 276578
rect 114071 276544 114100 276578
rect 113000 276538 114100 276544
rect 114178 276502 114226 276594
rect 112874 276458 114226 276502
rect 114324 276619 114396 276660
rect 114570 276652 114576 276686
rect 114610 276652 114616 276686
rect 114570 276629 114616 276652
rect 114898 276758 114944 276781
rect 114898 276724 114904 276758
rect 114938 276724 114944 276758
rect 114898 276686 114944 276724
rect 114898 276652 114904 276686
rect 114938 276652 114944 276686
rect 114898 276629 114944 276652
rect 115261 276758 115307 276781
rect 115261 276724 115267 276758
rect 115301 276724 115307 276758
rect 115261 276686 115307 276724
rect 115261 276652 115267 276686
rect 115301 276652 115307 276686
rect 115261 276629 115307 276652
rect 115589 276758 115635 276781
rect 115589 276724 115595 276758
rect 115629 276724 115635 276758
rect 115589 276686 115635 276724
rect 115862 276752 115897 276867
rect 116135 276860 117235 276866
rect 116135 276826 116164 276860
rect 116198 276826 116236 276860
rect 116270 276826 116308 276860
rect 116342 276826 116380 276860
rect 116414 276826 116452 276860
rect 116486 276826 116524 276860
rect 116558 276826 116596 276860
rect 116630 276826 116668 276860
rect 116702 276826 116740 276860
rect 116774 276826 116812 276860
rect 116846 276826 116884 276860
rect 116918 276826 116956 276860
rect 116990 276826 117028 276860
rect 117062 276826 117100 276860
rect 117134 276826 117172 276860
rect 117206 276826 117235 276860
rect 116135 276820 117235 276826
rect 117461 276764 117503 276970
rect 117581 276956 118681 276962
rect 117581 276922 117610 276956
rect 117644 276922 117682 276956
rect 117716 276922 117754 276956
rect 117788 276922 117826 276956
rect 117860 276922 117898 276956
rect 117932 276922 117970 276956
rect 118004 276922 118042 276956
rect 118076 276922 118114 276956
rect 118148 276922 118186 276956
rect 118220 276922 118258 276956
rect 118292 276922 118330 276956
rect 118364 276922 118402 276956
rect 118436 276922 118474 276956
rect 118508 276922 118546 276956
rect 118580 276922 118618 276956
rect 118652 276922 118681 276956
rect 117581 276916 118681 276922
rect 117581 276814 118681 276820
rect 117581 276780 117610 276814
rect 117644 276780 117682 276814
rect 117716 276780 117754 276814
rect 117788 276780 117826 276814
rect 117860 276780 117898 276814
rect 117932 276780 117970 276814
rect 118004 276780 118042 276814
rect 118076 276780 118114 276814
rect 118148 276780 118186 276814
rect 118220 276780 118258 276814
rect 118292 276780 118330 276814
rect 118364 276780 118402 276814
rect 118436 276780 118474 276814
rect 118508 276780 118546 276814
rect 118580 276780 118618 276814
rect 118652 276780 118681 276814
rect 117581 276774 118681 276780
rect 118759 276764 118801 276972
rect 115862 276722 116362 276752
rect 117461 276741 117549 276764
rect 115862 276716 117205 276722
rect 115862 276711 116134 276716
rect 115589 276652 115595 276686
rect 115629 276652 115635 276686
rect 116105 276682 116134 276711
rect 116168 276682 116206 276716
rect 116240 276682 116278 276716
rect 116312 276682 116350 276716
rect 116384 276682 116422 276716
rect 116456 276682 116494 276716
rect 116528 276682 116566 276716
rect 116600 276682 116638 276716
rect 116672 276682 116710 276716
rect 116744 276682 116782 276716
rect 116816 276682 116854 276716
rect 116888 276682 116926 276716
rect 116960 276682 116998 276716
rect 117032 276682 117070 276716
rect 117104 276682 117142 276716
rect 117176 276682 117205 276716
rect 116105 276676 117205 276682
rect 117461 276707 117509 276741
rect 117543 276707 117549 276741
rect 117461 276669 117549 276707
rect 115589 276629 115635 276652
rect 115809 276619 115881 276660
rect 114324 276585 114342 276619
rect 114376 276585 114396 276619
rect 114324 276529 114396 276585
rect 114657 276613 114857 276619
rect 114657 276579 114704 276613
rect 114738 276579 114776 276613
rect 114810 276579 114857 276613
rect 114657 276573 114857 276579
rect 115348 276613 115548 276619
rect 115348 276579 115395 276613
rect 115429 276579 115467 276613
rect 115501 276579 115548 276613
rect 115348 276573 115548 276579
rect 115809 276585 115828 276619
rect 115862 276585 115881 276619
rect 114843 276529 115030 276544
rect 114324 276484 114781 276529
rect 112874 276368 112922 276458
rect 113000 276418 114100 276424
rect 113000 276384 113029 276418
rect 113063 276384 113101 276418
rect 113135 276384 113173 276418
rect 113207 276384 113245 276418
rect 113279 276384 113317 276418
rect 113351 276384 113389 276418
rect 113423 276384 113461 276418
rect 113495 276384 113533 276418
rect 113567 276384 113605 276418
rect 113639 276384 113677 276418
rect 113711 276384 113749 276418
rect 113783 276384 113821 276418
rect 113855 276384 113893 276418
rect 113927 276384 113965 276418
rect 113999 276384 114037 276418
rect 114071 276384 114100 276418
rect 113000 276378 114100 276384
rect 114178 276368 114226 276458
rect 114737 276429 114781 276484
rect 114843 276477 114891 276529
rect 114943 276477 115030 276529
rect 114843 276459 115030 276477
rect 115175 276529 115362 276544
rect 115809 276529 115881 276585
rect 115175 276477 115262 276529
rect 115314 276477 115362 276529
rect 115175 276459 115362 276477
rect 115424 276484 115881 276529
rect 115979 276647 116073 276666
rect 115979 276613 116033 276647
rect 116067 276613 116073 276647
rect 115979 276594 116073 276613
rect 117237 276647 117331 276666
rect 117237 276613 117243 276647
rect 117277 276613 117331 276647
rect 117237 276594 117331 276613
rect 115979 276502 116027 276594
rect 116105 276578 117205 276584
rect 116105 276544 116134 276578
rect 116168 276544 116206 276578
rect 116240 276544 116278 276578
rect 116312 276544 116350 276578
rect 116384 276544 116422 276578
rect 116456 276544 116494 276578
rect 116528 276544 116566 276578
rect 116600 276544 116638 276578
rect 116672 276544 116710 276578
rect 116744 276544 116782 276578
rect 116816 276544 116854 276578
rect 116888 276544 116926 276578
rect 116960 276544 116998 276578
rect 117032 276544 117070 276578
rect 117104 276544 117142 276578
rect 117176 276544 117205 276578
rect 116105 276538 117205 276544
rect 117283 276502 117331 276594
rect 115424 276429 115468 276484
rect 115979 276458 117331 276502
rect 114657 276423 114857 276429
rect 114657 276389 114704 276423
rect 114738 276389 114776 276423
rect 114810 276389 114857 276423
rect 114657 276383 114857 276389
rect 115348 276423 115548 276429
rect 115348 276389 115395 276423
rect 115429 276389 115467 276423
rect 115501 276389 115548 276423
rect 115348 276383 115548 276389
rect 112874 276349 112968 276368
rect 112874 276315 112928 276349
rect 112962 276315 112968 276349
rect 112874 276296 112968 276315
rect 114132 276349 114226 276368
rect 114132 276315 114138 276349
rect 114172 276315 114226 276349
rect 114132 276296 114226 276315
rect 114570 276350 114616 276373
rect 114570 276316 114576 276350
rect 114610 276316 114616 276350
rect 111524 276236 112624 276242
rect 111524 276202 111553 276236
rect 111587 276202 111625 276236
rect 111659 276202 111697 276236
rect 111731 276202 111769 276236
rect 111803 276202 111841 276236
rect 111875 276202 111913 276236
rect 111947 276202 111985 276236
rect 112019 276202 112057 276236
rect 112091 276202 112129 276236
rect 112163 276202 112201 276236
rect 112235 276202 112273 276236
rect 112307 276202 112345 276236
rect 112379 276202 112417 276236
rect 112451 276202 112489 276236
rect 112523 276202 112561 276236
rect 112595 276202 112624 276236
rect 111524 276198 112624 276202
rect 112874 276202 112922 276296
rect 114327 276291 114395 276292
rect 114570 276291 114616 276316
rect 113000 276280 114100 276286
rect 113000 276246 113029 276280
rect 113063 276246 113101 276280
rect 113135 276246 113173 276280
rect 113207 276246 113245 276280
rect 113279 276246 113317 276280
rect 113351 276246 113389 276280
rect 113423 276246 113461 276280
rect 113495 276246 113533 276280
rect 113567 276246 113605 276280
rect 113639 276246 113677 276280
rect 113711 276246 113749 276280
rect 113783 276246 113821 276280
rect 113855 276246 113893 276280
rect 113927 276246 113965 276280
rect 113999 276246 114037 276280
rect 114071 276246 114100 276280
rect 113000 276240 114100 276246
rect 114327 276278 114616 276291
rect 114327 276244 114576 276278
rect 114610 276244 114616 276278
rect 114327 276231 114616 276244
rect 114327 276202 114395 276231
rect 114570 276221 114616 276231
rect 114898 276350 114944 276373
rect 114898 276316 114904 276350
rect 114938 276316 114944 276350
rect 114898 276278 114944 276316
rect 114898 276244 114904 276278
rect 114938 276244 114944 276278
rect 114898 276221 114944 276244
rect 115261 276350 115307 276373
rect 115261 276316 115267 276350
rect 115301 276316 115307 276350
rect 115261 276278 115307 276316
rect 115261 276244 115267 276278
rect 115301 276244 115307 276278
rect 115261 276221 115307 276244
rect 115589 276350 115635 276373
rect 115589 276316 115595 276350
rect 115629 276316 115635 276350
rect 115589 276291 115635 276316
rect 115979 276368 116027 276458
rect 116105 276418 117205 276424
rect 116105 276384 116134 276418
rect 116168 276384 116206 276418
rect 116240 276384 116278 276418
rect 116312 276384 116350 276418
rect 116384 276384 116422 276418
rect 116456 276384 116494 276418
rect 116528 276384 116566 276418
rect 116600 276384 116638 276418
rect 116672 276384 116710 276418
rect 116744 276384 116782 276418
rect 116816 276384 116854 276418
rect 116888 276384 116926 276418
rect 116960 276384 116998 276418
rect 117032 276384 117070 276418
rect 117104 276384 117142 276418
rect 117176 276384 117205 276418
rect 116105 276378 117205 276384
rect 117283 276368 117331 276458
rect 115979 276349 116073 276368
rect 115979 276315 116033 276349
rect 116067 276315 116073 276349
rect 115979 276296 116073 276315
rect 117237 276349 117331 276368
rect 117237 276315 117243 276349
rect 117277 276315 117331 276349
rect 117237 276296 117331 276315
rect 115810 276291 115878 276292
rect 115589 276278 115878 276291
rect 115589 276244 115595 276278
rect 115629 276244 115878 276278
rect 115589 276231 115878 276244
rect 116105 276280 117205 276286
rect 116105 276246 116134 276280
rect 116168 276246 116206 276280
rect 116240 276246 116278 276280
rect 116312 276246 116350 276280
rect 116384 276246 116422 276280
rect 116456 276246 116494 276280
rect 116528 276246 116566 276280
rect 116600 276246 116638 276280
rect 116672 276246 116710 276280
rect 116744 276246 116782 276280
rect 116816 276246 116854 276280
rect 116888 276246 116926 276280
rect 116960 276246 116998 276280
rect 117032 276246 117070 276280
rect 117104 276246 117142 276280
rect 117176 276246 117205 276280
rect 116105 276240 117205 276246
rect 115589 276221 115635 276231
rect 112874 276198 114395 276202
rect 111524 276196 114395 276198
rect 112044 276162 114395 276196
rect 114657 276205 114857 276211
rect 114657 276171 114704 276205
rect 114738 276171 114776 276205
rect 114810 276171 114857 276205
rect 114657 276165 114857 276171
rect 115348 276205 115548 276211
rect 115348 276171 115395 276205
rect 115429 276171 115467 276205
rect 115501 276171 115548 276205
rect 115348 276165 115548 276171
rect 115810 276202 115878 276231
rect 117283 276202 117331 276296
rect 117461 276635 117509 276669
rect 117543 276635 117549 276669
rect 117461 276612 117549 276635
rect 118713 276741 118801 276764
rect 118713 276707 118719 276741
rect 118753 276707 118801 276741
rect 118713 276669 118801 276707
rect 118713 276635 118719 276669
rect 118753 276635 118801 276669
rect 118713 276612 118801 276635
rect 120377 277100 120423 277117
rect 120377 277066 120383 277100
rect 120417 277066 120423 277100
rect 120377 277028 120423 277066
rect 120377 276994 120383 277028
rect 120417 276994 120423 277028
rect 120377 276956 120423 276994
rect 120377 276922 120383 276956
rect 120417 276922 120423 276956
rect 120377 276884 120423 276922
rect 120377 276850 120383 276884
rect 120417 276850 120423 276884
rect 120377 276812 120423 276850
rect 120377 276778 120383 276812
rect 120417 276778 120423 276812
rect 120377 276740 120423 276778
rect 120377 276706 120383 276740
rect 120417 276706 120423 276740
rect 120377 276668 120423 276706
rect 120377 276634 120383 276668
rect 120417 276634 120423 276668
rect 120377 276617 120423 276634
rect 120835 277100 120881 277117
rect 120835 277066 120841 277100
rect 120875 277066 120881 277100
rect 120835 277028 120881 277066
rect 120835 276994 120841 277028
rect 120875 276994 120881 277028
rect 120835 276956 120881 276994
rect 120835 276922 120841 276956
rect 120875 276928 120881 276956
rect 120953 277072 121018 277585
rect 121077 277562 121083 277585
rect 121117 277562 121123 277596
rect 121077 277524 121123 277562
rect 121077 277490 121083 277524
rect 121117 277490 121123 277524
rect 121077 277452 121123 277490
rect 121077 277418 121083 277452
rect 121117 277418 121123 277452
rect 121077 277401 121123 277418
rect 121535 277884 121605 277901
rect 121535 277850 121541 277884
rect 121575 277870 121605 277884
rect 121657 277870 121677 277922
rect 121575 277858 121677 277870
rect 121575 277850 121605 277858
rect 121535 277812 121605 277850
rect 121535 277778 121541 277812
rect 121575 277806 121605 277812
rect 121657 277806 121677 277858
rect 121575 277794 121677 277806
rect 121575 277778 121605 277794
rect 121535 277742 121605 277778
rect 121657 277742 121677 277794
rect 122362 278226 122408 278266
rect 122362 278192 122368 278226
rect 122402 278192 122408 278226
rect 122362 278154 122408 278192
rect 122362 278120 122368 278154
rect 122402 278120 122408 278154
rect 122362 278082 122408 278120
rect 122362 278048 122368 278082
rect 122402 278048 122408 278082
rect 122362 278010 122408 278048
rect 122362 277976 122368 278010
rect 122402 277976 122408 278010
rect 122362 277938 122408 277976
rect 122362 277904 122368 277938
rect 122402 277904 122408 277938
rect 122362 277866 122408 277904
rect 122362 277832 122368 277866
rect 122402 277832 122408 277866
rect 122362 277792 122408 277832
rect 123296 278226 123342 278266
rect 123296 278192 123302 278226
rect 123336 278192 123342 278226
rect 123296 278154 123342 278192
rect 123296 278120 123302 278154
rect 123336 278120 123342 278154
rect 123296 278082 123342 278120
rect 123296 278048 123302 278082
rect 123336 278048 123342 278082
rect 123296 278010 123342 278048
rect 123296 277976 123302 278010
rect 123336 277976 123342 278010
rect 123296 277938 123342 277976
rect 123296 277904 123302 277938
rect 123336 277904 123342 277938
rect 123296 277866 123342 277904
rect 123296 277832 123302 277866
rect 123336 277832 123342 277866
rect 123296 277792 123342 277832
rect 121535 277740 121677 277742
rect 121535 277706 121541 277740
rect 121575 277730 121677 277740
rect 121575 277706 121605 277730
rect 121535 277678 121605 277706
rect 121657 277678 121677 277730
rect 121535 277668 121677 277678
rect 122418 277745 123286 277751
rect 122418 277711 122439 277745
rect 122473 277711 122511 277745
rect 122545 277711 122583 277745
rect 122617 277711 122655 277745
rect 122689 277711 122727 277745
rect 122761 277711 122799 277745
rect 122833 277711 122871 277745
rect 122905 277711 122943 277745
rect 122977 277711 123015 277745
rect 123049 277711 123087 277745
rect 123121 277711 123159 277745
rect 123193 277711 123231 277745
rect 123265 277711 123286 277745
rect 122418 277707 123286 277711
rect 123440 277707 123477 278342
rect 123660 278161 124206 278167
rect 123660 278127 123700 278161
rect 123734 278127 123772 278161
rect 123806 278127 123844 278161
rect 123878 278127 123916 278161
rect 123950 278127 123988 278161
rect 124022 278127 124060 278161
rect 124094 278127 124132 278161
rect 124166 278127 124206 278161
rect 123660 278121 124206 278127
rect 122418 277670 123477 277707
rect 121535 277634 121541 277668
rect 121575 277666 121677 277668
rect 121575 277634 121605 277666
rect 121535 277614 121605 277634
rect 121657 277614 121677 277666
rect 121535 277602 121677 277614
rect 121535 277596 121605 277602
rect 121535 277562 121541 277596
rect 121575 277562 121605 277596
rect 121535 277550 121605 277562
rect 121657 277550 121677 277602
rect 121535 277538 121677 277550
rect 121535 277524 121605 277538
rect 121535 277490 121541 277524
rect 121575 277490 121605 277524
rect 121535 277486 121605 277490
rect 121657 277486 121677 277538
rect 121535 277452 121677 277486
rect 121535 277418 121541 277452
rect 121575 277418 121677 277452
rect 121535 277401 121677 277418
rect 122364 277581 123212 277587
rect 122364 277547 122439 277581
rect 122473 277547 122511 277581
rect 122545 277547 122583 277581
rect 122617 277547 122655 277581
rect 122689 277547 122727 277581
rect 122761 277547 122799 277581
rect 122833 277547 122871 277581
rect 122905 277547 122943 277581
rect 122977 277547 123015 277581
rect 123049 277547 123087 277581
rect 123121 277547 123159 277581
rect 123193 277547 123212 277581
rect 122364 277541 123212 277547
rect 122364 277500 122420 277541
rect 123440 277500 123477 277670
rect 123604 278042 123650 278080
rect 123604 278008 123610 278042
rect 123644 278008 123650 278042
rect 123604 277970 123650 278008
rect 123604 277936 123610 277970
rect 123644 277936 123650 277970
rect 123604 277898 123650 277936
rect 123604 277864 123610 277898
rect 123644 277864 123650 277898
rect 123604 277826 123650 277864
rect 123604 277792 123610 277826
rect 123644 277792 123650 277826
rect 123604 277754 123650 277792
rect 123604 277720 123610 277754
rect 123644 277720 123650 277754
rect 123604 277682 123650 277720
rect 123604 277648 123610 277682
rect 123644 277648 123650 277682
rect 123604 277610 123650 277648
rect 123604 277576 123610 277610
rect 123644 277576 123650 277610
rect 123604 277538 123650 277576
rect 123604 277504 123610 277538
rect 123644 277504 123650 277538
rect 123604 277500 123650 277504
rect 122364 277467 122410 277500
rect 122364 277433 122370 277467
rect 122404 277433 122410 277467
rect 121133 277354 121525 277360
rect 121133 277320 121168 277354
rect 121202 277320 121240 277354
rect 121274 277320 121312 277354
rect 121346 277320 121384 277354
rect 121418 277320 121456 277354
rect 121490 277320 121525 277354
rect 121133 277198 121525 277320
rect 121133 277164 121168 277198
rect 121202 277164 121240 277198
rect 121274 277164 121312 277198
rect 121346 277164 121384 277198
rect 121418 277164 121456 277198
rect 121490 277164 121525 277198
rect 121133 277158 121525 277164
rect 121581 277117 121624 277401
rect 122364 277400 122410 277433
rect 123222 277467 123650 277500
rect 123222 277433 123228 277467
rect 123262 277466 123650 277467
rect 123262 277433 123610 277466
rect 123222 277432 123610 277433
rect 123644 277432 123650 277466
rect 123222 277400 123650 277432
rect 122364 277359 122420 277400
rect 123604 277394 123650 277400
rect 124216 278042 124262 278080
rect 124216 278008 124222 278042
rect 124256 278008 124262 278042
rect 124216 277970 124262 278008
rect 124216 277936 124222 277970
rect 124256 277936 124262 277970
rect 124216 277898 124262 277936
rect 124216 277864 124222 277898
rect 124256 277864 124262 277898
rect 124216 277826 124262 277864
rect 124216 277792 124222 277826
rect 124256 277792 124262 277826
rect 124216 277754 124262 277792
rect 124216 277720 124222 277754
rect 124256 277720 124262 277754
rect 124216 277682 124262 277720
rect 124216 277648 124222 277682
rect 124256 277648 124262 277682
rect 124216 277610 124262 277648
rect 124216 277576 124222 277610
rect 124256 277576 124262 277610
rect 124216 277538 124262 277576
rect 124216 277504 124222 277538
rect 124256 277528 124262 277538
rect 124256 277504 124567 277528
rect 124216 277466 124567 277504
rect 124216 277432 124222 277466
rect 124256 277432 124567 277466
rect 124216 277394 124567 277432
rect 122364 277353 123212 277359
rect 122364 277319 122439 277353
rect 122473 277319 122511 277353
rect 122545 277319 122583 277353
rect 122617 277319 122655 277353
rect 122689 277319 122727 277353
rect 122761 277319 122799 277353
rect 122833 277319 122871 277353
rect 122905 277319 122943 277353
rect 122977 277319 123015 277353
rect 123049 277319 123087 277353
rect 123121 277319 123159 277353
rect 123193 277319 123212 277353
rect 122364 277313 123212 277319
rect 123660 277347 124206 277353
rect 123660 277313 123700 277347
rect 123734 277313 123772 277347
rect 123806 277313 123844 277347
rect 123878 277313 123916 277347
rect 123950 277313 123988 277347
rect 124022 277313 124060 277347
rect 124094 277313 124132 277347
rect 124166 277313 124206 277347
rect 123660 277307 124206 277313
rect 120953 277020 120959 277072
rect 121011 277020 121018 277072
rect 120953 277008 121018 277020
rect 120953 276956 120959 277008
rect 121011 276956 121018 277008
rect 120953 276944 121018 276956
rect 120953 276928 120959 276944
rect 120875 276922 120959 276928
rect 120835 276892 120959 276922
rect 121011 276928 121018 276944
rect 121077 277100 121123 277117
rect 121077 277066 121083 277100
rect 121117 277066 121123 277100
rect 121077 277028 121123 277066
rect 121077 276994 121083 277028
rect 121117 276994 121123 277028
rect 121077 276956 121123 276994
rect 121077 276928 121083 276956
rect 121011 276922 121083 276928
rect 121117 276922 121123 276956
rect 121011 276892 121123 276922
rect 120835 276884 121123 276892
rect 120835 276850 120841 276884
rect 120875 276880 121083 276884
rect 120875 276850 120959 276880
rect 120835 276828 120959 276850
rect 121011 276850 121083 276880
rect 121117 276850 121123 276884
rect 121011 276828 121123 276850
rect 120835 276812 121123 276828
rect 120835 276778 120841 276812
rect 120875 276801 121083 276812
rect 120875 276778 120881 276801
rect 120835 276740 120881 276778
rect 120835 276706 120841 276740
rect 120875 276706 120881 276740
rect 120835 276668 120881 276706
rect 120835 276634 120841 276668
rect 120875 276634 120881 276668
rect 120835 276617 120881 276634
rect 121077 276778 121083 276801
rect 121117 276778 121123 276812
rect 121077 276740 121123 276778
rect 121077 276706 121083 276740
rect 121117 276706 121123 276740
rect 121077 276668 121123 276706
rect 121077 276634 121083 276668
rect 121117 276634 121123 276668
rect 121077 276617 121123 276634
rect 121535 277100 121624 277117
rect 121535 277066 121541 277100
rect 121575 277066 121624 277100
rect 123792 277076 123945 277307
rect 121535 277028 121624 277066
rect 121535 276994 121541 277028
rect 121575 276994 121624 277028
rect 121535 276956 121624 276994
rect 121535 276922 121541 276956
rect 121575 276922 121624 276956
rect 121535 276884 121624 276922
rect 121535 276850 121541 276884
rect 121575 276850 121624 276884
rect 121535 276812 121624 276850
rect 123686 277010 123945 277076
rect 123686 276904 123771 277010
rect 123877 276904 123945 277010
rect 123686 276837 123945 276904
rect 121535 276778 121541 276812
rect 121575 276778 121624 276812
rect 121535 276740 121624 276778
rect 121535 276706 121541 276740
rect 121575 276706 121624 276740
rect 122442 276749 123828 276755
rect 122442 276715 122470 276749
rect 122504 276715 122542 276749
rect 122576 276715 122614 276749
rect 122648 276715 122686 276749
rect 122720 276715 122758 276749
rect 122792 276715 122830 276749
rect 122864 276715 122902 276749
rect 122936 276715 122974 276749
rect 123008 276715 123046 276749
rect 123080 276715 123118 276749
rect 123152 276715 123190 276749
rect 123224 276715 123262 276749
rect 123296 276715 123334 276749
rect 123368 276715 123406 276749
rect 123440 276715 123478 276749
rect 123512 276715 123550 276749
rect 123584 276715 123622 276749
rect 123656 276715 123694 276749
rect 123728 276715 123766 276749
rect 123800 276715 123828 276749
rect 122442 276709 123828 276715
rect 121535 276668 121624 276706
rect 121535 276634 121541 276668
rect 121575 276634 121624 276668
rect 121535 276617 121624 276634
rect 122386 276633 122432 276668
rect 117461 276404 117503 276612
rect 117581 276596 118681 276602
rect 117581 276562 117610 276596
rect 117644 276562 117682 276596
rect 117716 276562 117754 276596
rect 117788 276562 117826 276596
rect 117860 276562 117898 276596
rect 117932 276562 117970 276596
rect 118004 276562 118042 276596
rect 118076 276562 118114 276596
rect 118148 276562 118186 276596
rect 118220 276562 118258 276596
rect 118292 276562 118330 276596
rect 118364 276562 118402 276596
rect 118436 276562 118474 276596
rect 118508 276562 118546 276596
rect 118580 276562 118618 276596
rect 118652 276562 118681 276596
rect 117581 276556 118681 276562
rect 117581 276454 118681 276460
rect 117581 276420 117610 276454
rect 117644 276420 117682 276454
rect 117716 276420 117754 276454
rect 117788 276420 117826 276454
rect 117860 276420 117898 276454
rect 117932 276420 117970 276454
rect 118004 276420 118042 276454
rect 118076 276420 118114 276454
rect 118148 276420 118186 276454
rect 118220 276420 118258 276454
rect 118292 276420 118330 276454
rect 118364 276420 118402 276454
rect 118436 276420 118474 276454
rect 118508 276420 118546 276454
rect 118580 276420 118618 276454
rect 118652 276420 118681 276454
rect 117581 276414 118681 276420
rect 118759 276404 118801 276612
rect 122386 276599 122392 276633
rect 122426 276599 122432 276633
rect 117461 276381 117549 276404
rect 117461 276347 117509 276381
rect 117543 276347 117549 276381
rect 117461 276309 117549 276347
rect 117461 276275 117509 276309
rect 117543 276275 117549 276309
rect 117461 276252 117549 276275
rect 118713 276381 118801 276404
rect 118713 276347 118719 276381
rect 118753 276347 118801 276381
rect 120433 276570 120825 276576
rect 120433 276536 120468 276570
rect 120502 276536 120540 276570
rect 120574 276536 120612 276570
rect 120646 276536 120684 276570
rect 120718 276536 120756 276570
rect 120790 276536 120825 276570
rect 120433 276414 120825 276536
rect 120433 276380 120468 276414
rect 120502 276380 120540 276414
rect 120574 276380 120612 276414
rect 120646 276380 120684 276414
rect 120718 276380 120756 276414
rect 120790 276380 120825 276414
rect 120433 276374 120825 276380
rect 121133 276570 121525 276576
rect 121133 276536 121168 276570
rect 121202 276536 121240 276570
rect 121274 276536 121312 276570
rect 121346 276536 121384 276570
rect 121418 276536 121456 276570
rect 121490 276536 121525 276570
rect 121133 276414 121525 276536
rect 122386 276561 122432 276599
rect 122386 276527 122392 276561
rect 122426 276527 122432 276561
rect 122386 276492 122432 276527
rect 123838 276646 123884 276668
rect 123838 276633 124112 276646
rect 123838 276599 123844 276633
rect 123878 276599 124112 276633
rect 123838 276561 124112 276599
rect 123838 276527 123844 276561
rect 123878 276527 124112 276561
rect 123838 276514 124112 276527
rect 123838 276492 123884 276514
rect 121133 276380 121168 276414
rect 121202 276380 121240 276414
rect 121274 276380 121312 276414
rect 121346 276380 121384 276414
rect 121418 276380 121456 276414
rect 121490 276380 121525 276414
rect 122442 276445 123828 276451
rect 122442 276411 122470 276445
rect 122504 276411 122542 276445
rect 122576 276411 122614 276445
rect 122648 276411 122686 276445
rect 122720 276411 122758 276445
rect 122792 276411 122830 276445
rect 122864 276411 122902 276445
rect 122936 276411 122974 276445
rect 123008 276411 123046 276445
rect 123080 276411 123118 276445
rect 123152 276411 123190 276445
rect 123224 276411 123262 276445
rect 123296 276411 123334 276445
rect 123368 276411 123406 276445
rect 123440 276411 123478 276445
rect 123512 276411 123550 276445
rect 123584 276411 123622 276445
rect 123656 276411 123694 276445
rect 123728 276411 123766 276445
rect 123800 276411 123828 276445
rect 122442 276405 123828 276411
rect 121133 276374 121525 276380
rect 118713 276309 118801 276347
rect 118713 276275 118719 276309
rect 118753 276275 118801 276309
rect 118713 276252 118801 276275
rect 120377 276316 120423 276333
rect 120377 276282 120383 276316
rect 120417 276282 120423 276316
rect 120377 276244 120423 276282
rect 115810 276198 117331 276202
rect 117581 276236 118681 276242
rect 117581 276202 117610 276236
rect 117644 276202 117682 276236
rect 117716 276202 117754 276236
rect 117788 276202 117826 276236
rect 117860 276202 117898 276236
rect 117932 276202 117970 276236
rect 118004 276202 118042 276236
rect 118076 276202 118114 276236
rect 118148 276202 118186 276236
rect 118220 276202 118258 276236
rect 118292 276202 118330 276236
rect 118364 276202 118402 276236
rect 118436 276202 118474 276236
rect 118508 276202 118546 276236
rect 118580 276202 118618 276236
rect 118652 276202 118681 276236
rect 117581 276198 118681 276202
rect 115810 276196 118681 276198
rect 120377 276210 120383 276244
rect 120417 276210 120423 276244
rect 112719 276120 112924 276162
rect 113982 276088 114266 276098
rect 114724 276088 114783 276165
rect 113982 276067 114783 276088
rect 113982 276033 114034 276067
rect 114068 276033 114106 276067
rect 114140 276033 114178 276067
rect 114212 276033 114783 276067
rect 113982 275999 114783 276033
rect 115422 276088 115481 276165
rect 115810 276162 118161 276196
rect 120377 276172 120423 276210
rect 117281 276120 117486 276162
rect 120377 276138 120383 276172
rect 120417 276138 120423 276172
rect 120377 276100 120423 276138
rect 115939 276088 116223 276098
rect 115422 276067 116223 276088
rect 115422 276033 115992 276067
rect 116026 276033 116064 276067
rect 116098 276033 116136 276067
rect 116170 276033 116223 276067
rect 115422 275999 116223 276033
rect 113982 275998 114266 275999
rect 115939 275998 116223 275999
rect 120377 276066 120383 276100
rect 120417 276066 120423 276100
rect 120377 276028 120423 276066
rect 120377 275994 120383 276028
rect 120417 275994 120423 276028
rect 120377 275956 120423 275994
rect 120377 275922 120383 275956
rect 120417 275922 120423 275956
rect 120377 275884 120423 275922
rect 112970 275876 114070 275882
rect 111524 275868 112624 275874
rect 111524 275834 111553 275868
rect 111587 275834 111625 275868
rect 111659 275834 111697 275868
rect 111731 275834 111769 275868
rect 111803 275834 111841 275868
rect 111875 275834 111913 275868
rect 111947 275834 111985 275868
rect 112019 275834 112057 275868
rect 112091 275834 112129 275868
rect 112163 275834 112201 275868
rect 112235 275834 112273 275868
rect 112307 275834 112345 275868
rect 112379 275834 112417 275868
rect 112451 275834 112489 275868
rect 112523 275834 112561 275868
rect 112595 275834 112624 275868
rect 112970 275842 112999 275876
rect 113033 275842 113071 275876
rect 113105 275842 113143 275876
rect 113177 275842 113215 275876
rect 113249 275842 113287 275876
rect 113321 275842 113359 275876
rect 113393 275842 113431 275876
rect 113465 275842 113503 275876
rect 113537 275842 113575 275876
rect 113609 275842 113647 275876
rect 113681 275842 113719 275876
rect 113753 275842 113791 275876
rect 113825 275842 113863 275876
rect 113897 275842 113935 275876
rect 113969 275842 114007 275876
rect 114041 275842 114070 275876
rect 116135 275876 117235 275882
rect 112970 275836 114070 275842
rect 114657 275851 114857 275857
rect 111524 275828 112624 275834
rect 111404 275795 111492 275818
rect 111404 275761 111452 275795
rect 111486 275761 111492 275795
rect 111404 275723 111492 275761
rect 111404 275689 111452 275723
rect 111486 275689 111492 275723
rect 111404 275666 111492 275689
rect 112656 275795 112744 275818
rect 112656 275761 112662 275795
rect 112696 275761 112744 275795
rect 112656 275750 112744 275761
rect 112850 275783 112938 275826
rect 112850 275750 112898 275783
rect 112656 275749 112898 275750
rect 112932 275749 112938 275783
rect 112656 275723 112938 275749
rect 112656 275689 112662 275723
rect 112696 275711 112938 275723
rect 112696 275689 112898 275711
rect 112656 275688 112898 275689
rect 112656 275666 112744 275688
rect 111404 275458 111446 275666
rect 111524 275650 112624 275656
rect 111524 275616 111553 275650
rect 111587 275616 111625 275650
rect 111659 275616 111697 275650
rect 111731 275616 111769 275650
rect 111803 275616 111841 275650
rect 111875 275616 111913 275650
rect 111947 275616 111985 275650
rect 112019 275616 112057 275650
rect 112091 275616 112129 275650
rect 112163 275616 112201 275650
rect 112235 275616 112273 275650
rect 112307 275616 112345 275650
rect 112379 275616 112417 275650
rect 112451 275616 112489 275650
rect 112523 275616 112561 275650
rect 112595 275616 112624 275650
rect 111524 275610 112624 275616
rect 112702 275634 112744 275666
rect 112850 275677 112898 275688
rect 112932 275677 112938 275711
rect 112850 275634 112938 275677
rect 114102 275783 114190 275826
rect 114657 275817 114704 275851
rect 114738 275817 114776 275851
rect 114810 275817 114857 275851
rect 114657 275811 114857 275817
rect 115348 275851 115548 275857
rect 115348 275817 115395 275851
rect 115429 275817 115467 275851
rect 115501 275817 115548 275851
rect 116135 275842 116164 275876
rect 116198 275842 116236 275876
rect 116270 275842 116308 275876
rect 116342 275842 116380 275876
rect 116414 275842 116452 275876
rect 116486 275842 116524 275876
rect 116558 275842 116596 275876
rect 116630 275842 116668 275876
rect 116702 275842 116740 275876
rect 116774 275842 116812 275876
rect 116846 275842 116884 275876
rect 116918 275842 116956 275876
rect 116990 275842 117028 275876
rect 117062 275842 117100 275876
rect 117134 275842 117172 275876
rect 117206 275842 117235 275876
rect 116135 275836 117235 275842
rect 117581 275868 118681 275874
rect 117581 275834 117610 275868
rect 117644 275834 117682 275868
rect 117716 275834 117754 275868
rect 117788 275834 117826 275868
rect 117860 275834 117898 275868
rect 117932 275834 117970 275868
rect 118004 275834 118042 275868
rect 118076 275834 118114 275868
rect 118148 275834 118186 275868
rect 118220 275834 118258 275868
rect 118292 275834 118330 275868
rect 118364 275834 118402 275868
rect 118436 275834 118474 275868
rect 118508 275834 118546 275868
rect 118580 275834 118618 275868
rect 118652 275834 118681 275868
rect 117581 275828 118681 275834
rect 120377 275850 120383 275884
rect 120417 275850 120423 275884
rect 120377 275833 120423 275850
rect 120835 276316 120881 276333
rect 120835 276282 120841 276316
rect 120875 276282 120881 276316
rect 120835 276244 120881 276282
rect 120835 276210 120841 276244
rect 120875 276210 120881 276244
rect 120835 276172 120881 276210
rect 120835 276138 120841 276172
rect 120875 276139 120881 276172
rect 121077 276316 121123 276333
rect 121077 276282 121083 276316
rect 121117 276282 121123 276316
rect 121077 276244 121123 276282
rect 121077 276210 121083 276244
rect 121117 276210 121123 276244
rect 121077 276172 121123 276210
rect 121077 276139 121083 276172
rect 120875 276138 121083 276139
rect 121117 276138 121123 276172
rect 120835 276103 121123 276138
rect 120835 276100 120969 276103
rect 120835 276066 120841 276100
rect 120875 276069 120969 276100
rect 121003 276100 121123 276103
rect 121003 276069 121083 276100
rect 120875 276066 121083 276069
rect 121117 276066 121123 276100
rect 120835 276032 121123 276066
rect 120835 276028 120881 276032
rect 120835 275994 120841 276028
rect 120875 275994 120881 276028
rect 120835 275956 120881 275994
rect 120835 275922 120841 275956
rect 120875 275922 120881 275956
rect 120835 275884 120881 275922
rect 120835 275850 120841 275884
rect 120875 275850 120881 275884
rect 120835 275833 120881 275850
rect 115348 275811 115548 275817
rect 114102 275749 114108 275783
rect 114142 275760 114190 275783
rect 114570 275766 114616 275801
rect 114570 275760 114576 275766
rect 114142 275749 114576 275760
rect 114102 275732 114576 275749
rect 114610 275732 114616 275766
rect 114102 275711 114616 275732
rect 114102 275677 114108 275711
rect 114142 275694 114616 275711
rect 114142 275677 114576 275694
rect 114102 275660 114576 275677
rect 114610 275660 114616 275694
rect 114102 275634 114616 275660
rect 111524 275508 112624 275514
rect 111524 275474 111553 275508
rect 111587 275474 111625 275508
rect 111659 275474 111697 275508
rect 111731 275474 111769 275508
rect 111803 275474 111841 275508
rect 111875 275474 111913 275508
rect 111947 275474 111985 275508
rect 112019 275474 112057 275508
rect 112091 275474 112129 275508
rect 112163 275474 112201 275508
rect 112235 275474 112273 275508
rect 112307 275474 112345 275508
rect 112379 275474 112417 275508
rect 112451 275474 112489 275508
rect 112523 275474 112561 275508
rect 112595 275474 112624 275508
rect 111524 275468 112624 275474
rect 112702 275458 112746 275634
rect 111404 275435 111492 275458
rect 111404 275401 111452 275435
rect 111486 275401 111492 275435
rect 111404 275363 111492 275401
rect 111404 275329 111452 275363
rect 111486 275329 111492 275363
rect 111404 275306 111492 275329
rect 112656 275435 112746 275458
rect 112656 275401 112662 275435
rect 112696 275414 112746 275435
rect 112850 275534 112892 275634
rect 114148 275627 114616 275634
rect 112970 275618 114070 275624
rect 112970 275584 112999 275618
rect 113033 275584 113071 275618
rect 113105 275584 113143 275618
rect 113177 275584 113215 275618
rect 113249 275584 113287 275618
rect 113321 275584 113359 275618
rect 113393 275584 113431 275618
rect 113465 275584 113503 275618
rect 113537 275584 113575 275618
rect 113609 275584 113647 275618
rect 113681 275584 113719 275618
rect 113753 275584 113791 275618
rect 113825 275584 113863 275618
rect 113897 275584 113935 275618
rect 113969 275584 114007 275618
rect 114041 275584 114070 275618
rect 112970 275578 114070 275584
rect 114148 275534 114190 275627
rect 112850 275496 114190 275534
rect 112696 275401 112744 275414
rect 112656 275366 112744 275401
rect 112850 275402 112892 275496
rect 112970 275452 114070 275458
rect 112970 275418 112999 275452
rect 113033 275418 113071 275452
rect 113105 275418 113143 275452
rect 113177 275418 113215 275452
rect 113249 275418 113287 275452
rect 113321 275418 113359 275452
rect 113393 275418 113431 275452
rect 113465 275418 113503 275452
rect 113537 275418 113575 275452
rect 113609 275418 113647 275452
rect 113681 275418 113719 275452
rect 113753 275418 113791 275452
rect 113825 275418 113863 275452
rect 113897 275418 113935 275452
rect 113969 275418 114007 275452
rect 114041 275418 114070 275452
rect 112970 275412 114070 275418
rect 114148 275402 114190 275496
rect 114570 275622 114616 275627
rect 114570 275588 114576 275622
rect 114610 275588 114616 275622
rect 114570 275550 114616 275588
rect 114570 275516 114576 275550
rect 114610 275516 114616 275550
rect 114570 275478 114616 275516
rect 114570 275444 114576 275478
rect 114610 275444 114616 275478
rect 114570 275409 114616 275444
rect 114898 275766 114944 275801
rect 114898 275732 114904 275766
rect 114938 275732 114944 275766
rect 114898 275694 114944 275732
rect 114898 275660 114904 275694
rect 114938 275660 114944 275694
rect 114898 275622 114944 275660
rect 114898 275588 114904 275622
rect 114938 275588 114944 275622
rect 114898 275550 114944 275588
rect 114898 275516 114904 275550
rect 114938 275516 114944 275550
rect 114898 275478 114944 275516
rect 114898 275444 114904 275478
rect 114938 275444 114944 275478
rect 114898 275409 114944 275444
rect 115261 275766 115307 275801
rect 115261 275732 115267 275766
rect 115301 275732 115307 275766
rect 115261 275694 115307 275732
rect 115261 275660 115267 275694
rect 115301 275660 115307 275694
rect 115261 275622 115307 275660
rect 115261 275588 115267 275622
rect 115301 275588 115307 275622
rect 115261 275550 115307 275588
rect 115261 275516 115267 275550
rect 115301 275516 115307 275550
rect 115261 275478 115307 275516
rect 115261 275444 115267 275478
rect 115301 275444 115307 275478
rect 115261 275409 115307 275444
rect 115589 275766 115635 275801
rect 115589 275732 115595 275766
rect 115629 275760 115635 275766
rect 116015 275783 116103 275826
rect 116015 275760 116063 275783
rect 115629 275749 116063 275760
rect 116097 275749 116103 275783
rect 115629 275732 116103 275749
rect 115589 275711 116103 275732
rect 115589 275694 116063 275711
rect 115589 275660 115595 275694
rect 115629 275677 116063 275694
rect 116097 275677 116103 275711
rect 115629 275660 116103 275677
rect 115589 275634 116103 275660
rect 117267 275783 117355 275826
rect 117267 275749 117273 275783
rect 117307 275750 117355 275783
rect 117461 275795 117549 275818
rect 117461 275761 117509 275795
rect 117543 275761 117549 275795
rect 117461 275750 117549 275761
rect 117307 275749 117549 275750
rect 117267 275723 117549 275749
rect 117267 275711 117509 275723
rect 117267 275677 117273 275711
rect 117307 275689 117509 275711
rect 117543 275689 117549 275723
rect 117307 275688 117549 275689
rect 117307 275677 117355 275688
rect 117267 275634 117355 275677
rect 117461 275666 117549 275688
rect 118713 275795 118801 275818
rect 118713 275761 118719 275795
rect 118753 275761 118801 275795
rect 118713 275723 118801 275761
rect 118713 275689 118719 275723
rect 118753 275689 118801 275723
rect 118713 275666 118801 275689
rect 117461 275634 117503 275666
rect 115589 275627 116057 275634
rect 115589 275622 115635 275627
rect 115589 275588 115595 275622
rect 115629 275588 115635 275622
rect 115589 275550 115635 275588
rect 115589 275516 115595 275550
rect 115629 275516 115635 275550
rect 115589 275478 115635 275516
rect 115589 275444 115595 275478
rect 115629 275444 115635 275478
rect 115589 275409 115635 275444
rect 116015 275534 116057 275627
rect 116135 275618 117235 275624
rect 116135 275584 116164 275618
rect 116198 275584 116236 275618
rect 116270 275584 116308 275618
rect 116342 275584 116380 275618
rect 116414 275584 116452 275618
rect 116486 275584 116524 275618
rect 116558 275584 116596 275618
rect 116630 275584 116668 275618
rect 116702 275584 116740 275618
rect 116774 275584 116812 275618
rect 116846 275584 116884 275618
rect 116918 275584 116956 275618
rect 116990 275584 117028 275618
rect 117062 275584 117100 275618
rect 117134 275584 117172 275618
rect 117206 275584 117235 275618
rect 116135 275578 117235 275584
rect 117313 275534 117355 275634
rect 116015 275496 117355 275534
rect 112850 275366 112938 275402
rect 112656 275363 112938 275366
rect 112656 275329 112662 275363
rect 112696 275359 112938 275363
rect 112696 275329 112898 275359
rect 112656 275325 112898 275329
rect 112932 275325 112938 275359
rect 112656 275306 112938 275325
rect 111404 275098 111446 275306
rect 112702 275304 112938 275306
rect 111524 275290 112624 275296
rect 111524 275256 111553 275290
rect 111587 275256 111625 275290
rect 111659 275256 111697 275290
rect 111731 275256 111769 275290
rect 111803 275256 111841 275290
rect 111875 275256 111913 275290
rect 111947 275256 111985 275290
rect 112019 275256 112057 275290
rect 112091 275256 112129 275290
rect 112163 275256 112201 275290
rect 112235 275256 112273 275290
rect 112307 275256 112345 275290
rect 112379 275256 112417 275290
rect 112451 275256 112489 275290
rect 112523 275256 112561 275290
rect 112595 275256 112624 275290
rect 111524 275250 112624 275256
rect 111524 275148 112624 275154
rect 111524 275114 111553 275148
rect 111587 275114 111625 275148
rect 111659 275114 111697 275148
rect 111731 275114 111769 275148
rect 111803 275114 111841 275148
rect 111875 275114 111913 275148
rect 111947 275114 111985 275148
rect 112019 275114 112057 275148
rect 112091 275114 112129 275148
rect 112163 275114 112201 275148
rect 112235 275114 112273 275148
rect 112307 275114 112345 275148
rect 112379 275114 112417 275148
rect 112451 275114 112489 275148
rect 112523 275114 112561 275148
rect 112595 275114 112624 275148
rect 111524 275108 112624 275114
rect 112702 275098 112744 275304
rect 112850 275287 112938 275304
rect 112850 275253 112898 275287
rect 112932 275253 112938 275287
rect 112850 275210 112938 275253
rect 114102 275359 114190 275402
rect 116015 275402 116057 275496
rect 116135 275452 117235 275458
rect 116135 275418 116164 275452
rect 116198 275418 116236 275452
rect 116270 275418 116308 275452
rect 116342 275418 116380 275452
rect 116414 275418 116452 275452
rect 116486 275418 116524 275452
rect 116558 275418 116596 275452
rect 116630 275418 116668 275452
rect 116702 275418 116740 275452
rect 116774 275418 116812 275452
rect 116846 275418 116884 275452
rect 116918 275418 116956 275452
rect 116990 275418 117028 275452
rect 117062 275418 117100 275452
rect 117134 275418 117172 275452
rect 117206 275418 117235 275452
rect 116135 275412 117235 275418
rect 117313 275402 117355 275496
rect 117459 275458 117503 275634
rect 117581 275650 118681 275656
rect 117581 275616 117610 275650
rect 117644 275616 117682 275650
rect 117716 275616 117754 275650
rect 117788 275616 117826 275650
rect 117860 275616 117898 275650
rect 117932 275616 117970 275650
rect 118004 275616 118042 275650
rect 118076 275616 118114 275650
rect 118148 275616 118186 275650
rect 118220 275616 118258 275650
rect 118292 275616 118330 275650
rect 118364 275616 118402 275650
rect 118436 275616 118474 275650
rect 118508 275616 118546 275650
rect 118580 275616 118618 275650
rect 118652 275616 118681 275650
rect 117581 275610 118681 275616
rect 117581 275508 118681 275514
rect 117581 275474 117610 275508
rect 117644 275474 117682 275508
rect 117716 275474 117754 275508
rect 117788 275474 117826 275508
rect 117860 275474 117898 275508
rect 117932 275474 117970 275508
rect 118004 275474 118042 275508
rect 118076 275474 118114 275508
rect 118148 275474 118186 275508
rect 118220 275474 118258 275508
rect 118292 275474 118330 275508
rect 118364 275474 118402 275508
rect 118436 275474 118474 275508
rect 118508 275474 118546 275508
rect 118580 275474 118618 275508
rect 118652 275474 118681 275508
rect 117581 275468 118681 275474
rect 118759 275458 118801 275666
rect 120433 275786 120825 275792
rect 120433 275752 120468 275786
rect 120502 275752 120540 275786
rect 120574 275752 120612 275786
rect 120646 275752 120684 275786
rect 120718 275752 120756 275786
rect 120790 275752 120825 275786
rect 120433 275630 120825 275752
rect 120433 275596 120468 275630
rect 120502 275596 120540 275630
rect 120574 275596 120612 275630
rect 120646 275596 120684 275630
rect 120718 275596 120756 275630
rect 120790 275596 120825 275630
rect 120433 275590 120825 275596
rect 117459 275435 117549 275458
rect 117459 275414 117509 275435
rect 114102 275325 114108 275359
rect 114142 275325 114190 275359
rect 114657 275393 114857 275399
rect 114657 275359 114704 275393
rect 114738 275359 114776 275393
rect 114810 275359 114857 275393
rect 114657 275353 114857 275359
rect 115348 275393 115548 275399
rect 115348 275359 115395 275393
rect 115429 275359 115467 275393
rect 115501 275359 115548 275393
rect 115348 275353 115548 275359
rect 116015 275359 116103 275402
rect 114102 275287 114190 275325
rect 114102 275253 114108 275287
rect 114142 275253 114190 275287
rect 114720 275285 114790 275353
rect 114102 275210 114190 275253
rect 114308 275201 114790 275285
rect 114865 275288 114970 275313
rect 114865 275236 114890 275288
rect 114942 275236 114970 275288
rect 114865 275206 114970 275236
rect 115235 275288 115340 275313
rect 115235 275236 115262 275288
rect 115314 275236 115340 275288
rect 115235 275206 115340 275236
rect 115415 275285 115485 275353
rect 116015 275325 116063 275359
rect 116097 275325 116103 275359
rect 116015 275287 116103 275325
rect 112970 275194 114070 275200
rect 112970 275160 112999 275194
rect 113033 275160 113071 275194
rect 113105 275160 113143 275194
rect 113177 275160 113215 275194
rect 113249 275160 113287 275194
rect 113321 275160 113359 275194
rect 113393 275160 113431 275194
rect 113465 275160 113503 275194
rect 113537 275160 113575 275194
rect 113609 275160 113647 275194
rect 113681 275160 113719 275194
rect 113753 275160 113791 275194
rect 113825 275160 113863 275194
rect 113897 275160 113935 275194
rect 113969 275160 114007 275194
rect 114041 275160 114070 275194
rect 112970 275154 114070 275160
rect 111404 275075 111492 275098
rect 111404 275041 111452 275075
rect 111486 275041 111492 275075
rect 111404 275003 111492 275041
rect 111404 274969 111452 275003
rect 111486 274969 111492 275003
rect 111404 274946 111492 274969
rect 112656 275075 112744 275098
rect 114308 275086 114343 275201
rect 114720 275171 114790 275201
rect 115415 275201 115897 275285
rect 116015 275253 116063 275287
rect 116097 275253 116103 275287
rect 116015 275210 116103 275253
rect 117267 275366 117355 275402
rect 117461 275401 117509 275414
rect 117543 275401 117549 275435
rect 117461 275366 117549 275401
rect 117267 275363 117549 275366
rect 117267 275359 117509 275363
rect 117267 275325 117273 275359
rect 117307 275329 117509 275359
rect 117543 275329 117549 275363
rect 117307 275325 117549 275329
rect 117267 275306 117549 275325
rect 118713 275435 118801 275458
rect 118713 275401 118719 275435
rect 118753 275401 118801 275435
rect 118713 275363 118801 275401
rect 118713 275329 118719 275363
rect 118753 275329 118801 275363
rect 118713 275306 118801 275329
rect 117267 275304 117503 275306
rect 117267 275287 117355 275304
rect 117267 275253 117273 275287
rect 117307 275253 117355 275287
rect 117267 275210 117355 275253
rect 115415 275171 115485 275201
rect 114657 275165 114857 275171
rect 114657 275131 114704 275165
rect 114738 275131 114776 275165
rect 114810 275131 114857 275165
rect 114657 275125 114857 275131
rect 115348 275165 115548 275171
rect 115348 275131 115395 275165
rect 115429 275131 115467 275165
rect 115501 275131 115548 275165
rect 115348 275125 115548 275131
rect 112656 275041 112662 275075
rect 112696 275041 112744 275075
rect 113843 275056 114343 275086
rect 112656 275003 112744 275041
rect 113000 275050 114343 275056
rect 113000 275016 113029 275050
rect 113063 275016 113101 275050
rect 113135 275016 113173 275050
rect 113207 275016 113245 275050
rect 113279 275016 113317 275050
rect 113351 275016 113389 275050
rect 113423 275016 113461 275050
rect 113495 275016 113533 275050
rect 113567 275016 113605 275050
rect 113639 275016 113677 275050
rect 113711 275016 113749 275050
rect 113783 275016 113821 275050
rect 113855 275016 113893 275050
rect 113927 275016 113965 275050
rect 113999 275016 114037 275050
rect 114071 275045 114343 275050
rect 114570 275092 114616 275115
rect 114570 275058 114576 275092
rect 114610 275058 114616 275092
rect 114071 275016 114100 275045
rect 113000 275010 114100 275016
rect 114570 275020 114616 275058
rect 112656 274969 112662 275003
rect 112696 274969 112744 275003
rect 112656 274946 112744 274969
rect 111404 274738 111446 274946
rect 111524 274930 112624 274936
rect 111524 274896 111553 274930
rect 111587 274896 111625 274930
rect 111659 274896 111697 274930
rect 111731 274896 111769 274930
rect 111803 274896 111841 274930
rect 111875 274896 111913 274930
rect 111947 274896 111985 274930
rect 112019 274896 112057 274930
rect 112091 274896 112129 274930
rect 112163 274896 112201 274930
rect 112235 274896 112273 274930
rect 112307 274896 112345 274930
rect 112379 274896 112417 274930
rect 112451 274896 112489 274930
rect 112523 274896 112561 274930
rect 112595 274896 112624 274930
rect 111524 274890 112624 274896
rect 111524 274788 112624 274794
rect 111524 274754 111553 274788
rect 111587 274754 111625 274788
rect 111659 274754 111697 274788
rect 111731 274754 111769 274788
rect 111803 274754 111841 274788
rect 111875 274754 111913 274788
rect 111947 274754 111985 274788
rect 112019 274754 112057 274788
rect 112091 274754 112129 274788
rect 112163 274754 112201 274788
rect 112235 274754 112273 274788
rect 112307 274754 112345 274788
rect 112379 274754 112417 274788
rect 112451 274754 112489 274788
rect 112523 274754 112561 274788
rect 112595 274754 112624 274788
rect 111524 274748 112624 274754
rect 112702 274738 112744 274946
rect 111404 274715 111492 274738
rect 111404 274681 111452 274715
rect 111486 274681 111492 274715
rect 111404 274643 111492 274681
rect 111404 274609 111452 274643
rect 111486 274609 111492 274643
rect 111404 274586 111492 274609
rect 112656 274715 112744 274738
rect 112656 274681 112662 274715
rect 112696 274681 112744 274715
rect 112656 274643 112744 274681
rect 112656 274609 112662 274643
rect 112696 274609 112744 274643
rect 112656 274586 112744 274609
rect 112874 274981 112968 275000
rect 112874 274947 112928 274981
rect 112962 274947 112968 274981
rect 112874 274928 112968 274947
rect 114132 274981 114226 275000
rect 114132 274947 114138 274981
rect 114172 274947 114226 274981
rect 114132 274928 114226 274947
rect 112874 274836 112922 274928
rect 113000 274912 114100 274918
rect 113000 274878 113029 274912
rect 113063 274878 113101 274912
rect 113135 274878 113173 274912
rect 113207 274878 113245 274912
rect 113279 274878 113317 274912
rect 113351 274878 113389 274912
rect 113423 274878 113461 274912
rect 113495 274878 113533 274912
rect 113567 274878 113605 274912
rect 113639 274878 113677 274912
rect 113711 274878 113749 274912
rect 113783 274878 113821 274912
rect 113855 274878 113893 274912
rect 113927 274878 113965 274912
rect 113999 274878 114037 274912
rect 114071 274878 114100 274912
rect 113000 274872 114100 274878
rect 114178 274836 114226 274928
rect 112874 274792 114226 274836
rect 114324 274953 114396 274994
rect 114570 274986 114576 275020
rect 114610 274986 114616 275020
rect 114570 274963 114616 274986
rect 114898 275092 114944 275115
rect 114898 275058 114904 275092
rect 114938 275058 114944 275092
rect 114898 275020 114944 275058
rect 114898 274986 114904 275020
rect 114938 274986 114944 275020
rect 114898 274963 114944 274986
rect 115261 275092 115307 275115
rect 115261 275058 115267 275092
rect 115301 275058 115307 275092
rect 115261 275020 115307 275058
rect 115261 274986 115267 275020
rect 115301 274986 115307 275020
rect 115261 274963 115307 274986
rect 115589 275092 115635 275115
rect 115589 275058 115595 275092
rect 115629 275058 115635 275092
rect 115589 275020 115635 275058
rect 115862 275086 115897 275201
rect 116135 275194 117235 275200
rect 116135 275160 116164 275194
rect 116198 275160 116236 275194
rect 116270 275160 116308 275194
rect 116342 275160 116380 275194
rect 116414 275160 116452 275194
rect 116486 275160 116524 275194
rect 116558 275160 116596 275194
rect 116630 275160 116668 275194
rect 116702 275160 116740 275194
rect 116774 275160 116812 275194
rect 116846 275160 116884 275194
rect 116918 275160 116956 275194
rect 116990 275160 117028 275194
rect 117062 275160 117100 275194
rect 117134 275160 117172 275194
rect 117206 275160 117235 275194
rect 116135 275154 117235 275160
rect 117461 275098 117503 275304
rect 117581 275290 118681 275296
rect 117581 275256 117610 275290
rect 117644 275256 117682 275290
rect 117716 275256 117754 275290
rect 117788 275256 117826 275290
rect 117860 275256 117898 275290
rect 117932 275256 117970 275290
rect 118004 275256 118042 275290
rect 118076 275256 118114 275290
rect 118148 275256 118186 275290
rect 118220 275256 118258 275290
rect 118292 275256 118330 275290
rect 118364 275256 118402 275290
rect 118436 275256 118474 275290
rect 118508 275256 118546 275290
rect 118580 275256 118618 275290
rect 118652 275256 118681 275290
rect 117581 275250 118681 275256
rect 117581 275148 118681 275154
rect 117581 275114 117610 275148
rect 117644 275114 117682 275148
rect 117716 275114 117754 275148
rect 117788 275114 117826 275148
rect 117860 275114 117898 275148
rect 117932 275114 117970 275148
rect 118004 275114 118042 275148
rect 118076 275114 118114 275148
rect 118148 275114 118186 275148
rect 118220 275114 118258 275148
rect 118292 275114 118330 275148
rect 118364 275114 118402 275148
rect 118436 275114 118474 275148
rect 118508 275114 118546 275148
rect 118580 275114 118618 275148
rect 118652 275114 118681 275148
rect 117581 275108 118681 275114
rect 118759 275098 118801 275306
rect 115862 275056 116362 275086
rect 117461 275075 117549 275098
rect 115862 275050 117205 275056
rect 115862 275045 116134 275050
rect 115589 274986 115595 275020
rect 115629 274986 115635 275020
rect 116105 275016 116134 275045
rect 116168 275016 116206 275050
rect 116240 275016 116278 275050
rect 116312 275016 116350 275050
rect 116384 275016 116422 275050
rect 116456 275016 116494 275050
rect 116528 275016 116566 275050
rect 116600 275016 116638 275050
rect 116672 275016 116710 275050
rect 116744 275016 116782 275050
rect 116816 275016 116854 275050
rect 116888 275016 116926 275050
rect 116960 275016 116998 275050
rect 117032 275016 117070 275050
rect 117104 275016 117142 275050
rect 117176 275016 117205 275050
rect 116105 275010 117205 275016
rect 117461 275041 117509 275075
rect 117543 275041 117549 275075
rect 117461 275003 117549 275041
rect 115589 274963 115635 274986
rect 115809 274953 115881 274994
rect 114324 274919 114342 274953
rect 114376 274919 114396 274953
rect 114324 274863 114396 274919
rect 114657 274947 114857 274953
rect 114657 274913 114704 274947
rect 114738 274913 114776 274947
rect 114810 274913 114857 274947
rect 114657 274907 114857 274913
rect 115348 274947 115548 274953
rect 115348 274913 115395 274947
rect 115429 274913 115467 274947
rect 115501 274913 115548 274947
rect 115348 274907 115548 274913
rect 115809 274919 115828 274953
rect 115862 274919 115881 274953
rect 114843 274863 115030 274878
rect 114324 274818 114781 274863
rect 112874 274702 112922 274792
rect 113000 274752 114100 274758
rect 113000 274718 113029 274752
rect 113063 274718 113101 274752
rect 113135 274718 113173 274752
rect 113207 274718 113245 274752
rect 113279 274718 113317 274752
rect 113351 274718 113389 274752
rect 113423 274718 113461 274752
rect 113495 274718 113533 274752
rect 113567 274718 113605 274752
rect 113639 274718 113677 274752
rect 113711 274718 113749 274752
rect 113783 274718 113821 274752
rect 113855 274718 113893 274752
rect 113927 274718 113965 274752
rect 113999 274718 114037 274752
rect 114071 274718 114100 274752
rect 113000 274712 114100 274718
rect 114178 274702 114226 274792
rect 114737 274763 114781 274818
rect 114843 274811 114891 274863
rect 114943 274811 115030 274863
rect 114843 274793 115030 274811
rect 115175 274863 115362 274878
rect 115809 274863 115881 274919
rect 115175 274811 115262 274863
rect 115314 274811 115362 274863
rect 115175 274793 115362 274811
rect 115424 274818 115881 274863
rect 115979 274981 116073 275000
rect 115979 274947 116033 274981
rect 116067 274947 116073 274981
rect 115979 274928 116073 274947
rect 117237 274981 117331 275000
rect 117237 274947 117243 274981
rect 117277 274947 117331 274981
rect 117237 274928 117331 274947
rect 115979 274836 116027 274928
rect 116105 274912 117205 274918
rect 116105 274878 116134 274912
rect 116168 274878 116206 274912
rect 116240 274878 116278 274912
rect 116312 274878 116350 274912
rect 116384 274878 116422 274912
rect 116456 274878 116494 274912
rect 116528 274878 116566 274912
rect 116600 274878 116638 274912
rect 116672 274878 116710 274912
rect 116744 274878 116782 274912
rect 116816 274878 116854 274912
rect 116888 274878 116926 274912
rect 116960 274878 116998 274912
rect 117032 274878 117070 274912
rect 117104 274878 117142 274912
rect 117176 274878 117205 274912
rect 116105 274872 117205 274878
rect 117283 274836 117331 274928
rect 115424 274763 115468 274818
rect 115979 274792 117331 274836
rect 114657 274757 114857 274763
rect 114657 274723 114704 274757
rect 114738 274723 114776 274757
rect 114810 274723 114857 274757
rect 114657 274717 114857 274723
rect 115348 274757 115548 274763
rect 115348 274723 115395 274757
rect 115429 274723 115467 274757
rect 115501 274723 115548 274757
rect 115348 274717 115548 274723
rect 112874 274683 112968 274702
rect 112874 274649 112928 274683
rect 112962 274649 112968 274683
rect 112874 274630 112968 274649
rect 114132 274683 114226 274702
rect 114132 274649 114138 274683
rect 114172 274649 114226 274683
rect 114132 274630 114226 274649
rect 114570 274684 114616 274707
rect 114570 274650 114576 274684
rect 114610 274650 114616 274684
rect 111524 274570 112624 274576
rect 111524 274536 111553 274570
rect 111587 274536 111625 274570
rect 111659 274536 111697 274570
rect 111731 274536 111769 274570
rect 111803 274536 111841 274570
rect 111875 274536 111913 274570
rect 111947 274536 111985 274570
rect 112019 274536 112057 274570
rect 112091 274536 112129 274570
rect 112163 274536 112201 274570
rect 112235 274536 112273 274570
rect 112307 274536 112345 274570
rect 112379 274536 112417 274570
rect 112451 274536 112489 274570
rect 112523 274536 112561 274570
rect 112595 274536 112624 274570
rect 111524 274532 112624 274536
rect 112874 274536 112922 274630
rect 114327 274625 114395 274626
rect 114570 274625 114616 274650
rect 113000 274614 114100 274620
rect 113000 274580 113029 274614
rect 113063 274580 113101 274614
rect 113135 274580 113173 274614
rect 113207 274580 113245 274614
rect 113279 274580 113317 274614
rect 113351 274580 113389 274614
rect 113423 274580 113461 274614
rect 113495 274580 113533 274614
rect 113567 274580 113605 274614
rect 113639 274580 113677 274614
rect 113711 274580 113749 274614
rect 113783 274580 113821 274614
rect 113855 274580 113893 274614
rect 113927 274580 113965 274614
rect 113999 274580 114037 274614
rect 114071 274580 114100 274614
rect 113000 274574 114100 274580
rect 114327 274612 114616 274625
rect 114327 274578 114576 274612
rect 114610 274578 114616 274612
rect 114327 274565 114616 274578
rect 114327 274536 114395 274565
rect 114570 274555 114616 274565
rect 114898 274684 114944 274707
rect 114898 274650 114904 274684
rect 114938 274650 114944 274684
rect 114898 274612 114944 274650
rect 114898 274578 114904 274612
rect 114938 274578 114944 274612
rect 114898 274555 114944 274578
rect 115261 274684 115307 274707
rect 115261 274650 115267 274684
rect 115301 274650 115307 274684
rect 115261 274612 115307 274650
rect 115261 274578 115267 274612
rect 115301 274578 115307 274612
rect 115261 274555 115307 274578
rect 115589 274684 115635 274707
rect 115589 274650 115595 274684
rect 115629 274650 115635 274684
rect 115589 274625 115635 274650
rect 115979 274702 116027 274792
rect 116105 274752 117205 274758
rect 116105 274718 116134 274752
rect 116168 274718 116206 274752
rect 116240 274718 116278 274752
rect 116312 274718 116350 274752
rect 116384 274718 116422 274752
rect 116456 274718 116494 274752
rect 116528 274718 116566 274752
rect 116600 274718 116638 274752
rect 116672 274718 116710 274752
rect 116744 274718 116782 274752
rect 116816 274718 116854 274752
rect 116888 274718 116926 274752
rect 116960 274718 116998 274752
rect 117032 274718 117070 274752
rect 117104 274718 117142 274752
rect 117176 274718 117205 274752
rect 116105 274712 117205 274718
rect 117283 274702 117331 274792
rect 115979 274683 116073 274702
rect 115979 274649 116033 274683
rect 116067 274649 116073 274683
rect 115979 274630 116073 274649
rect 117237 274683 117331 274702
rect 117237 274649 117243 274683
rect 117277 274649 117331 274683
rect 117237 274630 117331 274649
rect 115810 274625 115878 274626
rect 115589 274612 115878 274625
rect 115589 274578 115595 274612
rect 115629 274578 115878 274612
rect 115589 274565 115878 274578
rect 116105 274614 117205 274620
rect 116105 274580 116134 274614
rect 116168 274580 116206 274614
rect 116240 274580 116278 274614
rect 116312 274580 116350 274614
rect 116384 274580 116422 274614
rect 116456 274580 116494 274614
rect 116528 274580 116566 274614
rect 116600 274580 116638 274614
rect 116672 274580 116710 274614
rect 116744 274580 116782 274614
rect 116816 274580 116854 274614
rect 116888 274580 116926 274614
rect 116960 274580 116998 274614
rect 117032 274580 117070 274614
rect 117104 274580 117142 274614
rect 117176 274580 117205 274614
rect 116105 274574 117205 274580
rect 115589 274555 115635 274565
rect 112874 274532 114395 274536
rect 111524 274530 114395 274532
rect 108355 274505 111012 274509
rect 106072 274503 111014 274505
rect 102557 274043 105283 274145
rect 102557 273799 102638 274043
rect 105186 273799 105283 274043
rect 106053 274267 111014 274503
rect 112044 274496 114395 274530
rect 114657 274539 114857 274545
rect 114657 274505 114704 274539
rect 114738 274505 114776 274539
rect 114810 274505 114857 274539
rect 114657 274499 114857 274505
rect 115348 274539 115548 274545
rect 115348 274505 115395 274539
rect 115429 274505 115467 274539
rect 115501 274505 115548 274539
rect 115348 274499 115548 274505
rect 115810 274536 115878 274565
rect 117283 274536 117331 274630
rect 117461 274969 117509 275003
rect 117543 274969 117549 275003
rect 117461 274946 117549 274969
rect 118713 275075 118801 275098
rect 118713 275041 118719 275075
rect 118753 275041 118801 275075
rect 120377 275532 120423 275549
rect 120377 275498 120383 275532
rect 120417 275498 120423 275532
rect 120377 275460 120423 275498
rect 120377 275426 120383 275460
rect 120417 275426 120423 275460
rect 120377 275388 120423 275426
rect 120377 275354 120383 275388
rect 120417 275354 120423 275388
rect 120377 275316 120423 275354
rect 120377 275282 120383 275316
rect 120417 275282 120423 275316
rect 120377 275244 120423 275282
rect 120377 275210 120383 275244
rect 120417 275210 120423 275244
rect 120377 275172 120423 275210
rect 120377 275138 120383 275172
rect 120417 275138 120423 275172
rect 120377 275100 120423 275138
rect 120377 275066 120383 275100
rect 120417 275066 120423 275100
rect 120377 275049 120423 275066
rect 120835 275532 120881 275549
rect 120835 275498 120841 275532
rect 120875 275498 120881 275532
rect 120835 275460 120881 275498
rect 120835 275426 120841 275460
rect 120875 275426 120881 275460
rect 120835 275388 120881 275426
rect 120835 275354 120841 275388
rect 120875 275354 120881 275388
rect 120835 275316 120881 275354
rect 120835 275282 120841 275316
rect 120875 275282 120881 275316
rect 120835 275244 120881 275282
rect 120835 275210 120841 275244
rect 120875 275210 120881 275244
rect 120835 275172 120881 275210
rect 120835 275138 120841 275172
rect 120875 275138 120881 275172
rect 120835 275100 120881 275138
rect 120835 275066 120841 275100
rect 120875 275066 120881 275100
rect 120835 275049 120881 275066
rect 118713 275003 118801 275041
rect 118713 274969 118719 275003
rect 118753 274969 118801 275003
rect 118713 274946 118801 274969
rect 117461 274738 117503 274946
rect 117581 274930 118681 274936
rect 117581 274896 117610 274930
rect 117644 274896 117682 274930
rect 117716 274896 117754 274930
rect 117788 274896 117826 274930
rect 117860 274896 117898 274930
rect 117932 274896 117970 274930
rect 118004 274896 118042 274930
rect 118076 274896 118114 274930
rect 118148 274896 118186 274930
rect 118220 274896 118258 274930
rect 118292 274896 118330 274930
rect 118364 274896 118402 274930
rect 118436 274896 118474 274930
rect 118508 274896 118546 274930
rect 118580 274896 118618 274930
rect 118652 274896 118681 274930
rect 117581 274890 118681 274896
rect 117581 274788 118681 274794
rect 117581 274754 117610 274788
rect 117644 274754 117682 274788
rect 117716 274754 117754 274788
rect 117788 274754 117826 274788
rect 117860 274754 117898 274788
rect 117932 274754 117970 274788
rect 118004 274754 118042 274788
rect 118076 274754 118114 274788
rect 118148 274754 118186 274788
rect 118220 274754 118258 274788
rect 118292 274754 118330 274788
rect 118364 274754 118402 274788
rect 118436 274754 118474 274788
rect 118508 274754 118546 274788
rect 118580 274754 118618 274788
rect 118652 274754 118681 274788
rect 117581 274748 118681 274754
rect 118759 274738 118801 274946
rect 120433 275002 120825 275008
rect 120433 274968 120468 275002
rect 120502 274968 120540 275002
rect 120574 274968 120612 275002
rect 120646 274968 120684 275002
rect 120718 274968 120756 275002
rect 120790 274968 120825 275002
rect 120433 274846 120825 274968
rect 120433 274812 120468 274846
rect 120502 274812 120540 274846
rect 120574 274812 120612 274846
rect 120646 274812 120684 274846
rect 120718 274812 120756 274846
rect 120790 274812 120825 274846
rect 120433 274806 120825 274812
rect 117461 274715 117549 274738
rect 117461 274681 117509 274715
rect 117543 274681 117549 274715
rect 117461 274643 117549 274681
rect 117461 274609 117509 274643
rect 117543 274609 117549 274643
rect 117461 274586 117549 274609
rect 118713 274715 118801 274738
rect 118713 274681 118719 274715
rect 118753 274681 118801 274715
rect 118713 274643 118801 274681
rect 118713 274609 118719 274643
rect 118753 274609 118801 274643
rect 118713 274586 118801 274609
rect 120377 274748 120423 274765
rect 120377 274714 120383 274748
rect 120417 274714 120423 274748
rect 120377 274676 120423 274714
rect 120377 274642 120383 274676
rect 120417 274642 120423 274676
rect 120377 274604 120423 274642
rect 115810 274532 117331 274536
rect 117581 274570 118681 274576
rect 117581 274536 117610 274570
rect 117644 274536 117682 274570
rect 117716 274536 117754 274570
rect 117788 274536 117826 274570
rect 117860 274536 117898 274570
rect 117932 274536 117970 274570
rect 118004 274536 118042 274570
rect 118076 274536 118114 274570
rect 118148 274536 118186 274570
rect 118220 274536 118258 274570
rect 118292 274536 118330 274570
rect 118364 274536 118402 274570
rect 118436 274536 118474 274570
rect 118508 274536 118546 274570
rect 118580 274536 118618 274570
rect 118652 274536 118681 274570
rect 117581 274532 118681 274536
rect 115810 274530 118681 274532
rect 120377 274570 120383 274604
rect 120417 274570 120423 274604
rect 120377 274532 120423 274570
rect 112719 274454 112924 274496
rect 113982 274422 114266 274432
rect 114724 274422 114783 274499
rect 113982 274401 114783 274422
rect 113982 274367 114034 274401
rect 114068 274367 114106 274401
rect 114140 274367 114178 274401
rect 114212 274367 114783 274401
rect 113982 274333 114783 274367
rect 115422 274422 115481 274499
rect 115810 274496 118161 274530
rect 120377 274498 120383 274532
rect 120417 274498 120423 274532
rect 117281 274454 117486 274496
rect 120377 274460 120423 274498
rect 115939 274422 116223 274432
rect 115422 274401 116223 274422
rect 115422 274367 115992 274401
rect 116026 274367 116064 274401
rect 116098 274367 116136 274401
rect 116170 274367 116223 274401
rect 115422 274333 116223 274367
rect 113982 274332 114266 274333
rect 115939 274332 116223 274333
rect 120377 274426 120383 274460
rect 120417 274426 120423 274460
rect 120377 274388 120423 274426
rect 120377 274354 120383 274388
rect 120417 274354 120423 274388
rect 120377 274316 120423 274354
rect 120377 274282 120383 274316
rect 120417 274282 120423 274316
rect 106053 273841 111015 274267
rect 120377 274265 120423 274282
rect 120835 274748 120881 274765
rect 120835 274714 120841 274748
rect 120875 274714 120881 274748
rect 120835 274676 120881 274714
rect 120835 274642 120841 274676
rect 120875 274642 120881 274676
rect 120835 274604 120881 274642
rect 120835 274570 120841 274604
rect 120875 274570 120881 274604
rect 120835 274532 120881 274570
rect 120835 274498 120841 274532
rect 120875 274498 120881 274532
rect 120835 274460 120881 274498
rect 120835 274426 120841 274460
rect 120875 274426 120881 274460
rect 120835 274388 120881 274426
rect 120835 274354 120841 274388
rect 120875 274354 120881 274388
rect 120835 274316 120881 274354
rect 120835 274282 120841 274316
rect 120875 274282 120881 274316
rect 120835 274265 120881 274282
rect 120433 274218 120825 274224
rect 112970 274210 114070 274216
rect 111524 274202 112624 274208
rect 111524 274168 111553 274202
rect 111587 274168 111625 274202
rect 111659 274168 111697 274202
rect 111731 274168 111769 274202
rect 111803 274168 111841 274202
rect 111875 274168 111913 274202
rect 111947 274168 111985 274202
rect 112019 274168 112057 274202
rect 112091 274168 112129 274202
rect 112163 274168 112201 274202
rect 112235 274168 112273 274202
rect 112307 274168 112345 274202
rect 112379 274168 112417 274202
rect 112451 274168 112489 274202
rect 112523 274168 112561 274202
rect 112595 274168 112624 274202
rect 112970 274176 112999 274210
rect 113033 274176 113071 274210
rect 113105 274176 113143 274210
rect 113177 274176 113215 274210
rect 113249 274176 113287 274210
rect 113321 274176 113359 274210
rect 113393 274176 113431 274210
rect 113465 274176 113503 274210
rect 113537 274176 113575 274210
rect 113609 274176 113647 274210
rect 113681 274176 113719 274210
rect 113753 274176 113791 274210
rect 113825 274176 113863 274210
rect 113897 274176 113935 274210
rect 113969 274176 114007 274210
rect 114041 274176 114070 274210
rect 116135 274210 117235 274216
rect 112970 274170 114070 274176
rect 114657 274185 114857 274191
rect 111524 274162 112624 274168
rect 111404 274129 111492 274152
rect 111404 274095 111452 274129
rect 111486 274095 111492 274129
rect 111404 274057 111492 274095
rect 111404 274023 111452 274057
rect 111486 274023 111492 274057
rect 111404 274000 111492 274023
rect 112656 274129 112744 274152
rect 112656 274095 112662 274129
rect 112696 274095 112744 274129
rect 112656 274084 112744 274095
rect 112850 274117 112938 274160
rect 112850 274084 112898 274117
rect 112656 274083 112898 274084
rect 112932 274083 112938 274117
rect 112656 274057 112938 274083
rect 112656 274023 112662 274057
rect 112696 274045 112938 274057
rect 112696 274023 112898 274045
rect 112656 274022 112898 274023
rect 112656 274000 112744 274022
rect 102557 273716 105283 273799
rect 108199 273428 108478 273841
rect 105964 273149 108478 273428
rect 111404 273792 111446 274000
rect 111524 273984 112624 273990
rect 111524 273950 111553 273984
rect 111587 273950 111625 273984
rect 111659 273950 111697 273984
rect 111731 273950 111769 273984
rect 111803 273950 111841 273984
rect 111875 273950 111913 273984
rect 111947 273950 111985 273984
rect 112019 273950 112057 273984
rect 112091 273950 112129 273984
rect 112163 273950 112201 273984
rect 112235 273950 112273 273984
rect 112307 273950 112345 273984
rect 112379 273950 112417 273984
rect 112451 273950 112489 273984
rect 112523 273950 112561 273984
rect 112595 273950 112624 273984
rect 111524 273944 112624 273950
rect 112702 273968 112744 274000
rect 112850 274011 112898 274022
rect 112932 274011 112938 274045
rect 112850 273968 112938 274011
rect 114102 274117 114190 274160
rect 114657 274151 114704 274185
rect 114738 274151 114776 274185
rect 114810 274151 114857 274185
rect 114657 274145 114857 274151
rect 115348 274185 115548 274191
rect 115348 274151 115395 274185
rect 115429 274151 115467 274185
rect 115501 274151 115548 274185
rect 116135 274176 116164 274210
rect 116198 274176 116236 274210
rect 116270 274176 116308 274210
rect 116342 274176 116380 274210
rect 116414 274176 116452 274210
rect 116486 274176 116524 274210
rect 116558 274176 116596 274210
rect 116630 274176 116668 274210
rect 116702 274176 116740 274210
rect 116774 274176 116812 274210
rect 116846 274176 116884 274210
rect 116918 274176 116956 274210
rect 116990 274176 117028 274210
rect 117062 274176 117100 274210
rect 117134 274176 117172 274210
rect 117206 274176 117235 274210
rect 116135 274170 117235 274176
rect 117581 274202 118681 274208
rect 117581 274168 117610 274202
rect 117644 274168 117682 274202
rect 117716 274168 117754 274202
rect 117788 274168 117826 274202
rect 117860 274168 117898 274202
rect 117932 274168 117970 274202
rect 118004 274168 118042 274202
rect 118076 274168 118114 274202
rect 118148 274168 118186 274202
rect 118220 274168 118258 274202
rect 118292 274168 118330 274202
rect 118364 274168 118402 274202
rect 118436 274168 118474 274202
rect 118508 274168 118546 274202
rect 118580 274168 118618 274202
rect 118652 274168 118681 274202
rect 117581 274162 118681 274168
rect 120433 274184 120468 274218
rect 120502 274184 120540 274218
rect 120574 274184 120612 274218
rect 120646 274184 120684 274218
rect 120718 274184 120756 274218
rect 120790 274184 120825 274218
rect 115348 274145 115548 274151
rect 114102 274083 114108 274117
rect 114142 274094 114190 274117
rect 114570 274100 114616 274135
rect 114570 274094 114576 274100
rect 114142 274083 114576 274094
rect 114102 274066 114576 274083
rect 114610 274066 114616 274100
rect 114102 274045 114616 274066
rect 114102 274011 114108 274045
rect 114142 274028 114616 274045
rect 114142 274011 114576 274028
rect 114102 273994 114576 274011
rect 114610 273994 114616 274028
rect 114102 273968 114616 273994
rect 111524 273842 112624 273848
rect 111524 273808 111553 273842
rect 111587 273808 111625 273842
rect 111659 273808 111697 273842
rect 111731 273808 111769 273842
rect 111803 273808 111841 273842
rect 111875 273808 111913 273842
rect 111947 273808 111985 273842
rect 112019 273808 112057 273842
rect 112091 273808 112129 273842
rect 112163 273808 112201 273842
rect 112235 273808 112273 273842
rect 112307 273808 112345 273842
rect 112379 273808 112417 273842
rect 112451 273808 112489 273842
rect 112523 273808 112561 273842
rect 112595 273808 112624 273842
rect 111524 273802 112624 273808
rect 112702 273792 112746 273968
rect 111404 273769 111492 273792
rect 111404 273735 111452 273769
rect 111486 273735 111492 273769
rect 111404 273697 111492 273735
rect 111404 273663 111452 273697
rect 111486 273663 111492 273697
rect 111404 273640 111492 273663
rect 112656 273769 112746 273792
rect 112656 273735 112662 273769
rect 112696 273748 112746 273769
rect 112850 273868 112892 273968
rect 114148 273961 114616 273968
rect 112970 273952 114070 273958
rect 112970 273918 112999 273952
rect 113033 273918 113071 273952
rect 113105 273918 113143 273952
rect 113177 273918 113215 273952
rect 113249 273918 113287 273952
rect 113321 273918 113359 273952
rect 113393 273918 113431 273952
rect 113465 273918 113503 273952
rect 113537 273918 113575 273952
rect 113609 273918 113647 273952
rect 113681 273918 113719 273952
rect 113753 273918 113791 273952
rect 113825 273918 113863 273952
rect 113897 273918 113935 273952
rect 113969 273918 114007 273952
rect 114041 273918 114070 273952
rect 112970 273912 114070 273918
rect 114148 273868 114190 273961
rect 112850 273830 114190 273868
rect 112696 273735 112744 273748
rect 112656 273700 112744 273735
rect 112850 273736 112892 273830
rect 112970 273786 114070 273792
rect 112970 273752 112999 273786
rect 113033 273752 113071 273786
rect 113105 273752 113143 273786
rect 113177 273752 113215 273786
rect 113249 273752 113287 273786
rect 113321 273752 113359 273786
rect 113393 273752 113431 273786
rect 113465 273752 113503 273786
rect 113537 273752 113575 273786
rect 113609 273752 113647 273786
rect 113681 273752 113719 273786
rect 113753 273752 113791 273786
rect 113825 273752 113863 273786
rect 113897 273752 113935 273786
rect 113969 273752 114007 273786
rect 114041 273752 114070 273786
rect 112970 273746 114070 273752
rect 114148 273736 114190 273830
rect 114570 273956 114616 273961
rect 114570 273922 114576 273956
rect 114610 273922 114616 273956
rect 114570 273884 114616 273922
rect 114570 273850 114576 273884
rect 114610 273850 114616 273884
rect 114570 273812 114616 273850
rect 114570 273778 114576 273812
rect 114610 273778 114616 273812
rect 114570 273743 114616 273778
rect 114898 274100 114944 274135
rect 114898 274066 114904 274100
rect 114938 274066 114944 274100
rect 114898 274028 114944 274066
rect 114898 273994 114904 274028
rect 114938 273994 114944 274028
rect 114898 273956 114944 273994
rect 114898 273922 114904 273956
rect 114938 273922 114944 273956
rect 114898 273884 114944 273922
rect 114898 273850 114904 273884
rect 114938 273850 114944 273884
rect 114898 273812 114944 273850
rect 114898 273778 114904 273812
rect 114938 273778 114944 273812
rect 114898 273743 114944 273778
rect 115261 274100 115307 274135
rect 115261 274066 115267 274100
rect 115301 274066 115307 274100
rect 115261 274028 115307 274066
rect 115261 273994 115267 274028
rect 115301 273994 115307 274028
rect 115261 273956 115307 273994
rect 115261 273922 115267 273956
rect 115301 273922 115307 273956
rect 115261 273884 115307 273922
rect 115261 273850 115267 273884
rect 115301 273850 115307 273884
rect 115261 273812 115307 273850
rect 115261 273778 115267 273812
rect 115301 273778 115307 273812
rect 115261 273743 115307 273778
rect 115589 274100 115635 274135
rect 115589 274066 115595 274100
rect 115629 274094 115635 274100
rect 116015 274117 116103 274160
rect 116015 274094 116063 274117
rect 115629 274083 116063 274094
rect 116097 274083 116103 274117
rect 115629 274066 116103 274083
rect 115589 274045 116103 274066
rect 115589 274028 116063 274045
rect 115589 273994 115595 274028
rect 115629 274011 116063 274028
rect 116097 274011 116103 274045
rect 115629 273994 116103 274011
rect 115589 273968 116103 273994
rect 117267 274117 117355 274160
rect 117267 274083 117273 274117
rect 117307 274084 117355 274117
rect 117461 274129 117549 274152
rect 117461 274095 117509 274129
rect 117543 274095 117549 274129
rect 117461 274084 117549 274095
rect 117307 274083 117549 274084
rect 117267 274057 117549 274083
rect 117267 274045 117509 274057
rect 117267 274011 117273 274045
rect 117307 274023 117509 274045
rect 117543 274023 117549 274057
rect 117307 274022 117549 274023
rect 117307 274011 117355 274022
rect 117267 273968 117355 274011
rect 117461 274000 117549 274022
rect 118713 274129 118801 274152
rect 118713 274095 118719 274129
rect 118753 274095 118801 274129
rect 118713 274057 118801 274095
rect 118713 274023 118719 274057
rect 118753 274023 118801 274057
rect 118713 274000 118801 274023
rect 120433 274062 120825 274184
rect 120433 274028 120468 274062
rect 120502 274028 120540 274062
rect 120574 274028 120612 274062
rect 120646 274028 120684 274062
rect 120718 274028 120756 274062
rect 120790 274028 120825 274062
rect 120433 274022 120825 274028
rect 117461 273968 117503 274000
rect 115589 273961 116057 273968
rect 115589 273956 115635 273961
rect 115589 273922 115595 273956
rect 115629 273922 115635 273956
rect 115589 273884 115635 273922
rect 115589 273850 115595 273884
rect 115629 273850 115635 273884
rect 115589 273812 115635 273850
rect 115589 273778 115595 273812
rect 115629 273778 115635 273812
rect 115589 273743 115635 273778
rect 116015 273868 116057 273961
rect 116135 273952 117235 273958
rect 116135 273918 116164 273952
rect 116198 273918 116236 273952
rect 116270 273918 116308 273952
rect 116342 273918 116380 273952
rect 116414 273918 116452 273952
rect 116486 273918 116524 273952
rect 116558 273918 116596 273952
rect 116630 273918 116668 273952
rect 116702 273918 116740 273952
rect 116774 273918 116812 273952
rect 116846 273918 116884 273952
rect 116918 273918 116956 273952
rect 116990 273918 117028 273952
rect 117062 273918 117100 273952
rect 117134 273918 117172 273952
rect 117206 273918 117235 273952
rect 116135 273912 117235 273918
rect 117313 273868 117355 273968
rect 116015 273830 117355 273868
rect 112850 273700 112938 273736
rect 112656 273697 112938 273700
rect 112656 273663 112662 273697
rect 112696 273693 112938 273697
rect 112696 273663 112898 273693
rect 112656 273659 112898 273663
rect 112932 273659 112938 273693
rect 112656 273640 112938 273659
rect 111404 273432 111446 273640
rect 112702 273638 112938 273640
rect 111524 273624 112624 273630
rect 111524 273590 111553 273624
rect 111587 273590 111625 273624
rect 111659 273590 111697 273624
rect 111731 273590 111769 273624
rect 111803 273590 111841 273624
rect 111875 273590 111913 273624
rect 111947 273590 111985 273624
rect 112019 273590 112057 273624
rect 112091 273590 112129 273624
rect 112163 273590 112201 273624
rect 112235 273590 112273 273624
rect 112307 273590 112345 273624
rect 112379 273590 112417 273624
rect 112451 273590 112489 273624
rect 112523 273590 112561 273624
rect 112595 273590 112624 273624
rect 111524 273584 112624 273590
rect 111524 273482 112624 273488
rect 111524 273448 111553 273482
rect 111587 273448 111625 273482
rect 111659 273448 111697 273482
rect 111731 273448 111769 273482
rect 111803 273448 111841 273482
rect 111875 273448 111913 273482
rect 111947 273448 111985 273482
rect 112019 273448 112057 273482
rect 112091 273448 112129 273482
rect 112163 273448 112201 273482
rect 112235 273448 112273 273482
rect 112307 273448 112345 273482
rect 112379 273448 112417 273482
rect 112451 273448 112489 273482
rect 112523 273448 112561 273482
rect 112595 273448 112624 273482
rect 111524 273442 112624 273448
rect 112702 273432 112744 273638
rect 112850 273621 112938 273638
rect 112850 273587 112898 273621
rect 112932 273587 112938 273621
rect 112850 273544 112938 273587
rect 114102 273693 114190 273736
rect 116015 273736 116057 273830
rect 116135 273786 117235 273792
rect 116135 273752 116164 273786
rect 116198 273752 116236 273786
rect 116270 273752 116308 273786
rect 116342 273752 116380 273786
rect 116414 273752 116452 273786
rect 116486 273752 116524 273786
rect 116558 273752 116596 273786
rect 116630 273752 116668 273786
rect 116702 273752 116740 273786
rect 116774 273752 116812 273786
rect 116846 273752 116884 273786
rect 116918 273752 116956 273786
rect 116990 273752 117028 273786
rect 117062 273752 117100 273786
rect 117134 273752 117172 273786
rect 117206 273752 117235 273786
rect 116135 273746 117235 273752
rect 117313 273736 117355 273830
rect 117459 273792 117503 273968
rect 117581 273984 118681 273990
rect 117581 273950 117610 273984
rect 117644 273950 117682 273984
rect 117716 273950 117754 273984
rect 117788 273950 117826 273984
rect 117860 273950 117898 273984
rect 117932 273950 117970 273984
rect 118004 273950 118042 273984
rect 118076 273950 118114 273984
rect 118148 273950 118186 273984
rect 118220 273950 118258 273984
rect 118292 273950 118330 273984
rect 118364 273950 118402 273984
rect 118436 273950 118474 273984
rect 118508 273950 118546 273984
rect 118580 273950 118618 273984
rect 118652 273950 118681 273984
rect 117581 273944 118681 273950
rect 117581 273842 118681 273848
rect 117581 273808 117610 273842
rect 117644 273808 117682 273842
rect 117716 273808 117754 273842
rect 117788 273808 117826 273842
rect 117860 273808 117898 273842
rect 117932 273808 117970 273842
rect 118004 273808 118042 273842
rect 118076 273808 118114 273842
rect 118148 273808 118186 273842
rect 118220 273808 118258 273842
rect 118292 273808 118330 273842
rect 118364 273808 118402 273842
rect 118436 273808 118474 273842
rect 118508 273808 118546 273842
rect 118580 273808 118618 273842
rect 118652 273808 118681 273842
rect 117581 273802 118681 273808
rect 118759 273792 118801 274000
rect 117459 273769 117549 273792
rect 117459 273748 117509 273769
rect 114102 273659 114108 273693
rect 114142 273659 114190 273693
rect 114657 273727 114857 273733
rect 114657 273693 114704 273727
rect 114738 273693 114776 273727
rect 114810 273693 114857 273727
rect 114657 273687 114857 273693
rect 115348 273727 115548 273733
rect 115348 273693 115395 273727
rect 115429 273693 115467 273727
rect 115501 273693 115548 273727
rect 115348 273687 115548 273693
rect 116015 273693 116103 273736
rect 114102 273621 114190 273659
rect 114102 273587 114108 273621
rect 114142 273587 114190 273621
rect 114720 273619 114790 273687
rect 114102 273544 114190 273587
rect 114308 273535 114790 273619
rect 114865 273622 114970 273647
rect 114865 273570 114890 273622
rect 114942 273570 114970 273622
rect 114865 273540 114970 273570
rect 115235 273622 115340 273647
rect 115235 273570 115262 273622
rect 115314 273570 115340 273622
rect 115235 273540 115340 273570
rect 115415 273619 115485 273687
rect 116015 273659 116063 273693
rect 116097 273659 116103 273693
rect 116015 273621 116103 273659
rect 112970 273528 114070 273534
rect 112970 273494 112999 273528
rect 113033 273494 113071 273528
rect 113105 273494 113143 273528
rect 113177 273494 113215 273528
rect 113249 273494 113287 273528
rect 113321 273494 113359 273528
rect 113393 273494 113431 273528
rect 113465 273494 113503 273528
rect 113537 273494 113575 273528
rect 113609 273494 113647 273528
rect 113681 273494 113719 273528
rect 113753 273494 113791 273528
rect 113825 273494 113863 273528
rect 113897 273494 113935 273528
rect 113969 273494 114007 273528
rect 114041 273494 114070 273528
rect 112970 273488 114070 273494
rect 111404 273409 111492 273432
rect 111404 273375 111452 273409
rect 111486 273375 111492 273409
rect 111404 273337 111492 273375
rect 111404 273303 111452 273337
rect 111486 273303 111492 273337
rect 111404 273280 111492 273303
rect 112656 273409 112744 273432
rect 114308 273420 114343 273535
rect 114720 273505 114790 273535
rect 115415 273535 115897 273619
rect 116015 273587 116063 273621
rect 116097 273587 116103 273621
rect 116015 273544 116103 273587
rect 117267 273700 117355 273736
rect 117461 273735 117509 273748
rect 117543 273735 117549 273769
rect 117461 273700 117549 273735
rect 117267 273697 117549 273700
rect 117267 273693 117509 273697
rect 117267 273659 117273 273693
rect 117307 273663 117509 273693
rect 117543 273663 117549 273697
rect 117307 273659 117549 273663
rect 117267 273640 117549 273659
rect 118713 273769 118801 273792
rect 118713 273735 118719 273769
rect 118753 273735 118801 273769
rect 118713 273697 118801 273735
rect 118713 273663 118719 273697
rect 118753 273663 118801 273697
rect 118713 273640 118801 273663
rect 117267 273638 117503 273640
rect 117267 273621 117355 273638
rect 117267 273587 117273 273621
rect 117307 273587 117355 273621
rect 117267 273544 117355 273587
rect 115415 273505 115485 273535
rect 114657 273499 114857 273505
rect 114657 273465 114704 273499
rect 114738 273465 114776 273499
rect 114810 273465 114857 273499
rect 114657 273459 114857 273465
rect 115348 273499 115548 273505
rect 115348 273465 115395 273499
rect 115429 273465 115467 273499
rect 115501 273465 115548 273499
rect 115348 273459 115548 273465
rect 112656 273375 112662 273409
rect 112696 273375 112744 273409
rect 113843 273390 114343 273420
rect 112656 273337 112744 273375
rect 113000 273384 114343 273390
rect 113000 273350 113029 273384
rect 113063 273350 113101 273384
rect 113135 273350 113173 273384
rect 113207 273350 113245 273384
rect 113279 273350 113317 273384
rect 113351 273350 113389 273384
rect 113423 273350 113461 273384
rect 113495 273350 113533 273384
rect 113567 273350 113605 273384
rect 113639 273350 113677 273384
rect 113711 273350 113749 273384
rect 113783 273350 113821 273384
rect 113855 273350 113893 273384
rect 113927 273350 113965 273384
rect 113999 273350 114037 273384
rect 114071 273379 114343 273384
rect 114570 273426 114616 273449
rect 114570 273392 114576 273426
rect 114610 273392 114616 273426
rect 114071 273350 114100 273379
rect 113000 273344 114100 273350
rect 114570 273354 114616 273392
rect 112656 273303 112662 273337
rect 112696 273303 112744 273337
rect 112656 273280 112744 273303
rect 105964 270099 106243 273149
rect 111404 273072 111446 273280
rect 111524 273264 112624 273270
rect 111524 273230 111553 273264
rect 111587 273230 111625 273264
rect 111659 273230 111697 273264
rect 111731 273230 111769 273264
rect 111803 273230 111841 273264
rect 111875 273230 111913 273264
rect 111947 273230 111985 273264
rect 112019 273230 112057 273264
rect 112091 273230 112129 273264
rect 112163 273230 112201 273264
rect 112235 273230 112273 273264
rect 112307 273230 112345 273264
rect 112379 273230 112417 273264
rect 112451 273230 112489 273264
rect 112523 273230 112561 273264
rect 112595 273230 112624 273264
rect 111524 273224 112624 273230
rect 111524 273122 112624 273128
rect 111524 273088 111553 273122
rect 111587 273088 111625 273122
rect 111659 273088 111697 273122
rect 111731 273088 111769 273122
rect 111803 273088 111841 273122
rect 111875 273088 111913 273122
rect 111947 273088 111985 273122
rect 112019 273088 112057 273122
rect 112091 273088 112129 273122
rect 112163 273088 112201 273122
rect 112235 273088 112273 273122
rect 112307 273088 112345 273122
rect 112379 273088 112417 273122
rect 112451 273088 112489 273122
rect 112523 273088 112561 273122
rect 112595 273088 112624 273122
rect 111524 273082 112624 273088
rect 112702 273072 112744 273280
rect 111404 273049 111492 273072
rect 111404 273015 111452 273049
rect 111486 273015 111492 273049
rect 111404 272977 111492 273015
rect 111404 272943 111452 272977
rect 111486 272943 111492 272977
rect 111404 272920 111492 272943
rect 112656 273049 112744 273072
rect 112656 273015 112662 273049
rect 112696 273015 112744 273049
rect 112656 272977 112744 273015
rect 112656 272943 112662 272977
rect 112696 272943 112744 272977
rect 112656 272920 112744 272943
rect 112874 273315 112968 273334
rect 112874 273281 112928 273315
rect 112962 273281 112968 273315
rect 112874 273262 112968 273281
rect 114132 273315 114226 273334
rect 114132 273281 114138 273315
rect 114172 273281 114226 273315
rect 114132 273262 114226 273281
rect 112874 273170 112922 273262
rect 113000 273246 114100 273252
rect 113000 273212 113029 273246
rect 113063 273212 113101 273246
rect 113135 273212 113173 273246
rect 113207 273212 113245 273246
rect 113279 273212 113317 273246
rect 113351 273212 113389 273246
rect 113423 273212 113461 273246
rect 113495 273212 113533 273246
rect 113567 273212 113605 273246
rect 113639 273212 113677 273246
rect 113711 273212 113749 273246
rect 113783 273212 113821 273246
rect 113855 273212 113893 273246
rect 113927 273212 113965 273246
rect 113999 273212 114037 273246
rect 114071 273212 114100 273246
rect 113000 273206 114100 273212
rect 114178 273170 114226 273262
rect 112874 273126 114226 273170
rect 114324 273287 114396 273328
rect 114570 273320 114576 273354
rect 114610 273320 114616 273354
rect 114570 273297 114616 273320
rect 114898 273426 114944 273449
rect 114898 273392 114904 273426
rect 114938 273392 114944 273426
rect 114898 273354 114944 273392
rect 114898 273320 114904 273354
rect 114938 273320 114944 273354
rect 114898 273297 114944 273320
rect 115261 273426 115307 273449
rect 115261 273392 115267 273426
rect 115301 273392 115307 273426
rect 115261 273354 115307 273392
rect 115261 273320 115267 273354
rect 115301 273320 115307 273354
rect 115261 273297 115307 273320
rect 115589 273426 115635 273449
rect 115589 273392 115595 273426
rect 115629 273392 115635 273426
rect 115589 273354 115635 273392
rect 115862 273420 115897 273535
rect 116135 273528 117235 273534
rect 116135 273494 116164 273528
rect 116198 273494 116236 273528
rect 116270 273494 116308 273528
rect 116342 273494 116380 273528
rect 116414 273494 116452 273528
rect 116486 273494 116524 273528
rect 116558 273494 116596 273528
rect 116630 273494 116668 273528
rect 116702 273494 116740 273528
rect 116774 273494 116812 273528
rect 116846 273494 116884 273528
rect 116918 273494 116956 273528
rect 116990 273494 117028 273528
rect 117062 273494 117100 273528
rect 117134 273494 117172 273528
rect 117206 273494 117235 273528
rect 116135 273488 117235 273494
rect 117461 273432 117503 273638
rect 117581 273624 118681 273630
rect 117581 273590 117610 273624
rect 117644 273590 117682 273624
rect 117716 273590 117754 273624
rect 117788 273590 117826 273624
rect 117860 273590 117898 273624
rect 117932 273590 117970 273624
rect 118004 273590 118042 273624
rect 118076 273590 118114 273624
rect 118148 273590 118186 273624
rect 118220 273590 118258 273624
rect 118292 273590 118330 273624
rect 118364 273590 118402 273624
rect 118436 273590 118474 273624
rect 118508 273590 118546 273624
rect 118580 273590 118618 273624
rect 118652 273590 118681 273624
rect 117581 273584 118681 273590
rect 117581 273482 118681 273488
rect 117581 273448 117610 273482
rect 117644 273448 117682 273482
rect 117716 273448 117754 273482
rect 117788 273448 117826 273482
rect 117860 273448 117898 273482
rect 117932 273448 117970 273482
rect 118004 273448 118042 273482
rect 118076 273448 118114 273482
rect 118148 273448 118186 273482
rect 118220 273448 118258 273482
rect 118292 273448 118330 273482
rect 118364 273448 118402 273482
rect 118436 273448 118474 273482
rect 118508 273448 118546 273482
rect 118580 273448 118618 273482
rect 118652 273448 118681 273482
rect 117581 273442 118681 273448
rect 118759 273432 118801 273640
rect 120377 273964 120423 273981
rect 120377 273930 120383 273964
rect 120417 273930 120423 273964
rect 120377 273892 120423 273930
rect 120377 273858 120383 273892
rect 120417 273858 120423 273892
rect 120377 273820 120423 273858
rect 120377 273786 120383 273820
rect 120417 273786 120423 273820
rect 120377 273748 120423 273786
rect 120377 273714 120383 273748
rect 120417 273714 120423 273748
rect 120377 273676 120423 273714
rect 120377 273642 120383 273676
rect 120417 273642 120423 273676
rect 120377 273604 120423 273642
rect 120377 273570 120383 273604
rect 120417 273570 120423 273604
rect 120377 273532 120423 273570
rect 120377 273498 120383 273532
rect 120417 273498 120423 273532
rect 120377 273481 120423 273498
rect 120835 273964 120881 273981
rect 120835 273930 120841 273964
rect 120875 273930 120881 273964
rect 120835 273892 120881 273930
rect 120835 273858 120841 273892
rect 120875 273858 120881 273892
rect 120835 273820 120881 273858
rect 120835 273786 120841 273820
rect 120875 273786 120881 273820
rect 120835 273778 120881 273786
rect 120950 273778 121028 276032
rect 121077 276028 121123 276032
rect 121077 275994 121083 276028
rect 121117 275994 121123 276028
rect 121077 275956 121123 275994
rect 121077 275922 121083 275956
rect 121117 275922 121123 275956
rect 121077 275884 121123 275922
rect 121077 275850 121083 275884
rect 121117 275850 121123 275884
rect 121077 275833 121123 275850
rect 121535 276316 121581 276333
rect 121535 276282 121541 276316
rect 121575 276282 121581 276316
rect 121535 276244 121581 276282
rect 121535 276210 121541 276244
rect 121575 276210 121581 276244
rect 121535 276172 121581 276210
rect 121802 276207 121933 276287
rect 121802 276172 121841 276207
rect 121535 276138 121541 276172
rect 121575 276138 121581 276172
rect 121535 276135 121581 276138
rect 121801 276155 121841 276172
rect 121893 276155 121933 276207
rect 121801 276143 121933 276155
rect 121801 276135 121841 276143
rect 121535 276100 121841 276135
rect 121535 276066 121541 276100
rect 121575 276091 121841 276100
rect 121893 276091 121933 276143
rect 121575 276079 121933 276091
rect 121575 276066 121841 276079
rect 121535 276028 121841 276066
rect 121535 275994 121541 276028
rect 121575 275994 121581 276028
rect 121535 275956 121581 275994
rect 121535 275922 121541 275956
rect 121575 275922 121581 275956
rect 121802 276027 121841 276028
rect 121893 276027 121933 276079
rect 122096 276118 122427 276154
rect 124055 276118 124112 276514
rect 122096 276112 124349 276118
rect 122096 276078 122137 276112
rect 122171 276078 122209 276112
rect 122243 276078 122281 276112
rect 122315 276078 122353 276112
rect 122387 276078 124349 276112
rect 122096 276049 124349 276078
rect 124445 276049 124567 277394
rect 122096 276035 122427 276049
rect 121802 275945 121933 276027
rect 121535 275884 121581 275922
rect 121535 275850 121541 275884
rect 121575 275850 121581 275884
rect 121535 275833 121581 275850
rect 122390 275807 122422 276035
rect 122629 275863 122686 276049
rect 122466 275857 122866 275863
rect 122466 275823 122505 275857
rect 122539 275823 122577 275857
rect 122611 275823 122649 275857
rect 122683 275823 122721 275857
rect 122755 275823 122793 275857
rect 122827 275823 122866 275857
rect 122466 275817 122866 275823
rect 122970 275807 123002 276049
rect 123272 275863 123329 276049
rect 123102 275857 123502 275863
rect 123102 275823 123141 275857
rect 123175 275823 123213 275857
rect 123247 275823 123285 275857
rect 123319 275823 123357 275857
rect 123391 275823 123429 275857
rect 123463 275823 123502 275857
rect 123102 275817 123502 275823
rect 123605 275807 123637 276049
rect 123915 275863 123972 276049
rect 124240 275863 124272 276049
rect 124445 276015 124490 276049
rect 124524 276015 124567 276049
rect 124445 275955 124567 276015
rect 123738 275857 124138 275863
rect 123738 275823 123777 275857
rect 123811 275823 123849 275857
rect 123883 275823 123921 275857
rect 123955 275823 123993 275857
rect 124027 275823 124065 275857
rect 124099 275823 124138 275857
rect 123738 275817 124138 275823
rect 124240 275857 124774 275863
rect 124240 275823 124413 275857
rect 124447 275823 124485 275857
rect 124519 275823 124557 275857
rect 124591 275823 124629 275857
rect 124663 275823 124701 275857
rect 124735 275823 124774 275857
rect 124240 275817 124774 275823
rect 124240 275807 124374 275817
rect 121133 275786 121525 275792
rect 121133 275752 121168 275786
rect 121202 275752 121240 275786
rect 121274 275752 121312 275786
rect 121346 275752 121384 275786
rect 121418 275752 121456 275786
rect 121490 275752 121525 275786
rect 121133 275630 121525 275752
rect 122379 275778 122425 275807
rect 122379 275744 122385 275778
rect 122419 275744 122425 275778
rect 122379 275715 122425 275744
rect 122907 275778 123061 275807
rect 122907 275744 122913 275778
rect 122947 275744 123021 275778
rect 123055 275744 123061 275778
rect 122907 275715 123061 275744
rect 123543 275778 123697 275807
rect 123543 275744 123549 275778
rect 123583 275744 123657 275778
rect 123691 275744 123697 275778
rect 123543 275715 123697 275744
rect 124179 275797 124374 275807
rect 124179 275778 124333 275797
rect 124179 275744 124185 275778
rect 124219 275744 124293 275778
rect 124327 275744 124333 275778
rect 124179 275715 124333 275744
rect 124815 275778 124861 275807
rect 124815 275744 124821 275778
rect 124855 275744 124861 275778
rect 124815 275715 124861 275744
rect 122466 275699 122866 275705
rect 122466 275665 122505 275699
rect 122539 275665 122577 275699
rect 122611 275665 122649 275699
rect 122683 275665 122721 275699
rect 122755 275665 122793 275699
rect 122827 275665 122866 275699
rect 122466 275659 122866 275665
rect 123102 275699 123502 275705
rect 123102 275665 123141 275699
rect 123175 275665 123213 275699
rect 123247 275665 123285 275699
rect 123319 275665 123357 275699
rect 123391 275665 123429 275699
rect 123463 275665 123502 275699
rect 123102 275659 123502 275665
rect 123738 275699 124138 275705
rect 123738 275665 123777 275699
rect 123811 275665 123849 275699
rect 123883 275665 123921 275699
rect 123955 275665 123993 275699
rect 124027 275665 124065 275699
rect 124099 275665 124138 275699
rect 123738 275659 124138 275665
rect 121133 275596 121168 275630
rect 121202 275596 121240 275630
rect 121274 275596 121312 275630
rect 121346 275596 121384 275630
rect 121418 275596 121456 275630
rect 121490 275596 121525 275630
rect 121133 275590 121525 275596
rect 121077 275532 121123 275549
rect 121077 275498 121083 275532
rect 121117 275498 121123 275532
rect 121077 275460 121123 275498
rect 121077 275426 121083 275460
rect 121117 275426 121123 275460
rect 121077 275388 121123 275426
rect 121077 275354 121083 275388
rect 121117 275354 121123 275388
rect 121077 275316 121123 275354
rect 121077 275282 121083 275316
rect 121117 275282 121123 275316
rect 121077 275244 121123 275282
rect 121077 275210 121083 275244
rect 121117 275210 121123 275244
rect 121077 275172 121123 275210
rect 121077 275138 121083 275172
rect 121117 275138 121123 275172
rect 121077 275100 121123 275138
rect 121077 275066 121083 275100
rect 121117 275066 121123 275100
rect 121077 275049 121123 275066
rect 121535 275532 121628 275549
rect 121535 275498 121541 275532
rect 121575 275498 121628 275532
rect 121535 275460 121628 275498
rect 121535 275426 121541 275460
rect 121575 275426 121628 275460
rect 124244 275475 124285 275715
rect 124374 275699 124774 275705
rect 124374 275665 124413 275699
rect 124447 275665 124485 275699
rect 124519 275665 124557 275699
rect 124591 275665 124629 275699
rect 124663 275665 124701 275699
rect 124735 275665 124774 275699
rect 124374 275659 124774 275665
rect 124818 275475 124859 275715
rect 124244 275432 124859 275475
rect 121535 275388 121628 275426
rect 121535 275354 121541 275388
rect 121575 275354 121628 275388
rect 121535 275316 121628 275354
rect 123213 275368 123457 275431
rect 121535 275282 121541 275316
rect 121575 275282 121628 275316
rect 121535 275244 121628 275282
rect 121535 275210 121541 275244
rect 121575 275210 121628 275244
rect 121535 275172 121628 275210
rect 121535 275138 121541 275172
rect 121575 275138 121628 275172
rect 121535 275100 121628 275138
rect 121535 275066 121541 275100
rect 121575 275070 121628 275100
rect 122354 275286 122587 275333
rect 122354 275070 122415 275286
rect 121575 275066 122415 275070
rect 121535 275049 122415 275066
rect 121133 275002 121525 275008
rect 121133 274968 121168 275002
rect 121202 274968 121240 275002
rect 121274 274968 121312 275002
rect 121346 274968 121384 275002
rect 121418 274968 121456 275002
rect 121490 274968 121525 275002
rect 121133 274846 121525 274968
rect 121133 274812 121168 274846
rect 121202 274812 121240 274846
rect 121274 274812 121312 274846
rect 121346 274812 121384 274846
rect 121418 274812 121456 274846
rect 121490 274812 121525 274846
rect 121133 274806 121525 274812
rect 121581 274786 122415 275049
rect 122531 274786 122587 275286
rect 123213 275190 123246 275368
rect 123424 275336 123457 275368
rect 123424 275231 124318 275336
rect 123424 275190 123457 275231
rect 123213 275140 123457 275190
rect 124132 274973 124318 275231
rect 123881 274943 124318 274973
rect 125452 275151 128452 275523
rect 125452 275136 125825 275151
rect 128019 275136 128452 275151
rect 123881 274940 124366 274943
rect 122956 274934 123948 274940
rect 122956 274900 123003 274934
rect 123037 274900 123075 274934
rect 123109 274900 123147 274934
rect 123181 274900 123219 274934
rect 123253 274900 123291 274934
rect 123325 274900 123363 274934
rect 123397 274900 123435 274934
rect 123469 274900 123507 274934
rect 123541 274900 123579 274934
rect 123613 274900 123651 274934
rect 123685 274900 123723 274934
rect 123757 274900 123795 274934
rect 123829 274900 123867 274934
rect 123901 274900 123948 274934
rect 122956 274894 123948 274900
rect 122900 274815 122946 274862
rect 122900 274807 122906 274815
rect 121581 274765 122587 274786
rect 121077 274748 121123 274765
rect 121077 274714 121083 274748
rect 121117 274714 121123 274748
rect 121077 274676 121123 274714
rect 121077 274642 121083 274676
rect 121117 274642 121123 274676
rect 121077 274604 121123 274642
rect 121077 274570 121083 274604
rect 121117 274570 121123 274604
rect 121077 274532 121123 274570
rect 121077 274498 121083 274532
rect 121117 274498 121123 274532
rect 121077 274460 121123 274498
rect 121077 274426 121083 274460
rect 121117 274426 121123 274460
rect 121077 274388 121123 274426
rect 121077 274354 121083 274388
rect 121117 274354 121123 274388
rect 121077 274316 121123 274354
rect 121077 274282 121083 274316
rect 121117 274282 121123 274316
rect 121077 274265 121123 274282
rect 121535 274748 122587 274765
rect 121535 274714 121541 274748
rect 121575 274736 122587 274748
rect 122706 274781 122906 274807
rect 122940 274781 122946 274815
rect 122706 274765 122946 274781
rect 121575 274714 121628 274736
rect 121535 274676 121628 274714
rect 121535 274642 121541 274676
rect 121575 274642 121628 274676
rect 121535 274604 121628 274642
rect 121535 274570 121541 274604
rect 121575 274570 121628 274604
rect 121535 274532 121628 274570
rect 121535 274498 121541 274532
rect 121575 274498 121628 274532
rect 121535 274460 121628 274498
rect 121535 274426 121541 274460
rect 121575 274426 121628 274460
rect 121535 274388 121628 274426
rect 122706 274454 122746 274765
rect 122900 274743 122946 274765
rect 122900 274709 122906 274743
rect 122940 274709 122946 274743
rect 122900 274662 122946 274709
rect 123958 274815 124004 274862
rect 123958 274781 123964 274815
rect 123998 274781 124004 274815
rect 123958 274743 124004 274781
rect 123958 274709 123964 274743
rect 123998 274709 124004 274743
rect 123958 274662 124004 274709
rect 122956 274624 123948 274630
rect 122956 274590 123003 274624
rect 123037 274590 123075 274624
rect 123109 274590 123147 274624
rect 123181 274590 123219 274624
rect 123253 274590 123291 274624
rect 123325 274590 123363 274624
rect 123397 274590 123435 274624
rect 123469 274590 123507 274624
rect 123541 274590 123579 274624
rect 123613 274590 123651 274624
rect 123685 274590 123723 274624
rect 123757 274590 123795 274624
rect 123829 274590 123867 274624
rect 123901 274590 123948 274624
rect 122956 274584 123948 274590
rect 124116 274584 124366 274940
rect 123879 274574 124366 274584
rect 123879 274551 124148 274574
rect 122706 274452 123624 274454
rect 122706 274443 123670 274452
rect 122706 274418 123534 274443
rect 123497 274409 123534 274418
rect 123568 274409 123606 274443
rect 123640 274409 123670 274443
rect 123497 274401 123670 274409
rect 121535 274354 121541 274388
rect 121575 274354 121628 274388
rect 124001 274397 124921 274447
rect 124001 274356 124100 274397
rect 121535 274316 121628 274354
rect 121535 274282 121541 274316
rect 121575 274282 121628 274316
rect 122281 274350 122477 274356
rect 122281 274316 122324 274350
rect 122358 274316 122396 274350
rect 122430 274316 122477 274350
rect 122281 274310 122477 274316
rect 122697 274350 124137 274356
rect 122697 274316 122740 274350
rect 122774 274316 122812 274350
rect 122846 274316 123156 274350
rect 123190 274316 123228 274350
rect 123262 274316 123572 274350
rect 123606 274316 123644 274350
rect 123678 274316 123988 274350
rect 124022 274316 124060 274350
rect 124094 274316 124137 274350
rect 122697 274310 124137 274316
rect 124357 274350 124553 274356
rect 124357 274316 124404 274350
rect 124438 274316 124476 274350
rect 124510 274316 124553 274350
rect 124357 274310 124553 274316
rect 121535 274265 121628 274282
rect 122225 274261 122271 274278
rect 122225 274227 122231 274261
rect 122265 274227 122271 274261
rect 121133 274218 121525 274224
rect 121133 274184 121168 274218
rect 121202 274184 121240 274218
rect 121274 274184 121312 274218
rect 121346 274184 121384 274218
rect 121418 274184 121456 274218
rect 121490 274184 121525 274218
rect 121133 274062 121525 274184
rect 121133 274028 121168 274062
rect 121202 274028 121240 274062
rect 121274 274028 121312 274062
rect 121346 274028 121384 274062
rect 121418 274028 121456 274062
rect 121490 274028 121525 274062
rect 121133 274022 121525 274028
rect 122225 274189 122271 274227
rect 122225 274155 122231 274189
rect 122265 274155 122271 274189
rect 122225 274117 122271 274155
rect 122225 274083 122231 274117
rect 122265 274083 122271 274117
rect 122225 274045 122271 274083
rect 122225 274011 122231 274045
rect 122265 274011 122271 274045
rect 121077 273964 121123 273981
rect 121077 273930 121083 273964
rect 121117 273930 121123 273964
rect 121077 273892 121123 273930
rect 121077 273858 121083 273892
rect 121117 273858 121123 273892
rect 121077 273820 121123 273858
rect 121077 273786 121083 273820
rect 121117 273786 121123 273820
rect 121077 273778 121123 273786
rect 120835 273748 121123 273778
rect 120835 273714 120841 273748
rect 120875 273741 121083 273748
rect 120875 273714 120972 273741
rect 120835 273707 120972 273714
rect 121006 273714 121083 273741
rect 121117 273714 121123 273748
rect 121006 273707 121123 273714
rect 120835 273676 121123 273707
rect 120835 273642 120841 273676
rect 120875 273671 121083 273676
rect 120875 273642 120881 273671
rect 120835 273604 120881 273642
rect 120835 273570 120841 273604
rect 120875 273570 120881 273604
rect 120835 273532 120881 273570
rect 120835 273498 120841 273532
rect 120875 273498 120881 273532
rect 120835 273481 120881 273498
rect 121077 273642 121083 273671
rect 121117 273642 121123 273676
rect 121077 273604 121123 273642
rect 121077 273570 121083 273604
rect 121117 273570 121123 273604
rect 121077 273532 121123 273570
rect 121077 273498 121083 273532
rect 121117 273498 121123 273532
rect 121077 273481 121123 273498
rect 121535 273964 121581 273981
rect 121535 273930 121541 273964
rect 121575 273930 121581 273964
rect 121535 273892 121581 273930
rect 121535 273858 121541 273892
rect 121575 273858 121581 273892
rect 122225 273973 122271 274011
rect 122225 273939 122231 273973
rect 122265 273939 122271 273973
rect 122225 273901 122271 273939
rect 121535 273820 121581 273858
rect 121535 273786 121541 273820
rect 121575 273786 121581 273820
rect 121535 273769 121581 273786
rect 121803 273805 121934 273885
rect 121803 273770 121842 273805
rect 121764 273769 121842 273770
rect 121535 273753 121842 273769
rect 121894 273753 121934 273805
rect 122225 273867 122231 273901
rect 122265 273867 122271 273901
rect 122225 273829 122271 273867
rect 122225 273795 122231 273829
rect 122265 273795 122271 273829
rect 122225 273778 122271 273795
rect 122483 274261 122529 274278
rect 122483 274227 122489 274261
rect 122523 274227 122529 274261
rect 122483 274189 122529 274227
rect 122483 274155 122489 274189
rect 122523 274155 122529 274189
rect 122483 274117 122529 274155
rect 122483 274083 122489 274117
rect 122523 274083 122529 274117
rect 122483 274045 122529 274083
rect 122483 274011 122489 274045
rect 122523 274011 122529 274045
rect 122641 274261 122687 274278
rect 122641 274227 122647 274261
rect 122681 274227 122687 274261
rect 122641 274189 122687 274227
rect 122641 274155 122647 274189
rect 122681 274155 122687 274189
rect 122641 274117 122687 274155
rect 122641 274083 122647 274117
rect 122681 274083 122687 274117
rect 122641 274045 122687 274083
rect 122641 274044 122647 274045
rect 122483 273973 122529 274011
rect 122483 273939 122489 273973
rect 122523 273939 122529 273973
rect 122483 273901 122529 273939
rect 122483 273867 122489 273901
rect 122523 273867 122529 273901
rect 122483 273829 122529 273867
rect 122483 273795 122489 273829
rect 122523 273795 122529 273829
rect 122483 273778 122529 273795
rect 122602 274011 122647 274044
rect 122681 274011 122687 274045
rect 122602 273973 122687 274011
rect 122602 273939 122647 273973
rect 122681 273939 122687 273973
rect 122602 273901 122687 273939
rect 122602 273867 122647 273901
rect 122681 273867 122687 273901
rect 122602 273829 122687 273867
rect 122602 273795 122647 273829
rect 122681 273795 122687 273829
rect 122602 273778 122687 273795
rect 122899 274261 122945 274278
rect 122899 274227 122905 274261
rect 122939 274227 122945 274261
rect 122899 274189 122945 274227
rect 122899 274155 122905 274189
rect 122939 274155 122945 274189
rect 122899 274117 122945 274155
rect 122899 274083 122905 274117
rect 122939 274083 122945 274117
rect 122899 274045 122945 274083
rect 122899 274011 122905 274045
rect 122939 274011 122945 274045
rect 123057 274261 123103 274278
rect 123057 274227 123063 274261
rect 123097 274227 123103 274261
rect 123057 274189 123103 274227
rect 123057 274155 123063 274189
rect 123097 274155 123103 274189
rect 123057 274117 123103 274155
rect 123057 274083 123063 274117
rect 123097 274083 123103 274117
rect 123057 274045 123103 274083
rect 123057 274044 123063 274045
rect 122899 273973 122945 274011
rect 122899 273939 122905 273973
rect 122939 273939 122945 273973
rect 122899 273901 122945 273939
rect 122899 273867 122905 273901
rect 122939 273867 122945 273901
rect 122899 273829 122945 273867
rect 122899 273795 122905 273829
rect 122939 273795 122945 273829
rect 122899 273778 122945 273795
rect 123018 274011 123063 274044
rect 123097 274011 123103 274045
rect 123018 273973 123103 274011
rect 123018 273939 123063 273973
rect 123097 273939 123103 273973
rect 123018 273901 123103 273939
rect 123018 273867 123063 273901
rect 123097 273867 123103 273901
rect 123018 273829 123103 273867
rect 123018 273795 123063 273829
rect 123097 273795 123103 273829
rect 123018 273778 123103 273795
rect 123315 274261 123361 274278
rect 123315 274227 123321 274261
rect 123355 274227 123361 274261
rect 123315 274189 123361 274227
rect 123315 274155 123321 274189
rect 123355 274155 123361 274189
rect 123315 274117 123361 274155
rect 123315 274083 123321 274117
rect 123355 274083 123361 274117
rect 123315 274045 123361 274083
rect 123315 274011 123321 274045
rect 123355 274011 123361 274045
rect 123473 274261 123519 274278
rect 123473 274227 123479 274261
rect 123513 274227 123519 274261
rect 123473 274189 123519 274227
rect 123473 274155 123479 274189
rect 123513 274155 123519 274189
rect 123473 274117 123519 274155
rect 123473 274083 123479 274117
rect 123513 274083 123519 274117
rect 123473 274045 123519 274083
rect 123473 274044 123479 274045
rect 123315 273973 123361 274011
rect 123315 273939 123321 273973
rect 123355 273939 123361 273973
rect 123315 273901 123361 273939
rect 123315 273867 123321 273901
rect 123355 273867 123361 273901
rect 123315 273829 123361 273867
rect 123315 273795 123321 273829
rect 123355 273795 123361 273829
rect 123315 273778 123361 273795
rect 123434 274011 123479 274044
rect 123513 274011 123519 274045
rect 123434 273973 123519 274011
rect 123434 273939 123479 273973
rect 123513 273939 123519 273973
rect 123434 273901 123519 273939
rect 123434 273867 123479 273901
rect 123513 273867 123519 273901
rect 123434 273829 123519 273867
rect 123434 273795 123479 273829
rect 123513 273795 123519 273829
rect 123434 273778 123519 273795
rect 123731 274261 123777 274278
rect 123731 274227 123737 274261
rect 123771 274227 123777 274261
rect 123731 274189 123777 274227
rect 123731 274155 123737 274189
rect 123771 274155 123777 274189
rect 123731 274117 123777 274155
rect 123731 274083 123737 274117
rect 123771 274083 123777 274117
rect 123731 274045 123777 274083
rect 123731 274011 123737 274045
rect 123771 274011 123777 274045
rect 123889 274261 123935 274278
rect 123889 274227 123895 274261
rect 123929 274227 123935 274261
rect 123889 274189 123935 274227
rect 123889 274155 123895 274189
rect 123929 274155 123935 274189
rect 123889 274117 123935 274155
rect 123889 274083 123895 274117
rect 123929 274083 123935 274117
rect 123889 274045 123935 274083
rect 123889 274044 123895 274045
rect 123731 273973 123777 274011
rect 123731 273939 123737 273973
rect 123771 273939 123777 273973
rect 123731 273901 123777 273939
rect 123731 273867 123737 273901
rect 123771 273867 123777 273901
rect 123731 273829 123777 273867
rect 123731 273795 123737 273829
rect 123771 273795 123777 273829
rect 123731 273778 123777 273795
rect 123850 274011 123895 274044
rect 123929 274011 123935 274045
rect 123850 273973 123935 274011
rect 123850 273939 123895 273973
rect 123929 273939 123935 273973
rect 123850 273901 123935 273939
rect 123850 273867 123895 273901
rect 123929 273867 123935 273901
rect 123850 273829 123935 273867
rect 123850 273795 123895 273829
rect 123929 273795 123935 273829
rect 123850 273778 123935 273795
rect 124147 274261 124193 274278
rect 124147 274227 124153 274261
rect 124187 274227 124193 274261
rect 124147 274189 124193 274227
rect 124147 274155 124153 274189
rect 124187 274155 124193 274189
rect 124147 274117 124193 274155
rect 124147 274083 124153 274117
rect 124187 274083 124193 274117
rect 124147 274045 124193 274083
rect 124147 274011 124153 274045
rect 124187 274011 124193 274045
rect 124147 273973 124193 274011
rect 124147 273939 124153 273973
rect 124187 273939 124193 273973
rect 124147 273901 124193 273939
rect 124147 273867 124153 273901
rect 124187 273867 124193 273901
rect 124147 273829 124193 273867
rect 124147 273795 124153 273829
rect 124187 273795 124193 273829
rect 124147 273778 124193 273795
rect 124305 274261 124351 274278
rect 124305 274227 124311 274261
rect 124345 274227 124351 274261
rect 124305 274189 124351 274227
rect 124305 274155 124311 274189
rect 124345 274155 124351 274189
rect 124305 274117 124351 274155
rect 124305 274083 124311 274117
rect 124345 274083 124351 274117
rect 124305 274045 124351 274083
rect 124305 274011 124311 274045
rect 124345 274011 124351 274045
rect 124305 273973 124351 274011
rect 124305 273939 124311 273973
rect 124345 273939 124351 273973
rect 124305 273901 124351 273939
rect 124305 273867 124311 273901
rect 124345 273867 124351 273901
rect 124305 273829 124351 273867
rect 124305 273795 124311 273829
rect 124345 273795 124351 273829
rect 124305 273778 124351 273795
rect 124563 274261 124609 274278
rect 124563 274227 124569 274261
rect 124603 274227 124609 274261
rect 124563 274189 124609 274227
rect 124563 274155 124569 274189
rect 124603 274155 124609 274189
rect 124563 274117 124609 274155
rect 124563 274083 124569 274117
rect 124603 274083 124609 274117
rect 124563 274045 124609 274083
rect 124563 274011 124569 274045
rect 124603 274011 124609 274045
rect 124563 273973 124609 274011
rect 124563 273939 124569 273973
rect 124603 273939 124609 273973
rect 124563 273901 124609 273939
rect 124563 273867 124569 273901
rect 124603 273867 124609 273901
rect 124563 273829 124609 273867
rect 124563 273795 124569 273829
rect 124603 273795 124609 273829
rect 124563 273778 124609 273795
rect 121535 273748 121934 273753
rect 121535 273714 121541 273748
rect 121575 273741 121934 273748
rect 121575 273714 121842 273741
rect 121535 273689 121842 273714
rect 121894 273689 121934 273741
rect 122281 273740 122473 273746
rect 122281 273706 122324 273740
rect 122358 273706 122396 273740
rect 122430 273706 122473 273740
rect 122281 273700 122473 273706
rect 121535 273677 121934 273689
rect 121535 273676 121842 273677
rect 121535 273642 121541 273676
rect 121575 273662 121842 273676
rect 121575 273642 121581 273662
rect 121764 273661 121842 273662
rect 121535 273604 121581 273642
rect 121535 273570 121541 273604
rect 121575 273570 121581 273604
rect 121535 273532 121581 273570
rect 121803 273625 121842 273661
rect 121894 273625 121934 273677
rect 121803 273543 121934 273625
rect 121535 273498 121541 273532
rect 121575 273498 121581 273532
rect 121535 273481 121581 273498
rect 122602 273468 122652 273778
rect 122697 273740 122889 273746
rect 122697 273706 122740 273740
rect 122774 273706 122812 273740
rect 122846 273706 122889 273740
rect 122697 273700 122889 273706
rect 123018 273477 123068 273778
rect 123113 273740 123305 273746
rect 123113 273706 123156 273740
rect 123190 273706 123228 273740
rect 123262 273706 123305 273740
rect 123113 273700 123305 273706
rect 123434 273477 123484 273778
rect 123529 273740 123721 273746
rect 123529 273706 123572 273740
rect 123606 273706 123644 273740
rect 123678 273706 123721 273740
rect 123529 273700 123721 273706
rect 122602 273449 122755 273468
rect 115862 273390 116362 273420
rect 117461 273409 117549 273432
rect 115862 273384 117205 273390
rect 115862 273379 116134 273384
rect 115589 273320 115595 273354
rect 115629 273320 115635 273354
rect 116105 273350 116134 273379
rect 116168 273350 116206 273384
rect 116240 273350 116278 273384
rect 116312 273350 116350 273384
rect 116384 273350 116422 273384
rect 116456 273350 116494 273384
rect 116528 273350 116566 273384
rect 116600 273350 116638 273384
rect 116672 273350 116710 273384
rect 116744 273350 116782 273384
rect 116816 273350 116854 273384
rect 116888 273350 116926 273384
rect 116960 273350 116998 273384
rect 117032 273350 117070 273384
rect 117104 273350 117142 273384
rect 117176 273350 117205 273384
rect 116105 273344 117205 273350
rect 117461 273375 117509 273409
rect 117543 273375 117549 273409
rect 117461 273337 117549 273375
rect 115589 273297 115635 273320
rect 115809 273287 115881 273328
rect 114324 273253 114342 273287
rect 114376 273253 114396 273287
rect 114324 273197 114396 273253
rect 114657 273281 114857 273287
rect 114657 273247 114704 273281
rect 114738 273247 114776 273281
rect 114810 273247 114857 273281
rect 114657 273241 114857 273247
rect 115348 273281 115548 273287
rect 115348 273247 115395 273281
rect 115429 273247 115467 273281
rect 115501 273247 115548 273281
rect 115348 273241 115548 273247
rect 115809 273253 115828 273287
rect 115862 273253 115881 273287
rect 114843 273197 115030 273212
rect 114324 273152 114781 273197
rect 112874 273036 112922 273126
rect 113000 273086 114100 273092
rect 113000 273052 113029 273086
rect 113063 273052 113101 273086
rect 113135 273052 113173 273086
rect 113207 273052 113245 273086
rect 113279 273052 113317 273086
rect 113351 273052 113389 273086
rect 113423 273052 113461 273086
rect 113495 273052 113533 273086
rect 113567 273052 113605 273086
rect 113639 273052 113677 273086
rect 113711 273052 113749 273086
rect 113783 273052 113821 273086
rect 113855 273052 113893 273086
rect 113927 273052 113965 273086
rect 113999 273052 114037 273086
rect 114071 273052 114100 273086
rect 113000 273046 114100 273052
rect 114178 273036 114226 273126
rect 114737 273097 114781 273152
rect 114843 273145 114891 273197
rect 114943 273145 115030 273197
rect 114843 273127 115030 273145
rect 115175 273197 115362 273212
rect 115809 273197 115881 273253
rect 115175 273145 115262 273197
rect 115314 273145 115362 273197
rect 115175 273127 115362 273145
rect 115424 273152 115881 273197
rect 115979 273315 116073 273334
rect 115979 273281 116033 273315
rect 116067 273281 116073 273315
rect 115979 273262 116073 273281
rect 117237 273315 117331 273334
rect 117237 273281 117243 273315
rect 117277 273281 117331 273315
rect 117237 273262 117331 273281
rect 115979 273170 116027 273262
rect 116105 273246 117205 273252
rect 116105 273212 116134 273246
rect 116168 273212 116206 273246
rect 116240 273212 116278 273246
rect 116312 273212 116350 273246
rect 116384 273212 116422 273246
rect 116456 273212 116494 273246
rect 116528 273212 116566 273246
rect 116600 273212 116638 273246
rect 116672 273212 116710 273246
rect 116744 273212 116782 273246
rect 116816 273212 116854 273246
rect 116888 273212 116926 273246
rect 116960 273212 116998 273246
rect 117032 273212 117070 273246
rect 117104 273212 117142 273246
rect 117176 273212 117205 273246
rect 116105 273206 117205 273212
rect 117283 273170 117331 273262
rect 115424 273097 115468 273152
rect 115979 273126 117331 273170
rect 114657 273091 114857 273097
rect 114657 273057 114704 273091
rect 114738 273057 114776 273091
rect 114810 273057 114857 273091
rect 114657 273051 114857 273057
rect 115348 273091 115548 273097
rect 115348 273057 115395 273091
rect 115429 273057 115467 273091
rect 115501 273057 115548 273091
rect 115348 273051 115548 273057
rect 112874 273017 112968 273036
rect 112874 272983 112928 273017
rect 112962 272983 112968 273017
rect 112874 272964 112968 272983
rect 114132 273017 114226 273036
rect 114132 272983 114138 273017
rect 114172 272983 114226 273017
rect 114132 272964 114226 272983
rect 114570 273018 114616 273041
rect 114570 272984 114576 273018
rect 114610 272984 114616 273018
rect 111524 272904 112624 272910
rect 111524 272870 111553 272904
rect 111587 272870 111625 272904
rect 111659 272870 111697 272904
rect 111731 272870 111769 272904
rect 111803 272870 111841 272904
rect 111875 272870 111913 272904
rect 111947 272870 111985 272904
rect 112019 272870 112057 272904
rect 112091 272870 112129 272904
rect 112163 272870 112201 272904
rect 112235 272870 112273 272904
rect 112307 272870 112345 272904
rect 112379 272870 112417 272904
rect 112451 272870 112489 272904
rect 112523 272870 112561 272904
rect 112595 272870 112624 272904
rect 111524 272866 112624 272870
rect 112874 272870 112922 272964
rect 114327 272959 114395 272960
rect 114570 272959 114616 272984
rect 113000 272948 114100 272954
rect 113000 272914 113029 272948
rect 113063 272914 113101 272948
rect 113135 272914 113173 272948
rect 113207 272914 113245 272948
rect 113279 272914 113317 272948
rect 113351 272914 113389 272948
rect 113423 272914 113461 272948
rect 113495 272914 113533 272948
rect 113567 272914 113605 272948
rect 113639 272914 113677 272948
rect 113711 272914 113749 272948
rect 113783 272914 113821 272948
rect 113855 272914 113893 272948
rect 113927 272914 113965 272948
rect 113999 272914 114037 272948
rect 114071 272914 114100 272948
rect 113000 272908 114100 272914
rect 114327 272946 114616 272959
rect 114327 272912 114576 272946
rect 114610 272912 114616 272946
rect 114327 272899 114616 272912
rect 114327 272870 114395 272899
rect 114570 272889 114616 272899
rect 114898 273018 114944 273041
rect 114898 272984 114904 273018
rect 114938 272984 114944 273018
rect 114898 272946 114944 272984
rect 114898 272912 114904 272946
rect 114938 272912 114944 272946
rect 114898 272889 114944 272912
rect 115261 273018 115307 273041
rect 115261 272984 115267 273018
rect 115301 272984 115307 273018
rect 115261 272946 115307 272984
rect 115261 272912 115267 272946
rect 115301 272912 115307 272946
rect 115261 272889 115307 272912
rect 115589 273018 115635 273041
rect 115589 272984 115595 273018
rect 115629 272984 115635 273018
rect 115589 272959 115635 272984
rect 115979 273036 116027 273126
rect 116105 273086 117205 273092
rect 116105 273052 116134 273086
rect 116168 273052 116206 273086
rect 116240 273052 116278 273086
rect 116312 273052 116350 273086
rect 116384 273052 116422 273086
rect 116456 273052 116494 273086
rect 116528 273052 116566 273086
rect 116600 273052 116638 273086
rect 116672 273052 116710 273086
rect 116744 273052 116782 273086
rect 116816 273052 116854 273086
rect 116888 273052 116926 273086
rect 116960 273052 116998 273086
rect 117032 273052 117070 273086
rect 117104 273052 117142 273086
rect 117176 273052 117205 273086
rect 116105 273046 117205 273052
rect 117283 273036 117331 273126
rect 115979 273017 116073 273036
rect 115979 272983 116033 273017
rect 116067 272983 116073 273017
rect 115979 272964 116073 272983
rect 117237 273017 117331 273036
rect 117237 272983 117243 273017
rect 117277 272983 117331 273017
rect 117237 272964 117331 272983
rect 115810 272959 115878 272960
rect 115589 272946 115878 272959
rect 115589 272912 115595 272946
rect 115629 272912 115878 272946
rect 115589 272899 115878 272912
rect 116105 272948 117205 272954
rect 116105 272914 116134 272948
rect 116168 272914 116206 272948
rect 116240 272914 116278 272948
rect 116312 272914 116350 272948
rect 116384 272914 116422 272948
rect 116456 272914 116494 272948
rect 116528 272914 116566 272948
rect 116600 272914 116638 272948
rect 116672 272914 116710 272948
rect 116744 272914 116782 272948
rect 116816 272914 116854 272948
rect 116888 272914 116926 272948
rect 116960 272914 116998 272948
rect 117032 272914 117070 272948
rect 117104 272914 117142 272948
rect 117176 272914 117205 272948
rect 116105 272908 117205 272914
rect 115589 272889 115635 272899
rect 112874 272866 114395 272870
rect 111524 272864 114395 272866
rect 112044 272830 114395 272864
rect 114657 272873 114857 272879
rect 114657 272839 114704 272873
rect 114738 272839 114776 272873
rect 114810 272839 114857 272873
rect 114657 272833 114857 272839
rect 115348 272873 115548 272879
rect 115348 272839 115395 272873
rect 115429 272839 115467 272873
rect 115501 272839 115548 272873
rect 115348 272833 115548 272839
rect 115810 272870 115878 272899
rect 117283 272870 117331 272964
rect 117461 273303 117509 273337
rect 117543 273303 117549 273337
rect 117461 273280 117549 273303
rect 118713 273409 118801 273432
rect 118713 273375 118719 273409
rect 118753 273375 118801 273409
rect 118713 273337 118801 273375
rect 118713 273303 118719 273337
rect 118753 273303 118801 273337
rect 118713 273280 118801 273303
rect 117461 273072 117503 273280
rect 117581 273264 118681 273270
rect 117581 273230 117610 273264
rect 117644 273230 117682 273264
rect 117716 273230 117754 273264
rect 117788 273230 117826 273264
rect 117860 273230 117898 273264
rect 117932 273230 117970 273264
rect 118004 273230 118042 273264
rect 118076 273230 118114 273264
rect 118148 273230 118186 273264
rect 118220 273230 118258 273264
rect 118292 273230 118330 273264
rect 118364 273230 118402 273264
rect 118436 273230 118474 273264
rect 118508 273230 118546 273264
rect 118580 273230 118618 273264
rect 118652 273230 118681 273264
rect 117581 273224 118681 273230
rect 117581 273122 118681 273128
rect 117581 273088 117610 273122
rect 117644 273088 117682 273122
rect 117716 273088 117754 273122
rect 117788 273088 117826 273122
rect 117860 273088 117898 273122
rect 117932 273088 117970 273122
rect 118004 273088 118042 273122
rect 118076 273088 118114 273122
rect 118148 273088 118186 273122
rect 118220 273088 118258 273122
rect 118292 273088 118330 273122
rect 118364 273088 118402 273122
rect 118436 273088 118474 273122
rect 118508 273088 118546 273122
rect 118580 273088 118618 273122
rect 118652 273088 118681 273122
rect 117581 273082 118681 273088
rect 118759 273072 118801 273280
rect 120433 273434 120825 273440
rect 120433 273400 120468 273434
rect 120502 273400 120540 273434
rect 120574 273400 120612 273434
rect 120646 273400 120684 273434
rect 120718 273400 120756 273434
rect 120790 273400 120825 273434
rect 120433 273278 120825 273400
rect 120433 273244 120468 273278
rect 120502 273244 120540 273278
rect 120574 273244 120612 273278
rect 120646 273244 120684 273278
rect 120718 273244 120756 273278
rect 120790 273244 120825 273278
rect 120433 273238 120825 273244
rect 121133 273434 121525 273440
rect 121133 273400 121168 273434
rect 121202 273400 121240 273434
rect 121274 273400 121312 273434
rect 121346 273400 121384 273434
rect 121418 273400 121456 273434
rect 121490 273400 121525 273434
rect 121133 273278 121525 273400
rect 122602 273397 122652 273449
rect 122704 273397 122755 273449
rect 122602 273371 122755 273397
rect 123018 273420 123484 273477
rect 123850 273468 123900 273778
rect 123945 273740 124137 273746
rect 123945 273706 123988 273740
rect 124022 273706 124060 273740
rect 124094 273706 124137 273740
rect 123945 273700 124137 273706
rect 124361 273740 124553 273746
rect 124361 273706 124404 273740
rect 124438 273706 124476 273740
rect 124510 273706 124553 273740
rect 124361 273700 124553 273706
rect 124865 273477 124921 274397
rect 123747 273449 123900 273468
rect 123018 273320 123689 273420
rect 123747 273397 123797 273449
rect 123849 273397 123900 273449
rect 123747 273371 123900 273397
rect 124396 273399 124921 273477
rect 121133 273244 121168 273278
rect 121202 273244 121240 273278
rect 121274 273244 121312 273278
rect 121346 273244 121384 273278
rect 121418 273244 121456 273278
rect 121490 273244 121525 273278
rect 121133 273238 121525 273244
rect 117461 273049 117549 273072
rect 117461 273015 117509 273049
rect 117543 273015 117549 273049
rect 117461 272977 117549 273015
rect 117461 272943 117509 272977
rect 117543 272943 117549 272977
rect 117461 272920 117549 272943
rect 118713 273049 118801 273072
rect 118713 273015 118719 273049
rect 118753 273015 118801 273049
rect 118713 272977 118801 273015
rect 118713 272943 118719 272977
rect 118753 272943 118801 272977
rect 118713 272920 118801 272943
rect 120377 273180 120423 273197
rect 120377 273146 120383 273180
rect 120417 273146 120423 273180
rect 120377 273108 120423 273146
rect 120377 273074 120383 273108
rect 120417 273074 120423 273108
rect 120377 273036 120423 273074
rect 120377 273002 120383 273036
rect 120417 273002 120423 273036
rect 120377 272964 120423 273002
rect 120377 272930 120383 272964
rect 120417 272930 120423 272964
rect 115810 272866 117331 272870
rect 117581 272904 118681 272910
rect 117581 272870 117610 272904
rect 117644 272870 117682 272904
rect 117716 272870 117754 272904
rect 117788 272870 117826 272904
rect 117860 272870 117898 272904
rect 117932 272870 117970 272904
rect 118004 272870 118042 272904
rect 118076 272870 118114 272904
rect 118148 272870 118186 272904
rect 118220 272870 118258 272904
rect 118292 272870 118330 272904
rect 118364 272870 118402 272904
rect 118436 272870 118474 272904
rect 118508 272870 118546 272904
rect 118580 272870 118618 272904
rect 118652 272870 118681 272904
rect 117581 272866 118681 272870
rect 115810 272864 118681 272866
rect 120377 272892 120423 272930
rect 112719 272788 112924 272830
rect 113982 272756 114266 272766
rect 114724 272756 114783 272833
rect 113982 272735 114783 272756
rect 113982 272701 114034 272735
rect 114068 272701 114106 272735
rect 114140 272701 114178 272735
rect 114212 272701 114783 272735
rect 113982 272667 114783 272701
rect 114928 272766 115275 272825
rect 113982 272666 114266 272667
rect 114928 272540 115016 272766
rect 109394 272507 109556 272513
rect 109394 272473 109458 272507
rect 109492 272473 109556 272507
rect 109394 272467 109556 272473
rect 110973 272444 115016 272540
rect 115194 272444 115275 272766
rect 115422 272756 115481 272833
rect 115810 272830 118161 272864
rect 120377 272858 120383 272892
rect 120417 272858 120423 272892
rect 117281 272788 117486 272830
rect 120377 272820 120423 272858
rect 120377 272786 120383 272820
rect 120417 272786 120423 272820
rect 115939 272756 116223 272766
rect 115422 272735 116223 272756
rect 115422 272701 115992 272735
rect 116026 272701 116064 272735
rect 116098 272701 116136 272735
rect 116170 272701 116223 272735
rect 115422 272667 116223 272701
rect 120377 272748 120423 272786
rect 120377 272714 120383 272748
rect 120417 272714 120423 272748
rect 120377 272697 120423 272714
rect 120835 273180 120881 273197
rect 120835 273146 120841 273180
rect 120875 273146 120881 273180
rect 120835 273108 120881 273146
rect 120835 273074 120841 273108
rect 120875 273074 120881 273108
rect 120835 273036 120881 273074
rect 120835 273002 120841 273036
rect 120875 273008 120881 273036
rect 121077 273180 121123 273197
rect 121077 273146 121083 273180
rect 121117 273146 121123 273180
rect 121077 273108 121123 273146
rect 121077 273074 121083 273108
rect 121117 273074 121123 273108
rect 121077 273036 121123 273074
rect 121077 273008 121083 273036
rect 120875 273002 121083 273008
rect 121117 273002 121123 273036
rect 120835 272981 121123 273002
rect 120835 272964 120959 272981
rect 120835 272930 120841 272964
rect 120875 272930 120959 272964
rect 120835 272929 120959 272930
rect 121011 272964 121123 272981
rect 121011 272930 121083 272964
rect 121117 272930 121123 272964
rect 121011 272929 121123 272930
rect 120835 272917 121123 272929
rect 120835 272892 120959 272917
rect 120835 272858 120841 272892
rect 120875 272881 120959 272892
rect 120875 272858 120881 272881
rect 120835 272820 120881 272858
rect 120835 272786 120841 272820
rect 120875 272786 120881 272820
rect 120835 272748 120881 272786
rect 120835 272714 120841 272748
rect 120875 272714 120881 272748
rect 120835 272697 120881 272714
rect 120953 272865 120959 272881
rect 121011 272892 121123 272917
rect 121011 272881 121083 272892
rect 121011 272865 121018 272881
rect 120953 272853 121018 272865
rect 120953 272801 120959 272853
rect 121011 272801 121018 272853
rect 120953 272789 121018 272801
rect 120953 272737 120959 272789
rect 121011 272737 121018 272789
rect 115939 272666 116223 272667
rect 120433 272650 120825 272656
rect 120433 272616 120468 272650
rect 120502 272616 120540 272650
rect 120574 272616 120612 272650
rect 120646 272616 120684 272650
rect 120718 272616 120756 272650
rect 120790 272616 120825 272650
rect 120433 272494 120825 272616
rect 120433 272460 120468 272494
rect 120502 272460 120540 272494
rect 120574 272460 120612 272494
rect 120646 272460 120684 272494
rect 120718 272460 120756 272494
rect 120790 272460 120825 272494
rect 120433 272454 120825 272460
rect 109388 272411 109434 272426
rect 109388 272377 109394 272411
rect 109428 272377 109434 272411
rect 109388 272339 109434 272377
rect 109388 272305 109394 272339
rect 109428 272305 109434 272339
rect 109388 272267 109434 272305
rect 109388 272233 109394 272267
rect 109428 272233 109434 272267
rect 106985 272157 108373 272215
rect 106985 272043 107187 272157
rect 107463 272151 108075 272157
rect 107463 272117 107500 272151
rect 107534 272117 107572 272151
rect 107606 272117 107644 272151
rect 107678 272117 107716 272151
rect 107750 272117 107788 272151
rect 107822 272117 107860 272151
rect 107894 272117 107932 272151
rect 107966 272117 108004 272151
rect 108038 272117 108075 272151
rect 107463 272111 108075 272117
rect 106985 272009 106997 272043
rect 107031 272009 107069 272043
rect 107103 272009 107141 272043
rect 107175 272009 107187 272043
rect 106985 272003 107187 272009
rect 107407 272032 107453 272079
rect 107407 271998 107413 272032
rect 107447 271998 107453 272032
rect 107407 271971 107453 271998
rect 106929 271942 106975 271971
rect 106929 271908 106935 271942
rect 106969 271908 106975 271942
rect 106929 271870 106975 271908
rect 106929 271836 106935 271870
rect 106969 271836 106975 271870
rect 106929 271807 106975 271836
rect 107197 271960 107453 271971
rect 107197 271949 107413 271960
rect 107197 271942 107300 271949
rect 107197 271908 107203 271942
rect 107237 271908 107300 271942
rect 107197 271897 107300 271908
rect 107352 271926 107413 271949
rect 107447 271926 107453 271960
rect 107352 271897 107453 271926
rect 107197 271888 107453 271897
rect 107197 271885 107413 271888
rect 107197 271870 107300 271885
rect 107197 271836 107203 271870
rect 107237 271836 107300 271870
rect 107197 271833 107300 271836
rect 107352 271854 107413 271885
rect 107447 271854 107453 271888
rect 107352 271833 107453 271854
rect 107197 271816 107453 271833
rect 107197 271807 107413 271816
rect 107407 271782 107413 271807
rect 107447 271782 107453 271816
rect 106951 271769 107187 271775
rect 106951 271735 106997 271769
rect 107031 271735 107069 271769
rect 107103 271735 107141 271769
rect 107175 271735 107187 271769
rect 107407 271735 107453 271782
rect 108085 272032 108131 272079
rect 108085 271998 108091 272032
rect 108125 271998 108131 272032
rect 108085 271985 108131 271998
rect 108243 271985 108373 272157
rect 109388 272195 109434 272233
rect 109388 272161 109394 272195
rect 109428 272161 109434 272195
rect 109388 272123 109434 272161
rect 108595 272088 108841 272113
rect 109388 272089 109394 272123
rect 109428 272089 109434 272123
rect 109388 272088 109434 272089
rect 108595 272078 109434 272088
rect 108595 272026 108651 272078
rect 108703 272026 108715 272078
rect 108767 272026 108779 272078
rect 108831 272051 109434 272078
rect 108831 272026 109394 272051
rect 108595 272017 109394 272026
rect 109428 272017 109434 272051
rect 108595 272010 109434 272017
rect 108595 271995 108841 272010
rect 108085 271960 108373 271985
rect 108085 271926 108091 271960
rect 108125 271926 108373 271960
rect 108085 271888 108373 271926
rect 108085 271854 108091 271888
rect 108125 271854 108373 271888
rect 108085 271821 108373 271854
rect 108085 271816 108131 271821
rect 108085 271782 108091 271816
rect 108125 271782 108131 271816
rect 108085 271735 108131 271782
rect 106951 271637 107187 271735
rect 107463 271697 108075 271703
rect 107463 271663 107500 271697
rect 107534 271663 107572 271697
rect 107606 271663 107644 271697
rect 107678 271663 107716 271697
rect 107750 271663 107788 271697
rect 107822 271663 107860 271697
rect 107894 271663 107932 271697
rect 107966 271663 108004 271697
rect 108038 271663 108075 271697
rect 107463 271637 108075 271663
rect 106951 271587 108075 271637
rect 106951 271485 107027 271587
rect 107463 271541 108075 271587
rect 108265 271659 108373 271821
rect 109388 271979 109434 272010
rect 109388 271945 109394 271979
rect 109428 271945 109434 271979
rect 109388 271907 109434 271945
rect 109388 271873 109394 271907
rect 109428 271873 109434 271907
rect 109388 271835 109434 271873
rect 109388 271801 109394 271835
rect 109428 271801 109434 271835
rect 109388 271763 109434 271801
rect 109388 271729 109394 271763
rect 109428 271729 109434 271763
rect 109388 271691 109434 271729
rect 108265 271611 108507 271659
rect 108265 271541 108373 271611
rect 107173 271535 108373 271541
rect 107173 271501 107216 271535
rect 107250 271501 107288 271535
rect 107322 271501 107360 271535
rect 107394 271501 107432 271535
rect 107466 271501 107504 271535
rect 107538 271501 107576 271535
rect 107610 271501 107648 271535
rect 107682 271501 107720 271535
rect 107754 271501 107792 271535
rect 107826 271501 107864 271535
rect 107898 271501 107936 271535
rect 107970 271501 108008 271535
rect 108042 271501 108080 271535
rect 108114 271501 108152 271535
rect 108186 271501 108224 271535
rect 108258 271501 108296 271535
rect 108330 271501 108373 271535
rect 107173 271495 108373 271501
rect 108465 271485 108507 271611
rect 106951 271458 107141 271485
rect 106951 271406 107049 271458
rect 107101 271453 107141 271458
rect 107135 271419 107141 271453
rect 107101 271406 107141 271419
rect 106951 271394 107141 271406
rect 106951 271342 107049 271394
rect 107101 271381 107141 271394
rect 107135 271347 107141 271381
rect 107101 271342 107141 271347
rect 106951 271315 107141 271342
rect 108405 271458 108507 271485
rect 108405 271453 108445 271458
rect 108405 271419 108411 271453
rect 108405 271406 108445 271419
rect 108497 271406 108507 271458
rect 108405 271394 108507 271406
rect 108405 271381 108445 271394
rect 108405 271347 108411 271381
rect 108405 271342 108445 271347
rect 108497 271342 108507 271394
rect 108405 271315 108507 271342
rect 109388 271657 109394 271691
rect 109428 271657 109434 271691
rect 109388 271619 109434 271657
rect 109388 271585 109394 271619
rect 109428 271585 109434 271619
rect 109388 271547 109434 271585
rect 109388 271513 109394 271547
rect 109428 271513 109434 271547
rect 109388 271475 109434 271513
rect 109388 271441 109394 271475
rect 109428 271441 109434 271475
rect 109388 271403 109434 271441
rect 109388 271369 109394 271403
rect 109428 271369 109434 271403
rect 109388 271331 109434 271369
rect 106951 271304 107039 271315
rect 106951 271252 106967 271304
rect 107019 271252 107039 271304
rect 107173 271299 108373 271305
rect 107173 271265 107216 271299
rect 107250 271265 107288 271299
rect 107322 271265 107360 271299
rect 107394 271265 107432 271299
rect 107466 271265 107504 271299
rect 107538 271265 107576 271299
rect 107610 271265 107648 271299
rect 107682 271265 107720 271299
rect 107754 271265 107792 271299
rect 107826 271265 107864 271299
rect 107898 271265 107936 271299
rect 107970 271265 108008 271299
rect 108042 271265 108080 271299
rect 108114 271265 108152 271299
rect 108186 271265 108224 271299
rect 108258 271265 108296 271299
rect 108330 271265 108373 271299
rect 107173 271259 108373 271265
rect 109388 271297 109394 271331
rect 109428 271297 109434 271331
rect 109388 271259 109434 271297
rect 106951 271240 107039 271252
rect 106951 271188 106967 271240
rect 107019 271213 107039 271240
rect 108103 271217 108697 271259
rect 107019 271188 107229 271213
rect 106951 271177 107229 271188
rect 106951 271176 107039 271177
rect 106951 271124 106967 271176
rect 107019 271124 107039 271176
rect 107173 271171 107229 271177
rect 107173 271165 108373 271171
rect 107173 271131 107216 271165
rect 107250 271131 107288 271165
rect 107322 271131 107360 271165
rect 107394 271131 107432 271165
rect 107466 271131 107504 271165
rect 107538 271131 107576 271165
rect 107610 271131 107648 271165
rect 107682 271131 107720 271165
rect 107754 271131 107792 271165
rect 107826 271131 107864 271165
rect 107898 271131 107936 271165
rect 107970 271131 108008 271165
rect 108042 271131 108080 271165
rect 108114 271131 108152 271165
rect 108186 271131 108224 271165
rect 108258 271131 108296 271165
rect 108330 271131 108373 271165
rect 107173 271125 108373 271131
rect 106951 271115 107039 271124
rect 106951 271088 107141 271115
rect 106951 271036 107049 271088
rect 107101 271083 107141 271088
rect 107135 271049 107141 271083
rect 107101 271036 107141 271049
rect 106951 271024 107141 271036
rect 106951 270972 107049 271024
rect 107101 271011 107141 271024
rect 107135 270977 107141 271011
rect 107101 270972 107141 270977
rect 106951 270945 107141 270972
rect 108405 271088 108507 271115
rect 108405 271083 108445 271088
rect 108405 271049 108411 271083
rect 108405 271036 108445 271049
rect 108497 271036 108507 271088
rect 108405 271024 108507 271036
rect 108405 271011 108445 271024
rect 108405 270977 108411 271011
rect 108405 270972 108445 270977
rect 108497 270972 108507 271024
rect 108405 270945 108507 270972
rect 108551 271029 108697 271217
rect 109388 271225 109394 271259
rect 109428 271225 109434 271259
rect 109388 271187 109434 271225
rect 109388 271153 109394 271187
rect 109428 271153 109434 271187
rect 109388 271115 109434 271153
rect 109388 271081 109394 271115
rect 109428 271081 109434 271115
rect 109388 271043 109434 271081
rect 108551 270974 109106 271029
rect 108551 270940 109009 270974
rect 109043 270940 109106 270974
rect 107173 270929 108373 270935
rect 107173 270895 107216 270929
rect 107250 270895 107288 270929
rect 107322 270895 107360 270929
rect 107394 270895 107432 270929
rect 107466 270895 107504 270929
rect 107538 270895 107576 270929
rect 107610 270895 107648 270929
rect 107682 270895 107720 270929
rect 107754 270895 107792 270929
rect 107826 270895 107864 270929
rect 107898 270895 107936 270929
rect 107970 270895 108008 270929
rect 108042 270895 108080 270929
rect 108114 270895 108152 270929
rect 108186 270895 108224 270929
rect 108258 270895 108296 270929
rect 108330 270895 108373 270929
rect 107173 270891 108373 270895
rect 108551 270902 109106 270940
rect 108551 270891 109009 270902
rect 107173 270889 109009 270891
rect 108103 270868 109009 270889
rect 109043 270868 109106 270902
rect 108103 270811 109106 270868
rect 109388 271009 109394 271043
rect 109428 271009 109434 271043
rect 109388 270971 109434 271009
rect 109388 270937 109394 270971
rect 109428 270937 109434 270971
rect 109388 270899 109434 270937
rect 109388 270865 109394 270899
rect 109428 270865 109434 270899
rect 109388 270827 109434 270865
rect 108776 270099 109055 270811
rect 109388 270793 109394 270827
rect 109428 270793 109434 270827
rect 109388 270755 109434 270793
rect 109388 270721 109394 270755
rect 109428 270721 109434 270755
rect 109388 270706 109434 270721
rect 109516 272411 109562 272426
rect 109516 272377 109522 272411
rect 109556 272377 109562 272411
rect 109516 272339 109562 272377
rect 109516 272305 109522 272339
rect 109556 272305 109562 272339
rect 109516 272267 109562 272305
rect 109516 272233 109522 272267
rect 109556 272233 109562 272267
rect 109516 272195 109562 272233
rect 109516 272161 109522 272195
rect 109556 272161 109562 272195
rect 109516 272123 109562 272161
rect 109516 272089 109522 272123
rect 109556 272089 109562 272123
rect 109516 272051 109562 272089
rect 109516 272017 109522 272051
rect 109556 272017 109562 272051
rect 109516 271979 109562 272017
rect 109516 271945 109522 271979
rect 109556 271945 109562 271979
rect 109516 271907 109562 271945
rect 109516 271873 109522 271907
rect 109556 271873 109562 271907
rect 109516 271835 109562 271873
rect 109516 271801 109522 271835
rect 109556 271801 109562 271835
rect 109516 271763 109562 271801
rect 109516 271729 109522 271763
rect 109556 271729 109562 271763
rect 109516 271691 109562 271729
rect 109516 271657 109522 271691
rect 109556 271657 109562 271691
rect 109516 271619 109562 271657
rect 109516 271585 109522 271619
rect 109556 271585 109562 271619
rect 109516 271547 109562 271585
rect 109516 271513 109522 271547
rect 109556 271513 109562 271547
rect 109516 271475 109562 271513
rect 109516 271441 109522 271475
rect 109556 271441 109562 271475
rect 109516 271403 109562 271441
rect 109516 271369 109522 271403
rect 109556 271369 109562 271403
rect 109516 271331 109562 271369
rect 109516 271297 109522 271331
rect 109556 271297 109562 271331
rect 109516 271259 109562 271297
rect 109516 271225 109522 271259
rect 109556 271225 109562 271259
rect 109516 271187 109562 271225
rect 109516 271153 109522 271187
rect 109556 271153 109562 271187
rect 109516 271115 109562 271153
rect 109516 271081 109522 271115
rect 109556 271081 109562 271115
rect 109516 271043 109562 271081
rect 109516 271009 109522 271043
rect 109556 271009 109562 271043
rect 109516 270971 109562 271009
rect 109516 270937 109522 270971
rect 109556 270937 109562 270971
rect 109516 270899 109562 270937
rect 109516 270865 109522 270899
rect 109556 270865 109562 270899
rect 109516 270827 109562 270865
rect 109516 270793 109522 270827
rect 109556 270793 109562 270827
rect 109516 270755 109562 270793
rect 109516 270721 109522 270755
rect 109556 270721 109562 270755
rect 109516 270706 109562 270721
rect 110973 272309 115275 272444
rect 120377 272396 120423 272413
rect 120377 272362 120383 272396
rect 120417 272362 120423 272396
rect 120377 272324 120423 272362
rect 110973 272303 115138 272309
rect 109444 270659 109506 270665
rect 109394 270625 109458 270659
rect 109492 270625 109556 270659
rect 109394 270609 109556 270625
rect 105964 269820 109055 270099
rect 110973 266766 111559 272303
rect 113799 272003 114103 272303
rect 120377 272290 120383 272324
rect 120417 272290 120423 272324
rect 120377 272252 120423 272290
rect 116590 272193 118192 272248
rect 116590 272159 116644 272193
rect 116678 272159 116716 272193
rect 116750 272159 116788 272193
rect 116822 272159 116860 272193
rect 116894 272159 116932 272193
rect 116966 272159 117004 272193
rect 117038 272159 117076 272193
rect 117110 272159 117148 272193
rect 117182 272159 117220 272193
rect 117254 272159 117292 272193
rect 117326 272159 117364 272193
rect 117398 272159 117436 272193
rect 117470 272159 117508 272193
rect 117542 272159 117580 272193
rect 117614 272159 117652 272193
rect 117686 272159 117724 272193
rect 117758 272159 117796 272193
rect 117830 272159 117868 272193
rect 117902 272159 117940 272193
rect 117974 272159 118012 272193
rect 118046 272159 118084 272193
rect 118118 272159 118192 272193
rect 116590 272129 118192 272159
rect 120377 272218 120383 272252
rect 120417 272218 120423 272252
rect 120377 272180 120423 272218
rect 120377 272146 120383 272180
rect 120417 272146 120423 272180
rect 115787 272096 118629 272129
rect 114761 272004 115601 272048
rect 113800 271981 114102 272003
rect 113800 271731 113863 271981
rect 114041 271731 114102 271981
rect 114761 271824 114830 272004
rect 115522 271984 115601 272004
rect 115522 271950 115523 271984
rect 115557 271950 115601 271984
rect 115522 271824 115601 271950
rect 114761 271763 115601 271824
rect 115787 271924 115829 272096
rect 115885 271996 116037 272002
rect 115885 271962 115908 271996
rect 115942 271962 115980 271996
rect 116014 271962 116037 271996
rect 115885 271956 116037 271962
rect 116187 271924 116229 272096
rect 116285 271996 116437 272002
rect 116285 271962 116308 271996
rect 116342 271962 116380 271996
rect 116414 271962 116437 271996
rect 116285 271956 116437 271962
rect 116587 271924 116629 272096
rect 116685 271996 116837 272002
rect 116685 271962 116708 271996
rect 116742 271962 116780 271996
rect 116814 271962 116837 271996
rect 116685 271956 116837 271962
rect 116987 271924 117029 272096
rect 117085 271996 117237 272002
rect 117085 271962 117108 271996
rect 117142 271962 117180 271996
rect 117214 271962 117237 271996
rect 117085 271956 117237 271962
rect 117387 271924 117429 272096
rect 117485 271996 117637 272002
rect 117485 271962 117508 271996
rect 117542 271962 117580 271996
rect 117614 271962 117637 271996
rect 117485 271956 117637 271962
rect 117787 271924 117829 272096
rect 117885 271996 118037 272002
rect 117885 271962 117908 271996
rect 117942 271962 117980 271996
rect 118014 271962 118037 271996
rect 117885 271956 118037 271962
rect 118187 271924 118229 272096
rect 118285 271996 118437 272002
rect 118285 271962 118308 271996
rect 118342 271962 118380 271996
rect 118414 271962 118437 271996
rect 118285 271956 118437 271962
rect 118587 271924 118629 272096
rect 120377 272108 120423 272146
rect 120377 272074 120383 272108
rect 120417 272074 120423 272108
rect 120377 272036 120423 272074
rect 120377 272002 120383 272036
rect 120417 272002 120423 272036
rect 118685 271996 118837 272002
rect 118685 271962 118708 271996
rect 118742 271962 118780 271996
rect 118814 271962 118837 271996
rect 118685 271956 118837 271962
rect 120377 271964 120423 272002
rect 120377 271930 120383 271964
rect 120417 271930 120423 271964
rect 115787 271895 115875 271924
rect 115787 271861 115835 271895
rect 115869 271861 115875 271895
rect 115787 271823 115875 271861
rect 115787 271789 115835 271823
rect 115869 271789 115875 271823
rect 113800 271668 114102 271731
rect 113068 271601 113461 271643
rect 113068 271567 113100 271601
rect 113134 271567 113172 271601
rect 113206 271567 113244 271601
rect 113278 271567 113316 271601
rect 113350 271567 113388 271601
rect 113422 271567 113461 271601
rect 113068 271540 113461 271567
rect 112790 271501 113726 271540
rect 112582 271387 112734 271393
rect 112582 271353 112605 271387
rect 112639 271353 112677 271387
rect 112711 271353 112734 271387
rect 112582 271347 112734 271353
rect 112790 271306 112840 271501
rect 112982 271387 113134 271393
rect 112982 271353 113005 271387
rect 113039 271353 113077 271387
rect 113111 271353 113134 271387
rect 112982 271347 113134 271353
rect 113233 271306 113283 271501
rect 113382 271387 113534 271393
rect 113382 271353 113405 271387
rect 113439 271353 113477 271387
rect 113511 271353 113534 271387
rect 113382 271347 113534 271353
rect 113676 271306 113726 271501
rect 113782 271387 114490 271393
rect 113782 271353 113805 271387
rect 113839 271353 113877 271387
rect 113911 271353 114490 271387
rect 115091 271364 115154 271763
rect 115787 271751 115875 271789
rect 115787 271717 115835 271751
rect 115869 271717 115875 271751
rect 115787 271679 115875 271717
rect 115787 271645 115835 271679
rect 115869 271645 115875 271679
rect 115787 271607 115875 271645
rect 115787 271573 115835 271607
rect 115869 271573 115875 271607
rect 115787 271535 115875 271573
rect 115787 271501 115835 271535
rect 115869 271501 115875 271535
rect 115787 271463 115875 271501
rect 115787 271429 115835 271463
rect 115869 271429 115875 271463
rect 115787 271391 115875 271429
rect 113782 271347 114490 271353
rect 113900 271346 114490 271347
rect 112484 271259 112572 271306
rect 112484 271225 112532 271259
rect 112566 271225 112572 271259
rect 112484 271187 112572 271225
rect 112484 271153 112532 271187
rect 112566 271153 112572 271187
rect 112484 271106 112572 271153
rect 112744 271259 112840 271306
rect 112744 271225 112750 271259
rect 112784 271225 112840 271259
rect 112744 271187 112840 271225
rect 112744 271153 112750 271187
rect 112784 271153 112840 271187
rect 112744 271106 112840 271153
rect 112884 271259 112972 271306
rect 112884 271225 112932 271259
rect 112966 271225 112972 271259
rect 112884 271187 112972 271225
rect 112884 271153 112932 271187
rect 112966 271153 112972 271187
rect 112884 271106 112972 271153
rect 113144 271259 113372 271306
rect 113144 271225 113150 271259
rect 113184 271247 113332 271259
rect 113184 271225 113190 271247
rect 113144 271187 113190 271225
rect 113144 271153 113150 271187
rect 113184 271153 113190 271187
rect 113144 271106 113190 271153
rect 113326 271225 113332 271247
rect 113366 271225 113372 271259
rect 113326 271187 113372 271225
rect 113326 271153 113332 271187
rect 113366 271153 113372 271187
rect 113326 271106 113372 271153
rect 113544 271259 113632 271306
rect 113544 271225 113550 271259
rect 113584 271225 113632 271259
rect 113544 271187 113632 271225
rect 113544 271153 113550 271187
rect 113584 271153 113632 271187
rect 113544 271106 113632 271153
rect 113676 271259 113772 271306
rect 113676 271225 113732 271259
rect 113766 271225 113772 271259
rect 113676 271187 113772 271225
rect 113676 271153 113732 271187
rect 113766 271153 113772 271187
rect 113676 271106 113772 271153
rect 113944 271259 114032 271306
rect 113944 271225 113950 271259
rect 113984 271225 114032 271259
rect 114425 271277 114490 271346
rect 114641 271358 115193 271364
rect 114641 271324 114664 271358
rect 114698 271324 114736 271358
rect 114770 271324 115064 271358
rect 115098 271324 115136 271358
rect 115170 271324 115193 271358
rect 114641 271318 115193 271324
rect 115787 271357 115835 271391
rect 115869 271357 115875 271391
rect 115787 271319 115875 271357
rect 115787 271285 115835 271319
rect 115869 271285 115875 271319
rect 114425 271230 114631 271277
rect 113944 271187 114032 271225
rect 113944 271153 113950 271187
rect 113984 271153 114032 271187
rect 113944 271106 114032 271153
rect 112484 270939 112526 271106
rect 112582 271059 112734 271065
rect 112582 271025 112605 271059
rect 112639 271025 112677 271059
rect 112711 271025 112734 271059
rect 112582 271019 112734 271025
rect 112884 270939 112926 271106
rect 112982 271059 113134 271065
rect 112982 271025 113005 271059
rect 113039 271025 113077 271059
rect 113111 271025 113134 271059
rect 112982 271019 113134 271025
rect 113382 271059 113534 271065
rect 113382 271025 113405 271059
rect 113439 271025 113477 271059
rect 113511 271025 113534 271059
rect 113382 271019 113534 271025
rect 113590 270939 113632 271106
rect 113782 271059 113934 271065
rect 113782 271025 113805 271059
rect 113839 271025 113877 271059
rect 113911 271025 113934 271059
rect 113782 271019 113934 271025
rect 113990 270939 114032 271106
rect 112484 270901 114032 270939
rect 114537 271196 114591 271230
rect 114625 271196 114631 271230
rect 114537 271158 114631 271196
rect 114537 271124 114591 271158
rect 114625 271124 114631 271158
rect 114537 271077 114631 271124
rect 114803 271230 114849 271277
rect 114803 271196 114809 271230
rect 114843 271196 114849 271230
rect 114803 271158 114849 271196
rect 114803 271124 114809 271158
rect 114843 271124 114849 271158
rect 114803 271077 114849 271124
rect 114985 271230 115031 271277
rect 114985 271196 114991 271230
rect 115025 271196 115031 271230
rect 114985 271158 115031 271196
rect 114985 271124 114991 271158
rect 115025 271124 115031 271158
rect 114985 271077 115031 271124
rect 115203 271230 115297 271277
rect 115203 271196 115209 271230
rect 115243 271196 115297 271230
rect 115203 271158 115297 271196
rect 115203 271124 115209 271158
rect 115243 271124 115297 271158
rect 115203 271077 115297 271124
rect 114537 270909 114585 271077
rect 114641 271030 114793 271036
rect 114641 270996 114664 271030
rect 114698 270996 114736 271030
rect 114770 270996 114793 271030
rect 114641 270990 114793 270996
rect 115041 271030 115193 271036
rect 115041 270996 115064 271030
rect 115098 270996 115136 271030
rect 115170 270996 115193 271030
rect 115041 270990 115193 270996
rect 115249 270909 115297 271077
rect 112676 270715 112792 270901
rect 114537 270869 115297 270909
rect 115787 271247 115875 271285
rect 115787 271213 115835 271247
rect 115869 271213 115875 271247
rect 115787 271175 115875 271213
rect 115787 271141 115835 271175
rect 115869 271141 115875 271175
rect 115787 271103 115875 271141
rect 115787 271069 115835 271103
rect 115869 271069 115875 271103
rect 115787 271031 115875 271069
rect 115787 270997 115835 271031
rect 115869 270997 115875 271031
rect 115787 270959 115875 270997
rect 115787 270925 115835 270959
rect 115869 270925 115875 270959
rect 115787 270887 115875 270925
rect 112194 270648 113508 270715
rect 112194 270468 112288 270648
rect 113428 270468 113508 270648
rect 114050 270657 114542 270693
rect 114850 270657 114976 270869
rect 115787 270853 115835 270887
rect 115869 270853 115875 270887
rect 115787 270824 115875 270853
rect 116047 271895 116135 271924
rect 116047 271861 116053 271895
rect 116087 271861 116135 271895
rect 116047 271823 116135 271861
rect 116047 271789 116053 271823
rect 116087 271789 116135 271823
rect 116047 271751 116135 271789
rect 116047 271717 116053 271751
rect 116087 271717 116135 271751
rect 116047 271679 116135 271717
rect 116047 271645 116053 271679
rect 116087 271645 116135 271679
rect 116047 271607 116135 271645
rect 116047 271573 116053 271607
rect 116087 271573 116135 271607
rect 116047 271535 116135 271573
rect 116047 271501 116053 271535
rect 116087 271501 116135 271535
rect 116047 271463 116135 271501
rect 116047 271429 116053 271463
rect 116087 271429 116135 271463
rect 116047 271391 116135 271429
rect 116047 271357 116053 271391
rect 116087 271357 116135 271391
rect 116047 271319 116135 271357
rect 116047 271285 116053 271319
rect 116087 271285 116135 271319
rect 116047 271247 116135 271285
rect 116047 271213 116053 271247
rect 116087 271213 116135 271247
rect 116047 271175 116135 271213
rect 116047 271141 116053 271175
rect 116087 271141 116135 271175
rect 116047 271103 116135 271141
rect 116047 271069 116053 271103
rect 116087 271069 116135 271103
rect 116047 271031 116135 271069
rect 116047 270997 116053 271031
rect 116087 270997 116135 271031
rect 116047 270959 116135 270997
rect 116047 270925 116053 270959
rect 116087 270925 116135 270959
rect 116047 270887 116135 270925
rect 116047 270853 116053 270887
rect 116087 270853 116135 270887
rect 116047 270824 116135 270853
rect 116187 271895 116275 271924
rect 116187 271861 116235 271895
rect 116269 271861 116275 271895
rect 116187 271823 116275 271861
rect 116187 271789 116235 271823
rect 116269 271789 116275 271823
rect 116187 271751 116275 271789
rect 116187 271717 116235 271751
rect 116269 271717 116275 271751
rect 116187 271679 116275 271717
rect 116187 271645 116235 271679
rect 116269 271645 116275 271679
rect 116187 271607 116275 271645
rect 116187 271573 116235 271607
rect 116269 271573 116275 271607
rect 116187 271535 116275 271573
rect 116187 271501 116235 271535
rect 116269 271501 116275 271535
rect 116187 271463 116275 271501
rect 116187 271429 116235 271463
rect 116269 271429 116275 271463
rect 116187 271391 116275 271429
rect 116187 271357 116235 271391
rect 116269 271357 116275 271391
rect 116187 271319 116275 271357
rect 116187 271285 116235 271319
rect 116269 271285 116275 271319
rect 116187 271247 116275 271285
rect 116187 271213 116235 271247
rect 116269 271213 116275 271247
rect 116187 271175 116275 271213
rect 116187 271141 116235 271175
rect 116269 271141 116275 271175
rect 116187 271103 116275 271141
rect 116187 271069 116235 271103
rect 116269 271069 116275 271103
rect 116187 271031 116275 271069
rect 116187 270997 116235 271031
rect 116269 270997 116275 271031
rect 116187 270959 116275 270997
rect 116187 270925 116235 270959
rect 116269 270925 116275 270959
rect 116187 270887 116275 270925
rect 116187 270853 116235 270887
rect 116269 270853 116275 270887
rect 116187 270824 116275 270853
rect 116447 271895 116535 271924
rect 116447 271861 116453 271895
rect 116487 271861 116535 271895
rect 116447 271823 116535 271861
rect 116447 271789 116453 271823
rect 116487 271789 116535 271823
rect 116447 271751 116535 271789
rect 116447 271717 116453 271751
rect 116487 271717 116535 271751
rect 116447 271679 116535 271717
rect 116447 271645 116453 271679
rect 116487 271645 116535 271679
rect 116447 271607 116535 271645
rect 116447 271573 116453 271607
rect 116487 271573 116535 271607
rect 116447 271535 116535 271573
rect 116447 271501 116453 271535
rect 116487 271501 116535 271535
rect 116447 271463 116535 271501
rect 116447 271429 116453 271463
rect 116487 271429 116535 271463
rect 116447 271391 116535 271429
rect 116447 271357 116453 271391
rect 116487 271357 116535 271391
rect 116447 271319 116535 271357
rect 116447 271285 116453 271319
rect 116487 271285 116535 271319
rect 116447 271247 116535 271285
rect 116447 271213 116453 271247
rect 116487 271213 116535 271247
rect 116447 271175 116535 271213
rect 116447 271141 116453 271175
rect 116487 271141 116535 271175
rect 116447 271103 116535 271141
rect 116447 271069 116453 271103
rect 116487 271069 116535 271103
rect 116447 271031 116535 271069
rect 116447 270997 116453 271031
rect 116487 270997 116535 271031
rect 116447 270959 116535 270997
rect 116447 270925 116453 270959
rect 116487 270925 116535 270959
rect 116447 270887 116535 270925
rect 116447 270853 116453 270887
rect 116487 270853 116535 270887
rect 116447 270824 116535 270853
rect 116587 271895 116675 271924
rect 116587 271861 116635 271895
rect 116669 271861 116675 271895
rect 116587 271823 116675 271861
rect 116587 271789 116635 271823
rect 116669 271789 116675 271823
rect 116587 271751 116675 271789
rect 116587 271717 116635 271751
rect 116669 271717 116675 271751
rect 116587 271679 116675 271717
rect 116587 271645 116635 271679
rect 116669 271645 116675 271679
rect 116587 271607 116675 271645
rect 116587 271573 116635 271607
rect 116669 271573 116675 271607
rect 116587 271535 116675 271573
rect 116587 271501 116635 271535
rect 116669 271501 116675 271535
rect 116587 271463 116675 271501
rect 116587 271429 116635 271463
rect 116669 271429 116675 271463
rect 116587 271391 116675 271429
rect 116587 271357 116635 271391
rect 116669 271357 116675 271391
rect 116587 271319 116675 271357
rect 116587 271285 116635 271319
rect 116669 271285 116675 271319
rect 116587 271247 116675 271285
rect 116587 271213 116635 271247
rect 116669 271213 116675 271247
rect 116587 271175 116675 271213
rect 116587 271141 116635 271175
rect 116669 271141 116675 271175
rect 116587 271103 116675 271141
rect 116587 271069 116635 271103
rect 116669 271069 116675 271103
rect 116587 271031 116675 271069
rect 116587 270997 116635 271031
rect 116669 270997 116675 271031
rect 116587 270959 116675 270997
rect 116587 270925 116635 270959
rect 116669 270925 116675 270959
rect 116587 270887 116675 270925
rect 116587 270853 116635 270887
rect 116669 270853 116675 270887
rect 116587 270824 116675 270853
rect 116847 271895 116935 271924
rect 116847 271861 116853 271895
rect 116887 271861 116935 271895
rect 116847 271823 116935 271861
rect 116847 271789 116853 271823
rect 116887 271789 116935 271823
rect 116847 271751 116935 271789
rect 116847 271717 116853 271751
rect 116887 271717 116935 271751
rect 116847 271679 116935 271717
rect 116847 271645 116853 271679
rect 116887 271645 116935 271679
rect 116847 271607 116935 271645
rect 116847 271573 116853 271607
rect 116887 271573 116935 271607
rect 116847 271535 116935 271573
rect 116847 271501 116853 271535
rect 116887 271501 116935 271535
rect 116847 271463 116935 271501
rect 116847 271429 116853 271463
rect 116887 271429 116935 271463
rect 116847 271391 116935 271429
rect 116847 271357 116853 271391
rect 116887 271357 116935 271391
rect 116847 271319 116935 271357
rect 116847 271285 116853 271319
rect 116887 271285 116935 271319
rect 116847 271247 116935 271285
rect 116847 271213 116853 271247
rect 116887 271213 116935 271247
rect 116847 271175 116935 271213
rect 116847 271141 116853 271175
rect 116887 271141 116935 271175
rect 116847 271103 116935 271141
rect 116847 271069 116853 271103
rect 116887 271069 116935 271103
rect 116847 271031 116935 271069
rect 116847 270997 116853 271031
rect 116887 270997 116935 271031
rect 116847 270959 116935 270997
rect 116847 270925 116853 270959
rect 116887 270925 116935 270959
rect 116847 270887 116935 270925
rect 116847 270853 116853 270887
rect 116887 270853 116935 270887
rect 116847 270824 116935 270853
rect 116987 271895 117075 271924
rect 116987 271861 117035 271895
rect 117069 271861 117075 271895
rect 116987 271823 117075 271861
rect 116987 271789 117035 271823
rect 117069 271789 117075 271823
rect 116987 271751 117075 271789
rect 116987 271717 117035 271751
rect 117069 271717 117075 271751
rect 116987 271679 117075 271717
rect 116987 271645 117035 271679
rect 117069 271645 117075 271679
rect 116987 271607 117075 271645
rect 116987 271573 117035 271607
rect 117069 271573 117075 271607
rect 116987 271535 117075 271573
rect 116987 271501 117035 271535
rect 117069 271501 117075 271535
rect 116987 271463 117075 271501
rect 116987 271429 117035 271463
rect 117069 271429 117075 271463
rect 116987 271391 117075 271429
rect 116987 271357 117035 271391
rect 117069 271357 117075 271391
rect 116987 271319 117075 271357
rect 116987 271285 117035 271319
rect 117069 271285 117075 271319
rect 116987 271247 117075 271285
rect 116987 271213 117035 271247
rect 117069 271213 117075 271247
rect 116987 271175 117075 271213
rect 116987 271141 117035 271175
rect 117069 271141 117075 271175
rect 116987 271103 117075 271141
rect 116987 271069 117035 271103
rect 117069 271069 117075 271103
rect 116987 271031 117075 271069
rect 116987 270997 117035 271031
rect 117069 270997 117075 271031
rect 116987 270959 117075 270997
rect 116987 270925 117035 270959
rect 117069 270925 117075 270959
rect 116987 270887 117075 270925
rect 116987 270853 117035 270887
rect 117069 270853 117075 270887
rect 116987 270824 117075 270853
rect 117247 271895 117335 271924
rect 117247 271861 117253 271895
rect 117287 271861 117335 271895
rect 117247 271823 117335 271861
rect 117247 271789 117253 271823
rect 117287 271789 117335 271823
rect 117247 271751 117335 271789
rect 117247 271717 117253 271751
rect 117287 271717 117335 271751
rect 117247 271679 117335 271717
rect 117247 271645 117253 271679
rect 117287 271645 117335 271679
rect 117247 271607 117335 271645
rect 117247 271573 117253 271607
rect 117287 271573 117335 271607
rect 117247 271535 117335 271573
rect 117247 271501 117253 271535
rect 117287 271501 117335 271535
rect 117247 271463 117335 271501
rect 117247 271429 117253 271463
rect 117287 271429 117335 271463
rect 117247 271391 117335 271429
rect 117247 271357 117253 271391
rect 117287 271357 117335 271391
rect 117247 271319 117335 271357
rect 117247 271285 117253 271319
rect 117287 271285 117335 271319
rect 117247 271247 117335 271285
rect 117247 271213 117253 271247
rect 117287 271213 117335 271247
rect 117247 271175 117335 271213
rect 117247 271141 117253 271175
rect 117287 271141 117335 271175
rect 117247 271103 117335 271141
rect 117247 271069 117253 271103
rect 117287 271069 117335 271103
rect 117247 271031 117335 271069
rect 117247 270997 117253 271031
rect 117287 270997 117335 271031
rect 117247 270959 117335 270997
rect 117247 270925 117253 270959
rect 117287 270925 117335 270959
rect 117247 270887 117335 270925
rect 117247 270853 117253 270887
rect 117287 270853 117335 270887
rect 117247 270824 117335 270853
rect 117387 271895 117475 271924
rect 117387 271861 117435 271895
rect 117469 271861 117475 271895
rect 117387 271823 117475 271861
rect 117387 271789 117435 271823
rect 117469 271789 117475 271823
rect 117387 271751 117475 271789
rect 117387 271717 117435 271751
rect 117469 271717 117475 271751
rect 117387 271679 117475 271717
rect 117387 271645 117435 271679
rect 117469 271645 117475 271679
rect 117387 271607 117475 271645
rect 117387 271573 117435 271607
rect 117469 271573 117475 271607
rect 117387 271535 117475 271573
rect 117387 271501 117435 271535
rect 117469 271501 117475 271535
rect 117387 271463 117475 271501
rect 117387 271429 117435 271463
rect 117469 271429 117475 271463
rect 117387 271391 117475 271429
rect 117387 271357 117435 271391
rect 117469 271357 117475 271391
rect 117387 271319 117475 271357
rect 117387 271285 117435 271319
rect 117469 271285 117475 271319
rect 117387 271247 117475 271285
rect 117387 271213 117435 271247
rect 117469 271213 117475 271247
rect 117387 271175 117475 271213
rect 117387 271141 117435 271175
rect 117469 271141 117475 271175
rect 117387 271103 117475 271141
rect 117387 271069 117435 271103
rect 117469 271069 117475 271103
rect 117387 271031 117475 271069
rect 117387 270997 117435 271031
rect 117469 270997 117475 271031
rect 117387 270959 117475 270997
rect 117387 270925 117435 270959
rect 117469 270925 117475 270959
rect 117387 270887 117475 270925
rect 117387 270853 117435 270887
rect 117469 270853 117475 270887
rect 117387 270824 117475 270853
rect 117647 271895 117735 271924
rect 117647 271861 117653 271895
rect 117687 271861 117735 271895
rect 117647 271823 117735 271861
rect 117647 271789 117653 271823
rect 117687 271789 117735 271823
rect 117647 271751 117735 271789
rect 117647 271717 117653 271751
rect 117687 271717 117735 271751
rect 117647 271679 117735 271717
rect 117647 271645 117653 271679
rect 117687 271645 117735 271679
rect 117647 271607 117735 271645
rect 117647 271573 117653 271607
rect 117687 271573 117735 271607
rect 117647 271535 117735 271573
rect 117647 271501 117653 271535
rect 117687 271501 117735 271535
rect 117647 271463 117735 271501
rect 117647 271429 117653 271463
rect 117687 271429 117735 271463
rect 117647 271391 117735 271429
rect 117647 271357 117653 271391
rect 117687 271357 117735 271391
rect 117647 271319 117735 271357
rect 117647 271285 117653 271319
rect 117687 271285 117735 271319
rect 117647 271247 117735 271285
rect 117647 271213 117653 271247
rect 117687 271213 117735 271247
rect 117647 271175 117735 271213
rect 117647 271141 117653 271175
rect 117687 271141 117735 271175
rect 117647 271103 117735 271141
rect 117647 271069 117653 271103
rect 117687 271069 117735 271103
rect 117647 271031 117735 271069
rect 117647 270997 117653 271031
rect 117687 270997 117735 271031
rect 117647 270959 117735 270997
rect 117647 270925 117653 270959
rect 117687 270925 117735 270959
rect 117647 270887 117735 270925
rect 117647 270853 117653 270887
rect 117687 270853 117735 270887
rect 117647 270824 117735 270853
rect 117787 271895 117875 271924
rect 117787 271861 117835 271895
rect 117869 271861 117875 271895
rect 117787 271823 117875 271861
rect 117787 271789 117835 271823
rect 117869 271789 117875 271823
rect 117787 271751 117875 271789
rect 117787 271717 117835 271751
rect 117869 271717 117875 271751
rect 117787 271679 117875 271717
rect 117787 271645 117835 271679
rect 117869 271645 117875 271679
rect 117787 271607 117875 271645
rect 117787 271573 117835 271607
rect 117869 271573 117875 271607
rect 117787 271535 117875 271573
rect 117787 271501 117835 271535
rect 117869 271501 117875 271535
rect 117787 271463 117875 271501
rect 117787 271429 117835 271463
rect 117869 271429 117875 271463
rect 117787 271391 117875 271429
rect 117787 271357 117835 271391
rect 117869 271357 117875 271391
rect 117787 271319 117875 271357
rect 117787 271285 117835 271319
rect 117869 271285 117875 271319
rect 117787 271247 117875 271285
rect 117787 271213 117835 271247
rect 117869 271213 117875 271247
rect 117787 271175 117875 271213
rect 117787 271141 117835 271175
rect 117869 271141 117875 271175
rect 117787 271103 117875 271141
rect 117787 271069 117835 271103
rect 117869 271069 117875 271103
rect 117787 271031 117875 271069
rect 117787 270997 117835 271031
rect 117869 270997 117875 271031
rect 117787 270959 117875 270997
rect 117787 270925 117835 270959
rect 117869 270925 117875 270959
rect 117787 270887 117875 270925
rect 117787 270853 117835 270887
rect 117869 270853 117875 270887
rect 117787 270824 117875 270853
rect 118047 271895 118135 271924
rect 118047 271861 118053 271895
rect 118087 271861 118135 271895
rect 118047 271823 118135 271861
rect 118047 271789 118053 271823
rect 118087 271789 118135 271823
rect 118047 271751 118135 271789
rect 118047 271717 118053 271751
rect 118087 271717 118135 271751
rect 118047 271679 118135 271717
rect 118047 271645 118053 271679
rect 118087 271645 118135 271679
rect 118047 271607 118135 271645
rect 118047 271573 118053 271607
rect 118087 271573 118135 271607
rect 118047 271535 118135 271573
rect 118047 271501 118053 271535
rect 118087 271501 118135 271535
rect 118047 271463 118135 271501
rect 118047 271429 118053 271463
rect 118087 271429 118135 271463
rect 118047 271391 118135 271429
rect 118047 271357 118053 271391
rect 118087 271357 118135 271391
rect 118047 271319 118135 271357
rect 118047 271285 118053 271319
rect 118087 271285 118135 271319
rect 118047 271247 118135 271285
rect 118047 271213 118053 271247
rect 118087 271213 118135 271247
rect 118047 271175 118135 271213
rect 118047 271141 118053 271175
rect 118087 271141 118135 271175
rect 118047 271103 118135 271141
rect 118047 271069 118053 271103
rect 118087 271069 118135 271103
rect 118047 271031 118135 271069
rect 118047 270997 118053 271031
rect 118087 270997 118135 271031
rect 118047 270959 118135 270997
rect 118047 270925 118053 270959
rect 118087 270925 118135 270959
rect 118047 270887 118135 270925
rect 118047 270853 118053 270887
rect 118087 270853 118135 270887
rect 118047 270824 118135 270853
rect 118187 271895 118275 271924
rect 118187 271861 118235 271895
rect 118269 271861 118275 271895
rect 118187 271823 118275 271861
rect 118187 271789 118235 271823
rect 118269 271789 118275 271823
rect 118187 271751 118275 271789
rect 118187 271717 118235 271751
rect 118269 271717 118275 271751
rect 118187 271679 118275 271717
rect 118187 271645 118235 271679
rect 118269 271645 118275 271679
rect 118187 271607 118275 271645
rect 118187 271573 118235 271607
rect 118269 271573 118275 271607
rect 118187 271535 118275 271573
rect 118187 271501 118235 271535
rect 118269 271501 118275 271535
rect 118187 271463 118275 271501
rect 118187 271429 118235 271463
rect 118269 271429 118275 271463
rect 118187 271391 118275 271429
rect 118187 271357 118235 271391
rect 118269 271357 118275 271391
rect 118187 271319 118275 271357
rect 118187 271285 118235 271319
rect 118269 271285 118275 271319
rect 118187 271247 118275 271285
rect 118187 271213 118235 271247
rect 118269 271213 118275 271247
rect 118187 271175 118275 271213
rect 118187 271141 118235 271175
rect 118269 271141 118275 271175
rect 118187 271103 118275 271141
rect 118187 271069 118235 271103
rect 118269 271069 118275 271103
rect 118187 271031 118275 271069
rect 118187 270997 118235 271031
rect 118269 270997 118275 271031
rect 118187 270959 118275 270997
rect 118187 270925 118235 270959
rect 118269 270925 118275 270959
rect 118187 270887 118275 270925
rect 118187 270853 118235 270887
rect 118269 270853 118275 270887
rect 118187 270824 118275 270853
rect 118447 271895 118535 271924
rect 118447 271861 118453 271895
rect 118487 271861 118535 271895
rect 118447 271823 118535 271861
rect 118447 271789 118453 271823
rect 118487 271789 118535 271823
rect 118447 271751 118535 271789
rect 118447 271717 118453 271751
rect 118487 271717 118535 271751
rect 118447 271679 118535 271717
rect 118447 271645 118453 271679
rect 118487 271645 118535 271679
rect 118447 271607 118535 271645
rect 118447 271573 118453 271607
rect 118487 271573 118535 271607
rect 118447 271535 118535 271573
rect 118447 271501 118453 271535
rect 118487 271501 118535 271535
rect 118447 271463 118535 271501
rect 118447 271429 118453 271463
rect 118487 271429 118535 271463
rect 118447 271391 118535 271429
rect 118447 271357 118453 271391
rect 118487 271357 118535 271391
rect 118447 271319 118535 271357
rect 118447 271285 118453 271319
rect 118487 271285 118535 271319
rect 118447 271247 118535 271285
rect 118447 271213 118453 271247
rect 118487 271213 118535 271247
rect 118447 271175 118535 271213
rect 118447 271141 118453 271175
rect 118487 271141 118535 271175
rect 118447 271103 118535 271141
rect 118447 271069 118453 271103
rect 118487 271069 118535 271103
rect 118447 271031 118535 271069
rect 118447 270997 118453 271031
rect 118487 270997 118535 271031
rect 118447 270959 118535 270997
rect 118447 270925 118453 270959
rect 118487 270925 118535 270959
rect 118447 270887 118535 270925
rect 118447 270853 118453 270887
rect 118487 270853 118535 270887
rect 118447 270824 118535 270853
rect 118587 271895 118675 271924
rect 118587 271861 118635 271895
rect 118669 271861 118675 271895
rect 118587 271823 118675 271861
rect 118587 271789 118635 271823
rect 118669 271789 118675 271823
rect 118587 271751 118675 271789
rect 118587 271717 118635 271751
rect 118669 271717 118675 271751
rect 118587 271679 118675 271717
rect 118587 271645 118635 271679
rect 118669 271645 118675 271679
rect 118587 271607 118675 271645
rect 118587 271573 118635 271607
rect 118669 271573 118675 271607
rect 118587 271535 118675 271573
rect 118587 271501 118635 271535
rect 118669 271501 118675 271535
rect 118587 271463 118675 271501
rect 118587 271429 118635 271463
rect 118669 271429 118675 271463
rect 118587 271391 118675 271429
rect 118587 271357 118635 271391
rect 118669 271357 118675 271391
rect 118587 271319 118675 271357
rect 118587 271285 118635 271319
rect 118669 271285 118675 271319
rect 118587 271247 118675 271285
rect 118587 271213 118635 271247
rect 118669 271213 118675 271247
rect 118587 271175 118675 271213
rect 118587 271141 118635 271175
rect 118669 271141 118675 271175
rect 118587 271103 118675 271141
rect 118587 271069 118635 271103
rect 118669 271069 118675 271103
rect 118587 271031 118675 271069
rect 118587 270997 118635 271031
rect 118669 270997 118675 271031
rect 118587 270959 118675 270997
rect 118587 270925 118635 270959
rect 118669 270925 118675 270959
rect 118587 270887 118675 270925
rect 118587 270853 118635 270887
rect 118669 270853 118675 270887
rect 118587 270824 118675 270853
rect 118847 271895 118935 271924
rect 120377 271913 120423 271930
rect 120835 272396 120881 272413
rect 120835 272362 120841 272396
rect 120875 272362 120881 272396
rect 120835 272324 120881 272362
rect 120835 272290 120841 272324
rect 120875 272290 120881 272324
rect 120835 272252 120881 272290
rect 120835 272218 120841 272252
rect 120875 272224 120881 272252
rect 120953 272224 121018 272737
rect 121077 272858 121083 272881
rect 121117 272858 121123 272892
rect 121077 272820 121123 272858
rect 121077 272786 121083 272820
rect 121117 272786 121123 272820
rect 121077 272748 121123 272786
rect 121077 272714 121083 272748
rect 121117 272714 121123 272748
rect 121077 272697 121123 272714
rect 121535 273180 121624 273197
rect 121535 273146 121541 273180
rect 121575 273146 121624 273180
rect 121535 273108 121624 273146
rect 121535 273074 121541 273108
rect 121575 273074 121624 273108
rect 121535 273036 121624 273074
rect 121535 273002 121541 273036
rect 121575 273002 121624 273036
rect 121535 272964 121624 273002
rect 121535 272930 121541 272964
rect 121575 272930 121624 272964
rect 121535 272892 121624 272930
rect 121535 272858 121541 272892
rect 121575 272858 121624 272892
rect 121535 272820 121624 272858
rect 121535 272786 121541 272820
rect 121575 272786 121624 272820
rect 121535 272748 121624 272786
rect 121535 272714 121541 272748
rect 121575 272714 121624 272748
rect 121535 272697 121624 272714
rect 121133 272650 121525 272656
rect 121133 272616 121168 272650
rect 121202 272616 121240 272650
rect 121274 272616 121312 272650
rect 121346 272616 121384 272650
rect 121418 272616 121456 272650
rect 121490 272616 121525 272650
rect 121133 272494 121525 272616
rect 121133 272460 121168 272494
rect 121202 272460 121240 272494
rect 121274 272460 121312 272494
rect 121346 272460 121384 272494
rect 121418 272460 121456 272494
rect 121490 272460 121525 272494
rect 121133 272454 121525 272460
rect 121581 272413 121624 272697
rect 121796 273059 123438 273127
rect 121077 272396 121123 272413
rect 121077 272362 121083 272396
rect 121117 272362 121123 272396
rect 121077 272324 121123 272362
rect 121077 272290 121083 272324
rect 121117 272290 121123 272324
rect 121077 272252 121123 272290
rect 121077 272224 121083 272252
rect 120875 272218 121083 272224
rect 121117 272218 121123 272252
rect 120835 272180 121123 272218
rect 120835 272146 120841 272180
rect 120875 272146 121083 272180
rect 121117 272146 121123 272180
rect 120835 272108 121123 272146
rect 120835 272074 120841 272108
rect 120875 272097 121083 272108
rect 120875 272074 120881 272097
rect 120835 272036 120881 272074
rect 120835 272002 120841 272036
rect 120875 272002 120881 272036
rect 120835 271964 120881 272002
rect 120835 271930 120841 271964
rect 120875 271930 120881 271964
rect 120835 271913 120881 271930
rect 118847 271861 118853 271895
rect 118887 271861 118935 271895
rect 118847 271823 118935 271861
rect 118847 271789 118853 271823
rect 118887 271789 118935 271823
rect 118847 271751 118935 271789
rect 118847 271717 118853 271751
rect 118887 271717 118935 271751
rect 118847 271679 118935 271717
rect 118847 271645 118853 271679
rect 118887 271645 118935 271679
rect 120433 271866 120825 271872
rect 120433 271832 120468 271866
rect 120502 271832 120540 271866
rect 120574 271832 120612 271866
rect 120646 271832 120684 271866
rect 120718 271832 120756 271866
rect 120790 271832 120825 271866
rect 120433 271710 120825 271832
rect 120433 271676 120468 271710
rect 120502 271676 120540 271710
rect 120574 271676 120612 271710
rect 120646 271676 120684 271710
rect 120718 271676 120756 271710
rect 120790 271676 120825 271710
rect 120433 271670 120825 271676
rect 118847 271607 118935 271645
rect 118847 271573 118853 271607
rect 118887 271573 118935 271607
rect 118847 271535 118935 271573
rect 118847 271501 118853 271535
rect 118887 271501 118935 271535
rect 118847 271463 118935 271501
rect 118847 271429 118853 271463
rect 118887 271429 118935 271463
rect 118847 271391 118935 271429
rect 118847 271357 118853 271391
rect 118887 271357 118935 271391
rect 118847 271319 118935 271357
rect 118847 271285 118853 271319
rect 118887 271285 118935 271319
rect 118847 271247 118935 271285
rect 118847 271213 118853 271247
rect 118887 271213 118935 271247
rect 118847 271175 118935 271213
rect 118847 271141 118853 271175
rect 118887 271141 118935 271175
rect 118847 271103 118935 271141
rect 120377 271612 120423 271629
rect 120377 271578 120383 271612
rect 120417 271578 120423 271612
rect 120377 271540 120423 271578
rect 120377 271506 120383 271540
rect 120417 271506 120423 271540
rect 120377 271468 120423 271506
rect 120377 271434 120383 271468
rect 120417 271434 120423 271468
rect 120377 271396 120423 271434
rect 120377 271362 120383 271396
rect 120417 271362 120423 271396
rect 120377 271324 120423 271362
rect 120377 271290 120383 271324
rect 120417 271290 120423 271324
rect 120377 271252 120423 271290
rect 120377 271218 120383 271252
rect 120417 271218 120423 271252
rect 120377 271180 120423 271218
rect 120377 271146 120383 271180
rect 120417 271146 120423 271180
rect 120377 271129 120423 271146
rect 120835 271612 120881 271629
rect 120835 271578 120841 271612
rect 120875 271578 120881 271612
rect 120835 271540 120881 271578
rect 120835 271506 120841 271540
rect 120875 271506 120881 271540
rect 120835 271468 120881 271506
rect 120835 271434 120841 271468
rect 120875 271440 120881 271468
rect 120953 271440 121018 272097
rect 121077 272074 121083 272097
rect 121117 272074 121123 272108
rect 121077 272036 121123 272074
rect 121077 272002 121083 272036
rect 121117 272002 121123 272036
rect 121077 271964 121123 272002
rect 121077 271930 121083 271964
rect 121117 271930 121123 271964
rect 121077 271913 121123 271930
rect 121535 272396 121677 272413
rect 121535 272362 121541 272396
rect 121575 272362 121677 272396
rect 121535 272338 121677 272362
rect 121535 272324 121605 272338
rect 121535 272290 121541 272324
rect 121575 272290 121605 272324
rect 121535 272286 121605 272290
rect 121657 272286 121677 272338
rect 121535 272274 121677 272286
rect 121535 272252 121605 272274
rect 121535 272218 121541 272252
rect 121575 272222 121605 272252
rect 121657 272222 121677 272274
rect 121575 272218 121677 272222
rect 121535 272210 121677 272218
rect 121535 272180 121605 272210
rect 121535 272146 121541 272180
rect 121575 272158 121605 272180
rect 121657 272158 121677 272210
rect 121575 272146 121677 272158
rect 121535 272108 121605 272146
rect 121535 272074 121541 272108
rect 121575 272094 121605 272108
rect 121657 272094 121677 272146
rect 121575 272082 121677 272094
rect 121575 272074 121605 272082
rect 121535 272036 121605 272074
rect 121535 272002 121541 272036
rect 121575 272030 121605 272036
rect 121657 272030 121677 272082
rect 121575 272018 121677 272030
rect 121575 272002 121605 272018
rect 121535 271966 121605 272002
rect 121657 271966 121677 272018
rect 121535 271964 121677 271966
rect 121535 271930 121541 271964
rect 121575 271954 121677 271964
rect 121575 271930 121605 271954
rect 121535 271913 121605 271930
rect 121581 271902 121605 271913
rect 121657 271902 121677 271954
rect 121581 271890 121677 271902
rect 121133 271866 121525 271872
rect 121133 271832 121168 271866
rect 121202 271832 121240 271866
rect 121274 271832 121312 271866
rect 121346 271832 121384 271866
rect 121418 271832 121456 271866
rect 121490 271832 121525 271866
rect 121133 271710 121525 271832
rect 121133 271676 121168 271710
rect 121202 271676 121240 271710
rect 121274 271676 121312 271710
rect 121346 271676 121384 271710
rect 121418 271676 121456 271710
rect 121490 271676 121525 271710
rect 121133 271670 121525 271676
rect 121581 271838 121605 271890
rect 121657 271838 121677 271890
rect 121581 271826 121677 271838
rect 121581 271774 121605 271826
rect 121657 271774 121677 271826
rect 121581 271762 121677 271774
rect 121581 271710 121605 271762
rect 121657 271710 121677 271762
rect 121581 271698 121677 271710
rect 121581 271646 121605 271698
rect 121657 271646 121677 271698
rect 121581 271634 121677 271646
rect 121581 271629 121605 271634
rect 121077 271612 121123 271629
rect 121077 271578 121083 271612
rect 121117 271578 121123 271612
rect 121077 271540 121123 271578
rect 121077 271506 121083 271540
rect 121117 271506 121123 271540
rect 121077 271468 121123 271506
rect 121077 271440 121083 271468
rect 120875 271434 121083 271440
rect 121117 271434 121123 271468
rect 120835 271396 121123 271434
rect 120835 271362 120841 271396
rect 120875 271362 121083 271396
rect 121117 271362 121123 271396
rect 120835 271324 121123 271362
rect 120835 271290 120841 271324
rect 120875 271313 121083 271324
rect 120875 271290 120881 271313
rect 120835 271252 120881 271290
rect 120835 271218 120841 271252
rect 120875 271218 120881 271252
rect 120835 271180 120881 271218
rect 120835 271146 120841 271180
rect 120875 271146 120881 271180
rect 120835 271129 120881 271146
rect 118847 271069 118853 271103
rect 118887 271069 118935 271103
rect 118847 271031 118935 271069
rect 118847 270997 118853 271031
rect 118887 270997 118935 271031
rect 118847 270959 118935 270997
rect 118847 270925 118853 270959
rect 118887 270925 118935 270959
rect 118847 270887 118935 270925
rect 118847 270853 118853 270887
rect 118887 270853 118935 270887
rect 120433 271082 120825 271088
rect 120433 271048 120468 271082
rect 120502 271048 120540 271082
rect 120574 271048 120612 271082
rect 120646 271048 120684 271082
rect 120718 271048 120756 271082
rect 120790 271048 120825 271082
rect 120433 270926 120825 271048
rect 120433 270892 120468 270926
rect 120502 270892 120540 270926
rect 120574 270892 120612 270926
rect 120646 270892 120684 270926
rect 120718 270892 120756 270926
rect 120790 270892 120825 270926
rect 120433 270886 120825 270892
rect 118847 270824 118935 270853
rect 115885 270786 116037 270792
rect 115885 270752 115908 270786
rect 115942 270752 115980 270786
rect 116014 270752 116037 270786
rect 115885 270746 116037 270752
rect 114050 270641 114976 270657
rect 114050 270607 114096 270641
rect 114130 270607 114168 270641
rect 114202 270607 114240 270641
rect 114274 270607 114312 270641
rect 114346 270607 114384 270641
rect 114418 270607 114456 270641
rect 114490 270617 114976 270641
rect 116093 270621 116135 270824
rect 116285 270786 116437 270792
rect 116285 270752 116308 270786
rect 116342 270752 116380 270786
rect 116414 270752 116437 270786
rect 116285 270746 116437 270752
rect 116493 270621 116535 270824
rect 116685 270786 116837 270792
rect 116685 270752 116708 270786
rect 116742 270752 116780 270786
rect 116814 270752 116837 270786
rect 116685 270746 116837 270752
rect 116893 270621 116935 270824
rect 117085 270786 117237 270792
rect 117085 270752 117108 270786
rect 117142 270752 117180 270786
rect 117214 270752 117237 270786
rect 117085 270746 117237 270752
rect 117293 270621 117335 270824
rect 117485 270786 117637 270792
rect 117485 270752 117508 270786
rect 117542 270752 117580 270786
rect 117614 270752 117637 270786
rect 117485 270746 117637 270752
rect 117693 270621 117735 270824
rect 117885 270786 118037 270792
rect 117885 270752 117908 270786
rect 117942 270752 117980 270786
rect 118014 270752 118037 270786
rect 117885 270746 118037 270752
rect 118093 270621 118135 270824
rect 118285 270786 118437 270792
rect 118285 270752 118308 270786
rect 118342 270752 118380 270786
rect 118414 270752 118437 270786
rect 118285 270746 118437 270752
rect 118493 270621 118535 270824
rect 118685 270786 118837 270792
rect 118685 270752 118708 270786
rect 118742 270752 118780 270786
rect 118814 270752 118837 270786
rect 118685 270746 118837 270752
rect 118893 270621 118935 270824
rect 116093 270617 118935 270621
rect 114490 270607 118935 270617
rect 114050 270588 118935 270607
rect 120377 270828 120423 270845
rect 120377 270794 120383 270828
rect 120417 270794 120423 270828
rect 120377 270756 120423 270794
rect 120377 270722 120383 270756
rect 120417 270722 120423 270756
rect 120377 270684 120423 270722
rect 120377 270650 120383 270684
rect 120417 270650 120423 270684
rect 120377 270612 120423 270650
rect 114050 270587 116771 270588
rect 114050 270586 114877 270587
rect 114050 270545 114542 270586
rect 120377 270578 120383 270612
rect 120417 270578 120423 270612
rect 112194 270429 113508 270468
rect 120377 270540 120423 270578
rect 120377 270506 120383 270540
rect 120417 270506 120423 270540
rect 120377 270468 120423 270506
rect 120377 270434 120383 270468
rect 120417 270434 120423 270468
rect 112194 270399 118508 270429
rect 112466 270396 118508 270399
rect 112466 270224 112508 270396
rect 112564 270296 112716 270302
rect 112564 270262 112587 270296
rect 112621 270262 112659 270296
rect 112693 270262 112716 270296
rect 112564 270256 112716 270262
rect 112866 270224 112908 270396
rect 112964 270296 113116 270302
rect 112964 270262 112987 270296
rect 113021 270262 113059 270296
rect 113093 270262 113116 270296
rect 112964 270256 113116 270262
rect 113266 270224 113308 270396
rect 113364 270296 113516 270302
rect 113364 270262 113387 270296
rect 113421 270262 113459 270296
rect 113493 270262 113516 270296
rect 113364 270256 113516 270262
rect 113666 270224 113708 270396
rect 113764 270296 113916 270302
rect 113764 270262 113787 270296
rect 113821 270262 113859 270296
rect 113893 270262 113916 270296
rect 113764 270256 113916 270262
rect 114066 270224 114108 270396
rect 114164 270296 114316 270302
rect 114164 270262 114187 270296
rect 114221 270262 114259 270296
rect 114293 270262 114316 270296
rect 114164 270256 114316 270262
rect 114466 270224 114508 270396
rect 114564 270296 114716 270302
rect 114564 270262 114587 270296
rect 114621 270262 114659 270296
rect 114693 270262 114716 270296
rect 114564 270256 114716 270262
rect 114866 270224 114908 270396
rect 114964 270296 115116 270302
rect 114964 270262 114987 270296
rect 115021 270262 115059 270296
rect 115093 270262 115116 270296
rect 114964 270256 115116 270262
rect 115266 270224 115308 270396
rect 115364 270296 115516 270302
rect 115364 270262 115387 270296
rect 115421 270262 115459 270296
rect 115493 270262 115516 270296
rect 115364 270256 115516 270262
rect 115666 270224 115708 270396
rect 115764 270296 115916 270302
rect 115764 270262 115787 270296
rect 115821 270262 115859 270296
rect 115893 270262 115916 270296
rect 115764 270256 115916 270262
rect 116066 270224 116108 270396
rect 116164 270296 116316 270302
rect 116164 270262 116187 270296
rect 116221 270262 116259 270296
rect 116293 270262 116316 270296
rect 116164 270256 116316 270262
rect 116466 270224 116508 270396
rect 116564 270296 116716 270302
rect 116564 270262 116587 270296
rect 116621 270262 116659 270296
rect 116693 270262 116716 270296
rect 116564 270256 116716 270262
rect 116866 270224 116908 270396
rect 116964 270296 117116 270302
rect 116964 270262 116987 270296
rect 117021 270262 117059 270296
rect 117093 270262 117116 270296
rect 116964 270256 117116 270262
rect 117266 270224 117308 270396
rect 117364 270296 117516 270302
rect 117364 270262 117387 270296
rect 117421 270262 117459 270296
rect 117493 270262 117516 270296
rect 117364 270256 117516 270262
rect 117666 270224 117708 270396
rect 117764 270296 117916 270302
rect 117764 270262 117787 270296
rect 117821 270262 117859 270296
rect 117893 270262 117916 270296
rect 117764 270256 117916 270262
rect 118066 270224 118108 270396
rect 118164 270296 118316 270302
rect 118164 270262 118187 270296
rect 118221 270262 118259 270296
rect 118293 270262 118316 270296
rect 118164 270256 118316 270262
rect 118466 270224 118508 270396
rect 120377 270396 120423 270434
rect 120377 270362 120383 270396
rect 120417 270362 120423 270396
rect 120377 270345 120423 270362
rect 120835 270828 120881 270845
rect 120835 270794 120841 270828
rect 120875 270794 120881 270828
rect 120835 270756 120881 270794
rect 120835 270722 120841 270756
rect 120875 270722 120881 270756
rect 120835 270684 120881 270722
rect 120835 270650 120841 270684
rect 120875 270656 120881 270684
rect 120953 270656 121018 271313
rect 121077 271290 121083 271313
rect 121117 271290 121123 271324
rect 121077 271252 121123 271290
rect 121077 271218 121083 271252
rect 121117 271218 121123 271252
rect 121077 271180 121123 271218
rect 121077 271146 121083 271180
rect 121117 271146 121123 271180
rect 121077 271129 121123 271146
rect 121535 271612 121605 271629
rect 121535 271578 121541 271612
rect 121575 271582 121605 271612
rect 121657 271582 121677 271634
rect 121575 271578 121677 271582
rect 121535 271570 121677 271578
rect 121535 271540 121605 271570
rect 121535 271506 121541 271540
rect 121575 271518 121605 271540
rect 121657 271518 121677 271570
rect 121575 271506 121677 271518
rect 121535 271468 121605 271506
rect 121535 271434 121541 271468
rect 121575 271454 121605 271468
rect 121657 271454 121677 271506
rect 121575 271442 121677 271454
rect 121575 271434 121605 271442
rect 121535 271396 121605 271434
rect 121535 271362 121541 271396
rect 121575 271390 121605 271396
rect 121657 271390 121677 271442
rect 121575 271378 121677 271390
rect 121575 271362 121605 271378
rect 121535 271326 121605 271362
rect 121657 271326 121677 271378
rect 121535 271324 121677 271326
rect 121535 271290 121541 271324
rect 121575 271314 121677 271324
rect 121575 271290 121605 271314
rect 121535 271262 121605 271290
rect 121657 271262 121677 271314
rect 121535 271252 121677 271262
rect 121535 271218 121541 271252
rect 121575 271250 121677 271252
rect 121575 271218 121605 271250
rect 121535 271198 121605 271218
rect 121657 271198 121677 271250
rect 121535 271186 121677 271198
rect 121535 271180 121605 271186
rect 121535 271146 121541 271180
rect 121575 271146 121605 271180
rect 121535 271134 121605 271146
rect 121657 271134 121677 271186
rect 121535 271129 121677 271134
rect 121581 271122 121677 271129
rect 121133 271082 121525 271088
rect 121133 271048 121168 271082
rect 121202 271048 121240 271082
rect 121274 271048 121312 271082
rect 121346 271048 121384 271082
rect 121418 271048 121456 271082
rect 121490 271048 121525 271082
rect 121133 270926 121525 271048
rect 121133 270892 121168 270926
rect 121202 270892 121240 270926
rect 121274 270892 121312 270926
rect 121346 270892 121384 270926
rect 121418 270892 121456 270926
rect 121490 270892 121525 270926
rect 121133 270886 121525 270892
rect 121581 271070 121605 271122
rect 121657 271070 121677 271122
rect 121581 271058 121677 271070
rect 121581 271006 121605 271058
rect 121657 271006 121677 271058
rect 121581 270994 121677 271006
rect 121581 270942 121605 270994
rect 121657 270942 121677 270994
rect 121581 270930 121677 270942
rect 121581 270878 121605 270930
rect 121657 270878 121677 270930
rect 121581 270866 121677 270878
rect 121581 270845 121605 270866
rect 121077 270828 121123 270845
rect 121077 270794 121083 270828
rect 121117 270794 121123 270828
rect 121077 270756 121123 270794
rect 121077 270722 121083 270756
rect 121117 270722 121123 270756
rect 121077 270684 121123 270722
rect 121077 270656 121083 270684
rect 120875 270650 121083 270656
rect 121117 270650 121123 270684
rect 120835 270612 121123 270650
rect 120835 270578 120841 270612
rect 120875 270578 121083 270612
rect 121117 270578 121123 270612
rect 120835 270540 121123 270578
rect 120835 270506 120841 270540
rect 120875 270529 121083 270540
rect 120875 270506 120881 270529
rect 120835 270468 120881 270506
rect 120835 270434 120841 270468
rect 120875 270434 120881 270468
rect 120835 270396 120881 270434
rect 120835 270362 120841 270396
rect 120875 270362 120881 270396
rect 120835 270345 120881 270362
rect 118564 270296 118716 270302
rect 118564 270262 118587 270296
rect 118621 270262 118659 270296
rect 118693 270262 118716 270296
rect 118564 270256 118716 270262
rect 120433 270298 120825 270304
rect 120433 270264 120468 270298
rect 120502 270264 120540 270298
rect 120574 270264 120612 270298
rect 120646 270264 120684 270298
rect 120718 270264 120756 270298
rect 120790 270264 120825 270298
rect 112466 270195 112554 270224
rect 112466 270161 112514 270195
rect 112548 270161 112554 270195
rect 112466 270123 112554 270161
rect 112466 270089 112514 270123
rect 112548 270089 112554 270123
rect 112466 270051 112554 270089
rect 112466 270017 112514 270051
rect 112548 270017 112554 270051
rect 112466 269979 112554 270017
rect 112466 269945 112514 269979
rect 112548 269945 112554 269979
rect 112466 269907 112554 269945
rect 112466 269873 112514 269907
rect 112548 269873 112554 269907
rect 112466 269835 112554 269873
rect 112466 269801 112514 269835
rect 112548 269801 112554 269835
rect 112466 269763 112554 269801
rect 112466 269729 112514 269763
rect 112548 269729 112554 269763
rect 112466 269691 112554 269729
rect 112466 269657 112514 269691
rect 112548 269657 112554 269691
rect 112466 269619 112554 269657
rect 112466 269585 112514 269619
rect 112548 269585 112554 269619
rect 112466 269547 112554 269585
rect 112466 269513 112514 269547
rect 112548 269513 112554 269547
rect 112466 269475 112554 269513
rect 112466 269441 112514 269475
rect 112548 269441 112554 269475
rect 112466 269403 112554 269441
rect 112466 269369 112514 269403
rect 112548 269369 112554 269403
rect 112466 269331 112554 269369
rect 112466 269297 112514 269331
rect 112548 269297 112554 269331
rect 112466 269259 112554 269297
rect 112466 269225 112514 269259
rect 112548 269225 112554 269259
rect 112466 269187 112554 269225
rect 112466 269153 112514 269187
rect 112548 269153 112554 269187
rect 112466 269124 112554 269153
rect 112726 270195 112814 270224
rect 112726 270161 112732 270195
rect 112766 270161 112814 270195
rect 112726 270123 112814 270161
rect 112726 270089 112732 270123
rect 112766 270089 112814 270123
rect 112726 270051 112814 270089
rect 112726 270017 112732 270051
rect 112766 270017 112814 270051
rect 112726 269979 112814 270017
rect 112726 269945 112732 269979
rect 112766 269945 112814 269979
rect 112726 269907 112814 269945
rect 112726 269873 112732 269907
rect 112766 269873 112814 269907
rect 112726 269835 112814 269873
rect 112726 269801 112732 269835
rect 112766 269801 112814 269835
rect 112726 269763 112814 269801
rect 112726 269729 112732 269763
rect 112766 269729 112814 269763
rect 112726 269691 112814 269729
rect 112726 269657 112732 269691
rect 112766 269657 112814 269691
rect 112726 269619 112814 269657
rect 112726 269585 112732 269619
rect 112766 269585 112814 269619
rect 112726 269547 112814 269585
rect 112726 269513 112732 269547
rect 112766 269513 112814 269547
rect 112726 269475 112814 269513
rect 112726 269441 112732 269475
rect 112766 269441 112814 269475
rect 112726 269403 112814 269441
rect 112726 269369 112732 269403
rect 112766 269369 112814 269403
rect 112726 269331 112814 269369
rect 112726 269297 112732 269331
rect 112766 269297 112814 269331
rect 112726 269259 112814 269297
rect 112726 269225 112732 269259
rect 112766 269225 112814 269259
rect 112726 269187 112814 269225
rect 112726 269153 112732 269187
rect 112766 269153 112814 269187
rect 112726 269124 112814 269153
rect 112866 270195 112954 270224
rect 112866 270161 112914 270195
rect 112948 270161 112954 270195
rect 112866 270123 112954 270161
rect 112866 270089 112914 270123
rect 112948 270089 112954 270123
rect 112866 270051 112954 270089
rect 112866 270017 112914 270051
rect 112948 270017 112954 270051
rect 112866 269979 112954 270017
rect 112866 269945 112914 269979
rect 112948 269945 112954 269979
rect 112866 269907 112954 269945
rect 112866 269873 112914 269907
rect 112948 269873 112954 269907
rect 112866 269835 112954 269873
rect 112866 269801 112914 269835
rect 112948 269801 112954 269835
rect 112866 269763 112954 269801
rect 112866 269729 112914 269763
rect 112948 269729 112954 269763
rect 112866 269691 112954 269729
rect 112866 269657 112914 269691
rect 112948 269657 112954 269691
rect 112866 269619 112954 269657
rect 112866 269585 112914 269619
rect 112948 269585 112954 269619
rect 112866 269547 112954 269585
rect 112866 269513 112914 269547
rect 112948 269513 112954 269547
rect 112866 269475 112954 269513
rect 112866 269441 112914 269475
rect 112948 269441 112954 269475
rect 112866 269403 112954 269441
rect 112866 269369 112914 269403
rect 112948 269369 112954 269403
rect 112866 269331 112954 269369
rect 112866 269297 112914 269331
rect 112948 269297 112954 269331
rect 112866 269259 112954 269297
rect 112866 269225 112914 269259
rect 112948 269225 112954 269259
rect 112866 269187 112954 269225
rect 112866 269153 112914 269187
rect 112948 269153 112954 269187
rect 112866 269124 112954 269153
rect 113126 270195 113214 270224
rect 113126 270161 113132 270195
rect 113166 270161 113214 270195
rect 113126 270123 113214 270161
rect 113126 270089 113132 270123
rect 113166 270089 113214 270123
rect 113126 270051 113214 270089
rect 113126 270017 113132 270051
rect 113166 270017 113214 270051
rect 113126 269979 113214 270017
rect 113126 269945 113132 269979
rect 113166 269945 113214 269979
rect 113126 269907 113214 269945
rect 113126 269873 113132 269907
rect 113166 269873 113214 269907
rect 113126 269835 113214 269873
rect 113126 269801 113132 269835
rect 113166 269801 113214 269835
rect 113126 269763 113214 269801
rect 113126 269729 113132 269763
rect 113166 269729 113214 269763
rect 113126 269691 113214 269729
rect 113126 269657 113132 269691
rect 113166 269657 113214 269691
rect 113126 269619 113214 269657
rect 113126 269585 113132 269619
rect 113166 269585 113214 269619
rect 113126 269547 113214 269585
rect 113126 269513 113132 269547
rect 113166 269513 113214 269547
rect 113126 269475 113214 269513
rect 113126 269441 113132 269475
rect 113166 269441 113214 269475
rect 113126 269403 113214 269441
rect 113126 269369 113132 269403
rect 113166 269369 113214 269403
rect 113126 269331 113214 269369
rect 113126 269297 113132 269331
rect 113166 269297 113214 269331
rect 113126 269259 113214 269297
rect 113126 269225 113132 269259
rect 113166 269225 113214 269259
rect 113126 269187 113214 269225
rect 113126 269153 113132 269187
rect 113166 269153 113214 269187
rect 113126 269124 113214 269153
rect 113266 270195 113354 270224
rect 113266 270161 113314 270195
rect 113348 270161 113354 270195
rect 113266 270123 113354 270161
rect 113266 270089 113314 270123
rect 113348 270089 113354 270123
rect 113266 270051 113354 270089
rect 113266 270017 113314 270051
rect 113348 270017 113354 270051
rect 113266 269979 113354 270017
rect 113266 269945 113314 269979
rect 113348 269945 113354 269979
rect 113266 269907 113354 269945
rect 113266 269873 113314 269907
rect 113348 269873 113354 269907
rect 113266 269835 113354 269873
rect 113266 269801 113314 269835
rect 113348 269801 113354 269835
rect 113266 269763 113354 269801
rect 113266 269729 113314 269763
rect 113348 269729 113354 269763
rect 113266 269691 113354 269729
rect 113266 269657 113314 269691
rect 113348 269657 113354 269691
rect 113266 269619 113354 269657
rect 113266 269585 113314 269619
rect 113348 269585 113354 269619
rect 113266 269547 113354 269585
rect 113266 269513 113314 269547
rect 113348 269513 113354 269547
rect 113266 269475 113354 269513
rect 113266 269441 113314 269475
rect 113348 269441 113354 269475
rect 113266 269403 113354 269441
rect 113266 269369 113314 269403
rect 113348 269369 113354 269403
rect 113266 269331 113354 269369
rect 113266 269297 113314 269331
rect 113348 269297 113354 269331
rect 113266 269259 113354 269297
rect 113266 269225 113314 269259
rect 113348 269225 113354 269259
rect 113266 269187 113354 269225
rect 113266 269153 113314 269187
rect 113348 269153 113354 269187
rect 113266 269124 113354 269153
rect 113526 270195 113614 270224
rect 113526 270161 113532 270195
rect 113566 270161 113614 270195
rect 113526 270123 113614 270161
rect 113526 270089 113532 270123
rect 113566 270089 113614 270123
rect 113526 270051 113614 270089
rect 113526 270017 113532 270051
rect 113566 270017 113614 270051
rect 113526 269979 113614 270017
rect 113526 269945 113532 269979
rect 113566 269945 113614 269979
rect 113526 269907 113614 269945
rect 113526 269873 113532 269907
rect 113566 269873 113614 269907
rect 113526 269835 113614 269873
rect 113526 269801 113532 269835
rect 113566 269801 113614 269835
rect 113526 269763 113614 269801
rect 113526 269729 113532 269763
rect 113566 269729 113614 269763
rect 113526 269691 113614 269729
rect 113526 269657 113532 269691
rect 113566 269657 113614 269691
rect 113526 269619 113614 269657
rect 113526 269585 113532 269619
rect 113566 269585 113614 269619
rect 113526 269547 113614 269585
rect 113526 269513 113532 269547
rect 113566 269513 113614 269547
rect 113526 269475 113614 269513
rect 113526 269441 113532 269475
rect 113566 269441 113614 269475
rect 113526 269403 113614 269441
rect 113526 269369 113532 269403
rect 113566 269369 113614 269403
rect 113526 269331 113614 269369
rect 113526 269297 113532 269331
rect 113566 269297 113614 269331
rect 113526 269259 113614 269297
rect 113526 269225 113532 269259
rect 113566 269225 113614 269259
rect 113526 269187 113614 269225
rect 113526 269153 113532 269187
rect 113566 269153 113614 269187
rect 113526 269124 113614 269153
rect 113666 270195 113754 270224
rect 113666 270161 113714 270195
rect 113748 270161 113754 270195
rect 113666 270123 113754 270161
rect 113666 270089 113714 270123
rect 113748 270089 113754 270123
rect 113666 270051 113754 270089
rect 113666 270017 113714 270051
rect 113748 270017 113754 270051
rect 113666 269979 113754 270017
rect 113666 269945 113714 269979
rect 113748 269945 113754 269979
rect 113666 269907 113754 269945
rect 113666 269873 113714 269907
rect 113748 269873 113754 269907
rect 113666 269835 113754 269873
rect 113666 269801 113714 269835
rect 113748 269801 113754 269835
rect 113666 269763 113754 269801
rect 113666 269729 113714 269763
rect 113748 269729 113754 269763
rect 113666 269691 113754 269729
rect 113666 269657 113714 269691
rect 113748 269657 113754 269691
rect 113666 269619 113754 269657
rect 113666 269585 113714 269619
rect 113748 269585 113754 269619
rect 113666 269547 113754 269585
rect 113666 269513 113714 269547
rect 113748 269513 113754 269547
rect 113666 269475 113754 269513
rect 113666 269441 113714 269475
rect 113748 269441 113754 269475
rect 113666 269403 113754 269441
rect 113666 269369 113714 269403
rect 113748 269369 113754 269403
rect 113666 269331 113754 269369
rect 113666 269297 113714 269331
rect 113748 269297 113754 269331
rect 113666 269259 113754 269297
rect 113666 269225 113714 269259
rect 113748 269225 113754 269259
rect 113666 269187 113754 269225
rect 113666 269153 113714 269187
rect 113748 269153 113754 269187
rect 113666 269124 113754 269153
rect 113926 270195 114014 270224
rect 113926 270161 113932 270195
rect 113966 270161 114014 270195
rect 113926 270123 114014 270161
rect 113926 270089 113932 270123
rect 113966 270089 114014 270123
rect 113926 270051 114014 270089
rect 113926 270017 113932 270051
rect 113966 270017 114014 270051
rect 113926 269979 114014 270017
rect 113926 269945 113932 269979
rect 113966 269945 114014 269979
rect 113926 269907 114014 269945
rect 113926 269873 113932 269907
rect 113966 269873 114014 269907
rect 113926 269835 114014 269873
rect 113926 269801 113932 269835
rect 113966 269801 114014 269835
rect 113926 269763 114014 269801
rect 113926 269729 113932 269763
rect 113966 269729 114014 269763
rect 113926 269691 114014 269729
rect 113926 269657 113932 269691
rect 113966 269657 114014 269691
rect 113926 269619 114014 269657
rect 113926 269585 113932 269619
rect 113966 269585 114014 269619
rect 113926 269547 114014 269585
rect 113926 269513 113932 269547
rect 113966 269513 114014 269547
rect 113926 269475 114014 269513
rect 113926 269441 113932 269475
rect 113966 269441 114014 269475
rect 113926 269403 114014 269441
rect 113926 269369 113932 269403
rect 113966 269369 114014 269403
rect 113926 269331 114014 269369
rect 113926 269297 113932 269331
rect 113966 269297 114014 269331
rect 113926 269259 114014 269297
rect 113926 269225 113932 269259
rect 113966 269225 114014 269259
rect 113926 269187 114014 269225
rect 113926 269153 113932 269187
rect 113966 269153 114014 269187
rect 113926 269124 114014 269153
rect 114066 270195 114154 270224
rect 114066 270161 114114 270195
rect 114148 270161 114154 270195
rect 114066 270123 114154 270161
rect 114066 270089 114114 270123
rect 114148 270089 114154 270123
rect 114066 270051 114154 270089
rect 114066 270017 114114 270051
rect 114148 270017 114154 270051
rect 114066 269979 114154 270017
rect 114066 269945 114114 269979
rect 114148 269945 114154 269979
rect 114066 269907 114154 269945
rect 114066 269873 114114 269907
rect 114148 269873 114154 269907
rect 114066 269835 114154 269873
rect 114066 269801 114114 269835
rect 114148 269801 114154 269835
rect 114066 269763 114154 269801
rect 114066 269729 114114 269763
rect 114148 269729 114154 269763
rect 114066 269691 114154 269729
rect 114066 269657 114114 269691
rect 114148 269657 114154 269691
rect 114066 269619 114154 269657
rect 114066 269585 114114 269619
rect 114148 269585 114154 269619
rect 114066 269547 114154 269585
rect 114066 269513 114114 269547
rect 114148 269513 114154 269547
rect 114066 269475 114154 269513
rect 114066 269441 114114 269475
rect 114148 269441 114154 269475
rect 114066 269403 114154 269441
rect 114066 269369 114114 269403
rect 114148 269369 114154 269403
rect 114066 269331 114154 269369
rect 114066 269297 114114 269331
rect 114148 269297 114154 269331
rect 114066 269259 114154 269297
rect 114066 269225 114114 269259
rect 114148 269225 114154 269259
rect 114066 269187 114154 269225
rect 114066 269153 114114 269187
rect 114148 269153 114154 269187
rect 114066 269124 114154 269153
rect 114326 270195 114414 270224
rect 114326 270161 114332 270195
rect 114366 270161 114414 270195
rect 114326 270123 114414 270161
rect 114326 270089 114332 270123
rect 114366 270089 114414 270123
rect 114326 270051 114414 270089
rect 114326 270017 114332 270051
rect 114366 270017 114414 270051
rect 114326 269979 114414 270017
rect 114326 269945 114332 269979
rect 114366 269945 114414 269979
rect 114326 269907 114414 269945
rect 114326 269873 114332 269907
rect 114366 269873 114414 269907
rect 114326 269835 114414 269873
rect 114326 269801 114332 269835
rect 114366 269801 114414 269835
rect 114326 269763 114414 269801
rect 114326 269729 114332 269763
rect 114366 269729 114414 269763
rect 114326 269691 114414 269729
rect 114326 269657 114332 269691
rect 114366 269657 114414 269691
rect 114326 269619 114414 269657
rect 114326 269585 114332 269619
rect 114366 269585 114414 269619
rect 114326 269547 114414 269585
rect 114326 269513 114332 269547
rect 114366 269513 114414 269547
rect 114326 269475 114414 269513
rect 114326 269441 114332 269475
rect 114366 269441 114414 269475
rect 114326 269403 114414 269441
rect 114326 269369 114332 269403
rect 114366 269369 114414 269403
rect 114326 269331 114414 269369
rect 114326 269297 114332 269331
rect 114366 269297 114414 269331
rect 114326 269259 114414 269297
rect 114326 269225 114332 269259
rect 114366 269225 114414 269259
rect 114326 269187 114414 269225
rect 114326 269153 114332 269187
rect 114366 269153 114414 269187
rect 114326 269124 114414 269153
rect 114466 270195 114554 270224
rect 114466 270161 114514 270195
rect 114548 270161 114554 270195
rect 114466 270123 114554 270161
rect 114466 270089 114514 270123
rect 114548 270089 114554 270123
rect 114466 270051 114554 270089
rect 114466 270017 114514 270051
rect 114548 270017 114554 270051
rect 114466 269979 114554 270017
rect 114466 269945 114514 269979
rect 114548 269945 114554 269979
rect 114466 269907 114554 269945
rect 114466 269873 114514 269907
rect 114548 269873 114554 269907
rect 114466 269835 114554 269873
rect 114466 269801 114514 269835
rect 114548 269801 114554 269835
rect 114466 269763 114554 269801
rect 114466 269729 114514 269763
rect 114548 269729 114554 269763
rect 114466 269691 114554 269729
rect 114466 269657 114514 269691
rect 114548 269657 114554 269691
rect 114466 269619 114554 269657
rect 114466 269585 114514 269619
rect 114548 269585 114554 269619
rect 114466 269547 114554 269585
rect 114466 269513 114514 269547
rect 114548 269513 114554 269547
rect 114466 269475 114554 269513
rect 114466 269441 114514 269475
rect 114548 269441 114554 269475
rect 114466 269403 114554 269441
rect 114466 269369 114514 269403
rect 114548 269369 114554 269403
rect 114466 269331 114554 269369
rect 114466 269297 114514 269331
rect 114548 269297 114554 269331
rect 114466 269259 114554 269297
rect 114466 269225 114514 269259
rect 114548 269225 114554 269259
rect 114466 269187 114554 269225
rect 114466 269153 114514 269187
rect 114548 269153 114554 269187
rect 114466 269124 114554 269153
rect 114726 270195 114814 270224
rect 114726 270161 114732 270195
rect 114766 270161 114814 270195
rect 114726 270123 114814 270161
rect 114726 270089 114732 270123
rect 114766 270089 114814 270123
rect 114726 270051 114814 270089
rect 114726 270017 114732 270051
rect 114766 270017 114814 270051
rect 114726 269979 114814 270017
rect 114726 269945 114732 269979
rect 114766 269945 114814 269979
rect 114726 269907 114814 269945
rect 114726 269873 114732 269907
rect 114766 269873 114814 269907
rect 114726 269835 114814 269873
rect 114726 269801 114732 269835
rect 114766 269801 114814 269835
rect 114726 269763 114814 269801
rect 114726 269729 114732 269763
rect 114766 269729 114814 269763
rect 114726 269691 114814 269729
rect 114726 269657 114732 269691
rect 114766 269657 114814 269691
rect 114726 269619 114814 269657
rect 114726 269585 114732 269619
rect 114766 269585 114814 269619
rect 114726 269547 114814 269585
rect 114726 269513 114732 269547
rect 114766 269513 114814 269547
rect 114726 269475 114814 269513
rect 114726 269441 114732 269475
rect 114766 269441 114814 269475
rect 114726 269403 114814 269441
rect 114726 269369 114732 269403
rect 114766 269369 114814 269403
rect 114726 269331 114814 269369
rect 114726 269297 114732 269331
rect 114766 269297 114814 269331
rect 114726 269259 114814 269297
rect 114726 269225 114732 269259
rect 114766 269225 114814 269259
rect 114726 269187 114814 269225
rect 114726 269153 114732 269187
rect 114766 269153 114814 269187
rect 114726 269124 114814 269153
rect 114866 270195 114954 270224
rect 114866 270161 114914 270195
rect 114948 270161 114954 270195
rect 114866 270123 114954 270161
rect 114866 270089 114914 270123
rect 114948 270089 114954 270123
rect 114866 270051 114954 270089
rect 114866 270017 114914 270051
rect 114948 270017 114954 270051
rect 114866 269979 114954 270017
rect 114866 269945 114914 269979
rect 114948 269945 114954 269979
rect 114866 269907 114954 269945
rect 114866 269873 114914 269907
rect 114948 269873 114954 269907
rect 114866 269835 114954 269873
rect 114866 269801 114914 269835
rect 114948 269801 114954 269835
rect 114866 269763 114954 269801
rect 114866 269729 114914 269763
rect 114948 269729 114954 269763
rect 114866 269691 114954 269729
rect 114866 269657 114914 269691
rect 114948 269657 114954 269691
rect 114866 269619 114954 269657
rect 114866 269585 114914 269619
rect 114948 269585 114954 269619
rect 114866 269547 114954 269585
rect 114866 269513 114914 269547
rect 114948 269513 114954 269547
rect 114866 269475 114954 269513
rect 114866 269441 114914 269475
rect 114948 269441 114954 269475
rect 114866 269403 114954 269441
rect 114866 269369 114914 269403
rect 114948 269369 114954 269403
rect 114866 269331 114954 269369
rect 114866 269297 114914 269331
rect 114948 269297 114954 269331
rect 114866 269259 114954 269297
rect 114866 269225 114914 269259
rect 114948 269225 114954 269259
rect 114866 269187 114954 269225
rect 114866 269153 114914 269187
rect 114948 269153 114954 269187
rect 114866 269124 114954 269153
rect 115126 270195 115214 270224
rect 115126 270161 115132 270195
rect 115166 270161 115214 270195
rect 115126 270123 115214 270161
rect 115126 270089 115132 270123
rect 115166 270089 115214 270123
rect 115126 270051 115214 270089
rect 115126 270017 115132 270051
rect 115166 270017 115214 270051
rect 115126 269979 115214 270017
rect 115126 269945 115132 269979
rect 115166 269945 115214 269979
rect 115126 269907 115214 269945
rect 115126 269873 115132 269907
rect 115166 269873 115214 269907
rect 115126 269835 115214 269873
rect 115126 269801 115132 269835
rect 115166 269801 115214 269835
rect 115126 269763 115214 269801
rect 115126 269729 115132 269763
rect 115166 269729 115214 269763
rect 115126 269691 115214 269729
rect 115126 269657 115132 269691
rect 115166 269657 115214 269691
rect 115126 269619 115214 269657
rect 115126 269585 115132 269619
rect 115166 269585 115214 269619
rect 115126 269547 115214 269585
rect 115126 269513 115132 269547
rect 115166 269513 115214 269547
rect 115126 269475 115214 269513
rect 115126 269441 115132 269475
rect 115166 269441 115214 269475
rect 115126 269403 115214 269441
rect 115126 269369 115132 269403
rect 115166 269369 115214 269403
rect 115126 269331 115214 269369
rect 115126 269297 115132 269331
rect 115166 269297 115214 269331
rect 115126 269259 115214 269297
rect 115126 269225 115132 269259
rect 115166 269225 115214 269259
rect 115126 269187 115214 269225
rect 115126 269153 115132 269187
rect 115166 269153 115214 269187
rect 115126 269124 115214 269153
rect 115266 270195 115354 270224
rect 115266 270161 115314 270195
rect 115348 270161 115354 270195
rect 115266 270123 115354 270161
rect 115266 270089 115314 270123
rect 115348 270089 115354 270123
rect 115266 270051 115354 270089
rect 115266 270017 115314 270051
rect 115348 270017 115354 270051
rect 115266 269979 115354 270017
rect 115266 269945 115314 269979
rect 115348 269945 115354 269979
rect 115266 269907 115354 269945
rect 115266 269873 115314 269907
rect 115348 269873 115354 269907
rect 115266 269835 115354 269873
rect 115266 269801 115314 269835
rect 115348 269801 115354 269835
rect 115266 269763 115354 269801
rect 115266 269729 115314 269763
rect 115348 269729 115354 269763
rect 115266 269691 115354 269729
rect 115266 269657 115314 269691
rect 115348 269657 115354 269691
rect 115266 269619 115354 269657
rect 115266 269585 115314 269619
rect 115348 269585 115354 269619
rect 115266 269547 115354 269585
rect 115266 269513 115314 269547
rect 115348 269513 115354 269547
rect 115266 269475 115354 269513
rect 115266 269441 115314 269475
rect 115348 269441 115354 269475
rect 115266 269403 115354 269441
rect 115266 269369 115314 269403
rect 115348 269369 115354 269403
rect 115266 269331 115354 269369
rect 115266 269297 115314 269331
rect 115348 269297 115354 269331
rect 115266 269259 115354 269297
rect 115266 269225 115314 269259
rect 115348 269225 115354 269259
rect 115266 269187 115354 269225
rect 115266 269153 115314 269187
rect 115348 269153 115354 269187
rect 115266 269124 115354 269153
rect 115526 270195 115614 270224
rect 115526 270161 115532 270195
rect 115566 270161 115614 270195
rect 115526 270123 115614 270161
rect 115526 270089 115532 270123
rect 115566 270089 115614 270123
rect 115526 270051 115614 270089
rect 115526 270017 115532 270051
rect 115566 270017 115614 270051
rect 115526 269979 115614 270017
rect 115526 269945 115532 269979
rect 115566 269945 115614 269979
rect 115526 269907 115614 269945
rect 115526 269873 115532 269907
rect 115566 269873 115614 269907
rect 115526 269835 115614 269873
rect 115526 269801 115532 269835
rect 115566 269801 115614 269835
rect 115526 269763 115614 269801
rect 115526 269729 115532 269763
rect 115566 269729 115614 269763
rect 115526 269691 115614 269729
rect 115526 269657 115532 269691
rect 115566 269657 115614 269691
rect 115526 269619 115614 269657
rect 115526 269585 115532 269619
rect 115566 269585 115614 269619
rect 115526 269547 115614 269585
rect 115526 269513 115532 269547
rect 115566 269513 115614 269547
rect 115526 269475 115614 269513
rect 115526 269441 115532 269475
rect 115566 269441 115614 269475
rect 115526 269403 115614 269441
rect 115526 269369 115532 269403
rect 115566 269369 115614 269403
rect 115526 269331 115614 269369
rect 115526 269297 115532 269331
rect 115566 269297 115614 269331
rect 115526 269259 115614 269297
rect 115526 269225 115532 269259
rect 115566 269225 115614 269259
rect 115526 269187 115614 269225
rect 115526 269153 115532 269187
rect 115566 269153 115614 269187
rect 115526 269124 115614 269153
rect 115666 270195 115754 270224
rect 115666 270161 115714 270195
rect 115748 270161 115754 270195
rect 115666 270123 115754 270161
rect 115666 270089 115714 270123
rect 115748 270089 115754 270123
rect 115666 270051 115754 270089
rect 115666 270017 115714 270051
rect 115748 270017 115754 270051
rect 115666 269979 115754 270017
rect 115666 269945 115714 269979
rect 115748 269945 115754 269979
rect 115666 269907 115754 269945
rect 115666 269873 115714 269907
rect 115748 269873 115754 269907
rect 115666 269835 115754 269873
rect 115666 269801 115714 269835
rect 115748 269801 115754 269835
rect 115666 269763 115754 269801
rect 115666 269729 115714 269763
rect 115748 269729 115754 269763
rect 115666 269691 115754 269729
rect 115666 269657 115714 269691
rect 115748 269657 115754 269691
rect 115666 269619 115754 269657
rect 115666 269585 115714 269619
rect 115748 269585 115754 269619
rect 115666 269547 115754 269585
rect 115666 269513 115714 269547
rect 115748 269513 115754 269547
rect 115666 269475 115754 269513
rect 115666 269441 115714 269475
rect 115748 269441 115754 269475
rect 115666 269403 115754 269441
rect 115666 269369 115714 269403
rect 115748 269369 115754 269403
rect 115666 269331 115754 269369
rect 115666 269297 115714 269331
rect 115748 269297 115754 269331
rect 115666 269259 115754 269297
rect 115666 269225 115714 269259
rect 115748 269225 115754 269259
rect 115666 269187 115754 269225
rect 115666 269153 115714 269187
rect 115748 269153 115754 269187
rect 115666 269124 115754 269153
rect 115926 270195 116014 270224
rect 115926 270161 115932 270195
rect 115966 270161 116014 270195
rect 115926 270123 116014 270161
rect 115926 270089 115932 270123
rect 115966 270089 116014 270123
rect 115926 270051 116014 270089
rect 115926 270017 115932 270051
rect 115966 270017 116014 270051
rect 115926 269979 116014 270017
rect 115926 269945 115932 269979
rect 115966 269945 116014 269979
rect 115926 269907 116014 269945
rect 115926 269873 115932 269907
rect 115966 269873 116014 269907
rect 115926 269835 116014 269873
rect 115926 269801 115932 269835
rect 115966 269801 116014 269835
rect 115926 269763 116014 269801
rect 115926 269729 115932 269763
rect 115966 269729 116014 269763
rect 115926 269691 116014 269729
rect 115926 269657 115932 269691
rect 115966 269657 116014 269691
rect 115926 269619 116014 269657
rect 115926 269585 115932 269619
rect 115966 269585 116014 269619
rect 115926 269547 116014 269585
rect 115926 269513 115932 269547
rect 115966 269513 116014 269547
rect 115926 269475 116014 269513
rect 115926 269441 115932 269475
rect 115966 269441 116014 269475
rect 115926 269403 116014 269441
rect 115926 269369 115932 269403
rect 115966 269369 116014 269403
rect 115926 269331 116014 269369
rect 115926 269297 115932 269331
rect 115966 269297 116014 269331
rect 115926 269259 116014 269297
rect 115926 269225 115932 269259
rect 115966 269225 116014 269259
rect 115926 269187 116014 269225
rect 115926 269153 115932 269187
rect 115966 269153 116014 269187
rect 115926 269124 116014 269153
rect 116066 270195 116154 270224
rect 116066 270161 116114 270195
rect 116148 270161 116154 270195
rect 116066 270123 116154 270161
rect 116066 270089 116114 270123
rect 116148 270089 116154 270123
rect 116066 270051 116154 270089
rect 116066 270017 116114 270051
rect 116148 270017 116154 270051
rect 116066 269979 116154 270017
rect 116066 269945 116114 269979
rect 116148 269945 116154 269979
rect 116066 269907 116154 269945
rect 116066 269873 116114 269907
rect 116148 269873 116154 269907
rect 116066 269835 116154 269873
rect 116066 269801 116114 269835
rect 116148 269801 116154 269835
rect 116066 269763 116154 269801
rect 116066 269729 116114 269763
rect 116148 269729 116154 269763
rect 116066 269691 116154 269729
rect 116066 269657 116114 269691
rect 116148 269657 116154 269691
rect 116066 269619 116154 269657
rect 116066 269585 116114 269619
rect 116148 269585 116154 269619
rect 116066 269547 116154 269585
rect 116066 269513 116114 269547
rect 116148 269513 116154 269547
rect 116066 269475 116154 269513
rect 116066 269441 116114 269475
rect 116148 269441 116154 269475
rect 116066 269403 116154 269441
rect 116066 269369 116114 269403
rect 116148 269369 116154 269403
rect 116066 269331 116154 269369
rect 116066 269297 116114 269331
rect 116148 269297 116154 269331
rect 116066 269259 116154 269297
rect 116066 269225 116114 269259
rect 116148 269225 116154 269259
rect 116066 269187 116154 269225
rect 116066 269153 116114 269187
rect 116148 269153 116154 269187
rect 116066 269124 116154 269153
rect 116326 270195 116414 270224
rect 116326 270161 116332 270195
rect 116366 270161 116414 270195
rect 116326 270123 116414 270161
rect 116326 270089 116332 270123
rect 116366 270089 116414 270123
rect 116326 270051 116414 270089
rect 116326 270017 116332 270051
rect 116366 270017 116414 270051
rect 116326 269979 116414 270017
rect 116326 269945 116332 269979
rect 116366 269945 116414 269979
rect 116326 269907 116414 269945
rect 116326 269873 116332 269907
rect 116366 269873 116414 269907
rect 116326 269835 116414 269873
rect 116326 269801 116332 269835
rect 116366 269801 116414 269835
rect 116326 269763 116414 269801
rect 116326 269729 116332 269763
rect 116366 269729 116414 269763
rect 116326 269691 116414 269729
rect 116326 269657 116332 269691
rect 116366 269657 116414 269691
rect 116326 269619 116414 269657
rect 116326 269585 116332 269619
rect 116366 269585 116414 269619
rect 116326 269547 116414 269585
rect 116326 269513 116332 269547
rect 116366 269513 116414 269547
rect 116326 269475 116414 269513
rect 116326 269441 116332 269475
rect 116366 269441 116414 269475
rect 116326 269403 116414 269441
rect 116326 269369 116332 269403
rect 116366 269369 116414 269403
rect 116326 269331 116414 269369
rect 116326 269297 116332 269331
rect 116366 269297 116414 269331
rect 116326 269259 116414 269297
rect 116326 269225 116332 269259
rect 116366 269225 116414 269259
rect 116326 269187 116414 269225
rect 116326 269153 116332 269187
rect 116366 269153 116414 269187
rect 116326 269124 116414 269153
rect 116466 270195 116554 270224
rect 116466 270161 116514 270195
rect 116548 270161 116554 270195
rect 116466 270123 116554 270161
rect 116466 270089 116514 270123
rect 116548 270089 116554 270123
rect 116466 270051 116554 270089
rect 116466 270017 116514 270051
rect 116548 270017 116554 270051
rect 116466 269979 116554 270017
rect 116466 269945 116514 269979
rect 116548 269945 116554 269979
rect 116466 269907 116554 269945
rect 116466 269873 116514 269907
rect 116548 269873 116554 269907
rect 116466 269835 116554 269873
rect 116466 269801 116514 269835
rect 116548 269801 116554 269835
rect 116466 269763 116554 269801
rect 116466 269729 116514 269763
rect 116548 269729 116554 269763
rect 116466 269691 116554 269729
rect 116466 269657 116514 269691
rect 116548 269657 116554 269691
rect 116466 269619 116554 269657
rect 116466 269585 116514 269619
rect 116548 269585 116554 269619
rect 116466 269547 116554 269585
rect 116466 269513 116514 269547
rect 116548 269513 116554 269547
rect 116466 269475 116554 269513
rect 116466 269441 116514 269475
rect 116548 269441 116554 269475
rect 116466 269403 116554 269441
rect 116466 269369 116514 269403
rect 116548 269369 116554 269403
rect 116466 269331 116554 269369
rect 116466 269297 116514 269331
rect 116548 269297 116554 269331
rect 116466 269259 116554 269297
rect 116466 269225 116514 269259
rect 116548 269225 116554 269259
rect 116466 269187 116554 269225
rect 116466 269153 116514 269187
rect 116548 269153 116554 269187
rect 116466 269124 116554 269153
rect 116726 270195 116814 270224
rect 116726 270161 116732 270195
rect 116766 270161 116814 270195
rect 116726 270123 116814 270161
rect 116726 270089 116732 270123
rect 116766 270089 116814 270123
rect 116726 270051 116814 270089
rect 116726 270017 116732 270051
rect 116766 270017 116814 270051
rect 116726 269979 116814 270017
rect 116726 269945 116732 269979
rect 116766 269945 116814 269979
rect 116726 269907 116814 269945
rect 116726 269873 116732 269907
rect 116766 269873 116814 269907
rect 116726 269835 116814 269873
rect 116726 269801 116732 269835
rect 116766 269801 116814 269835
rect 116726 269763 116814 269801
rect 116726 269729 116732 269763
rect 116766 269729 116814 269763
rect 116726 269691 116814 269729
rect 116726 269657 116732 269691
rect 116766 269657 116814 269691
rect 116726 269619 116814 269657
rect 116726 269585 116732 269619
rect 116766 269585 116814 269619
rect 116726 269547 116814 269585
rect 116726 269513 116732 269547
rect 116766 269513 116814 269547
rect 116726 269475 116814 269513
rect 116726 269441 116732 269475
rect 116766 269441 116814 269475
rect 116726 269403 116814 269441
rect 116726 269369 116732 269403
rect 116766 269369 116814 269403
rect 116726 269331 116814 269369
rect 116726 269297 116732 269331
rect 116766 269297 116814 269331
rect 116726 269259 116814 269297
rect 116726 269225 116732 269259
rect 116766 269225 116814 269259
rect 116726 269187 116814 269225
rect 116726 269153 116732 269187
rect 116766 269153 116814 269187
rect 116726 269124 116814 269153
rect 116866 270195 116954 270224
rect 116866 270161 116914 270195
rect 116948 270161 116954 270195
rect 116866 270123 116954 270161
rect 116866 270089 116914 270123
rect 116948 270089 116954 270123
rect 116866 270051 116954 270089
rect 116866 270017 116914 270051
rect 116948 270017 116954 270051
rect 116866 269979 116954 270017
rect 116866 269945 116914 269979
rect 116948 269945 116954 269979
rect 116866 269907 116954 269945
rect 116866 269873 116914 269907
rect 116948 269873 116954 269907
rect 116866 269835 116954 269873
rect 116866 269801 116914 269835
rect 116948 269801 116954 269835
rect 116866 269763 116954 269801
rect 116866 269729 116914 269763
rect 116948 269729 116954 269763
rect 116866 269691 116954 269729
rect 116866 269657 116914 269691
rect 116948 269657 116954 269691
rect 116866 269619 116954 269657
rect 116866 269585 116914 269619
rect 116948 269585 116954 269619
rect 116866 269547 116954 269585
rect 116866 269513 116914 269547
rect 116948 269513 116954 269547
rect 116866 269475 116954 269513
rect 116866 269441 116914 269475
rect 116948 269441 116954 269475
rect 116866 269403 116954 269441
rect 116866 269369 116914 269403
rect 116948 269369 116954 269403
rect 116866 269331 116954 269369
rect 116866 269297 116914 269331
rect 116948 269297 116954 269331
rect 116866 269259 116954 269297
rect 116866 269225 116914 269259
rect 116948 269225 116954 269259
rect 116866 269187 116954 269225
rect 116866 269153 116914 269187
rect 116948 269153 116954 269187
rect 116866 269124 116954 269153
rect 117126 270195 117214 270224
rect 117126 270161 117132 270195
rect 117166 270161 117214 270195
rect 117126 270123 117214 270161
rect 117126 270089 117132 270123
rect 117166 270089 117214 270123
rect 117126 270051 117214 270089
rect 117126 270017 117132 270051
rect 117166 270017 117214 270051
rect 117126 269979 117214 270017
rect 117126 269945 117132 269979
rect 117166 269945 117214 269979
rect 117126 269907 117214 269945
rect 117126 269873 117132 269907
rect 117166 269873 117214 269907
rect 117126 269835 117214 269873
rect 117126 269801 117132 269835
rect 117166 269801 117214 269835
rect 117126 269763 117214 269801
rect 117126 269729 117132 269763
rect 117166 269729 117214 269763
rect 117126 269691 117214 269729
rect 117126 269657 117132 269691
rect 117166 269657 117214 269691
rect 117126 269619 117214 269657
rect 117126 269585 117132 269619
rect 117166 269585 117214 269619
rect 117126 269547 117214 269585
rect 117126 269513 117132 269547
rect 117166 269513 117214 269547
rect 117126 269475 117214 269513
rect 117126 269441 117132 269475
rect 117166 269441 117214 269475
rect 117126 269403 117214 269441
rect 117126 269369 117132 269403
rect 117166 269369 117214 269403
rect 117126 269331 117214 269369
rect 117126 269297 117132 269331
rect 117166 269297 117214 269331
rect 117126 269259 117214 269297
rect 117126 269225 117132 269259
rect 117166 269225 117214 269259
rect 117126 269187 117214 269225
rect 117126 269153 117132 269187
rect 117166 269153 117214 269187
rect 117126 269124 117214 269153
rect 117266 270195 117354 270224
rect 117266 270161 117314 270195
rect 117348 270161 117354 270195
rect 117266 270123 117354 270161
rect 117266 270089 117314 270123
rect 117348 270089 117354 270123
rect 117266 270051 117354 270089
rect 117266 270017 117314 270051
rect 117348 270017 117354 270051
rect 117266 269979 117354 270017
rect 117266 269945 117314 269979
rect 117348 269945 117354 269979
rect 117266 269907 117354 269945
rect 117266 269873 117314 269907
rect 117348 269873 117354 269907
rect 117266 269835 117354 269873
rect 117266 269801 117314 269835
rect 117348 269801 117354 269835
rect 117266 269763 117354 269801
rect 117266 269729 117314 269763
rect 117348 269729 117354 269763
rect 117266 269691 117354 269729
rect 117266 269657 117314 269691
rect 117348 269657 117354 269691
rect 117266 269619 117354 269657
rect 117266 269585 117314 269619
rect 117348 269585 117354 269619
rect 117266 269547 117354 269585
rect 117266 269513 117314 269547
rect 117348 269513 117354 269547
rect 117266 269475 117354 269513
rect 117266 269441 117314 269475
rect 117348 269441 117354 269475
rect 117266 269403 117354 269441
rect 117266 269369 117314 269403
rect 117348 269369 117354 269403
rect 117266 269331 117354 269369
rect 117266 269297 117314 269331
rect 117348 269297 117354 269331
rect 117266 269259 117354 269297
rect 117266 269225 117314 269259
rect 117348 269225 117354 269259
rect 117266 269187 117354 269225
rect 117266 269153 117314 269187
rect 117348 269153 117354 269187
rect 117266 269124 117354 269153
rect 117526 270195 117614 270224
rect 117526 270161 117532 270195
rect 117566 270161 117614 270195
rect 117526 270123 117614 270161
rect 117526 270089 117532 270123
rect 117566 270089 117614 270123
rect 117526 270051 117614 270089
rect 117526 270017 117532 270051
rect 117566 270017 117614 270051
rect 117526 269979 117614 270017
rect 117526 269945 117532 269979
rect 117566 269945 117614 269979
rect 117526 269907 117614 269945
rect 117526 269873 117532 269907
rect 117566 269873 117614 269907
rect 117526 269835 117614 269873
rect 117526 269801 117532 269835
rect 117566 269801 117614 269835
rect 117526 269763 117614 269801
rect 117526 269729 117532 269763
rect 117566 269729 117614 269763
rect 117526 269691 117614 269729
rect 117526 269657 117532 269691
rect 117566 269657 117614 269691
rect 117526 269619 117614 269657
rect 117526 269585 117532 269619
rect 117566 269585 117614 269619
rect 117526 269547 117614 269585
rect 117526 269513 117532 269547
rect 117566 269513 117614 269547
rect 117526 269475 117614 269513
rect 117526 269441 117532 269475
rect 117566 269441 117614 269475
rect 117526 269403 117614 269441
rect 117526 269369 117532 269403
rect 117566 269369 117614 269403
rect 117526 269331 117614 269369
rect 117526 269297 117532 269331
rect 117566 269297 117614 269331
rect 117526 269259 117614 269297
rect 117526 269225 117532 269259
rect 117566 269225 117614 269259
rect 117526 269187 117614 269225
rect 117526 269153 117532 269187
rect 117566 269153 117614 269187
rect 117526 269124 117614 269153
rect 117666 270195 117754 270224
rect 117666 270161 117714 270195
rect 117748 270161 117754 270195
rect 117666 270123 117754 270161
rect 117666 270089 117714 270123
rect 117748 270089 117754 270123
rect 117666 270051 117754 270089
rect 117666 270017 117714 270051
rect 117748 270017 117754 270051
rect 117666 269979 117754 270017
rect 117666 269945 117714 269979
rect 117748 269945 117754 269979
rect 117666 269907 117754 269945
rect 117666 269873 117714 269907
rect 117748 269873 117754 269907
rect 117666 269835 117754 269873
rect 117666 269801 117714 269835
rect 117748 269801 117754 269835
rect 117666 269763 117754 269801
rect 117666 269729 117714 269763
rect 117748 269729 117754 269763
rect 117666 269691 117754 269729
rect 117666 269657 117714 269691
rect 117748 269657 117754 269691
rect 117666 269619 117754 269657
rect 117666 269585 117714 269619
rect 117748 269585 117754 269619
rect 117666 269547 117754 269585
rect 117666 269513 117714 269547
rect 117748 269513 117754 269547
rect 117666 269475 117754 269513
rect 117666 269441 117714 269475
rect 117748 269441 117754 269475
rect 117666 269403 117754 269441
rect 117666 269369 117714 269403
rect 117748 269369 117754 269403
rect 117666 269331 117754 269369
rect 117666 269297 117714 269331
rect 117748 269297 117754 269331
rect 117666 269259 117754 269297
rect 117666 269225 117714 269259
rect 117748 269225 117754 269259
rect 117666 269187 117754 269225
rect 117666 269153 117714 269187
rect 117748 269153 117754 269187
rect 117666 269124 117754 269153
rect 117926 270195 118014 270224
rect 117926 270161 117932 270195
rect 117966 270161 118014 270195
rect 117926 270123 118014 270161
rect 117926 270089 117932 270123
rect 117966 270089 118014 270123
rect 117926 270051 118014 270089
rect 117926 270017 117932 270051
rect 117966 270017 118014 270051
rect 117926 269979 118014 270017
rect 117926 269945 117932 269979
rect 117966 269945 118014 269979
rect 117926 269907 118014 269945
rect 117926 269873 117932 269907
rect 117966 269873 118014 269907
rect 117926 269835 118014 269873
rect 117926 269801 117932 269835
rect 117966 269801 118014 269835
rect 117926 269763 118014 269801
rect 117926 269729 117932 269763
rect 117966 269729 118014 269763
rect 117926 269691 118014 269729
rect 117926 269657 117932 269691
rect 117966 269657 118014 269691
rect 117926 269619 118014 269657
rect 117926 269585 117932 269619
rect 117966 269585 118014 269619
rect 117926 269547 118014 269585
rect 117926 269513 117932 269547
rect 117966 269513 118014 269547
rect 117926 269475 118014 269513
rect 117926 269441 117932 269475
rect 117966 269441 118014 269475
rect 117926 269403 118014 269441
rect 117926 269369 117932 269403
rect 117966 269369 118014 269403
rect 117926 269331 118014 269369
rect 117926 269297 117932 269331
rect 117966 269297 118014 269331
rect 117926 269259 118014 269297
rect 117926 269225 117932 269259
rect 117966 269225 118014 269259
rect 117926 269187 118014 269225
rect 117926 269153 117932 269187
rect 117966 269153 118014 269187
rect 117926 269124 118014 269153
rect 118066 270195 118154 270224
rect 118066 270161 118114 270195
rect 118148 270161 118154 270195
rect 118066 270123 118154 270161
rect 118066 270089 118114 270123
rect 118148 270089 118154 270123
rect 118066 270051 118154 270089
rect 118066 270017 118114 270051
rect 118148 270017 118154 270051
rect 118066 269979 118154 270017
rect 118066 269945 118114 269979
rect 118148 269945 118154 269979
rect 118066 269907 118154 269945
rect 118066 269873 118114 269907
rect 118148 269873 118154 269907
rect 118066 269835 118154 269873
rect 118066 269801 118114 269835
rect 118148 269801 118154 269835
rect 118066 269763 118154 269801
rect 118066 269729 118114 269763
rect 118148 269729 118154 269763
rect 118066 269691 118154 269729
rect 118066 269657 118114 269691
rect 118148 269657 118154 269691
rect 118066 269619 118154 269657
rect 118066 269585 118114 269619
rect 118148 269585 118154 269619
rect 118066 269547 118154 269585
rect 118066 269513 118114 269547
rect 118148 269513 118154 269547
rect 118066 269475 118154 269513
rect 118066 269441 118114 269475
rect 118148 269441 118154 269475
rect 118066 269403 118154 269441
rect 118066 269369 118114 269403
rect 118148 269369 118154 269403
rect 118066 269331 118154 269369
rect 118066 269297 118114 269331
rect 118148 269297 118154 269331
rect 118066 269259 118154 269297
rect 118066 269225 118114 269259
rect 118148 269225 118154 269259
rect 118066 269187 118154 269225
rect 118066 269153 118114 269187
rect 118148 269153 118154 269187
rect 118066 269124 118154 269153
rect 118326 270195 118414 270224
rect 118326 270161 118332 270195
rect 118366 270161 118414 270195
rect 118326 270123 118414 270161
rect 118326 270089 118332 270123
rect 118366 270089 118414 270123
rect 118326 270051 118414 270089
rect 118326 270017 118332 270051
rect 118366 270017 118414 270051
rect 118326 269979 118414 270017
rect 118326 269945 118332 269979
rect 118366 269945 118414 269979
rect 118326 269907 118414 269945
rect 118326 269873 118332 269907
rect 118366 269873 118414 269907
rect 118326 269835 118414 269873
rect 118326 269801 118332 269835
rect 118366 269801 118414 269835
rect 118326 269763 118414 269801
rect 118326 269729 118332 269763
rect 118366 269729 118414 269763
rect 118326 269691 118414 269729
rect 118326 269657 118332 269691
rect 118366 269657 118414 269691
rect 118326 269619 118414 269657
rect 118326 269585 118332 269619
rect 118366 269585 118414 269619
rect 118326 269547 118414 269585
rect 118326 269513 118332 269547
rect 118366 269513 118414 269547
rect 118326 269475 118414 269513
rect 118326 269441 118332 269475
rect 118366 269441 118414 269475
rect 118326 269403 118414 269441
rect 118326 269369 118332 269403
rect 118366 269369 118414 269403
rect 118326 269331 118414 269369
rect 118326 269297 118332 269331
rect 118366 269297 118414 269331
rect 118326 269259 118414 269297
rect 118326 269225 118332 269259
rect 118366 269225 118414 269259
rect 118326 269187 118414 269225
rect 118326 269153 118332 269187
rect 118366 269153 118414 269187
rect 118326 269124 118414 269153
rect 118466 270195 118554 270224
rect 118466 270161 118514 270195
rect 118548 270161 118554 270195
rect 118466 270123 118554 270161
rect 118466 270089 118514 270123
rect 118548 270089 118554 270123
rect 118466 270051 118554 270089
rect 118466 270017 118514 270051
rect 118548 270017 118554 270051
rect 118466 269979 118554 270017
rect 118466 269945 118514 269979
rect 118548 269945 118554 269979
rect 118466 269907 118554 269945
rect 118466 269873 118514 269907
rect 118548 269873 118554 269907
rect 118466 269835 118554 269873
rect 118466 269801 118514 269835
rect 118548 269801 118554 269835
rect 118466 269763 118554 269801
rect 118466 269729 118514 269763
rect 118548 269729 118554 269763
rect 118466 269691 118554 269729
rect 118466 269657 118514 269691
rect 118548 269657 118554 269691
rect 118466 269619 118554 269657
rect 118466 269585 118514 269619
rect 118548 269585 118554 269619
rect 118466 269547 118554 269585
rect 118466 269513 118514 269547
rect 118548 269513 118554 269547
rect 118466 269475 118554 269513
rect 118466 269441 118514 269475
rect 118548 269441 118554 269475
rect 118466 269403 118554 269441
rect 118466 269369 118514 269403
rect 118548 269369 118554 269403
rect 118466 269331 118554 269369
rect 118466 269297 118514 269331
rect 118548 269297 118554 269331
rect 118466 269259 118554 269297
rect 118466 269225 118514 269259
rect 118548 269225 118554 269259
rect 118466 269187 118554 269225
rect 118466 269153 118514 269187
rect 118548 269153 118554 269187
rect 118466 269124 118554 269153
rect 118726 270195 118814 270224
rect 118726 270161 118732 270195
rect 118766 270161 118814 270195
rect 118726 270123 118814 270161
rect 118726 270089 118732 270123
rect 118766 270089 118814 270123
rect 120433 270142 120825 270264
rect 120433 270108 120468 270142
rect 120502 270108 120540 270142
rect 120574 270108 120612 270142
rect 120646 270108 120684 270142
rect 120718 270108 120756 270142
rect 120790 270108 120825 270142
rect 120433 270102 120825 270108
rect 118726 270051 118814 270089
rect 118726 270017 118732 270051
rect 118766 270017 118814 270051
rect 118726 269979 118814 270017
rect 118726 269945 118732 269979
rect 118766 269945 118814 269979
rect 118726 269907 118814 269945
rect 118726 269873 118732 269907
rect 118766 269873 118814 269907
rect 118726 269835 118814 269873
rect 118726 269801 118732 269835
rect 118766 269801 118814 269835
rect 118726 269763 118814 269801
rect 118726 269729 118732 269763
rect 118766 269729 118814 269763
rect 118726 269691 118814 269729
rect 118726 269657 118732 269691
rect 118766 269657 118814 269691
rect 118726 269619 118814 269657
rect 118726 269585 118732 269619
rect 118766 269585 118814 269619
rect 118726 269547 118814 269585
rect 120377 270044 120423 270061
rect 120377 270010 120383 270044
rect 120417 270010 120423 270044
rect 120377 269972 120423 270010
rect 120377 269938 120383 269972
rect 120417 269938 120423 269972
rect 120377 269900 120423 269938
rect 120377 269866 120383 269900
rect 120417 269866 120423 269900
rect 120377 269828 120423 269866
rect 120377 269794 120383 269828
rect 120417 269794 120423 269828
rect 120377 269756 120423 269794
rect 120377 269722 120383 269756
rect 120417 269722 120423 269756
rect 120377 269684 120423 269722
rect 120377 269650 120383 269684
rect 120417 269650 120423 269684
rect 120377 269612 120423 269650
rect 120377 269578 120383 269612
rect 120417 269578 120423 269612
rect 120377 269561 120423 269578
rect 120835 270044 120881 270061
rect 120835 270010 120841 270044
rect 120875 270010 120881 270044
rect 120835 269972 120881 270010
rect 120835 269938 120841 269972
rect 120875 269938 120881 269972
rect 120835 269900 120881 269938
rect 120835 269866 120841 269900
rect 120875 269872 120881 269900
rect 120953 269872 121018 270529
rect 121077 270506 121083 270529
rect 121117 270506 121123 270540
rect 121077 270468 121123 270506
rect 121077 270434 121083 270468
rect 121117 270434 121123 270468
rect 121077 270396 121123 270434
rect 121077 270362 121083 270396
rect 121117 270362 121123 270396
rect 121077 270345 121123 270362
rect 121535 270828 121605 270845
rect 121535 270794 121541 270828
rect 121575 270814 121605 270828
rect 121657 270814 121677 270866
rect 121575 270802 121677 270814
rect 121575 270794 121605 270802
rect 121535 270756 121605 270794
rect 121535 270722 121541 270756
rect 121575 270750 121605 270756
rect 121657 270750 121677 270802
rect 121575 270738 121677 270750
rect 121575 270722 121605 270738
rect 121535 270686 121605 270722
rect 121657 270686 121677 270738
rect 121535 270684 121677 270686
rect 121535 270650 121541 270684
rect 121575 270674 121677 270684
rect 121575 270650 121605 270674
rect 121535 270622 121605 270650
rect 121657 270622 121677 270674
rect 121535 270612 121677 270622
rect 121535 270578 121541 270612
rect 121575 270610 121677 270612
rect 121575 270578 121605 270610
rect 121535 270558 121605 270578
rect 121657 270558 121677 270610
rect 121535 270546 121677 270558
rect 121535 270540 121605 270546
rect 121535 270506 121541 270540
rect 121575 270506 121605 270540
rect 121535 270494 121605 270506
rect 121657 270494 121677 270546
rect 121535 270482 121677 270494
rect 121535 270468 121605 270482
rect 121535 270434 121541 270468
rect 121575 270434 121605 270468
rect 121535 270430 121605 270434
rect 121657 270430 121677 270482
rect 121535 270396 121677 270430
rect 121535 270362 121541 270396
rect 121575 270362 121677 270396
rect 121535 270345 121677 270362
rect 121133 270298 121525 270304
rect 121133 270264 121168 270298
rect 121202 270264 121240 270298
rect 121274 270264 121312 270298
rect 121346 270264 121384 270298
rect 121418 270264 121456 270298
rect 121490 270264 121525 270298
rect 121133 270142 121525 270264
rect 121133 270108 121168 270142
rect 121202 270108 121240 270142
rect 121274 270108 121312 270142
rect 121346 270108 121384 270142
rect 121418 270108 121456 270142
rect 121490 270108 121525 270142
rect 121133 270102 121525 270108
rect 121581 270061 121624 270345
rect 121077 270044 121123 270061
rect 121077 270010 121083 270044
rect 121117 270010 121123 270044
rect 121077 269972 121123 270010
rect 121077 269938 121083 269972
rect 121117 269938 121123 269972
rect 121077 269900 121123 269938
rect 121077 269872 121083 269900
rect 120875 269866 121083 269872
rect 121117 269866 121123 269900
rect 120835 269828 121123 269866
rect 120835 269794 120841 269828
rect 120875 269794 121083 269828
rect 121117 269794 121123 269828
rect 120835 269756 121123 269794
rect 120835 269722 120841 269756
rect 120875 269745 121083 269756
rect 120875 269722 120881 269745
rect 120835 269684 120881 269722
rect 120835 269650 120841 269684
rect 120875 269650 120881 269684
rect 120835 269612 120881 269650
rect 120835 269578 120841 269612
rect 120875 269578 120881 269612
rect 120835 269561 120881 269578
rect 121077 269722 121083 269745
rect 121117 269722 121123 269756
rect 121077 269684 121123 269722
rect 121077 269650 121083 269684
rect 121117 269650 121123 269684
rect 121077 269612 121123 269650
rect 121077 269578 121083 269612
rect 121117 269578 121123 269612
rect 121077 269561 121123 269578
rect 121535 270044 121624 270061
rect 121535 270010 121541 270044
rect 121575 270010 121624 270044
rect 121535 269972 121624 270010
rect 121535 269938 121541 269972
rect 121575 269938 121624 269972
rect 121535 269900 121624 269938
rect 121535 269866 121541 269900
rect 121575 269866 121624 269900
rect 121535 269828 121624 269866
rect 121535 269794 121541 269828
rect 121575 269794 121624 269828
rect 121535 269756 121624 269794
rect 121535 269722 121541 269756
rect 121575 269722 121624 269756
rect 121535 269684 121624 269722
rect 121535 269650 121541 269684
rect 121575 269650 121624 269684
rect 121535 269612 121624 269650
rect 121535 269578 121541 269612
rect 121575 269578 121624 269612
rect 121535 269561 121624 269578
rect 118726 269513 118732 269547
rect 118766 269513 118814 269547
rect 118726 269475 118814 269513
rect 118726 269441 118732 269475
rect 118766 269441 118814 269475
rect 120433 269514 120825 269520
rect 120433 269480 120468 269514
rect 120502 269480 120540 269514
rect 120574 269480 120612 269514
rect 120646 269480 120684 269514
rect 120718 269480 120756 269514
rect 120790 269480 120825 269514
rect 121133 269514 121525 269520
rect 121133 269496 121168 269514
rect 120433 269474 120825 269480
rect 121132 269480 121168 269496
rect 121202 269480 121240 269514
rect 121274 269480 121312 269514
rect 121346 269480 121384 269514
rect 121418 269480 121456 269514
rect 121490 269496 121525 269514
rect 121796 269496 121864 273059
rect 122129 272894 122521 272900
rect 122129 272860 122164 272894
rect 122198 272860 122236 272894
rect 122270 272860 122308 272894
rect 122342 272860 122380 272894
rect 122414 272860 122452 272894
rect 122486 272860 122521 272894
rect 122129 272854 122521 272860
rect 122829 272894 123221 272900
rect 122829 272860 122864 272894
rect 122898 272860 122936 272894
rect 122970 272860 123008 272894
rect 123042 272860 123080 272894
rect 123114 272860 123152 272894
rect 123186 272860 123221 272894
rect 122829 272854 123221 272860
rect 122073 272780 122119 272813
rect 122073 272746 122079 272780
rect 122113 272746 122119 272780
rect 122073 272713 122119 272746
rect 122531 272780 122577 272813
rect 122531 272746 122537 272780
rect 122571 272746 122577 272780
rect 122531 272713 122577 272746
rect 122773 272780 122819 272813
rect 122773 272746 122779 272780
rect 122813 272746 122819 272780
rect 122773 272713 122819 272746
rect 123231 272780 123277 272813
rect 123231 272746 123237 272780
rect 123271 272746 123277 272780
rect 123231 272713 123277 272746
rect 122129 272666 122521 272672
rect 122129 272632 122164 272666
rect 122198 272632 122236 272666
rect 122270 272632 122308 272666
rect 122342 272632 122380 272666
rect 122414 272632 122452 272666
rect 122486 272632 122521 272666
rect 122129 272626 122521 272632
rect 122829 272666 123221 272672
rect 122829 272632 122864 272666
rect 122898 272632 122936 272666
rect 122970 272632 123008 272666
rect 123042 272632 123080 272666
rect 123114 272632 123152 272666
rect 123186 272632 123221 272666
rect 123368 272656 123438 273059
rect 122829 272626 123221 272632
rect 123333 272625 123462 272656
rect 123333 272591 123382 272625
rect 123416 272591 123462 272625
rect 123333 272553 123462 272591
rect 123333 272519 123382 272553
rect 123416 272519 123462 272553
rect 121490 269480 121864 269496
rect 118726 269403 118814 269441
rect 121132 269436 121864 269480
rect 121991 272510 122521 272516
rect 121991 272476 122164 272510
rect 122198 272476 122236 272510
rect 122270 272476 122308 272510
rect 122342 272476 122380 272510
rect 122414 272476 122452 272510
rect 122486 272476 122521 272510
rect 121991 272470 122521 272476
rect 122829 272510 123221 272516
rect 122829 272476 122864 272510
rect 122898 272476 122936 272510
rect 122970 272476 123008 272510
rect 123042 272476 123080 272510
rect 123114 272476 123152 272510
rect 123186 272476 123221 272510
rect 122829 272470 123221 272476
rect 123333 272481 123462 272519
rect 121991 271888 122023 272470
rect 123333 272447 123382 272481
rect 123416 272447 123462 272481
rect 122073 272412 122119 272429
rect 122073 272378 122079 272412
rect 122113 272378 122119 272412
rect 122073 272340 122119 272378
rect 122073 272306 122079 272340
rect 122113 272306 122119 272340
rect 122073 272268 122119 272306
rect 122073 272234 122079 272268
rect 122113 272234 122119 272268
rect 122073 272196 122119 272234
rect 122073 272162 122079 272196
rect 122113 272162 122119 272196
rect 122073 272124 122119 272162
rect 122073 272090 122079 272124
rect 122113 272090 122119 272124
rect 122073 272052 122119 272090
rect 122073 272018 122079 272052
rect 122113 272018 122119 272052
rect 122073 271980 122119 272018
rect 122073 271946 122079 271980
rect 122113 271946 122119 271980
rect 122073 271929 122119 271946
rect 122531 272412 122577 272429
rect 122531 272378 122537 272412
rect 122571 272378 122577 272412
rect 122531 272340 122577 272378
rect 122531 272306 122537 272340
rect 122571 272306 122577 272340
rect 122531 272268 122577 272306
rect 122531 272234 122537 272268
rect 122571 272235 122577 272268
rect 122773 272412 122819 272429
rect 122773 272378 122779 272412
rect 122813 272378 122819 272412
rect 122773 272340 122819 272378
rect 122773 272306 122779 272340
rect 122813 272306 122819 272340
rect 122773 272268 122819 272306
rect 122773 272235 122779 272268
rect 122571 272234 122779 272235
rect 122813 272234 122819 272268
rect 122531 272199 122819 272234
rect 122531 272196 122665 272199
rect 122531 272162 122537 272196
rect 122571 272165 122665 272196
rect 122699 272196 122819 272199
rect 122699 272165 122779 272196
rect 122571 272162 122779 272165
rect 122813 272162 122819 272196
rect 122531 272128 122819 272162
rect 122531 272124 122577 272128
rect 122531 272090 122537 272124
rect 122571 272090 122577 272124
rect 122531 272052 122577 272090
rect 122531 272018 122537 272052
rect 122571 272018 122577 272052
rect 122531 271980 122577 272018
rect 122531 271946 122537 271980
rect 122571 271946 122577 271980
rect 122531 271929 122577 271946
rect 121991 271882 122521 271888
rect 121991 271848 122164 271882
rect 122198 271848 122236 271882
rect 122270 271848 122308 271882
rect 122342 271848 122380 271882
rect 122414 271848 122452 271882
rect 122486 271848 122521 271882
rect 121991 271842 122521 271848
rect 121991 271732 122023 271842
rect 121991 271726 122521 271732
rect 121991 271692 122164 271726
rect 122198 271692 122236 271726
rect 122270 271692 122308 271726
rect 122342 271692 122380 271726
rect 122414 271692 122452 271726
rect 122486 271692 122521 271726
rect 121991 271686 122521 271692
rect 121991 271104 122023 271686
rect 122073 271628 122119 271645
rect 122073 271594 122079 271628
rect 122113 271594 122119 271628
rect 122073 271556 122119 271594
rect 122073 271522 122079 271556
rect 122113 271522 122119 271556
rect 122073 271484 122119 271522
rect 122073 271450 122079 271484
rect 122113 271450 122119 271484
rect 122073 271412 122119 271450
rect 122073 271378 122079 271412
rect 122113 271378 122119 271412
rect 122073 271340 122119 271378
rect 122073 271306 122079 271340
rect 122113 271306 122119 271340
rect 122073 271268 122119 271306
rect 122073 271234 122079 271268
rect 122113 271234 122119 271268
rect 122073 271196 122119 271234
rect 122073 271162 122079 271196
rect 122113 271162 122119 271196
rect 122073 271145 122119 271162
rect 122531 271628 122577 271645
rect 122531 271594 122537 271628
rect 122571 271594 122577 271628
rect 122531 271556 122577 271594
rect 122531 271522 122537 271556
rect 122571 271522 122577 271556
rect 122531 271484 122577 271522
rect 122531 271450 122537 271484
rect 122571 271450 122577 271484
rect 122531 271412 122577 271450
rect 122531 271378 122537 271412
rect 122571 271378 122577 271412
rect 122531 271340 122577 271378
rect 122531 271306 122537 271340
rect 122571 271306 122577 271340
rect 122531 271268 122577 271306
rect 122531 271234 122537 271268
rect 122571 271234 122577 271268
rect 122531 271196 122577 271234
rect 122531 271162 122537 271196
rect 122571 271162 122577 271196
rect 122531 271145 122577 271162
rect 121991 271098 122521 271104
rect 121991 271064 122164 271098
rect 122198 271064 122236 271098
rect 122270 271064 122308 271098
rect 122342 271064 122380 271098
rect 122414 271064 122452 271098
rect 122486 271064 122521 271098
rect 121991 271058 122521 271064
rect 121991 270948 122023 271058
rect 121991 270942 122521 270948
rect 121991 270908 122164 270942
rect 122198 270908 122236 270942
rect 122270 270908 122308 270942
rect 122342 270908 122380 270942
rect 122414 270908 122452 270942
rect 122486 270908 122521 270942
rect 121991 270902 122521 270908
rect 121991 270320 122023 270902
rect 122073 270844 122119 270861
rect 122073 270810 122079 270844
rect 122113 270810 122119 270844
rect 122073 270772 122119 270810
rect 122073 270738 122079 270772
rect 122113 270738 122119 270772
rect 122073 270700 122119 270738
rect 122073 270666 122079 270700
rect 122113 270666 122119 270700
rect 122073 270628 122119 270666
rect 122073 270594 122079 270628
rect 122113 270594 122119 270628
rect 122073 270556 122119 270594
rect 122073 270522 122079 270556
rect 122113 270522 122119 270556
rect 122073 270484 122119 270522
rect 122073 270450 122079 270484
rect 122113 270450 122119 270484
rect 122073 270412 122119 270450
rect 122073 270378 122079 270412
rect 122113 270378 122119 270412
rect 122073 270361 122119 270378
rect 122531 270844 122577 270861
rect 122531 270810 122537 270844
rect 122571 270810 122577 270844
rect 122531 270772 122577 270810
rect 122531 270738 122537 270772
rect 122571 270738 122577 270772
rect 122531 270700 122577 270738
rect 122531 270666 122537 270700
rect 122571 270666 122577 270700
rect 122531 270628 122577 270666
rect 122531 270594 122537 270628
rect 122571 270594 122577 270628
rect 122531 270556 122577 270594
rect 122531 270522 122537 270556
rect 122571 270522 122577 270556
rect 122531 270484 122577 270522
rect 122531 270450 122537 270484
rect 122571 270450 122577 270484
rect 122531 270412 122577 270450
rect 122531 270378 122537 270412
rect 122571 270378 122577 270412
rect 122531 270361 122577 270378
rect 121991 270314 122521 270320
rect 121991 270280 122164 270314
rect 122198 270280 122236 270314
rect 122270 270280 122308 270314
rect 122342 270280 122380 270314
rect 122414 270280 122452 270314
rect 122486 270280 122521 270314
rect 121991 270274 122521 270280
rect 121991 270164 122023 270274
rect 121991 270158 122521 270164
rect 121991 270124 122164 270158
rect 122198 270124 122236 270158
rect 122270 270124 122308 270158
rect 122342 270124 122380 270158
rect 122414 270124 122452 270158
rect 122486 270124 122521 270158
rect 121991 270118 122521 270124
rect 121991 269536 122023 270118
rect 122073 270060 122119 270077
rect 122073 270026 122079 270060
rect 122113 270026 122119 270060
rect 122073 269988 122119 270026
rect 122073 269954 122079 269988
rect 122113 269954 122119 269988
rect 122073 269916 122119 269954
rect 122073 269882 122079 269916
rect 122113 269882 122119 269916
rect 122073 269844 122119 269882
rect 122073 269810 122079 269844
rect 122113 269810 122119 269844
rect 122073 269772 122119 269810
rect 122073 269738 122079 269772
rect 122113 269738 122119 269772
rect 122073 269700 122119 269738
rect 122073 269666 122079 269700
rect 122113 269666 122119 269700
rect 122073 269628 122119 269666
rect 122073 269594 122079 269628
rect 122113 269594 122119 269628
rect 122073 269577 122119 269594
rect 122531 270060 122577 270077
rect 122531 270026 122537 270060
rect 122571 270026 122577 270060
rect 122531 269988 122577 270026
rect 122531 269954 122537 269988
rect 122571 269954 122577 269988
rect 122531 269916 122577 269954
rect 122531 269882 122537 269916
rect 122571 269882 122577 269916
rect 122531 269874 122577 269882
rect 122646 269874 122724 272128
rect 122773 272124 122819 272128
rect 122773 272090 122779 272124
rect 122813 272090 122819 272124
rect 122773 272052 122819 272090
rect 122773 272018 122779 272052
rect 122813 272018 122819 272052
rect 122773 271980 122819 272018
rect 122773 271946 122779 271980
rect 122813 271946 122819 271980
rect 122773 271929 122819 271946
rect 123231 272412 123277 272429
rect 123333 272427 123462 272447
rect 123231 272378 123237 272412
rect 123271 272378 123277 272412
rect 123231 272340 123277 272378
rect 123231 272306 123237 272340
rect 123271 272306 123277 272340
rect 123231 272268 123277 272306
rect 123231 272234 123237 272268
rect 123271 272234 123277 272268
rect 123231 272231 123277 272234
rect 123362 272231 123476 272233
rect 123231 272196 123476 272231
rect 123231 272162 123237 272196
rect 123271 272194 123476 272196
rect 123595 272194 123689 273320
rect 124396 273110 124462 273399
rect 123271 272178 123689 272194
rect 123271 272162 123395 272178
rect 123231 272126 123395 272162
rect 123447 272126 123689 272178
rect 123231 272125 123689 272126
rect 123231 272124 123329 272125
rect 123231 272090 123237 272124
rect 123271 272090 123277 272124
rect 123231 272052 123277 272090
rect 123231 272018 123237 272052
rect 123271 272018 123277 272052
rect 123231 271980 123277 272018
rect 123362 272114 123689 272125
rect 123362 272062 123395 272114
rect 123447 272083 123689 272114
rect 123774 273024 124462 273110
rect 124634 273033 124956 273071
rect 123447 272062 123476 272083
rect 123362 272007 123476 272062
rect 123231 271946 123237 271980
rect 123271 271946 123277 271980
rect 123231 271929 123277 271946
rect 122829 271882 123221 271888
rect 122829 271848 122864 271882
rect 122898 271848 122936 271882
rect 122970 271848 123008 271882
rect 123042 271848 123080 271882
rect 123114 271848 123152 271882
rect 123186 271848 123221 271882
rect 122829 271726 123221 271848
rect 122829 271692 122864 271726
rect 122898 271692 122936 271726
rect 122970 271692 123008 271726
rect 123042 271692 123080 271726
rect 123114 271692 123152 271726
rect 123186 271692 123221 271726
rect 122829 271686 123221 271692
rect 122773 271628 122819 271645
rect 122773 271594 122779 271628
rect 122813 271594 122819 271628
rect 122773 271556 122819 271594
rect 122773 271522 122779 271556
rect 122813 271522 122819 271556
rect 122773 271484 122819 271522
rect 122773 271450 122779 271484
rect 122813 271450 122819 271484
rect 122773 271412 122819 271450
rect 122773 271378 122779 271412
rect 122813 271378 122819 271412
rect 122773 271340 122819 271378
rect 122773 271306 122779 271340
rect 122813 271306 122819 271340
rect 122773 271268 122819 271306
rect 122773 271234 122779 271268
rect 122813 271234 122819 271268
rect 122773 271196 122819 271234
rect 122773 271162 122779 271196
rect 122813 271162 122819 271196
rect 122773 271145 122819 271162
rect 123231 271628 123337 271645
rect 123231 271594 123237 271628
rect 123271 271594 123337 271628
rect 123231 271556 123337 271594
rect 123231 271522 123237 271556
rect 123271 271522 123337 271556
rect 123231 271484 123337 271522
rect 123231 271450 123237 271484
rect 123271 271450 123337 271484
rect 123231 271412 123337 271450
rect 123231 271378 123237 271412
rect 123271 271378 123337 271412
rect 123231 271340 123337 271378
rect 123231 271306 123237 271340
rect 123271 271306 123337 271340
rect 123231 271268 123337 271306
rect 123231 271234 123237 271268
rect 123271 271234 123337 271268
rect 123231 271196 123337 271234
rect 123231 271162 123237 271196
rect 123271 271162 123337 271196
rect 123231 271145 123337 271162
rect 122829 271098 123221 271104
rect 122829 271064 122864 271098
rect 122898 271064 122936 271098
rect 122970 271064 123008 271098
rect 123042 271064 123080 271098
rect 123114 271064 123152 271098
rect 123186 271064 123221 271098
rect 122829 270942 123221 271064
rect 122829 270908 122864 270942
rect 122898 270908 122936 270942
rect 122970 270908 123008 270942
rect 123042 270908 123080 270942
rect 123114 270908 123152 270942
rect 123186 270908 123221 270942
rect 122829 270902 123221 270908
rect 123277 271065 123337 271145
rect 123774 271440 123842 273024
rect 124634 272915 124676 273033
rect 123930 272853 124676 272915
rect 124920 272853 124956 273033
rect 123930 272816 124956 272853
rect 123930 271856 123993 272816
rect 124634 272811 124956 272816
rect 124192 272566 124692 272572
rect 124192 272532 124209 272566
rect 124243 272532 124281 272566
rect 124315 272532 124353 272566
rect 124387 272532 124425 272566
rect 124459 272532 124497 272566
rect 124531 272532 124569 272566
rect 124603 272532 124641 272566
rect 124675 272532 124692 272566
rect 124192 272526 124692 272532
rect 124114 272473 124160 272516
rect 124114 272439 124120 272473
rect 124154 272439 124160 272473
rect 124114 272401 124160 272439
rect 124114 272367 124120 272401
rect 124154 272367 124160 272401
rect 124114 272324 124160 272367
rect 124724 272473 124770 272516
rect 124724 272439 124730 272473
rect 124764 272439 124770 272473
rect 124724 272401 124770 272439
rect 124724 272367 124730 272401
rect 124764 272367 124770 272401
rect 124724 272320 124770 272367
rect 124192 272308 124692 272314
rect 124192 272274 124209 272308
rect 124243 272274 124281 272308
rect 124315 272274 124353 272308
rect 124387 272274 124425 272308
rect 124459 272274 124497 272308
rect 124531 272274 124569 272308
rect 124603 272274 124641 272308
rect 124675 272274 124692 272308
rect 124192 272268 124692 272274
rect 124192 272150 124692 272156
rect 124192 272116 124209 272150
rect 124243 272116 124281 272150
rect 124315 272116 124353 272150
rect 124387 272116 124425 272150
rect 124459 272116 124497 272150
rect 124531 272116 124569 272150
rect 124603 272116 124641 272150
rect 124675 272116 124692 272150
rect 124192 272110 124692 272116
rect 124114 272057 124160 272100
rect 124114 272023 124120 272057
rect 124154 272023 124160 272057
rect 124114 271985 124160 272023
rect 124114 271951 124120 271985
rect 124154 271951 124160 271985
rect 124114 271908 124160 271951
rect 124724 272057 124770 272104
rect 124724 272023 124730 272057
rect 124764 272023 124770 272057
rect 124724 271985 124770 272023
rect 124724 271951 124730 271985
rect 124764 271951 124770 271985
rect 124192 271892 124692 271898
rect 124192 271858 124209 271892
rect 124243 271858 124281 271892
rect 124315 271858 124353 271892
rect 124387 271858 124425 271892
rect 124459 271858 124497 271892
rect 124531 271858 124569 271892
rect 124603 271858 124641 271892
rect 124675 271858 124692 271892
rect 124192 271856 124692 271858
rect 123930 271806 124692 271856
rect 123930 271804 123993 271806
rect 124192 271734 124692 271740
rect 124192 271700 124209 271734
rect 124243 271700 124281 271734
rect 124315 271700 124353 271734
rect 124387 271700 124425 271734
rect 124459 271700 124497 271734
rect 124531 271700 124569 271734
rect 124603 271700 124641 271734
rect 124675 271700 124692 271734
rect 124192 271694 124692 271700
rect 124114 271641 124160 271684
rect 124114 271607 124120 271641
rect 124154 271607 124160 271641
rect 124114 271569 124160 271607
rect 124114 271535 124120 271569
rect 124154 271535 124160 271569
rect 124114 271492 124160 271535
rect 124724 271641 124770 271951
rect 124724 271607 124730 271641
rect 124764 271607 124770 271641
rect 124724 271569 124770 271607
rect 124724 271535 124730 271569
rect 124764 271535 124770 271569
rect 124192 271476 124692 271482
rect 124192 271442 124209 271476
rect 124243 271442 124281 271476
rect 124315 271442 124353 271476
rect 124387 271442 124425 271476
rect 124459 271442 124497 271476
rect 124531 271442 124569 271476
rect 124603 271442 124641 271476
rect 124675 271442 124692 271476
rect 124192 271440 124692 271442
rect 123774 271390 124692 271440
rect 123774 271065 123847 271390
rect 124192 271318 124692 271324
rect 124192 271284 124209 271318
rect 124243 271284 124281 271318
rect 124315 271284 124353 271318
rect 124387 271284 124425 271318
rect 124459 271284 124497 271318
rect 124531 271284 124569 271318
rect 124603 271284 124641 271318
rect 124675 271284 124692 271318
rect 124192 271278 124692 271284
rect 124068 271225 124160 271268
rect 124068 271191 124120 271225
rect 124154 271191 124160 271225
rect 124068 271153 124160 271191
rect 124068 271119 124120 271153
rect 124154 271119 124160 271153
rect 124068 271093 124160 271119
rect 123277 270918 123847 271065
rect 123277 270861 123337 270918
rect 122773 270844 122819 270861
rect 122773 270810 122779 270844
rect 122813 270810 122819 270844
rect 122773 270772 122819 270810
rect 122773 270738 122779 270772
rect 122813 270738 122819 270772
rect 122773 270700 122819 270738
rect 122773 270666 122779 270700
rect 122813 270666 122819 270700
rect 122773 270628 122819 270666
rect 122773 270594 122779 270628
rect 122813 270594 122819 270628
rect 122773 270556 122819 270594
rect 122773 270522 122779 270556
rect 122813 270522 122819 270556
rect 122773 270484 122819 270522
rect 122773 270450 122779 270484
rect 122813 270450 122819 270484
rect 122773 270412 122819 270450
rect 122773 270378 122779 270412
rect 122813 270378 122819 270412
rect 122773 270361 122819 270378
rect 123231 270844 123337 270861
rect 123231 270810 123237 270844
rect 123271 270810 123337 270844
rect 123231 270772 123337 270810
rect 123231 270738 123237 270772
rect 123271 270738 123337 270772
rect 123231 270700 123337 270738
rect 123231 270666 123237 270700
rect 123271 270666 123337 270700
rect 123231 270628 123337 270666
rect 123231 270594 123237 270628
rect 123271 270594 123337 270628
rect 123231 270556 123337 270594
rect 123231 270522 123237 270556
rect 123271 270522 123337 270556
rect 123231 270484 123337 270522
rect 123231 270450 123237 270484
rect 123271 270450 123337 270484
rect 123231 270412 123337 270450
rect 123231 270378 123237 270412
rect 123271 270378 123337 270412
rect 123231 270361 123337 270378
rect 122829 270314 123221 270320
rect 122829 270280 122864 270314
rect 122898 270280 122936 270314
rect 122970 270280 123008 270314
rect 123042 270280 123080 270314
rect 123114 270280 123152 270314
rect 123186 270280 123221 270314
rect 122829 270158 123221 270280
rect 122829 270124 122864 270158
rect 122898 270124 122936 270158
rect 122970 270124 123008 270158
rect 123042 270124 123080 270158
rect 123114 270124 123152 270158
rect 123186 270124 123221 270158
rect 123774 270192 123847 270918
rect 123931 271076 124160 271093
rect 124724 271225 124770 271535
rect 124724 271191 124730 271225
rect 124764 271191 124770 271225
rect 124724 271153 124770 271191
rect 124724 271119 124730 271153
rect 124764 271119 124770 271153
rect 123931 271031 124114 271076
rect 123931 270979 123986 271031
rect 124038 271024 124114 271031
rect 124192 271060 124692 271066
rect 124192 271026 124209 271060
rect 124243 271026 124281 271060
rect 124315 271026 124353 271060
rect 124387 271026 124425 271060
rect 124459 271026 124497 271060
rect 124531 271026 124569 271060
rect 124603 271026 124641 271060
rect 124675 271026 124692 271060
rect 124192 271024 124692 271026
rect 124038 270979 124692 271024
rect 123931 270974 124692 270979
rect 123931 270967 124114 270974
rect 123931 270915 123986 270967
rect 124038 270915 124114 270967
rect 123931 270903 124114 270915
rect 123931 270851 123986 270903
rect 124038 270852 124114 270903
rect 124192 270902 124692 270908
rect 124192 270868 124209 270902
rect 124243 270868 124281 270902
rect 124315 270868 124353 270902
rect 124387 270868 124425 270902
rect 124459 270868 124497 270902
rect 124531 270868 124569 270902
rect 124603 270868 124641 270902
rect 124675 270868 124692 270902
rect 124192 270862 124692 270868
rect 124038 270851 124160 270852
rect 123931 270839 124160 270851
rect 123931 270787 123986 270839
rect 124038 270809 124160 270839
rect 124038 270787 124120 270809
rect 123931 270775 124120 270787
rect 124154 270775 124160 270809
rect 123931 270737 124160 270775
rect 123931 270717 124120 270737
rect 124068 270703 124120 270717
rect 124154 270703 124160 270737
rect 124068 270660 124160 270703
rect 124724 270809 124770 271119
rect 124724 270775 124730 270809
rect 124764 270775 124770 270809
rect 124724 270737 124770 270775
rect 124724 270703 124730 270737
rect 124764 270703 124770 270737
rect 124068 270608 124114 270660
rect 124192 270644 124692 270650
rect 124192 270610 124209 270644
rect 124243 270610 124281 270644
rect 124315 270610 124353 270644
rect 124387 270610 124425 270644
rect 124459 270610 124497 270644
rect 124531 270610 124569 270644
rect 124603 270610 124641 270644
rect 124675 270610 124692 270644
rect 124192 270608 124692 270610
rect 124068 270558 124692 270608
rect 124192 270486 124692 270492
rect 124192 270452 124209 270486
rect 124243 270452 124281 270486
rect 124315 270452 124353 270486
rect 124387 270452 124425 270486
rect 124459 270452 124497 270486
rect 124531 270452 124569 270486
rect 124603 270452 124641 270486
rect 124675 270452 124692 270486
rect 124192 270446 124692 270452
rect 124114 270393 124160 270436
rect 124114 270359 124120 270393
rect 124154 270359 124160 270393
rect 124114 270321 124160 270359
rect 124114 270287 124120 270321
rect 124154 270287 124160 270321
rect 124114 270244 124160 270287
rect 124724 270393 124770 270703
rect 124724 270359 124730 270393
rect 124764 270359 124770 270393
rect 124724 270321 124770 270359
rect 124724 270287 124730 270321
rect 124764 270287 124770 270321
rect 124192 270228 124692 270234
rect 124192 270194 124209 270228
rect 124243 270194 124281 270228
rect 124315 270194 124353 270228
rect 124387 270194 124425 270228
rect 124459 270194 124497 270228
rect 124531 270194 124569 270228
rect 124603 270194 124641 270228
rect 124675 270194 124692 270228
rect 124192 270192 124692 270194
rect 123774 270142 124692 270192
rect 122829 270118 123221 270124
rect 122773 270060 122819 270077
rect 122773 270026 122779 270060
rect 122813 270026 122819 270060
rect 122773 269988 122819 270026
rect 122773 269954 122779 269988
rect 122813 269954 122819 269988
rect 122773 269916 122819 269954
rect 122773 269882 122779 269916
rect 122813 269882 122819 269916
rect 122773 269874 122819 269882
rect 122531 269844 122819 269874
rect 122531 269810 122537 269844
rect 122571 269837 122779 269844
rect 122571 269810 122668 269837
rect 122531 269803 122668 269810
rect 122702 269810 122779 269837
rect 122813 269810 122819 269844
rect 122702 269803 122819 269810
rect 122531 269772 122819 269803
rect 122531 269738 122537 269772
rect 122571 269767 122779 269772
rect 122571 269738 122577 269767
rect 122531 269700 122577 269738
rect 122531 269666 122537 269700
rect 122571 269666 122577 269700
rect 122531 269628 122577 269666
rect 122531 269594 122537 269628
rect 122571 269594 122577 269628
rect 122531 269577 122577 269594
rect 122773 269738 122779 269767
rect 122813 269738 122819 269772
rect 122773 269700 122819 269738
rect 122773 269666 122779 269700
rect 122813 269666 122819 269700
rect 122773 269628 122819 269666
rect 122773 269594 122779 269628
rect 122813 269594 122819 269628
rect 122773 269577 122819 269594
rect 123231 270060 123277 270077
rect 123231 270026 123237 270060
rect 123271 270026 123277 270060
rect 124192 270070 124692 270076
rect 124192 270036 124209 270070
rect 124243 270036 124281 270070
rect 124315 270036 124353 270070
rect 124387 270036 124425 270070
rect 124459 270036 124497 270070
rect 124531 270036 124569 270070
rect 124603 270036 124641 270070
rect 124675 270036 124692 270070
rect 124192 270030 124692 270036
rect 123231 269988 123277 270026
rect 123231 269954 123237 269988
rect 123271 269954 123277 269988
rect 123231 269916 123277 269954
rect 123231 269882 123237 269916
rect 123271 269882 123277 269916
rect 123231 269865 123277 269882
rect 124114 269977 124160 270020
rect 124114 269943 124120 269977
rect 124154 269943 124160 269977
rect 124114 269905 124160 269943
rect 124114 269871 124120 269905
rect 124154 269871 124160 269905
rect 123231 269864 123411 269865
rect 123231 269844 123474 269864
rect 123231 269810 123237 269844
rect 123271 269811 123474 269844
rect 124114 269828 124160 269871
rect 124724 269977 124770 270287
rect 124724 269943 124730 269977
rect 124764 269943 124770 269977
rect 124724 269905 124770 269943
rect 124724 269871 124730 269905
rect 124764 269871 124770 269905
rect 124724 269824 124770 269871
rect 123271 269810 123392 269811
rect 123231 269772 123392 269810
rect 123231 269738 123237 269772
rect 123271 269759 123392 269772
rect 123444 269759 123474 269811
rect 123271 269758 123474 269759
rect 123271 269738 123277 269758
rect 123231 269700 123277 269738
rect 123231 269666 123237 269700
rect 123271 269666 123277 269700
rect 123231 269628 123277 269666
rect 123231 269594 123237 269628
rect 123271 269594 123277 269628
rect 123231 269577 123277 269594
rect 123360 269747 123474 269758
rect 123360 269695 123392 269747
rect 123444 269695 123474 269747
rect 124192 269812 124692 269818
rect 124192 269778 124209 269812
rect 124243 269778 124281 269812
rect 124315 269778 124353 269812
rect 124387 269778 124425 269812
rect 124459 269778 124497 269812
rect 124531 269778 124569 269812
rect 124603 269778 124641 269812
rect 124675 269790 124692 269812
rect 124878 269790 124944 272811
rect 124675 269778 124944 269790
rect 124192 269769 124944 269778
rect 124192 269737 124943 269769
rect 123360 269638 123474 269695
rect 124192 269654 124692 269660
rect 121991 269530 122521 269536
rect 121991 269496 122164 269530
rect 122198 269496 122236 269530
rect 122270 269496 122308 269530
rect 122342 269496 122380 269530
rect 122414 269496 122452 269530
rect 122486 269496 122521 269530
rect 121991 269490 122521 269496
rect 122829 269530 123221 269536
rect 122829 269496 122864 269530
rect 122898 269496 122936 269530
rect 122970 269496 123008 269530
rect 123042 269496 123080 269530
rect 123114 269496 123152 269530
rect 123186 269496 123221 269530
rect 122829 269490 123221 269496
rect 118726 269369 118732 269403
rect 118766 269369 118814 269403
rect 118726 269331 118814 269369
rect 118726 269297 118732 269331
rect 118766 269297 118814 269331
rect 120433 269358 120825 269364
rect 120433 269324 120468 269358
rect 120502 269324 120540 269358
rect 120574 269324 120612 269358
rect 120646 269324 120684 269358
rect 120718 269324 120756 269358
rect 120790 269324 120825 269358
rect 120433 269318 120825 269324
rect 121133 269358 121525 269364
rect 121133 269324 121168 269358
rect 121202 269324 121240 269358
rect 121274 269324 121312 269358
rect 121346 269324 121384 269358
rect 121418 269324 121456 269358
rect 121490 269324 121525 269358
rect 121133 269318 121525 269324
rect 118726 269259 118814 269297
rect 118726 269225 118732 269259
rect 118766 269225 118814 269259
rect 118726 269187 118814 269225
rect 118726 269153 118732 269187
rect 118766 269153 118814 269187
rect 120377 269244 120423 269277
rect 120377 269210 120383 269244
rect 120417 269210 120423 269244
rect 120377 269177 120423 269210
rect 120835 269244 120881 269277
rect 120835 269210 120841 269244
rect 120875 269210 120881 269244
rect 120835 269177 120881 269210
rect 121077 269244 121123 269277
rect 121077 269210 121083 269244
rect 121117 269210 121123 269244
rect 121077 269177 121123 269210
rect 121535 269244 121581 269277
rect 121535 269210 121541 269244
rect 121575 269210 121581 269244
rect 121535 269177 121581 269210
rect 118726 269124 118814 269153
rect 112564 269086 112716 269092
rect 112564 269052 112587 269086
rect 112621 269052 112659 269086
rect 112693 269052 112716 269086
rect 112564 269046 112716 269052
rect 112772 268921 112814 269124
rect 112964 269086 113116 269092
rect 112964 269052 112987 269086
rect 113021 269052 113059 269086
rect 113093 269052 113116 269086
rect 112964 269046 113116 269052
rect 113172 268921 113214 269124
rect 113364 269086 113516 269092
rect 113364 269052 113387 269086
rect 113421 269052 113459 269086
rect 113493 269052 113516 269086
rect 113364 269046 113516 269052
rect 113572 268921 113614 269124
rect 113764 269086 113916 269092
rect 113764 269052 113787 269086
rect 113821 269052 113859 269086
rect 113893 269052 113916 269086
rect 113764 269046 113916 269052
rect 113972 268921 114014 269124
rect 114164 269086 114316 269092
rect 114164 269052 114187 269086
rect 114221 269052 114259 269086
rect 114293 269052 114316 269086
rect 114164 269046 114316 269052
rect 114372 268921 114414 269124
rect 114564 269086 114716 269092
rect 114564 269052 114587 269086
rect 114621 269052 114659 269086
rect 114693 269052 114716 269086
rect 114564 269046 114716 269052
rect 114772 268921 114814 269124
rect 114964 269086 115116 269092
rect 114964 269052 114987 269086
rect 115021 269052 115059 269086
rect 115093 269052 115116 269086
rect 114964 269046 115116 269052
rect 115172 268921 115214 269124
rect 115364 269086 115516 269092
rect 115364 269052 115387 269086
rect 115421 269052 115459 269086
rect 115493 269052 115516 269086
rect 115364 269046 115516 269052
rect 115572 268921 115614 269124
rect 115764 269086 115916 269092
rect 115764 269052 115787 269086
rect 115821 269052 115859 269086
rect 115893 269052 115916 269086
rect 115764 269046 115916 269052
rect 115972 268921 116014 269124
rect 116164 269086 116316 269092
rect 116164 269052 116187 269086
rect 116221 269052 116259 269086
rect 116293 269052 116316 269086
rect 116164 269046 116316 269052
rect 116372 268921 116414 269124
rect 116564 269086 116716 269092
rect 116564 269052 116587 269086
rect 116621 269052 116659 269086
rect 116693 269052 116716 269086
rect 116564 269046 116716 269052
rect 116772 268921 116814 269124
rect 116964 269086 117116 269092
rect 116964 269052 116987 269086
rect 117021 269052 117059 269086
rect 117093 269052 117116 269086
rect 116964 269046 117116 269052
rect 117172 268921 117214 269124
rect 117364 269086 117516 269092
rect 117364 269052 117387 269086
rect 117421 269052 117459 269086
rect 117493 269052 117516 269086
rect 117364 269046 117516 269052
rect 117572 268921 117614 269124
rect 117764 269086 117916 269092
rect 117764 269052 117787 269086
rect 117821 269052 117859 269086
rect 117893 269052 117916 269086
rect 117764 269046 117916 269052
rect 117972 268921 118014 269124
rect 118164 269086 118316 269092
rect 118164 269052 118187 269086
rect 118221 269052 118259 269086
rect 118293 269052 118316 269086
rect 118164 269046 118316 269052
rect 118372 268921 118414 269124
rect 118564 269086 118716 269092
rect 118564 269052 118587 269086
rect 118621 269052 118659 269086
rect 118693 269052 118716 269086
rect 118564 269046 118716 269052
rect 118772 268921 118814 269124
rect 120433 269130 120825 269136
rect 120433 269096 120468 269130
rect 120502 269096 120540 269130
rect 120574 269096 120612 269130
rect 120646 269096 120684 269130
rect 120718 269096 120756 269130
rect 120790 269096 120825 269130
rect 120433 269090 120825 269096
rect 121133 269130 121525 269136
rect 121133 269096 121168 269130
rect 121202 269096 121240 269130
rect 121274 269096 121312 269130
rect 121346 269096 121384 269130
rect 121418 269096 121456 269130
rect 121490 269096 121525 269130
rect 121133 269090 121525 269096
rect 112772 268888 118814 268921
rect 121991 268966 122023 269490
rect 122129 269374 122521 269380
rect 122129 269340 122164 269374
rect 122198 269340 122236 269374
rect 122270 269340 122308 269374
rect 122342 269340 122380 269374
rect 122414 269340 122452 269374
rect 122486 269340 122521 269374
rect 122129 269334 122521 269340
rect 122829 269374 123221 269380
rect 122829 269340 122864 269374
rect 122898 269340 122936 269374
rect 122970 269340 123008 269374
rect 123042 269340 123080 269374
rect 123114 269340 123152 269374
rect 123186 269340 123221 269374
rect 122829 269334 123221 269340
rect 122073 269260 122119 269293
rect 122073 269226 122079 269260
rect 122113 269226 122119 269260
rect 122073 269193 122119 269226
rect 122531 269260 122577 269293
rect 122531 269226 122537 269260
rect 122571 269226 122577 269260
rect 122531 269193 122577 269226
rect 122773 269260 122819 269293
rect 122773 269226 122779 269260
rect 122813 269226 122819 269260
rect 122773 269193 122819 269226
rect 123231 269260 123277 269293
rect 123231 269226 123237 269260
rect 123271 269226 123277 269260
rect 123231 269193 123277 269226
rect 122129 269146 122521 269152
rect 122129 269112 122164 269146
rect 122198 269112 122236 269146
rect 122270 269112 122308 269146
rect 122342 269112 122380 269146
rect 122414 269112 122452 269146
rect 122486 269112 122521 269146
rect 122129 269106 122521 269112
rect 122829 269146 123221 269152
rect 122829 269112 122864 269146
rect 122898 269112 122936 269146
rect 122970 269112 123008 269146
rect 123042 269112 123080 269146
rect 123114 269112 123152 269146
rect 123186 269112 123221 269146
rect 122829 269106 123221 269112
rect 123360 268966 123413 269638
rect 124192 269620 124209 269654
rect 124243 269620 124281 269654
rect 124315 269620 124353 269654
rect 124387 269620 124425 269654
rect 124459 269620 124497 269654
rect 124531 269620 124569 269654
rect 124603 269620 124641 269654
rect 124675 269620 124692 269654
rect 124192 269614 124692 269620
rect 124114 269561 124160 269604
rect 124114 269527 124120 269561
rect 124154 269527 124160 269561
rect 124114 269489 124160 269527
rect 124114 269455 124120 269489
rect 124154 269455 124160 269489
rect 124114 269412 124160 269455
rect 124724 269561 124770 269608
rect 124724 269527 124730 269561
rect 124764 269527 124770 269561
rect 124724 269489 124770 269527
rect 124724 269455 124730 269489
rect 124764 269455 124770 269489
rect 124724 269412 124770 269455
rect 124192 269396 124692 269402
rect 124192 269362 124209 269396
rect 124243 269362 124281 269396
rect 124315 269362 124353 269396
rect 124387 269362 124425 269396
rect 124459 269362 124497 269396
rect 124531 269362 124569 269396
rect 124603 269362 124641 269396
rect 124675 269362 124692 269396
rect 124192 269356 124692 269362
rect 121991 268908 123413 268966
rect 121991 268901 123412 268908
rect 114230 268868 117626 268888
rect 114230 268762 114345 268868
rect 117475 268762 117626 268868
rect 114230 268711 117626 268762
rect 125452 268364 125808 275136
rect 128036 268364 128452 275136
rect 125452 268349 125825 268364
rect 128019 268349 128452 268364
rect 125452 268022 128452 268349
rect 104286 266548 111587 266766
rect 104286 265536 104489 266548
rect 111325 265536 111587 266548
rect 104286 265368 111587 265536
<< via1 >>
rect 106167 282446 113387 283650
rect 102272 280872 103092 281628
rect 107449 279529 107501 279581
rect 107513 279529 107565 279581
rect 107577 279529 107629 279581
rect 107641 279529 107693 279581
rect 108759 279529 108811 279581
rect 108823 279529 108875 279581
rect 108887 279529 108939 279581
rect 108951 279529 109003 279581
rect 107409 279115 107525 279231
rect 102266 275701 103086 276457
rect 107033 277478 107469 277722
rect 107795 277053 107847 277105
rect 107795 276989 107847 277041
rect 107795 276925 107847 276977
rect 107795 276861 107847 276913
rect 107987 276074 108039 276126
rect 107987 276010 108039 276062
rect 109692 278833 109744 278850
rect 109692 278799 109731 278833
rect 109731 278799 109744 278833
rect 109692 278798 109744 278799
rect 109692 278761 109744 278786
rect 109692 278734 109731 278761
rect 109731 278734 109744 278761
rect 109692 278689 109744 278722
rect 109692 278670 109731 278689
rect 109731 278670 109744 278689
rect 109692 278655 109731 278658
rect 109731 278655 109744 278658
rect 109692 278617 109744 278655
rect 109692 278606 109731 278617
rect 109731 278606 109744 278617
rect 109692 278583 109731 278594
rect 109731 278583 109744 278594
rect 109692 278545 109744 278583
rect 109692 278542 109731 278545
rect 109731 278542 109744 278545
rect 109692 278511 109731 278530
rect 109731 278511 109744 278530
rect 109692 278478 109744 278511
rect 109692 278439 109731 278466
rect 109731 278439 109744 278466
rect 109692 278414 109744 278439
rect 109692 278401 109744 278402
rect 109692 278367 109731 278401
rect 109731 278367 109744 278401
rect 109692 278350 109744 278367
rect 109692 278329 109744 278338
rect 109692 278295 109731 278329
rect 109731 278295 109744 278329
rect 109692 278286 109744 278295
rect 109692 278257 109744 278274
rect 109692 278223 109731 278257
rect 109731 278223 109744 278257
rect 109692 278222 109744 278223
rect 109692 278185 109744 278210
rect 109692 278158 109731 278185
rect 109731 278158 109744 278185
rect 109692 278113 109744 278146
rect 109692 278094 109731 278113
rect 109731 278094 109744 278113
rect 109692 278079 109731 278082
rect 109731 278079 109744 278082
rect 109692 278041 109744 278079
rect 109692 278030 109731 278041
rect 109731 278030 109744 278041
rect 109466 277223 109518 277275
rect 109466 277159 109518 277211
rect 109466 277095 109518 277147
rect 109466 277031 109518 277083
rect 109466 276967 109518 277019
rect 109466 276903 109518 276955
rect 109466 276839 109518 276891
rect 109466 276775 109518 276827
rect 109687 277687 109731 277696
rect 109731 277687 109739 277696
rect 109687 277649 109739 277687
rect 109687 277644 109731 277649
rect 109731 277644 109739 277649
rect 109687 277615 109731 277632
rect 109731 277615 109739 277632
rect 109687 277580 109739 277615
rect 109687 277543 109731 277568
rect 109731 277543 109739 277568
rect 109687 277516 109739 277543
rect 109687 277471 109731 277504
rect 109731 277471 109739 277504
rect 109687 277452 109739 277471
rect 109687 277433 109739 277440
rect 109687 277399 109731 277433
rect 109731 277399 109739 277433
rect 109687 277388 109739 277399
rect 109687 277361 109739 277376
rect 109687 277327 109731 277361
rect 109731 277327 109739 277361
rect 109687 277324 109739 277327
rect 109687 277289 109739 277312
rect 109687 277260 109731 277289
rect 109731 277260 109739 277289
rect 109687 277217 109739 277248
rect 109687 277196 109731 277217
rect 109731 277196 109739 277217
rect 109687 277183 109731 277184
rect 109731 277183 109739 277184
rect 109687 277145 109739 277183
rect 109687 277132 109731 277145
rect 109731 277132 109739 277145
rect 109687 277111 109731 277120
rect 109731 277111 109739 277120
rect 109687 277073 109739 277111
rect 109687 277068 109731 277073
rect 109731 277068 109739 277073
rect 109687 277039 109731 277056
rect 109731 277039 109739 277056
rect 109687 277004 109739 277039
rect 109687 276967 109731 276992
rect 109731 276967 109739 276992
rect 109687 276940 109739 276967
rect 109687 276895 109731 276928
rect 109731 276895 109739 276928
rect 109687 276876 109739 276895
rect 109466 276711 109518 276763
rect 109466 276647 109518 276699
rect 109927 276167 110171 276347
rect 109263 275878 109315 275930
rect 109327 275878 109379 275930
rect 109391 275878 109443 275930
rect 109455 275878 109507 275930
rect 109519 275878 109571 275930
rect 109583 275878 109635 275930
rect 108232 275593 108348 275709
rect 114890 280277 114942 280286
rect 114890 280243 114899 280277
rect 114899 280243 114933 280277
rect 114933 280243 114942 280277
rect 114890 280234 114942 280243
rect 115262 280277 115314 280286
rect 115262 280243 115271 280277
rect 115271 280243 115305 280277
rect 115305 280243 115314 280277
rect 115262 280234 115314 280243
rect 114891 279854 114943 279861
rect 114891 279820 114899 279854
rect 114899 279820 114933 279854
rect 114933 279820 114943 279854
rect 114891 279809 114943 279820
rect 115262 279854 115314 279861
rect 115262 279820 115271 279854
rect 115271 279820 115305 279854
rect 115305 279820 115314 279854
rect 115262 279809 115314 279820
rect 114890 278611 114942 278620
rect 114890 278577 114899 278611
rect 114899 278577 114933 278611
rect 114933 278577 114942 278611
rect 114890 278568 114942 278577
rect 115262 278611 115314 278620
rect 115262 278577 115271 278611
rect 115271 278577 115305 278611
rect 115305 278577 115314 278611
rect 115262 278568 115314 278577
rect 119363 278720 119735 281140
rect 124573 280587 124881 280767
rect 120529 279584 120581 279636
rect 120593 279584 120645 279636
rect 120657 279584 120709 279636
rect 114891 278188 114943 278195
rect 114891 278154 114899 278188
rect 114899 278154 114933 278188
rect 114933 278154 114943 278188
rect 114891 278143 114943 278154
rect 115262 278188 115314 278195
rect 115262 278154 115271 278188
rect 115271 278154 115305 278188
rect 115305 278154 115314 278188
rect 115262 278143 115314 278154
rect 121605 279342 121657 279394
rect 121605 279278 121657 279330
rect 121605 279214 121657 279266
rect 121866 279299 122174 279863
rect 121605 279150 121657 279202
rect 121605 279086 121657 279138
rect 121605 279022 121657 279074
rect 121605 278958 121657 279010
rect 121605 278894 121657 278946
rect 121605 278830 121657 278882
rect 121605 278766 121657 278818
rect 121605 278702 121657 278754
rect 121605 278638 121657 278690
rect 121605 278574 121657 278626
rect 121605 278510 121657 278562
rect 121605 278446 121657 278498
rect 121605 278382 121657 278434
rect 121605 278318 121657 278370
rect 121605 278254 121657 278306
rect 121605 278190 121657 278242
rect 121605 278126 121657 278178
rect 121605 278062 121657 278114
rect 121605 277998 121657 278050
rect 121605 277934 121657 277986
rect 114890 276945 114942 276954
rect 114890 276911 114899 276945
rect 114899 276911 114933 276945
rect 114933 276911 114942 276945
rect 114890 276902 114942 276911
rect 115262 276945 115314 276954
rect 115262 276911 115271 276945
rect 115271 276911 115305 276945
rect 115305 276911 115314 276945
rect 115262 276902 115314 276911
rect 114891 276522 114943 276529
rect 114891 276488 114899 276522
rect 114899 276488 114933 276522
rect 114933 276488 114943 276522
rect 114891 276477 114943 276488
rect 115262 276522 115314 276529
rect 115262 276488 115271 276522
rect 115271 276488 115305 276522
rect 115305 276488 115314 276522
rect 115262 276477 115314 276488
rect 121605 277870 121657 277922
rect 121605 277806 121657 277858
rect 121605 277742 121657 277794
rect 121605 277678 121657 277730
rect 121605 277614 121657 277666
rect 121605 277550 121657 277602
rect 121605 277486 121657 277538
rect 120959 277020 121011 277072
rect 120959 276956 121011 277008
rect 120959 276892 121011 276944
rect 120959 276828 121011 276880
rect 114890 275279 114942 275288
rect 114890 275245 114899 275279
rect 114899 275245 114933 275279
rect 114933 275245 114942 275279
rect 114890 275236 114942 275245
rect 115262 275279 115314 275288
rect 115262 275245 115271 275279
rect 115271 275245 115305 275279
rect 115305 275245 115314 275279
rect 115262 275236 115314 275245
rect 114891 274856 114943 274863
rect 114891 274822 114899 274856
rect 114899 274822 114933 274856
rect 114933 274822 114943 274856
rect 114891 274811 114943 274822
rect 115262 274856 115314 274863
rect 115262 274822 115271 274856
rect 115271 274822 115305 274856
rect 115305 274822 115314 274856
rect 115262 274811 115314 274822
rect 102638 273799 105186 274043
rect 114890 273613 114942 273622
rect 114890 273579 114899 273613
rect 114899 273579 114933 273613
rect 114933 273579 114942 273613
rect 114890 273570 114942 273579
rect 115262 273613 115314 273622
rect 115262 273579 115271 273613
rect 115271 273579 115305 273613
rect 115305 273579 115314 273613
rect 115262 273570 115314 273579
rect 121841 276155 121893 276207
rect 121841 276091 121893 276143
rect 121841 276027 121893 276079
rect 122415 274786 122531 275286
rect 121842 273753 121894 273805
rect 121842 273689 121894 273741
rect 121842 273625 121894 273677
rect 114891 273190 114943 273197
rect 114891 273156 114899 273190
rect 114899 273156 114933 273190
rect 114933 273156 114943 273190
rect 114891 273145 114943 273156
rect 115262 273190 115314 273197
rect 115262 273156 115271 273190
rect 115271 273156 115305 273190
rect 115305 273156 115314 273190
rect 115262 273145 115314 273156
rect 122652 273397 122704 273449
rect 123797 273397 123849 273449
rect 120959 272929 121011 272981
rect 120959 272865 121011 272917
rect 120959 272801 121011 272853
rect 120959 272737 121011 272789
rect 107300 271897 107352 271949
rect 107300 271833 107352 271885
rect 108651 272026 108703 272078
rect 108715 272026 108767 272078
rect 108779 272026 108831 272078
rect 107049 271406 107101 271458
rect 107049 271342 107101 271394
rect 108445 271406 108497 271458
rect 108445 271342 108497 271394
rect 106967 271252 107019 271304
rect 106967 271188 107019 271240
rect 106967 271124 107019 271176
rect 107049 271036 107101 271088
rect 107049 270972 107101 271024
rect 108445 271036 108497 271088
rect 108445 270972 108497 271024
rect 114830 271984 115522 272004
rect 114830 271950 115019 271984
rect 115019 271950 115053 271984
rect 115053 271950 115091 271984
rect 115091 271950 115125 271984
rect 115125 271950 115163 271984
rect 115163 271950 115197 271984
rect 115197 271950 115235 271984
rect 115235 271950 115269 271984
rect 115269 271950 115307 271984
rect 115307 271950 115341 271984
rect 115341 271950 115379 271984
rect 115379 271950 115413 271984
rect 115413 271950 115451 271984
rect 115451 271950 115485 271984
rect 115485 271950 115522 271984
rect 114830 271824 115522 271950
rect 112288 270468 113428 270648
rect 121605 272286 121657 272338
rect 121605 272222 121657 272274
rect 121605 272158 121657 272210
rect 121605 272094 121657 272146
rect 121605 272030 121657 272082
rect 121605 271966 121657 272018
rect 121605 271902 121657 271954
rect 121605 271838 121657 271890
rect 121605 271774 121657 271826
rect 121605 271710 121657 271762
rect 121605 271646 121657 271698
rect 121605 271582 121657 271634
rect 121605 271518 121657 271570
rect 121605 271454 121657 271506
rect 121605 271390 121657 271442
rect 121605 271326 121657 271378
rect 121605 271262 121657 271314
rect 121605 271198 121657 271250
rect 121605 271134 121657 271186
rect 121605 271070 121657 271122
rect 121605 271006 121657 271058
rect 121605 270942 121657 270994
rect 121605 270878 121657 270930
rect 121605 270814 121657 270866
rect 121605 270750 121657 270802
rect 121605 270686 121657 270738
rect 121605 270622 121657 270674
rect 121605 270558 121657 270610
rect 121605 270494 121657 270546
rect 121605 270430 121657 270482
rect 123395 272126 123447 272178
rect 123395 272062 123447 272114
rect 124676 272853 124920 273033
rect 123986 270979 124038 271031
rect 123986 270915 124038 270967
rect 123986 270851 124038 270903
rect 123986 270787 124038 270839
rect 123392 269759 123444 269811
rect 123392 269695 123444 269747
rect 125808 268364 125825 275136
rect 125825 268364 128019 275136
rect 128019 268364 128036 275136
rect 104489 265536 111325 266548
<< metal2 >>
rect 105796 283650 113672 283895
rect 105796 283636 106167 283650
rect 113387 283636 113672 283650
rect 105796 282460 106149 283636
rect 113405 282460 113672 283636
rect 105796 282446 106167 282460
rect 113387 282446 113672 282460
rect 105796 282251 113672 282446
rect 102098 281638 103259 281810
rect 102098 280862 102254 281638
rect 103110 280862 103259 281638
rect 119257 281148 119845 281225
rect 121769 281148 122109 281149
rect 119257 281140 122109 281148
rect 102098 280720 103259 280862
rect 114322 281007 115149 281071
rect 114322 279876 114413 281007
rect 114865 280288 114970 280311
rect 114865 280232 114888 280288
rect 114944 280232 114970 280288
rect 114865 280204 114970 280232
rect 115069 280265 115149 281007
rect 115235 280288 115340 280311
rect 115235 280265 115260 280288
rect 115069 280232 115260 280265
rect 115316 280232 115340 280288
rect 115069 280213 115340 280232
rect 115235 280204 115340 280213
rect 114322 279861 115030 279876
rect 114322 279805 114891 279861
rect 114947 279805 115030 279861
rect 114322 279791 115030 279805
rect 115175 279861 115900 279876
rect 115175 279805 115257 279861
rect 115314 279809 115900 279861
rect 115313 279805 115900 279809
rect 115175 279791 115900 279805
rect 107341 279581 107796 279642
rect 107341 279529 107449 279581
rect 107501 279529 107513 279581
rect 107565 279529 107577 279581
rect 107629 279529 107641 279581
rect 107693 279529 107796 279581
rect 107341 279471 107796 279529
rect 108650 279581 109105 279641
rect 108650 279529 108759 279581
rect 108811 279529 108823 279581
rect 108875 279529 108887 279581
rect 108939 279529 108951 279581
rect 109003 279554 109105 279581
rect 109003 279529 109575 279554
rect 108650 279491 109575 279529
rect 108650 279471 109576 279491
rect 107341 279231 107584 279471
rect 108978 279470 109576 279471
rect 107341 279115 107409 279231
rect 107525 279115 107584 279231
rect 107341 279074 107584 279115
rect 109441 278052 109576 279470
rect 109659 278850 109771 278903
rect 109659 278798 109692 278850
rect 109744 278798 109771 278850
rect 109659 278786 109771 278798
rect 109659 278734 109692 278786
rect 109744 278734 109771 278786
rect 109659 278722 109771 278734
rect 109659 278670 109692 278722
rect 109744 278670 109771 278722
rect 109659 278658 109771 278670
rect 109659 278606 109692 278658
rect 109744 278606 109771 278658
rect 114865 278628 114970 278645
rect 109659 278594 109771 278606
rect 109659 278542 109692 278594
rect 109744 278542 109771 278594
rect 109659 278530 109771 278542
rect 109659 278478 109692 278530
rect 109744 278478 109771 278530
rect 109659 278466 109771 278478
rect 109659 278414 109692 278466
rect 109744 278414 109771 278466
rect 109659 278402 109771 278414
rect 109659 278350 109692 278402
rect 109744 278350 109771 278402
rect 109659 278338 109771 278350
rect 109659 278286 109692 278338
rect 109744 278286 109771 278338
rect 109659 278274 109771 278286
rect 109659 278222 109692 278274
rect 109744 278222 109771 278274
rect 109659 278210 109771 278222
rect 109659 278158 109692 278210
rect 109744 278158 109771 278210
rect 109659 278146 109771 278158
rect 109659 278094 109692 278146
rect 109744 278094 109771 278146
rect 109659 278082 109771 278094
rect 109659 278052 109692 278082
rect 109441 278030 109692 278052
rect 109744 278030 109771 278082
rect 109441 277973 109771 278030
rect 114303 278622 114970 278628
rect 114303 278566 114888 278622
rect 114944 278566 114970 278622
rect 114303 278543 114970 278566
rect 106957 277748 107553 277799
rect 106957 277452 107023 277748
rect 107479 277452 107553 277748
rect 109441 277755 109709 277973
rect 109441 277696 109771 277755
rect 109441 277695 109687 277696
rect 106957 277403 107553 277452
rect 109659 277644 109687 277695
rect 109739 277644 109771 277696
rect 109659 277632 109771 277644
rect 109659 277580 109687 277632
rect 109739 277580 109771 277632
rect 109659 277568 109771 277580
rect 109659 277516 109687 277568
rect 109739 277516 109771 277568
rect 109659 277504 109771 277516
rect 109659 277452 109687 277504
rect 109739 277452 109771 277504
rect 109659 277440 109771 277452
rect 109659 277388 109687 277440
rect 109739 277388 109771 277440
rect 109659 277376 109771 277388
rect 109276 277275 109568 277341
rect 109276 277262 109466 277275
rect 107754 277105 107889 277153
rect 107754 277053 107795 277105
rect 107847 277053 107889 277105
rect 107754 277041 107889 277053
rect 107754 276989 107795 277041
rect 107847 276989 107889 277041
rect 107754 276977 107889 276989
rect 107754 276925 107795 276977
rect 107847 276925 107889 276977
rect 107754 276913 107889 276925
rect 107754 276861 107795 276913
rect 107847 276861 107889 276913
rect 107754 276808 107889 276861
rect 102098 276467 103259 276621
rect 102098 276457 102288 276467
rect 103064 276457 103259 276467
rect 102098 275701 102266 276457
rect 103086 275701 103259 276457
rect 107789 276165 107889 276808
rect 109276 276726 109356 277262
rect 109518 277223 109568 277275
rect 109492 277211 109568 277223
rect 109518 277159 109568 277211
rect 109492 277147 109568 277159
rect 109518 277095 109568 277147
rect 109492 277083 109568 277095
rect 109518 277031 109568 277083
rect 109492 277019 109568 277031
rect 109518 276967 109568 277019
rect 109492 276955 109568 276967
rect 109518 276903 109568 276955
rect 109492 276891 109568 276903
rect 109518 276839 109568 276891
rect 109492 276827 109568 276839
rect 109518 276775 109568 276827
rect 109659 277324 109687 277376
rect 109739 277324 109771 277376
rect 109659 277312 109771 277324
rect 109659 277260 109687 277312
rect 109739 277260 109771 277312
rect 109659 277248 109771 277260
rect 109659 277196 109687 277248
rect 109739 277196 109771 277248
rect 109659 277184 109771 277196
rect 109659 277132 109687 277184
rect 109739 277132 109771 277184
rect 109659 277120 109771 277132
rect 109659 277068 109687 277120
rect 109739 277068 109771 277120
rect 109659 277056 109771 277068
rect 109659 277004 109687 277056
rect 109739 277004 109771 277056
rect 109659 276992 109771 277004
rect 109659 276940 109687 276992
rect 109739 276940 109771 276992
rect 109659 276928 109771 276940
rect 109659 276876 109687 276928
rect 109739 276876 109771 276928
rect 109659 276825 109771 276876
rect 109492 276763 109568 276775
rect 109276 276711 109466 276726
rect 109518 276711 109568 276763
rect 109276 276699 109568 276711
rect 109276 276647 109466 276699
rect 109518 276647 109568 276699
rect 109276 276633 109568 276647
rect 109413 276577 109568 276633
rect 114303 276544 114407 278543
rect 114865 278538 114970 278543
rect 115235 278632 115340 278645
rect 115788 278632 115900 279791
rect 115235 278622 115900 278632
rect 119257 278720 119363 281140
rect 119735 280610 122109 281140
rect 119735 278720 119845 280610
rect 121747 280609 122109 280610
rect 121899 279937 122109 280609
rect 124495 280767 124958 280846
rect 124495 280587 124573 280767
rect 124881 280587 124958 280767
rect 124495 280498 124958 280587
rect 121797 279863 122235 279937
rect 120433 279654 120825 279712
rect 120433 279636 121677 279654
rect 120433 279584 120529 279636
rect 120581 279584 120593 279636
rect 120645 279584 120657 279636
rect 120709 279584 121677 279636
rect 120433 279559 121677 279584
rect 120433 279510 120825 279559
rect 119257 278631 119845 278720
rect 121587 279394 121677 279559
rect 121587 279342 121605 279394
rect 121657 279342 121677 279394
rect 121587 279330 121677 279342
rect 121587 279278 121605 279330
rect 121657 279278 121677 279330
rect 121587 279266 121677 279278
rect 121587 279214 121605 279266
rect 121657 279214 121677 279266
rect 121797 279299 121866 279863
rect 122174 279299 122235 279863
rect 121797 279225 122235 279299
rect 121587 279202 121677 279214
rect 121587 279150 121605 279202
rect 121657 279150 121677 279202
rect 121587 279138 121677 279150
rect 121587 279086 121605 279138
rect 121657 279086 121677 279138
rect 121587 279074 121677 279086
rect 121587 279022 121605 279074
rect 121657 279022 121677 279074
rect 121587 279010 121677 279022
rect 121587 278958 121605 279010
rect 121657 278958 121677 279010
rect 121587 278946 121677 278958
rect 121587 278894 121605 278946
rect 121657 278894 121677 278946
rect 121587 278882 121677 278894
rect 121587 278830 121605 278882
rect 121657 278830 121677 278882
rect 121587 278818 121677 278830
rect 121587 278766 121605 278818
rect 121657 278766 121677 278818
rect 121587 278754 121677 278766
rect 121587 278702 121605 278754
rect 121657 278702 121677 278754
rect 121587 278690 121677 278702
rect 121587 278638 121605 278690
rect 121657 278638 121677 278690
rect 115235 278566 115260 278622
rect 115316 278566 115900 278622
rect 115235 278547 115900 278566
rect 121587 278626 121677 278638
rect 121587 278574 121605 278626
rect 121657 278574 121677 278626
rect 121587 278562 121677 278574
rect 115235 278538 115340 278547
rect 121587 278510 121605 278562
rect 121657 278510 121677 278562
rect 121587 278498 121677 278510
rect 121587 278446 121605 278498
rect 121657 278446 121677 278498
rect 121587 278434 121677 278446
rect 121587 278382 121605 278434
rect 121657 278382 121677 278434
rect 121587 278370 121677 278382
rect 121587 278318 121605 278370
rect 121657 278318 121677 278370
rect 121587 278306 121677 278318
rect 121587 278254 121605 278306
rect 121657 278254 121677 278306
rect 121587 278242 121677 278254
rect 114843 278195 115030 278210
rect 114843 278139 114891 278195
rect 114947 278139 115030 278195
rect 114843 278125 115030 278139
rect 115175 278195 115362 278210
rect 115175 278139 115257 278195
rect 115314 278143 115362 278195
rect 115313 278139 115362 278143
rect 115175 278125 115362 278139
rect 121587 278190 121605 278242
rect 121657 278190 121677 278242
rect 121587 278178 121677 278190
rect 121587 278126 121605 278178
rect 121657 278126 121677 278178
rect 121587 278114 121677 278126
rect 121587 278062 121605 278114
rect 121657 278062 121677 278114
rect 121587 278050 121677 278062
rect 121587 277998 121605 278050
rect 121657 277998 121677 278050
rect 121587 277986 121677 277998
rect 121587 277934 121605 277986
rect 121657 277934 121677 277986
rect 121587 277922 121677 277934
rect 121587 277870 121605 277922
rect 121657 277870 121677 277922
rect 121587 277858 121677 277870
rect 121587 277806 121605 277858
rect 121657 277814 121677 277858
rect 121657 277806 121972 277814
rect 121587 277794 121972 277806
rect 121587 277742 121605 277794
rect 121657 277742 121972 277794
rect 121587 277730 121972 277742
rect 121587 277678 121605 277730
rect 121657 277718 121972 277730
rect 121657 277717 122169 277718
rect 121657 277678 122191 277717
rect 121587 277666 122191 277678
rect 121587 277614 121605 277666
rect 121657 277614 122191 277666
rect 121587 277602 122191 277614
rect 121587 277550 121605 277602
rect 121657 277550 122191 277602
rect 121587 277538 122191 277550
rect 121587 277486 121605 277538
rect 121657 277504 122191 277538
rect 121657 277486 121677 277504
rect 121908 277503 122191 277504
rect 120953 277072 121018 277099
rect 120953 277020 120959 277072
rect 121011 277020 121018 277072
rect 120953 277008 121018 277020
rect 114865 276956 114970 276979
rect 114865 276900 114888 276956
rect 114944 276900 114970 276956
rect 114865 276872 114970 276900
rect 115235 276956 115340 276979
rect 115235 276900 115260 276956
rect 115316 276900 115340 276956
rect 115235 276872 115340 276900
rect 120953 276956 120959 277008
rect 121011 276956 121018 277008
rect 120953 276944 121018 276956
rect 120953 276892 120959 276944
rect 121011 276892 121018 276944
rect 120953 276880 121018 276892
rect 120953 276828 120959 276880
rect 121011 276828 121018 276880
rect 114303 276529 115030 276544
rect 114303 276473 114891 276529
rect 114947 276473 115030 276529
rect 114303 276460 115030 276473
rect 114324 276459 115030 276460
rect 115175 276529 115900 276544
rect 115175 276473 115257 276529
rect 115314 276477 115900 276529
rect 115313 276473 115900 276477
rect 115175 276459 115900 276473
rect 109383 276316 109700 276394
rect 109383 276180 109475 276316
rect 109611 276180 109700 276316
rect 109383 276165 109700 276180
rect 109824 276347 110271 276420
rect 109824 276167 109927 276347
rect 110171 276167 110271 276347
rect 109824 276165 110271 276167
rect 107789 276126 110271 276165
rect 107789 276091 107987 276126
rect 107947 276074 107987 276091
rect 108039 276093 110271 276126
rect 108039 276091 109879 276093
rect 108039 276074 108079 276091
rect 107947 276062 108079 276074
rect 107947 276010 107987 276062
rect 108039 276010 108079 276062
rect 107947 275970 108079 276010
rect 108280 275968 109712 275969
rect 108216 275930 109712 275968
rect 108216 275878 109263 275930
rect 109315 275878 109327 275930
rect 109379 275878 109391 275930
rect 109443 275878 109455 275930
rect 109507 275878 109519 275930
rect 109571 275878 109583 275930
rect 109635 275878 109712 275930
rect 108216 275837 109712 275878
rect 108216 275765 108359 275837
rect 109193 275836 109712 275837
rect 102098 275691 102288 275701
rect 103064 275691 103259 275701
rect 102098 275531 103259 275691
rect 108187 275709 108393 275765
rect 108187 275593 108232 275709
rect 108348 275593 108393 275709
rect 108187 275522 108393 275593
rect 114865 275296 114970 275313
rect 114303 275290 114970 275296
rect 114303 275234 114888 275290
rect 114944 275234 114970 275290
rect 114303 275211 114970 275234
rect 102557 274069 105283 274145
rect 102557 274043 102644 274069
rect 105180 274043 105283 274069
rect 102557 273799 102638 274043
rect 105186 273799 105283 274043
rect 102557 273773 102644 273799
rect 105180 273773 105283 273799
rect 102557 273716 105283 273773
rect 114303 273212 114407 275211
rect 114865 275206 114970 275211
rect 115235 275304 115340 275313
rect 115788 275304 115900 276459
rect 115235 275290 115900 275304
rect 115235 275234 115260 275290
rect 115316 275234 115900 275290
rect 115235 275219 115900 275234
rect 115235 275206 115340 275219
rect 114843 274863 115030 274878
rect 114843 274807 114891 274863
rect 114947 274807 115030 274863
rect 114843 274793 115030 274807
rect 115175 274863 115362 274878
rect 115175 274807 115257 274863
rect 115314 274811 115362 274863
rect 115313 274807 115362 274811
rect 115175 274793 115362 274807
rect 114865 273632 114970 273647
rect 115235 273632 115340 273647
rect 114865 273624 115340 273632
rect 114865 273568 114888 273624
rect 114944 273568 115260 273624
rect 115316 273568 115340 273624
rect 114865 273554 115340 273568
rect 114865 273540 114970 273554
rect 115235 273540 115340 273554
rect 115209 273212 115899 273221
rect 114303 273197 115030 273212
rect 114303 273141 114891 273197
rect 114947 273141 115030 273197
rect 114303 273128 115030 273141
rect 114324 273127 115030 273128
rect 115175 273197 115899 273212
rect 115175 273141 115257 273197
rect 115314 273145 115899 273197
rect 115313 273141 115899 273145
rect 115175 273127 115899 273141
rect 115209 273107 115899 273127
rect 104687 272547 108128 272685
rect 115759 272659 115899 273107
rect 120953 272981 121018 276828
rect 120953 272929 120959 272981
rect 121011 272929 121018 272981
rect 120953 272917 121018 272929
rect 120953 272865 120959 272917
rect 121011 272865 121018 272917
rect 120953 272853 121018 272865
rect 120953 272801 120959 272853
rect 121011 272801 121018 272853
rect 120953 272789 121018 272801
rect 120953 272737 120959 272789
rect 121011 272737 121018 272789
rect 120953 272710 121018 272737
rect 115433 272645 115899 272659
rect 115433 272602 115898 272645
rect 104687 272454 108129 272547
rect 102092 271602 103253 271773
rect 102092 270826 102274 271602
rect 103050 271447 103253 271602
rect 104687 271447 104918 272454
rect 107985 272277 108129 272454
rect 107249 272207 108611 272277
rect 107249 271971 107351 272207
rect 108553 272113 108611 272207
rect 108553 272078 108841 272113
rect 108553 272026 108651 272078
rect 108703 272026 108715 272078
rect 108767 272026 108779 272078
rect 108831 272026 108841 272078
rect 115433 272048 115559 272602
rect 121587 272338 121677 277486
rect 121801 276207 121931 276287
rect 121801 276155 121841 276207
rect 121893 276155 121931 276207
rect 121801 276145 121931 276155
rect 121801 276143 121932 276145
rect 121801 276091 121841 276143
rect 121893 276091 121932 276143
rect 121801 276079 121932 276091
rect 121801 276027 121841 276079
rect 121893 276027 121932 276079
rect 121801 275945 121932 276027
rect 121802 273805 121932 275945
rect 121802 273753 121842 273805
rect 121894 273753 121932 273805
rect 121802 273741 121932 273753
rect 121802 273689 121842 273741
rect 121894 273689 121932 273741
rect 121802 273677 121932 273689
rect 121802 273625 121842 273677
rect 121894 273625 121932 273677
rect 121802 273253 121932 273625
rect 122077 273466 122191 277503
rect 122326 275317 122757 275386
rect 122326 274781 122402 275317
rect 122698 274781 122757 275317
rect 122326 274706 122757 274781
rect 122602 273466 122755 273468
rect 122077 273449 122755 273466
rect 123747 273449 123900 273468
rect 122077 273397 122652 273449
rect 122704 273402 123797 273449
rect 122704 273397 122755 273402
rect 122077 273390 122755 273397
rect 122602 273371 122755 273390
rect 123747 273397 123797 273402
rect 123849 273397 123900 273449
rect 123747 273371 123900 273397
rect 121802 273151 123740 273253
rect 121587 272286 121605 272338
rect 121657 272286 121677 272338
rect 121587 272274 121677 272286
rect 121587 272222 121605 272274
rect 121657 272222 121677 272274
rect 121587 272210 121677 272222
rect 121587 272158 121605 272210
rect 121657 272158 121677 272210
rect 121587 272146 121677 272158
rect 121587 272094 121605 272146
rect 121657 272094 121677 272146
rect 121587 272082 121677 272094
rect 108553 271995 108841 272026
rect 114761 272004 115601 272048
rect 107249 271949 107401 271971
rect 107249 271897 107300 271949
rect 107352 271897 107401 271949
rect 107249 271885 107401 271897
rect 107249 271833 107300 271885
rect 107352 271833 107401 271885
rect 107249 271807 107401 271833
rect 114761 271824 114830 272004
rect 115522 271824 115601 272004
rect 114761 271763 115601 271824
rect 121587 272030 121605 272082
rect 121657 272030 121677 272082
rect 121587 272018 121677 272030
rect 121587 271966 121605 272018
rect 121657 271966 121677 272018
rect 123362 272178 123476 272233
rect 123362 272126 123395 272178
rect 123447 272126 123476 272178
rect 123362 272114 123476 272126
rect 123362 272062 123395 272114
rect 123447 272062 123476 272114
rect 123362 272007 123476 272062
rect 121587 271954 121677 271966
rect 121587 271902 121605 271954
rect 121657 271902 121677 271954
rect 121587 271890 121677 271902
rect 121587 271838 121605 271890
rect 121657 271838 121677 271890
rect 121587 271826 121677 271838
rect 121587 271774 121605 271826
rect 121657 271774 121677 271826
rect 121587 271762 121677 271774
rect 121587 271710 121605 271762
rect 121657 271710 121677 271762
rect 121587 271698 121677 271710
rect 121587 271646 121605 271698
rect 121657 271646 121677 271698
rect 121587 271634 121677 271646
rect 121587 271582 121605 271634
rect 121657 271582 121677 271634
rect 121587 271570 121677 271582
rect 121587 271518 121605 271570
rect 121657 271518 121677 271570
rect 121587 271506 121677 271518
rect 103050 271216 104918 271447
rect 106951 271458 107141 271485
rect 106951 271406 107049 271458
rect 107101 271406 107141 271458
rect 106951 271394 107141 271406
rect 106951 271342 107049 271394
rect 107101 271342 107141 271394
rect 106951 271315 107141 271342
rect 108405 271458 108507 271485
rect 108405 271406 108445 271458
rect 108497 271406 108507 271458
rect 108405 271394 108507 271406
rect 108405 271342 108445 271394
rect 108497 271342 108507 271394
rect 108405 271315 108507 271342
rect 106951 271304 107095 271315
rect 106951 271252 106967 271304
rect 107019 271252 107095 271304
rect 106951 271240 107095 271252
rect 103050 270826 103253 271216
rect 106951 271188 106967 271240
rect 107019 271188 107095 271240
rect 106951 271176 107095 271188
rect 106951 271124 106967 271176
rect 107019 271124 107095 271176
rect 106951 271115 107095 271124
rect 108451 271115 108507 271315
rect 106951 271088 107141 271115
rect 106951 271036 107049 271088
rect 107101 271036 107141 271088
rect 106951 271024 107141 271036
rect 106951 270972 107049 271024
rect 107101 270972 107141 271024
rect 106951 270945 107141 270972
rect 108405 271088 108507 271115
rect 108405 271036 108445 271088
rect 108497 271036 108507 271088
rect 108405 271024 108507 271036
rect 108405 270972 108445 271024
rect 108497 270972 108507 271024
rect 108405 270945 108507 270972
rect 121587 271454 121605 271506
rect 121657 271454 121677 271506
rect 121587 271442 121677 271454
rect 121587 271390 121605 271442
rect 121657 271390 121677 271442
rect 121587 271378 121677 271390
rect 121587 271326 121605 271378
rect 121657 271326 121677 271378
rect 121587 271314 121677 271326
rect 121587 271262 121605 271314
rect 121657 271262 121677 271314
rect 121587 271250 121677 271262
rect 121587 271198 121605 271250
rect 121657 271198 121677 271250
rect 121587 271186 121677 271198
rect 121587 271134 121605 271186
rect 121657 271134 121677 271186
rect 121587 271122 121677 271134
rect 121587 271070 121605 271122
rect 121657 271070 121677 271122
rect 121587 271058 121677 271070
rect 121587 271006 121605 271058
rect 121657 271006 121677 271058
rect 121587 270994 121677 271006
rect 102092 270683 103253 270826
rect 121587 270942 121605 270994
rect 121657 270942 121677 270994
rect 121587 270930 121677 270942
rect 121587 270878 121605 270930
rect 121657 270878 121677 270930
rect 121587 270866 121677 270878
rect 121587 270814 121605 270866
rect 121657 270814 121677 270866
rect 121587 270802 121677 270814
rect 121587 270750 121605 270802
rect 121657 270750 121677 270802
rect 121587 270738 121677 270750
rect 112194 270648 113508 270715
rect 112194 270468 112288 270648
rect 113428 270468 113508 270648
rect 112194 270399 113508 270468
rect 121587 270686 121605 270738
rect 121657 270686 121677 270738
rect 121587 270674 121677 270686
rect 121587 270622 121605 270674
rect 121657 270622 121677 270674
rect 121587 270610 121677 270622
rect 121587 270558 121605 270610
rect 121657 270558 121677 270610
rect 121587 270546 121677 270558
rect 121587 270494 121605 270546
rect 121657 270494 121677 270546
rect 121587 270482 121677 270494
rect 121587 270430 121605 270482
rect 121657 270430 121677 270482
rect 112198 267513 112378 270399
rect 121587 270345 121677 270430
rect 123381 269864 123456 272007
rect 123629 271620 123739 273151
rect 124813 273071 124957 280498
rect 124634 273033 124957 273071
rect 124634 272853 124676 273033
rect 124920 272853 124957 273033
rect 124634 272849 124957 272853
rect 125452 275138 128452 275523
rect 125452 275136 125814 275138
rect 128030 275136 128452 275138
rect 124634 272811 124956 272849
rect 123629 271526 124017 271620
rect 123629 271524 123739 271526
rect 123940 271093 124017 271526
rect 123931 271031 124081 271093
rect 123931 270979 123986 271031
rect 124038 270979 124081 271031
rect 123931 270967 124081 270979
rect 123931 270915 123986 270967
rect 124038 270915 124081 270967
rect 123931 270903 124081 270915
rect 123931 270851 123986 270903
rect 124038 270851 124081 270903
rect 123931 270839 124081 270851
rect 123931 270787 123986 270839
rect 124038 270787 124081 270839
rect 123931 270717 124081 270787
rect 123360 269811 123474 269864
rect 123360 269759 123392 269811
rect 123444 269759 123474 269811
rect 123360 269747 123474 269759
rect 123360 269695 123392 269747
rect 123444 269695 123474 269747
rect 123360 269638 123474 269695
rect 125452 268364 125808 275136
rect 128036 268364 128452 275136
rect 125452 268362 125814 268364
rect 128030 268362 128452 268364
rect 125452 268022 128452 268362
rect 112198 267440 116858 267513
rect 112198 267384 112256 267440
rect 112312 267384 112336 267440
rect 112392 267384 112416 267440
rect 112472 267384 112496 267440
rect 112552 267384 112576 267440
rect 112632 267384 112656 267440
rect 112712 267384 112736 267440
rect 112792 267384 112816 267440
rect 112872 267384 112896 267440
rect 112952 267384 112976 267440
rect 113032 267384 113056 267440
rect 113112 267384 113136 267440
rect 113192 267384 113216 267440
rect 113272 267384 113296 267440
rect 113352 267384 113376 267440
rect 113432 267384 113456 267440
rect 113512 267384 113536 267440
rect 113592 267384 113616 267440
rect 113672 267384 113696 267440
rect 113752 267384 113776 267440
rect 113832 267384 113856 267440
rect 113912 267384 113936 267440
rect 113992 267384 114016 267440
rect 114072 267384 114096 267440
rect 114152 267384 114176 267440
rect 114232 267384 114256 267440
rect 114312 267384 114336 267440
rect 114392 267384 114416 267440
rect 114472 267384 114496 267440
rect 114552 267384 114576 267440
rect 114632 267384 114656 267440
rect 114712 267384 114736 267440
rect 114792 267384 114816 267440
rect 114872 267384 114896 267440
rect 114952 267384 114976 267440
rect 115032 267384 115056 267440
rect 115112 267384 115136 267440
rect 115192 267384 115216 267440
rect 115272 267384 115296 267440
rect 115352 267384 115376 267440
rect 115432 267384 115456 267440
rect 115512 267384 115536 267440
rect 115592 267384 115616 267440
rect 115672 267384 115696 267440
rect 115752 267384 115776 267440
rect 115832 267384 115856 267440
rect 115912 267384 115936 267440
rect 115992 267384 116016 267440
rect 116072 267384 116096 267440
rect 116152 267384 116176 267440
rect 116232 267384 116256 267440
rect 116312 267384 116336 267440
rect 116392 267384 116416 267440
rect 116472 267384 116496 267440
rect 116552 267384 116576 267440
rect 116632 267384 116656 267440
rect 116712 267384 116736 267440
rect 116792 267384 116858 267440
rect 112198 267333 116858 267384
rect 104286 266550 111587 266766
rect 104286 265534 104479 266550
rect 111335 265534 111587 266550
rect 104286 265368 111587 265534
<< via2 >>
rect 106149 282460 106167 283636
rect 106167 282460 113387 283636
rect 113387 282460 113405 283636
rect 102254 281628 103110 281638
rect 102254 280872 102272 281628
rect 102272 280872 103092 281628
rect 103092 280872 103110 281628
rect 102254 280862 103110 280872
rect 114888 280286 114944 280288
rect 114888 280234 114890 280286
rect 114890 280234 114942 280286
rect 114942 280234 114944 280286
rect 114888 280232 114944 280234
rect 115260 280286 115316 280288
rect 115260 280234 115262 280286
rect 115262 280234 115314 280286
rect 115314 280234 115316 280286
rect 115260 280232 115316 280234
rect 114891 279809 114943 279861
rect 114943 279809 114947 279861
rect 114891 279805 114947 279809
rect 115257 279809 115262 279861
rect 115262 279809 115313 279861
rect 115257 279805 115313 279809
rect 114888 278620 114944 278622
rect 114888 278568 114890 278620
rect 114890 278568 114942 278620
rect 114942 278568 114944 278620
rect 114888 278566 114944 278568
rect 107023 277722 107479 277748
rect 107023 277478 107033 277722
rect 107033 277478 107469 277722
rect 107469 277478 107479 277722
rect 107023 277452 107479 277478
rect 102288 276457 103064 276467
rect 102288 275701 103064 276457
rect 109356 277223 109466 277262
rect 109466 277223 109492 277262
rect 109356 277211 109492 277223
rect 109356 277159 109466 277211
rect 109466 277159 109492 277211
rect 109356 277147 109492 277159
rect 109356 277095 109466 277147
rect 109466 277095 109492 277147
rect 109356 277083 109492 277095
rect 109356 277031 109466 277083
rect 109466 277031 109492 277083
rect 109356 277019 109492 277031
rect 109356 276967 109466 277019
rect 109466 276967 109492 277019
rect 109356 276955 109492 276967
rect 109356 276903 109466 276955
rect 109466 276903 109492 276955
rect 109356 276891 109492 276903
rect 109356 276839 109466 276891
rect 109466 276839 109492 276891
rect 109356 276827 109492 276839
rect 109356 276775 109466 276827
rect 109466 276775 109492 276827
rect 109356 276763 109492 276775
rect 109356 276726 109466 276763
rect 109466 276726 109492 276763
rect 115260 278620 115316 278622
rect 115260 278568 115262 278620
rect 115262 278568 115314 278620
rect 115314 278568 115316 278620
rect 115260 278566 115316 278568
rect 114891 278143 114943 278195
rect 114943 278143 114947 278195
rect 114891 278139 114947 278143
rect 115257 278143 115262 278195
rect 115262 278143 115313 278195
rect 115257 278139 115313 278143
rect 114888 276954 114944 276956
rect 114888 276902 114890 276954
rect 114890 276902 114942 276954
rect 114942 276902 114944 276954
rect 114888 276900 114944 276902
rect 115260 276954 115316 276956
rect 115260 276902 115262 276954
rect 115262 276902 115314 276954
rect 115314 276902 115316 276954
rect 115260 276900 115316 276902
rect 114891 276477 114943 276529
rect 114943 276477 114947 276529
rect 114891 276473 114947 276477
rect 115257 276477 115262 276529
rect 115262 276477 115313 276529
rect 115257 276473 115313 276477
rect 109475 276180 109611 276316
rect 102288 275691 103064 275701
rect 114888 275288 114944 275290
rect 114888 275236 114890 275288
rect 114890 275236 114942 275288
rect 114942 275236 114944 275288
rect 114888 275234 114944 275236
rect 102644 274043 105180 274069
rect 102644 273799 105180 274043
rect 102644 273773 105180 273799
rect 115260 275288 115316 275290
rect 115260 275236 115262 275288
rect 115262 275236 115314 275288
rect 115314 275236 115316 275288
rect 115260 275234 115316 275236
rect 114891 274811 114943 274863
rect 114943 274811 114947 274863
rect 114891 274807 114947 274811
rect 115257 274811 115262 274863
rect 115262 274811 115313 274863
rect 115257 274807 115313 274811
rect 114888 273622 114944 273624
rect 114888 273570 114890 273622
rect 114890 273570 114942 273622
rect 114942 273570 114944 273622
rect 114888 273568 114944 273570
rect 115260 273622 115316 273624
rect 115260 273570 115262 273622
rect 115262 273570 115314 273622
rect 115314 273570 115316 273622
rect 115260 273568 115316 273570
rect 114891 273145 114943 273197
rect 114943 273145 114947 273197
rect 114891 273141 114947 273145
rect 115257 273145 115262 273197
rect 115262 273145 115313 273197
rect 115257 273141 115313 273145
rect 102274 270826 103050 271602
rect 122402 275286 122698 275317
rect 122402 274786 122415 275286
rect 122415 274786 122531 275286
rect 122531 274786 122698 275286
rect 122402 274781 122698 274786
rect 125814 275136 128030 275138
rect 125814 268364 128030 275136
rect 125814 268362 128030 268364
rect 112256 267384 112312 267440
rect 112336 267384 112392 267440
rect 112416 267384 112472 267440
rect 112496 267384 112552 267440
rect 112576 267384 112632 267440
rect 112656 267384 112712 267440
rect 112736 267384 112792 267440
rect 112816 267384 112872 267440
rect 112896 267384 112952 267440
rect 112976 267384 113032 267440
rect 113056 267384 113112 267440
rect 113136 267384 113192 267440
rect 113216 267384 113272 267440
rect 113296 267384 113352 267440
rect 113376 267384 113432 267440
rect 113456 267384 113512 267440
rect 113536 267384 113592 267440
rect 113616 267384 113672 267440
rect 113696 267384 113752 267440
rect 113776 267384 113832 267440
rect 113856 267384 113912 267440
rect 113936 267384 113992 267440
rect 114016 267384 114072 267440
rect 114096 267384 114152 267440
rect 114176 267384 114232 267440
rect 114256 267384 114312 267440
rect 114336 267384 114392 267440
rect 114416 267384 114472 267440
rect 114496 267384 114552 267440
rect 114576 267384 114632 267440
rect 114656 267384 114712 267440
rect 114736 267384 114792 267440
rect 114816 267384 114872 267440
rect 114896 267384 114952 267440
rect 114976 267384 115032 267440
rect 115056 267384 115112 267440
rect 115136 267384 115192 267440
rect 115216 267384 115272 267440
rect 115296 267384 115352 267440
rect 115376 267384 115432 267440
rect 115456 267384 115512 267440
rect 115536 267384 115592 267440
rect 115616 267384 115672 267440
rect 115696 267384 115752 267440
rect 115776 267384 115832 267440
rect 115856 267384 115912 267440
rect 115936 267384 115992 267440
rect 116016 267384 116072 267440
rect 116096 267384 116152 267440
rect 116176 267384 116232 267440
rect 116256 267384 116312 267440
rect 116336 267384 116392 267440
rect 116416 267384 116472 267440
rect 116496 267384 116552 267440
rect 116576 267384 116632 267440
rect 116656 267384 116712 267440
rect 116736 267384 116792 267440
rect 104479 266548 111335 266550
rect 104479 265536 104489 266548
rect 104489 265536 111325 266548
rect 111325 265536 111335 266548
rect 104479 265534 111335 265536
<< metal3 >>
rect 572176 406600 582975 406686
rect 572176 406488 583606 406600
rect 572176 406300 582975 406488
rect 572176 374237 572562 406300
rect 154704 373851 572562 374237
rect 5373 337581 128286 337911
rect 344 337472 128286 337581
rect 5373 336821 128286 337472
rect 2990 294360 109888 295024
rect 342 294248 109888 294360
rect 2990 293144 109888 294248
rect 106790 283895 109888 293144
rect 105796 283636 113672 283895
rect 105796 282460 106149 283636
rect 113405 282460 113672 283636
rect 105796 282251 113672 282460
rect 127196 281912 128286 336821
rect 102098 281808 103259 281810
rect 6645 281638 103259 281808
rect 6645 280862 102254 281638
rect 103110 280862 103259 281638
rect 6645 280720 103259 280862
rect 127196 280822 128357 281912
rect 6645 280718 102170 280720
rect 6645 251338 7735 280718
rect 101936 280716 102170 280718
rect 114841 280294 114994 280329
rect 114303 280288 114994 280294
rect 114303 280232 114888 280288
rect 114944 280232 114994 280288
rect 114303 280209 114994 280232
rect 106368 279497 109401 279505
rect 102586 279375 109401 279497
rect 102586 279266 106453 279375
rect 102586 279087 102817 279266
rect 107943 279238 109115 279266
rect 107943 279174 107963 279238
rect 108027 279174 109115 279238
rect 107943 279158 109115 279174
rect 107943 279094 107963 279158
rect 108027 279094 109115 279158
rect 342 251226 7735 251338
rect 6645 251087 7735 251226
rect 31331 277997 103259 279087
rect 107943 279078 109115 279094
rect 107943 279014 107963 279078
rect 108027 279014 109115 279078
rect 107943 278998 109115 279014
rect 107943 278934 107963 278998
rect 108027 278934 109115 278998
rect 107943 278918 109115 278934
rect 107943 278854 107963 278918
rect 108027 278854 109115 278918
rect 107943 278838 109115 278854
rect 107943 278774 107963 278838
rect 108027 278774 109115 278838
rect 107943 278758 109115 278774
rect 107943 278694 107963 278758
rect 108027 278694 109115 278758
rect 107943 278678 109115 278694
rect 107943 278614 107963 278678
rect 108027 278614 109115 278678
rect 107943 278598 109115 278614
rect 107943 278534 107963 278598
rect 108027 278534 109115 278598
rect 107943 278518 109115 278534
rect 107943 278454 107963 278518
rect 108027 278454 109115 278518
rect 107943 278438 109115 278454
rect 107943 278374 107963 278438
rect 108027 278374 109115 278438
rect 107943 278358 109115 278374
rect 107943 278294 107963 278358
rect 108027 278294 109115 278358
rect 107943 278278 109115 278294
rect 107943 278214 107963 278278
rect 108027 278214 109115 278278
rect 107943 278198 109115 278214
rect 107943 278134 107963 278198
rect 108027 278134 109115 278198
rect 107943 278118 109115 278134
rect 107943 278054 107963 278118
rect 108027 278054 109115 278118
rect 107943 278038 109115 278054
rect 31331 124117 32421 277997
rect 107943 277974 107963 278038
rect 108027 277974 109115 278038
rect 107943 277958 109115 277974
rect 107943 277894 107963 277958
rect 108027 277894 109115 277958
rect 107943 277878 109115 277894
rect 107943 277814 107963 277878
rect 108027 277814 109115 277878
rect 106957 277748 107553 277799
rect 106957 277712 107023 277748
rect 107479 277712 107553 277748
rect 106957 277488 107019 277712
rect 107483 277488 107553 277712
rect 106957 277452 107023 277488
rect 107479 277452 107553 277488
rect 106957 277403 107553 277452
rect 107943 277798 109115 277814
rect 107943 277734 107963 277798
rect 108027 277734 109115 277798
rect 107943 277718 109115 277734
rect 107943 277654 107963 277718
rect 108027 277654 109115 277718
rect 107943 277638 109115 277654
rect 107943 277574 107963 277638
rect 108027 277574 109115 277638
rect 107943 277558 109115 277574
rect 107943 277494 107963 277558
rect 108027 277494 109115 277558
rect 107943 277478 109115 277494
rect 107943 277414 107963 277478
rect 108027 277414 109115 277478
rect 107943 277398 109115 277414
rect 107943 277334 107963 277398
rect 108027 277334 109115 277398
rect 107943 277318 109115 277334
rect 107943 277254 107963 277318
rect 108027 277254 109115 277318
rect 107943 277238 109115 277254
rect 107943 277174 107963 277238
rect 108027 277174 109115 277238
rect 107943 277158 109115 277174
rect 107943 277094 107963 277158
rect 108027 277094 109115 277158
rect 107943 277078 109115 277094
rect 107943 277014 107963 277078
rect 108027 277014 109115 277078
rect 107943 276998 109115 277014
rect 107943 276934 107963 276998
rect 108027 276934 109115 276998
rect 107943 276918 109115 276934
rect 107943 276854 107963 276918
rect 108027 276854 109115 276918
rect 107943 276838 109115 276854
rect 107943 276774 107963 276838
rect 108027 276774 109115 276838
rect 107943 276758 109115 276774
rect 107943 276694 107963 276758
rect 108027 276694 109115 276758
rect 107943 276678 109115 276694
rect 102098 276620 103259 276621
rect 3945 123716 32421 124117
rect 326 123604 32421 123716
rect 3945 123027 32421 123604
rect 61553 276467 103259 276620
rect 61553 275691 102288 276467
rect 103064 275691 103259 276467
rect 107943 276614 107963 276678
rect 108027 276614 109115 276678
rect 109276 277341 109401 279375
rect 114303 278210 114407 280209
rect 114841 280178 114994 280209
rect 115211 280288 115364 280329
rect 115211 280232 115260 280288
rect 115316 280232 115364 280288
rect 115211 280178 115364 280232
rect 123842 279968 124731 280304
rect 127248 279968 127999 280822
rect 114843 279861 115030 279876
rect 114843 279805 114891 279861
rect 114947 279805 115030 279861
rect 114843 279791 115030 279805
rect 115175 279861 115362 279876
rect 115175 279805 115257 279861
rect 115313 279805 115362 279861
rect 115175 279791 115362 279805
rect 123842 279217 127999 279968
rect 123842 278876 124731 279217
rect 114841 278622 114994 278663
rect 114841 278566 114888 278622
rect 114944 278566 114994 278622
rect 114841 278512 114994 278566
rect 115211 278622 115364 278663
rect 115211 278566 115260 278622
rect 115316 278566 115364 278622
rect 115211 278512 115364 278566
rect 114303 278195 115030 278210
rect 114303 278139 114891 278195
rect 114947 278139 115030 278195
rect 114303 278126 115030 278139
rect 114324 278125 115030 278126
rect 115175 278195 115903 278210
rect 115175 278139 115257 278195
rect 115313 278139 115903 278195
rect 115175 278125 115903 278139
rect 109276 277262 109568 277341
rect 109276 276726 109356 277262
rect 109492 276726 109568 277262
rect 114841 276962 114994 276997
rect 109276 276633 109568 276726
rect 114303 276956 114994 276962
rect 114303 276900 114888 276956
rect 114944 276900 114994 276956
rect 114303 276877 114994 276900
rect 107943 276598 109115 276614
rect 107943 276534 107963 276598
rect 108027 276534 109115 276598
rect 107943 276518 109115 276534
rect 107943 276454 107963 276518
rect 108027 276454 109115 276518
rect 107943 276438 109115 276454
rect 107943 276374 107963 276438
rect 108027 276374 109115 276438
rect 107943 276358 109115 276374
rect 107943 276294 107963 276358
rect 108027 276294 109115 276358
rect 107943 276278 109115 276294
rect 107943 276214 107963 276278
rect 108027 276214 109115 276278
rect 107943 276186 109115 276214
rect 109383 276320 109700 276394
rect 109383 276176 109471 276320
rect 109615 276176 109700 276320
rect 109383 276091 109700 276176
rect 61553 275531 103259 275691
rect 61553 275530 102104 275531
rect 61553 80603 62643 275530
rect 114303 274878 114407 276877
rect 114841 276846 114994 276877
rect 115211 276972 115364 276997
rect 115791 276972 115903 278125
rect 124547 278165 124731 278876
rect 124547 277887 125086 278165
rect 115211 276956 115903 276972
rect 115211 276900 115260 276956
rect 115316 276900 115903 276956
rect 115211 276887 115903 276900
rect 115211 276846 115364 276887
rect 114843 276529 115030 276544
rect 114843 276473 114891 276529
rect 114947 276473 115030 276529
rect 114843 276459 115030 276473
rect 115175 276529 115362 276544
rect 115175 276473 115257 276529
rect 115313 276473 115362 276529
rect 115175 276459 115362 276473
rect 122326 275377 122757 275386
rect 124892 275377 125086 277887
rect 114841 275290 114994 275331
rect 114841 275234 114888 275290
rect 114944 275234 114994 275290
rect 114841 275180 114994 275234
rect 115211 275290 115364 275331
rect 115211 275234 115260 275290
rect 115316 275234 115364 275290
rect 115211 275180 115364 275234
rect 122326 275317 125086 275377
rect 114303 274863 115030 274878
rect 114303 274807 114891 274863
rect 114947 274807 115030 274863
rect 114303 274794 115030 274807
rect 114324 274793 115030 274794
rect 115175 274877 115362 274878
rect 115175 274863 115902 274877
rect 115175 274807 115257 274863
rect 115313 274807 115902 274863
rect 115175 274793 115902 274807
rect 115214 274792 115902 274793
rect 1853 80494 62643 80603
rect 342 80382 62643 80494
rect 1853 79513 62643 80382
rect 74033 274145 102558 274146
rect 74033 274069 105283 274145
rect 74033 273773 102644 274069
rect 105180 273773 105283 274069
rect 74033 273716 105283 273773
rect 1115 37272 4017 37406
rect 342 37245 4017 37272
rect 74033 37245 74463 273716
rect 114841 273624 114994 273665
rect 114841 273568 114888 273624
rect 114944 273568 114994 273624
rect 114841 273514 114994 273568
rect 115211 273635 115364 273665
rect 115790 273635 115902 274792
rect 122326 274781 122402 275317
rect 122698 275090 125086 275317
rect 125452 275138 128452 275523
rect 122698 274781 122757 275090
rect 122326 274706 122757 274781
rect 115211 273624 115902 273635
rect 115211 273568 115260 273624
rect 115316 273568 115902 273624
rect 115211 273550 115902 273568
rect 115211 273514 115364 273550
rect 114843 273197 115030 273212
rect 114843 273141 114891 273197
rect 114947 273141 115030 273197
rect 114843 273127 115030 273141
rect 115175 273197 115362 273212
rect 115175 273141 115257 273197
rect 115313 273141 115362 273197
rect 115175 273127 115362 273141
rect 342 37160 74463 37245
rect 1115 36815 74463 37160
rect 87083 271602 103253 271773
rect 87083 270826 102274 271602
rect 103050 270826 103253 271602
rect 87083 270683 103253 270826
rect 1115 36682 4017 36815
rect 87083 16181 88173 270683
rect 125452 268362 125814 275138
rect 128030 274476 128452 275138
rect 134328 274476 139500 350418
rect 128030 269304 139500 274476
rect 128030 268362 128452 269304
rect 125452 268022 128452 268362
rect 112198 267440 116858 267513
rect 112198 267384 112256 267440
rect 112312 267384 112336 267440
rect 112392 267384 112416 267440
rect 112472 267384 112496 267440
rect 112552 267384 112576 267440
rect 112632 267384 112656 267440
rect 112712 267384 112736 267440
rect 112792 267384 112816 267440
rect 112872 267384 112896 267440
rect 112952 267384 112976 267440
rect 113032 267384 113056 267440
rect 113112 267384 113136 267440
rect 113192 267384 113216 267440
rect 113272 267384 113296 267440
rect 113352 267384 113376 267440
rect 113432 267384 113456 267440
rect 113512 267384 113536 267440
rect 113592 267384 113616 267440
rect 113672 267384 113696 267440
rect 113752 267384 113776 267440
rect 113832 267384 113856 267440
rect 113912 267384 113936 267440
rect 113992 267384 114016 267440
rect 114072 267384 114096 267440
rect 114152 267384 114176 267440
rect 114232 267384 114256 267440
rect 114312 267384 114336 267440
rect 114392 267384 114416 267440
rect 114472 267384 114496 267440
rect 114552 267384 114576 267440
rect 114632 267384 114656 267440
rect 114712 267384 114736 267440
rect 114792 267384 114816 267440
rect 114872 267384 114896 267440
rect 114952 267384 114976 267440
rect 115032 267384 115056 267440
rect 115112 267384 115136 267440
rect 115192 267384 115216 267440
rect 115272 267384 115296 267440
rect 115352 267384 115376 267440
rect 115432 267384 115456 267440
rect 115512 267384 115536 267440
rect 115592 267384 115616 267440
rect 115672 267384 115696 267440
rect 115752 267384 115776 267440
rect 115832 267384 115856 267440
rect 115912 267384 115936 267440
rect 115992 267384 116016 267440
rect 116072 267384 116096 267440
rect 116152 267384 116176 267440
rect 116232 267384 116256 267440
rect 116312 267384 116336 267440
rect 116392 267384 116416 267440
rect 116472 267384 116496 267440
rect 116552 267384 116576 267440
rect 116632 267384 116656 267440
rect 116712 267384 116736 267440
rect 116792 267384 116858 267440
rect 112198 267333 116858 267384
rect 104286 266550 111587 266766
rect 104286 265534 104479 266550
rect 111335 265534 111587 266550
rect 104286 265368 111587 265534
rect 106618 236639 109716 265368
rect 115987 257334 116373 267333
rect 154704 257334 155090 373851
rect 115987 256948 155090 257334
rect 162337 364696 578379 366371
rect 162337 364584 581142 364696
rect 162337 363273 578379 364584
rect 162337 236639 165435 363273
rect 581030 360178 581142 364584
rect 581030 360066 583606 360178
rect 106618 233541 165435 236639
rect 1455 15850 88173 16181
rect 342 15738 88173 15850
rect 1455 15091 88173 15738
<< via3 >>
rect 107963 279174 108027 279238
rect 107963 279094 108027 279158
rect 107963 279014 108027 279078
rect 107963 278934 108027 278998
rect 107963 278854 108027 278918
rect 107963 278774 108027 278838
rect 107963 278694 108027 278758
rect 107963 278614 108027 278678
rect 107963 278534 108027 278598
rect 107963 278454 108027 278518
rect 107963 278374 108027 278438
rect 107963 278294 108027 278358
rect 107963 278214 108027 278278
rect 107963 278134 108027 278198
rect 107963 278054 108027 278118
rect 107963 277974 108027 278038
rect 107963 277894 108027 277958
rect 107963 277814 108027 277878
rect 107019 277488 107023 277712
rect 107023 277488 107479 277712
rect 107479 277488 107483 277712
rect 107963 277734 108027 277798
rect 107963 277654 108027 277718
rect 107963 277574 108027 277638
rect 107963 277494 108027 277558
rect 107963 277414 108027 277478
rect 107963 277334 108027 277398
rect 107963 277254 108027 277318
rect 107963 277174 108027 277238
rect 107963 277094 108027 277158
rect 107963 277014 108027 277078
rect 107963 276934 108027 276998
rect 107963 276854 108027 276918
rect 107963 276774 108027 276838
rect 107963 276694 108027 276758
rect 107963 276614 108027 276678
rect 107963 276534 108027 276598
rect 107963 276454 108027 276518
rect 107963 276374 108027 276438
rect 107963 276294 108027 276358
rect 107963 276214 108027 276278
rect 109471 276316 109615 276320
rect 109471 276180 109475 276316
rect 109475 276180 109611 276316
rect 109611 276180 109615 276316
rect 109471 276176 109615 276180
<< mimcap >>
rect 108275 279158 109075 279226
rect 108275 276294 108323 279158
rect 109027 276294 109075 279158
rect 108275 276226 109075 276294
<< mimcapcontact >>
rect 108323 276294 109027 279158
<< metal4 >>
rect 107947 279238 108043 279254
rect 107947 279174 107963 279238
rect 108027 279174 108043 279238
rect 107947 279158 108043 279174
rect 107947 279094 107963 279158
rect 108027 279094 108043 279158
rect 107947 279078 108043 279094
rect 107947 279014 107963 279078
rect 108027 279014 108043 279078
rect 107947 278998 108043 279014
rect 107947 278934 107963 278998
rect 108027 278934 108043 278998
rect 107947 278918 108043 278934
rect 107947 278854 107963 278918
rect 108027 278854 108043 278918
rect 107947 278838 108043 278854
rect 107947 278774 107963 278838
rect 108027 278774 108043 278838
rect 107947 278758 108043 278774
rect 107947 278694 107963 278758
rect 108027 278694 108043 278758
rect 107947 278678 108043 278694
rect 107947 278614 107963 278678
rect 108027 278614 108043 278678
rect 107947 278598 108043 278614
rect 107947 278534 107963 278598
rect 108027 278534 108043 278598
rect 107947 278518 108043 278534
rect 107947 278454 107963 278518
rect 108027 278454 108043 278518
rect 107947 278438 108043 278454
rect 107947 278374 107963 278438
rect 108027 278374 108043 278438
rect 107947 278358 108043 278374
rect 107947 278294 107963 278358
rect 108027 278294 108043 278358
rect 107947 278278 108043 278294
rect 107947 278214 107963 278278
rect 108027 278214 108043 278278
rect 107947 278198 108043 278214
rect 107947 278134 107963 278198
rect 108027 278134 108043 278198
rect 107947 278118 108043 278134
rect 107947 278054 107963 278118
rect 108027 278054 108043 278118
rect 107947 278038 108043 278054
rect 107947 277974 107963 278038
rect 108027 277974 108043 278038
rect 107947 277958 108043 277974
rect 107947 277894 107963 277958
rect 108027 277894 108043 277958
rect 107947 277878 108043 277894
rect 107947 277814 107963 277878
rect 108027 277814 108043 277878
rect 106957 277737 107553 277799
rect 107947 277798 108043 277814
rect 107947 277737 107963 277798
rect 106957 277734 107963 277737
rect 108027 277734 108043 277798
rect 106957 277718 108043 277734
rect 106957 277712 107963 277718
rect 106957 277488 107019 277712
rect 107483 277654 107963 277712
rect 108027 277654 108043 277718
rect 107483 277638 108043 277654
rect 107483 277574 107963 277638
rect 108027 277574 108043 277638
rect 107483 277558 108043 277574
rect 107483 277494 107963 277558
rect 108027 277494 108043 277558
rect 107483 277488 108043 277494
rect 106957 277478 108043 277488
rect 106957 277477 107963 277478
rect 106957 277403 107553 277477
rect 107947 277414 107963 277477
rect 108027 277414 108043 277478
rect 107947 277398 108043 277414
rect 107947 277334 107963 277398
rect 108027 277334 108043 277398
rect 107947 277318 108043 277334
rect 107947 277254 107963 277318
rect 108027 277254 108043 277318
rect 107947 277238 108043 277254
rect 107947 277174 107963 277238
rect 108027 277174 108043 277238
rect 107947 277158 108043 277174
rect 107947 277094 107963 277158
rect 108027 277094 108043 277158
rect 107947 277078 108043 277094
rect 107947 277014 107963 277078
rect 108027 277014 108043 277078
rect 107947 276998 108043 277014
rect 107947 276934 107963 276998
rect 108027 276934 108043 276998
rect 107947 276918 108043 276934
rect 107947 276854 107963 276918
rect 108027 276854 108043 276918
rect 107947 276838 108043 276854
rect 107947 276774 107963 276838
rect 108027 276774 108043 276838
rect 107947 276758 108043 276774
rect 107947 276694 107963 276758
rect 108027 276694 108043 276758
rect 107947 276678 108043 276694
rect 107947 276614 107963 276678
rect 108027 276614 108043 276678
rect 107947 276598 108043 276614
rect 107947 276534 107963 276598
rect 108027 276534 108043 276598
rect 107947 276518 108043 276534
rect 107947 276454 107963 276518
rect 108027 276454 108043 276518
rect 107947 276438 108043 276454
rect 107947 276374 107963 276438
rect 108027 276374 108043 276438
rect 107947 276358 108043 276374
rect 107947 276294 107963 276358
rect 108027 276294 108043 276358
rect 107947 276278 108043 276294
rect 107947 276214 107963 276278
rect 108027 276214 108043 276278
rect 108314 279158 109036 279187
rect 108314 276294 108323 279158
rect 109027 276394 109036 279158
rect 109027 276320 109700 276394
rect 109027 276294 109471 276320
rect 108314 276265 109471 276294
rect 107947 276198 108043 276214
rect 109383 276176 109471 276265
rect 109615 276176 109700 276320
rect 109383 276091 109700 276176
<< labels >>
flabel metal2 s 112229 267697 112349 267811 0 FreeSans 4000 90 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ring_out
port 1 nsew
flabel metal1 s 111201 267695 111321 267809 0 FreeSans 4000 90 0 0 pmu_circuits_top_level_0/pmu_circuits_0.dd_02
port 2 nsew
flabel metal2 s 106605 272511 106725 272625 0 FreeSans 4000 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.vref
port 3 nsew
flabel metal1 s 106117 277553 106237 277667 0 FreeSans 4000 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ldo_out
port 4 nsew
flabel metal1 s 105863 278241 105937 278329 0 FreeSans 4000 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ldo_vs
port 5 nsew
flabel metal3 s 105859 279345 105933 279433 0 FreeSans 4000 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ldo_vb
port 6 nsew
flabel metal1 s 105821 281133 105895 281221 0 FreeSans 4000 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ldo_iref
port 7 nsew
flabel metal1 s 106163 282527 106237 282615 0 FreeSans 4000 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.dd_01
port 8 nsew
flabel locali s 125137 281485 125329 281667 0 FreeSans 4000 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ss
port 9 nsew
flabel metal3 s 125259 279535 125451 279717 0 FreeSans 4000 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.iref
port 10 nsew
flabel metal2 s 108523 272221 108591 272269 0 FreeSans 2000 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.vref01_0.VREF
port 11 nsew
flabel metal1 s 108587 270871 108655 270919 0 FreeSans 2000 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.vref01_0.DD
port 12 nsew
flabel locali s 106809 271879 106877 271927 0 FreeSans 2000 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.vref01_0.SS
port 13 nsew
flabel locali s 118007 272352 118355 272604 0 FreeSans 2000 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.SS
port 14 nsew
flabel metal1 s 113347 272304 113553 272494 0 FreeSans 2000 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.DD
port 15 nsew
flabel metal1 s 112489 270487 112617 270591 0 FreeSans 2000 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.ring_100mV_buffer_0.OUT
port 16 nsew
flabel metal2 s 114788 271797 114916 271901 0 FreeSans 2000 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.ring_100mV_buffer_0.IN
port 17 nsew
flabel metal1 s 113883 271822 114011 271926 0 FreeSans 2000 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.ring_100mV_buffer_0.DD
port 18 nsew
flabel locali s 119001 272134 119129 272238 0 FreeSans 2000 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.ring_100mV_buffer_0.SS
port 19 nsew
rlabel metal1 s 114297 279009 114372 279073 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_9.IN
port 20 nsew
rlabel locali s 113345 277680 113420 277744 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_9.SS
port 21 nsew
rlabel locali s 114959 277764 114997 277798 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_9.DD
port 22 nsew
rlabel metal1 s 112782 277799 112826 277838 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_9.OUT
port 23 nsew
rlabel metal1 s 115833 279009 115908 279073 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_8.IN
port 24 nsew
rlabel locali s 116785 277680 116860 277744 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_8.SS
port 25 nsew
rlabel locali s 115208 277764 115246 277798 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_8.DD
port 26 nsew
rlabel metal1 s 117379 277799 117423 277838 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_8.OUT
port 27 nsew
rlabel metal1 s 114297 277343 114372 277407 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_7.IN
port 28 nsew
rlabel locali s 113345 276014 113420 276078 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_7.SS
port 29 nsew
rlabel locali s 114959 276098 114997 276132 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_7.DD
port 30 nsew
rlabel metal1 s 112782 276133 112826 276172 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_7.OUT
port 31 nsew
rlabel metal1 s 115833 277343 115908 277407 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_6.IN
port 32 nsew
rlabel locali s 116785 276014 116860 276078 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_6.SS
port 33 nsew
rlabel locali s 115208 276098 115246 276132 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_6.DD
port 34 nsew
rlabel metal1 s 117379 276133 117423 276172 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_6.OUT
port 35 nsew
rlabel metal1 s 114297 275677 114372 275741 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_5.IN
port 36 nsew
rlabel locali s 113345 274348 113420 274412 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_5.SS
port 37 nsew
rlabel locali s 114959 274432 114997 274466 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_5.DD
port 38 nsew
rlabel metal1 s 112782 274467 112826 274506 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_5.OUT
port 39 nsew
rlabel metal1 s 115833 275677 115908 275741 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_4.IN
port 40 nsew
rlabel locali s 116785 274348 116860 274412 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_4.SS
port 41 nsew
rlabel locali s 115208 274432 115246 274466 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_4.DD
port 42 nsew
rlabel metal1 s 117379 274467 117423 274506 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_4.OUT
port 43 nsew
rlabel metal1 s 115833 274011 115908 274075 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_3.IN
port 44 nsew
rlabel locali s 116785 272682 116860 272746 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_3.SS
port 45 nsew
rlabel locali s 115208 272766 115246 272800 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_3.DD
port 46 nsew
rlabel metal1 s 117379 272801 117423 272840 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_3.OUT
port 47 nsew
rlabel metal1 s 114297 274011 114372 274075 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_2.IN
port 48 nsew
rlabel locali s 113345 272682 113420 272746 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_2.SS
port 49 nsew
rlabel locali s 114959 272766 114997 272800 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_2.DD
port 50 nsew
rlabel metal1 s 112782 272801 112826 272840 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_2.OUT
port 51 nsew
rlabel metal1 s 115833 280675 115908 280739 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_1.IN
port 52 nsew
rlabel locali s 116785 279346 116860 279410 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_1.SS
port 53 nsew
rlabel locali s 115208 279430 115246 279464 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_1.DD
port 54 nsew
rlabel metal1 s 117379 279465 117423 279504 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_1.OUT
port 55 nsew
rlabel metal1 s 114297 280675 114372 280739 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_0.IN
port 56 nsew
rlabel locali s 113345 279346 113420 279410 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_0.SS
port 57 nsew
rlabel locali s 114959 279430 114997 279464 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_0.DD
port 58 nsew
rlabel metal1 s 112782 279465 112826 279504 4 pmu_circuits_top_level_0/pmu_circuits_0.ring_100mV_0.mdls_inv_0.OUT
port 59 nsew
flabel metal1 s 108183 280591 108259 280679 0 FreeSans 2000 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ldo_0.Iref
port 60 nsew
flabel locali s 109921 279361 109997 279449 0 FreeSans 2000 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ldo_0.SS
port 61 nsew
flabel metal3 s 106173 279327 106347 279459 0 FreeSans 2000 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ldo_0.VB
port 62 nsew
flabel metal1 s 106071 278255 106121 278309 0 FreeSans 2000 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ldo_0.VS
port 63 nsew
flabel metal1 s 106327 277543 106527 277719 0 FreeSans 2000 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ldo_0.OUT
port 64 nsew
flabel metal1 s 106143 274775 106235 274891 0 FreeSans 2000 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.ldo_0.DD
port 65 nsew
flabel metal2 s 120471 280709 120701 280913 0 FreeSans 2000 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.iref_2nA_0.DD
port 66 nsew
flabel metal3 s 124171 279421 124401 279625 0 FreeSans 2000 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.iref_2nA_0.IREF
port 67 nsew
flabel locali s 123893 268977 124041 269141 0 FreeSans 2000 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.iref_2nA_0.SS
port 68 nsew
flabel locali s 122378 278528 122456 278606 0 FreeSans 2000 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.iref_2nA_0.iref_2nA_vref_0.DD
port 69 nsew
flabel locali s 122060 276558 122134 276644 0 FreeSans 2000 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.iref_2nA_0.iref_2nA_vref_0.SS
port 70 nsew
flabel metal1 s 124468 276546 124542 276632 0 FreeSans 2000 0 0 0 pmu_circuits_top_level_0/pmu_circuits_0.iref_2nA_0.iref_2nA_vref_0.VREF
port 71 nsew
rlabel metal2 s 121796 277545 121931 277755 4 pmu_circuits_top_level_0/pmu_circuits_0.iref_2nA_0.iref_2nA_mirrors_0.Ip2
port 72 nsew
rlabel metal1 s 121951 274874 122001 274947 4 pmu_circuits_top_level_0/pmu_circuits_0.iref_2nA_0.iref_2nA_mirrors_0.Iref
port 73 nsew
rlabel metal1 s 123719 270947 123769 271020 4 pmu_circuits_top_level_0/pmu_circuits_0.iref_2nA_0.iref_2nA_mirrors_0.Vg
port 74 nsew
rlabel metal2 s 123405 269727 123455 269800 4 pmu_circuits_top_level_0/pmu_circuits_0.iref_2nA_0.iref_2nA_mirrors_0.Ip1
port 75 nsew
rlabel locali s 124373 269012 124499 269117 4 pmu_circuits_top_level_0/pmu_circuits_0.iref_2nA_0.iref_2nA_mirrors_0.SS
port 76 nsew
rlabel locali s 121944 279849 122032 279923 4 pmu_circuits_top_level_0/pmu_circuits_0.iref_2nA_0.iref_2nA_mirrors_0.DD
port 77 nsew
rlabel metal1 s 124871 273456 124913 273514 4 pmu_circuits_top_level_0/pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Vg
port 78 nsew
rlabel metal1 s 123437 273648 123479 273706 4 pmu_circuits_top_level_0/pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip1
port 79 nsew
rlabel metal1 s 123851 273648 123893 273706 4 pmu_circuits_top_level_0/pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.Ip2
port 80 nsew
rlabel locali s 124019 274734 124061 274792 4 pmu_circuits_top_level_0/pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.SS
port 81 nsew
rlabel metal1 s 124223 274754 124265 274812 4 pmu_circuits_top_level_0/pmu_circuits_0.iref_2nA_0.iref_2nA_igenerator_0.VCTAT
port 82 nsew
flabel metal3 s 10028 336906 11894 337768 0 FreeSans 10000 0 0 0 gpio_noesd[11]
port 83 nsew
flabel metal3 s 9412 293530 11278 294392 0 FreeSans 10000 0 0 0 gpio_noesd[12]
port 84 nsew
flabel metal3 s 6760 251254 7466 251912 0 FreeSans 10000 0 0 0 gpio_noesd[13]
port 85 nsew
flabel metal3 s 7748 123292 8454 123950 0 FreeSans 10000 0 0 0 gpio_noesd[14]
port 86 nsew
flabel metal3 s 7280 79630 7986 80288 0 FreeSans 10000 0 0 0 gpio_noesd[15]
port 87 nsew
flabel metal3 s 6896 36870 8062 37110 0 FreeSans 10000 0 0 0 gpio_noesd[16]
port 88 nsew
flabel metal3 s 6686 15490 7852 15730 0 FreeSans 10000 0 0 0 gpio_noesd[17]
port 89 nsew
flabel metal3 s 573308 364318 574122 364838 0 FreeSans 10000 0 0 0 gpio_noesd[2]
port 90 nsew
flabel metal3 s 575802 406322 576204 406584 0 FreeSans 10000 0 0 0 gpio_noesd[3]
port 91 nsew
flabel metal3 s 135612 346104 138678 348766 0 FreeSans 16000 0 0 0 vssa1
port 92 nsew
<< end >>

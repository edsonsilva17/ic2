magic
tech sky130A
magscale 1 2
timestamp 1699064461
<< nwell >>
rect 164480 538267 166680 539827
rect 168280 538267 170480 539827
rect 171980 538267 174180 539827
rect 175480 538267 177680 539827
rect 179080 538267 181280 539827
rect 182380 538267 184580 539827
rect 185680 538267 187880 539827
rect 188980 538267 191180 539827
rect 157550 535677 162910 537917
rect 172172 529784 187520 530350
rect 172172 528696 187520 529262
rect 172172 527608 187520 528174
rect 172172 526520 187520 527086
rect 172172 525432 187520 525998
rect 172172 524344 187520 524910
rect 172172 523256 187520 523822
rect 172172 522168 187520 522734
rect 172172 521080 187520 521646
rect 172172 519992 187520 520558
rect 172172 518904 187520 519470
rect 172172 517816 187520 518382
rect 172172 516728 187520 517294
rect 172172 515640 187520 516206
<< pwell >>
rect 164500 539827 166680 541347
rect 168300 539827 170480 541347
rect 172000 539827 174180 541347
rect 175500 539827 177680 541347
rect 179100 539827 181280 541347
rect 182400 539827 184580 541347
rect 185700 539827 187880 541347
rect 189000 539827 191180 541347
rect 157550 537927 162910 538857
rect 164152 535867 166780 538147
rect 167924 535867 169280 538147
rect 171660 535867 172380 538147
rect 175178 535867 175580 538147
rect 178778 536427 179180 538147
rect 182078 536707 182480 538147
rect 185378 536847 185780 538147
rect 188678 536751 189080 538147
rect 164122 533527 166750 535807
rect 172239 530590 172273 530628
rect 172975 530590 173009 530628
rect 173067 530590 173101 530628
rect 174171 530590 174205 530628
rect 174722 530600 174746 530622
rect 175367 530590 175401 530628
rect 175458 530600 175482 530622
rect 177299 530590 177333 530628
rect 177485 530599 177517 530621
rect 178311 530590 178345 530628
rect 178587 530590 178621 530628
rect 179139 530590 179173 530628
rect 179231 530590 179265 530628
rect 179785 530599 179817 530621
rect 180061 530599 180093 530621
rect 180298 530590 180332 530628
rect 181070 530600 181094 530622
rect 181844 530590 181878 530628
rect 181991 530590 182025 530628
rect 182635 530590 182669 530628
rect 183002 530600 183026 530622
rect 183095 530590 183129 530628
rect 183647 530590 183681 530628
rect 184751 530590 184785 530628
rect 185211 530590 185245 530628
rect 185763 530590 185797 530628
rect 186866 530600 186890 530622
rect 186959 530594 186993 530628
rect 187419 530590 187453 530628
rect 172211 530428 172485 530590
rect 172489 530454 173037 530590
rect 173039 530428 174141 530590
rect 174143 530428 174693 530590
rect 174789 530416 174875 530573
rect 174881 530454 175429 530590
rect 175523 530454 177361 530590
rect 175523 530408 175707 530454
rect 176273 530410 176459 530454
rect 177365 530416 177451 530573
rect 177658 530454 178351 530590
rect 177658 530408 177842 530454
rect 178375 530434 178649 530590
rect 178653 530454 179201 530590
rect 179203 530454 179751 530590
rect 179941 530416 180027 530573
rect 180215 530454 180995 530590
rect 181181 530454 181961 530590
rect 181963 530454 182511 530590
rect 180215 530408 180401 530454
rect 181775 530408 181961 530454
rect 182517 530416 182603 530573
rect 182607 530428 182973 530590
rect 183067 530454 183615 530590
rect 183619 530428 184721 530590
rect 184723 530428 185089 530590
rect 185093 530416 185179 530573
rect 185183 530454 185731 530590
rect 185735 530428 186837 530590
rect 187207 530428 187481 530590
rect 172211 529544 172485 529706
rect 172487 529544 173589 529706
rect 173591 529544 174693 529706
rect 175318 529680 175502 529726
rect 176425 529680 176611 529724
rect 177177 529680 177361 529726
rect 174809 529544 175502 529680
rect 175523 529544 177361 529680
rect 177365 529561 177451 529718
rect 178187 529680 178373 529726
rect 177593 529544 178373 529680
rect 178375 529680 178559 529726
rect 179125 529680 179311 529724
rect 181117 529680 181303 529724
rect 181869 529680 182053 529726
rect 178375 529544 180213 529680
rect 180215 529544 182053 529680
rect 182055 529544 182421 529706
rect 182517 529561 182603 529718
rect 182626 529680 182810 529726
rect 182626 529544 183319 529680
rect 183343 529544 184445 529706
rect 184447 529544 185549 529706
rect 185551 529544 186653 529706
rect 186655 529544 187205 529706
rect 187207 529544 187481 529706
rect 172239 529502 172273 529544
rect 172515 529502 172549 529544
rect 173619 529502 173653 529544
rect 174722 529512 174746 529534
rect 174815 529506 174849 529544
rect 174909 529511 174941 529533
rect 175551 529506 175585 529544
rect 175772 529502 175806 529540
rect 177482 529512 177506 529534
rect 177667 529502 177701 529540
rect 177759 529502 177793 529540
rect 178256 529506 178290 529544
rect 179598 529512 179622 529534
rect 179691 529502 179725 529540
rect 180059 529502 180093 529540
rect 180151 529506 180185 529544
rect 180243 529506 180277 529544
rect 180610 529512 180634 529534
rect 180703 529502 180737 529540
rect 182083 529506 182117 529544
rect 182450 529512 182474 529534
rect 182727 529502 182761 529540
rect 182819 529502 182853 529540
rect 183279 529506 183313 529544
rect 183371 529506 183405 529544
rect 183923 529502 183957 529540
rect 184475 529506 184509 529544
rect 185026 529512 185050 529534
rect 185211 529502 185245 529540
rect 185579 529506 185613 529544
rect 186315 529502 186349 529540
rect 186683 529506 186717 529544
rect 187053 529511 187085 529533
rect 187419 529502 187453 529544
rect 172211 529340 172485 529502
rect 172487 529340 173589 529502
rect 173591 529340 174693 529502
rect 174789 529328 174875 529485
rect 175109 529366 175889 529502
rect 175908 529366 177729 529502
rect 177731 529366 179569 529502
rect 175703 529320 175889 529366
rect 178633 529322 178819 529366
rect 179385 529320 179569 529366
rect 179663 529346 179937 529502
rect 179941 529328 180027 529485
rect 180031 529340 180581 529502
rect 180675 529366 182496 529502
rect 182515 529346 182789 529502
rect 182791 529340 183893 529502
rect 183895 529340 184997 529502
rect 185093 529328 185179 529485
rect 185183 529340 186285 529502
rect 186287 529340 187021 529502
rect 187207 529340 187481 529502
rect 172211 528456 172485 528618
rect 172487 528456 173589 528618
rect 173591 528456 174693 528618
rect 174695 528456 175797 528618
rect 175891 528456 176165 528612
rect 176167 528456 176441 528612
rect 177083 528592 177269 528638
rect 176489 528456 177269 528592
rect 177365 528473 177451 528630
rect 177474 528592 177658 528638
rect 177474 528456 178167 528592
rect 178375 528456 180196 528592
rect 180215 528456 180489 528612
rect 181393 528592 181579 528636
rect 182145 528592 182329 528638
rect 180491 528456 182329 528592
rect 182517 528473 182603 528630
rect 182607 528456 183709 528618
rect 183711 528456 184813 528618
rect 184815 528456 185917 528618
rect 185919 528456 187021 528618
rect 187207 528456 187481 528618
rect 172239 528414 172273 528456
rect 172515 528414 172549 528456
rect 173619 528414 173653 528456
rect 174723 528446 174757 528456
rect 174722 528424 174757 528446
rect 174723 528418 174757 528424
rect 174907 528414 174941 528452
rect 175826 528424 175850 528446
rect 175919 528418 175953 528456
rect 176010 528424 176034 528446
rect 176103 528414 176137 528452
rect 176195 528418 176229 528456
rect 177152 528418 177186 528456
rect 177298 528424 177322 528446
rect 178127 528414 178161 528456
rect 178219 528414 178253 528452
rect 178403 528418 178437 528456
rect 179010 528414 179044 528452
rect 179785 528423 179817 528445
rect 180059 528414 180093 528452
rect 180243 528418 180277 528456
rect 180519 528418 180553 528456
rect 180797 528423 180829 528445
rect 181034 528414 181068 528452
rect 181807 528414 181841 528452
rect 182361 528425 182393 528447
rect 182635 528418 182669 528456
rect 182911 528414 182945 528452
rect 183739 528418 183773 528456
rect 184015 528414 184049 528452
rect 184843 528418 184877 528456
rect 185211 528414 185245 528452
rect 185947 528418 185981 528456
rect 186315 528414 186349 528452
rect 187053 528423 187085 528447
rect 187419 528414 187453 528456
rect 172211 528252 172485 528414
rect 172487 528252 173589 528414
rect 173591 528252 174693 528414
rect 174789 528240 174875 528397
rect 174879 528252 175981 528414
rect 176075 528278 177913 528414
rect 176977 528234 177163 528278
rect 177729 528232 177913 528278
rect 177915 528258 178189 528414
rect 178191 528252 178925 528414
rect 178927 528278 179707 528414
rect 178927 528232 179113 528278
rect 179941 528240 180027 528397
rect 180031 528252 180765 528414
rect 180951 528278 181731 528414
rect 180951 528232 181137 528278
rect 181779 528252 182881 528414
rect 182883 528252 183985 528414
rect 183987 528252 185089 528414
rect 185093 528240 185179 528397
rect 185183 528252 186285 528414
rect 186287 528252 187021 528414
rect 187207 528252 187481 528414
rect 172211 527368 172485 527530
rect 172487 527368 173589 527530
rect 173591 527368 174693 527530
rect 174695 527368 175797 527530
rect 175799 527368 176349 527530
rect 176370 527504 176554 527550
rect 176370 527368 177063 527504
rect 177087 527368 177361 527530
rect 177365 527385 177451 527542
rect 177455 527368 178557 527530
rect 178559 527368 178925 527530
rect 178946 527504 179130 527550
rect 178946 527368 179639 527504
rect 179663 527368 180765 527530
rect 180767 527368 181869 527530
rect 181871 527368 182421 527530
rect 182517 527385 182603 527542
rect 182607 527368 183709 527530
rect 183711 527368 184813 527530
rect 184815 527368 185917 527530
rect 185919 527368 187021 527530
rect 187207 527368 187481 527530
rect 172239 527326 172273 527368
rect 172515 527326 172549 527368
rect 173619 527326 173653 527368
rect 174723 527358 174757 527368
rect 174722 527336 174757 527358
rect 174723 527330 174757 527336
rect 174907 527326 174941 527364
rect 175827 527330 175861 527368
rect 176011 527326 176045 527364
rect 177023 527330 177057 527368
rect 177115 527326 177149 527368
rect 177483 527330 177517 527368
rect 178219 527326 178253 527364
rect 178587 527330 178621 527368
rect 179323 527326 179357 527364
rect 179599 527330 179633 527368
rect 179691 527330 179725 527368
rect 179874 527336 179898 527358
rect 180059 527326 180093 527364
rect 180795 527330 180829 527368
rect 181163 527326 181197 527364
rect 181899 527330 181933 527368
rect 182267 527326 182301 527364
rect 182450 527336 182474 527358
rect 182635 527330 182669 527368
rect 183371 527326 183405 527364
rect 183739 527330 183773 527368
rect 184475 527326 184509 527364
rect 184843 527330 184877 527368
rect 185026 527336 185050 527358
rect 185211 527326 185245 527364
rect 185947 527330 185981 527368
rect 186315 527326 186349 527364
rect 187053 527335 187085 527359
rect 187419 527326 187453 527368
rect 172211 527164 172485 527326
rect 172487 527164 173589 527326
rect 173591 527164 174693 527326
rect 174789 527152 174875 527309
rect 174879 527164 175981 527326
rect 175983 527164 177085 527326
rect 177087 527164 178189 527326
rect 178191 527164 179293 527326
rect 179295 527164 179845 527326
rect 179941 527152 180027 527309
rect 180031 527164 181133 527326
rect 181135 527164 182237 527326
rect 182239 527164 183341 527326
rect 183343 527164 184445 527326
rect 184447 527164 184997 527326
rect 185093 527152 185179 527309
rect 185183 527164 186285 527326
rect 186287 527164 187021 527326
rect 187207 527164 187481 527326
rect 172211 526280 172485 526442
rect 172487 526280 173589 526442
rect 173591 526280 174693 526442
rect 174695 526280 175797 526442
rect 175799 526280 176901 526442
rect 176903 526280 177269 526442
rect 177365 526297 177451 526454
rect 177455 526280 178557 526442
rect 178559 526280 179661 526442
rect 179663 526280 180765 526442
rect 180767 526280 181869 526442
rect 181871 526280 182421 526442
rect 182517 526297 182603 526454
rect 182607 526280 183709 526442
rect 183711 526280 184813 526442
rect 184815 526280 185917 526442
rect 185919 526280 187021 526442
rect 187207 526280 187481 526442
rect 172239 526238 172273 526280
rect 172515 526238 172549 526280
rect 173619 526238 173653 526280
rect 174723 526270 174757 526280
rect 174722 526248 174757 526270
rect 174723 526242 174757 526248
rect 174907 526238 174941 526276
rect 175827 526242 175861 526280
rect 176011 526238 176045 526276
rect 176931 526242 176965 526280
rect 177115 526238 177149 526276
rect 177298 526248 177322 526270
rect 177483 526242 177517 526280
rect 178219 526238 178253 526276
rect 178587 526242 178621 526280
rect 179323 526238 179357 526276
rect 179691 526242 179725 526280
rect 179874 526248 179898 526270
rect 180059 526238 180093 526276
rect 180795 526242 180829 526280
rect 181163 526238 181197 526276
rect 181899 526242 181933 526280
rect 182267 526238 182301 526276
rect 182450 526248 182474 526270
rect 182635 526242 182669 526280
rect 183371 526238 183405 526276
rect 183739 526242 183773 526280
rect 184475 526238 184509 526276
rect 184843 526242 184877 526280
rect 185026 526248 185050 526270
rect 185211 526238 185245 526276
rect 185947 526242 185981 526280
rect 186315 526238 186349 526276
rect 187053 526247 187085 526271
rect 187419 526238 187453 526280
rect 172211 526076 172485 526238
rect 172487 526076 173589 526238
rect 173591 526076 174693 526238
rect 174789 526064 174875 526221
rect 174879 526076 175981 526238
rect 175983 526076 177085 526238
rect 177087 526076 178189 526238
rect 178191 526076 179293 526238
rect 179295 526076 179845 526238
rect 179941 526064 180027 526221
rect 180031 526076 181133 526238
rect 181135 526076 182237 526238
rect 182239 526076 183341 526238
rect 183343 526076 184445 526238
rect 184447 526076 184997 526238
rect 185093 526064 185179 526221
rect 185183 526076 186285 526238
rect 186287 526076 187021 526238
rect 187207 526076 187481 526238
rect 172211 525192 172485 525354
rect 172487 525192 173589 525354
rect 173591 525192 174693 525354
rect 174695 525192 175797 525354
rect 175799 525192 176901 525354
rect 176903 525192 177269 525354
rect 177365 525209 177451 525366
rect 177455 525192 178557 525354
rect 178559 525192 179661 525354
rect 179663 525192 180765 525354
rect 180767 525192 181869 525354
rect 181871 525192 182421 525354
rect 182517 525209 182603 525366
rect 182607 525192 183709 525354
rect 183711 525192 184813 525354
rect 184815 525192 185917 525354
rect 185919 525192 187021 525354
rect 187207 525192 187481 525354
rect 172239 525150 172273 525192
rect 172515 525150 172549 525192
rect 173619 525150 173653 525192
rect 174723 525182 174757 525192
rect 174722 525160 174757 525182
rect 174723 525154 174757 525160
rect 174907 525150 174941 525188
rect 175827 525154 175861 525192
rect 176011 525150 176045 525188
rect 176931 525154 176965 525192
rect 177115 525150 177149 525188
rect 177298 525160 177322 525182
rect 177483 525154 177517 525192
rect 178219 525150 178253 525188
rect 178587 525154 178621 525192
rect 179323 525150 179357 525188
rect 179691 525154 179725 525192
rect 179874 525160 179898 525182
rect 180059 525150 180093 525188
rect 180795 525154 180829 525192
rect 181163 525150 181197 525188
rect 181899 525154 181933 525192
rect 182267 525150 182301 525188
rect 182450 525160 182474 525182
rect 182635 525154 182669 525192
rect 183371 525150 183405 525188
rect 183739 525154 183773 525192
rect 184475 525150 184509 525188
rect 184843 525154 184877 525192
rect 185026 525160 185050 525182
rect 185211 525150 185245 525188
rect 185947 525154 185981 525192
rect 186315 525150 186349 525188
rect 187053 525159 187085 525183
rect 187419 525150 187453 525192
rect 172211 524988 172485 525150
rect 172487 524988 173589 525150
rect 173591 524988 174693 525150
rect 174789 524976 174875 525133
rect 174879 524988 175981 525150
rect 175983 524988 177085 525150
rect 177087 524988 178189 525150
rect 178191 524988 179293 525150
rect 179295 524988 179845 525150
rect 179941 524976 180027 525133
rect 180031 524988 181133 525150
rect 181135 524988 182237 525150
rect 182239 524988 183341 525150
rect 183343 524988 184445 525150
rect 184447 524988 184997 525150
rect 185093 524976 185179 525133
rect 185183 524988 186285 525150
rect 186287 524988 187021 525150
rect 187207 524988 187481 525150
rect 172211 524104 172485 524266
rect 172487 524104 173589 524266
rect 173591 524104 174693 524266
rect 174695 524104 175797 524266
rect 175799 524104 176901 524266
rect 176903 524104 177269 524266
rect 177365 524121 177451 524278
rect 177455 524104 178557 524266
rect 178559 524104 179661 524266
rect 179663 524104 180765 524266
rect 180767 524104 181869 524266
rect 181871 524104 182421 524266
rect 182517 524121 182603 524278
rect 182607 524104 183709 524266
rect 183711 524104 184813 524266
rect 184815 524104 185917 524266
rect 185919 524104 187021 524266
rect 187207 524104 187481 524266
rect 172239 524062 172273 524104
rect 172515 524062 172549 524104
rect 173619 524062 173653 524104
rect 174723 524094 174757 524104
rect 174722 524072 174757 524094
rect 174723 524066 174757 524072
rect 174907 524062 174941 524100
rect 175827 524066 175861 524104
rect 176011 524062 176045 524100
rect 176931 524066 176965 524104
rect 177115 524062 177149 524100
rect 177298 524072 177322 524094
rect 177483 524066 177517 524104
rect 178219 524062 178253 524100
rect 178587 524066 178621 524104
rect 179323 524062 179357 524100
rect 179691 524066 179725 524104
rect 179874 524072 179898 524094
rect 180059 524062 180093 524100
rect 180795 524066 180829 524104
rect 181163 524062 181197 524100
rect 181899 524066 181933 524104
rect 182267 524062 182301 524100
rect 182450 524072 182474 524094
rect 182635 524066 182669 524104
rect 183371 524062 183405 524100
rect 183739 524066 183773 524104
rect 184475 524062 184509 524100
rect 184843 524066 184877 524104
rect 185026 524072 185050 524094
rect 185211 524062 185245 524100
rect 185947 524066 185981 524104
rect 186315 524062 186349 524100
rect 187053 524071 187085 524095
rect 187419 524062 187453 524104
rect 172211 523900 172485 524062
rect 172487 523900 173589 524062
rect 173591 523900 174693 524062
rect 174789 523888 174875 524045
rect 174879 523900 175981 524062
rect 175983 523900 177085 524062
rect 177087 523900 178189 524062
rect 178191 523900 179293 524062
rect 179295 523900 179845 524062
rect 179941 523888 180027 524045
rect 180031 523900 181133 524062
rect 181135 523900 182237 524062
rect 182239 523900 183341 524062
rect 183343 523900 184445 524062
rect 184447 523900 184997 524062
rect 185093 523888 185179 524045
rect 185183 523900 186285 524062
rect 186287 523900 187021 524062
rect 187207 523900 187481 524062
rect 172211 523016 172485 523178
rect 172487 523016 173589 523178
rect 173591 523016 174693 523178
rect 174695 523016 175797 523178
rect 175799 523016 176901 523178
rect 176903 523016 177269 523178
rect 177365 523033 177451 523190
rect 177455 523016 178557 523178
rect 178559 523016 179661 523178
rect 179663 523016 180765 523178
rect 180767 523016 181869 523178
rect 181871 523016 182421 523178
rect 182517 523033 182603 523190
rect 182607 523016 183709 523178
rect 183711 523016 184813 523178
rect 184815 523016 185917 523178
rect 185919 523016 187021 523178
rect 187207 523016 187481 523178
rect 172239 522974 172273 523016
rect 172515 522974 172549 523016
rect 173619 522974 173653 523016
rect 174723 523006 174757 523016
rect 174722 522984 174757 523006
rect 174723 522978 174757 522984
rect 174907 522974 174941 523012
rect 175827 522978 175861 523016
rect 176011 522974 176045 523012
rect 176931 522978 176965 523016
rect 177115 522974 177149 523012
rect 177298 522984 177322 523006
rect 177483 522978 177517 523016
rect 178219 522974 178253 523012
rect 178587 522978 178621 523016
rect 179323 522974 179357 523012
rect 179691 522978 179725 523016
rect 179874 522984 179898 523006
rect 180059 522974 180093 523012
rect 180795 522978 180829 523016
rect 181163 522974 181197 523012
rect 181899 522978 181933 523016
rect 182267 522974 182301 523012
rect 182450 522984 182474 523006
rect 182635 522978 182669 523016
rect 183371 522974 183405 523012
rect 183739 522978 183773 523016
rect 184475 522974 184509 523012
rect 184843 522978 184877 523016
rect 185026 522984 185050 523006
rect 185211 522974 185245 523012
rect 185947 522978 185981 523016
rect 186315 522974 186349 523012
rect 187053 522983 187085 523007
rect 187419 522974 187453 523016
rect 172211 522812 172485 522974
rect 172487 522812 173589 522974
rect 173591 522812 174693 522974
rect 174789 522800 174875 522957
rect 174879 522812 175981 522974
rect 175983 522812 177085 522974
rect 177087 522812 178189 522974
rect 178191 522812 179293 522974
rect 179295 522812 179845 522974
rect 179941 522800 180027 522957
rect 180031 522812 181133 522974
rect 181135 522812 182237 522974
rect 182239 522812 183341 522974
rect 183343 522812 184445 522974
rect 184447 522812 184997 522974
rect 185093 522800 185179 522957
rect 185183 522812 186285 522974
rect 186287 522812 187021 522974
rect 187207 522812 187481 522974
rect 172211 521928 172485 522090
rect 172487 521928 173589 522090
rect 173591 521928 174693 522090
rect 174695 521928 175797 522090
rect 175799 521928 176901 522090
rect 176903 521928 177269 522090
rect 177365 521945 177451 522102
rect 177455 521928 178557 522090
rect 178559 521928 179661 522090
rect 179663 521928 180765 522090
rect 180767 521928 181869 522090
rect 181871 521928 182421 522090
rect 182517 521945 182603 522102
rect 182607 521928 183709 522090
rect 183711 521928 184813 522090
rect 184815 521928 185917 522090
rect 185919 521928 187021 522090
rect 187207 521928 187481 522090
rect 172239 521886 172273 521928
rect 172515 521886 172549 521928
rect 173619 521886 173653 521928
rect 174723 521918 174757 521928
rect 174722 521896 174757 521918
rect 174723 521890 174757 521896
rect 174907 521886 174941 521924
rect 175827 521890 175861 521928
rect 176011 521886 176045 521924
rect 176931 521890 176965 521928
rect 177115 521886 177149 521924
rect 177298 521896 177322 521918
rect 177483 521890 177517 521928
rect 178219 521886 178253 521924
rect 178587 521890 178621 521928
rect 179323 521886 179357 521924
rect 179691 521890 179725 521928
rect 179874 521896 179898 521918
rect 180059 521886 180093 521924
rect 180795 521890 180829 521928
rect 181163 521886 181197 521924
rect 181899 521890 181933 521928
rect 182267 521886 182301 521924
rect 182450 521896 182474 521918
rect 182635 521890 182669 521928
rect 183371 521886 183405 521924
rect 183739 521890 183773 521928
rect 184475 521886 184509 521924
rect 184843 521890 184877 521928
rect 185026 521896 185050 521918
rect 185211 521886 185245 521924
rect 185947 521890 185981 521928
rect 186315 521886 186349 521924
rect 187053 521895 187085 521919
rect 187419 521886 187453 521928
rect 172211 521724 172485 521886
rect 172487 521724 173589 521886
rect 173591 521724 174693 521886
rect 174789 521712 174875 521869
rect 174879 521724 175981 521886
rect 175983 521724 177085 521886
rect 177087 521724 178189 521886
rect 178191 521724 179293 521886
rect 179295 521724 179845 521886
rect 179941 521712 180027 521869
rect 180031 521724 181133 521886
rect 181135 521724 182237 521886
rect 182239 521724 183341 521886
rect 183343 521724 184445 521886
rect 184447 521724 184997 521886
rect 185093 521712 185179 521869
rect 185183 521724 186285 521886
rect 186287 521724 187021 521886
rect 187207 521724 187481 521886
rect 172211 520840 172485 521002
rect 172487 520840 173589 521002
rect 173591 520840 174693 521002
rect 174695 520840 175797 521002
rect 175799 520840 176901 521002
rect 176903 520840 177269 521002
rect 177365 520857 177451 521014
rect 177455 520840 178557 521002
rect 178559 520840 179661 521002
rect 179663 520840 180765 521002
rect 180767 520840 181869 521002
rect 181871 520840 182421 521002
rect 182517 520857 182603 521014
rect 182607 520840 183709 521002
rect 183711 520840 184813 521002
rect 184815 520840 185917 521002
rect 185919 520840 187021 521002
rect 187207 520840 187481 521002
rect 172239 520798 172273 520840
rect 172515 520798 172549 520840
rect 173619 520798 173653 520840
rect 174723 520830 174757 520840
rect 174722 520808 174757 520830
rect 174723 520802 174757 520808
rect 174907 520798 174941 520836
rect 175827 520802 175861 520840
rect 176011 520798 176045 520836
rect 176931 520802 176965 520840
rect 177115 520798 177149 520836
rect 177298 520808 177322 520830
rect 177483 520802 177517 520840
rect 178219 520798 178253 520836
rect 178587 520802 178621 520840
rect 179323 520798 179357 520836
rect 179691 520802 179725 520840
rect 179874 520808 179898 520830
rect 180059 520798 180093 520836
rect 180795 520802 180829 520840
rect 181163 520798 181197 520836
rect 181899 520802 181933 520840
rect 182267 520798 182301 520836
rect 182450 520808 182474 520830
rect 182635 520802 182669 520840
rect 183371 520798 183405 520836
rect 183739 520802 183773 520840
rect 184475 520798 184509 520836
rect 184843 520802 184877 520840
rect 185026 520808 185050 520830
rect 185211 520798 185245 520836
rect 185947 520802 185981 520840
rect 186315 520798 186349 520836
rect 187053 520807 187085 520831
rect 187419 520798 187453 520840
rect 172211 520636 172485 520798
rect 172487 520636 173589 520798
rect 173591 520636 174693 520798
rect 174789 520624 174875 520781
rect 174879 520636 175981 520798
rect 175983 520636 177085 520798
rect 177087 520636 178189 520798
rect 178191 520636 179293 520798
rect 179295 520636 179845 520798
rect 179941 520624 180027 520781
rect 180031 520636 181133 520798
rect 181135 520636 182237 520798
rect 182239 520636 183341 520798
rect 183343 520636 184445 520798
rect 184447 520636 184997 520798
rect 185093 520624 185179 520781
rect 185183 520636 186285 520798
rect 186287 520636 187021 520798
rect 187207 520636 187481 520798
rect 172211 519752 172485 519914
rect 172487 519752 173589 519914
rect 173591 519752 174693 519914
rect 174695 519752 175797 519914
rect 175799 519752 176901 519914
rect 176903 519752 177269 519914
rect 177365 519769 177451 519926
rect 177455 519752 178557 519914
rect 178559 519752 179661 519914
rect 179663 519752 180765 519914
rect 180767 519752 181869 519914
rect 181871 519752 182421 519914
rect 182517 519769 182603 519926
rect 182607 519752 183709 519914
rect 183711 519752 184813 519914
rect 184815 519752 185917 519914
rect 185919 519752 187021 519914
rect 187207 519752 187481 519914
rect 172239 519710 172273 519752
rect 172515 519710 172549 519752
rect 173619 519710 173653 519752
rect 174723 519742 174757 519752
rect 174722 519720 174757 519742
rect 174723 519714 174757 519720
rect 174907 519710 174941 519748
rect 175827 519714 175861 519752
rect 176011 519710 176045 519748
rect 176931 519714 176965 519752
rect 177115 519710 177149 519748
rect 177298 519720 177322 519742
rect 177483 519714 177517 519752
rect 178219 519710 178253 519748
rect 178587 519714 178621 519752
rect 179323 519710 179357 519748
rect 179691 519714 179725 519752
rect 179874 519720 179898 519742
rect 180059 519710 180093 519748
rect 180795 519714 180829 519752
rect 181163 519710 181197 519748
rect 181899 519714 181933 519752
rect 182267 519710 182301 519748
rect 182450 519720 182474 519742
rect 182635 519714 182669 519752
rect 183371 519710 183405 519748
rect 183739 519714 183773 519752
rect 184475 519710 184509 519748
rect 184843 519714 184877 519752
rect 185026 519720 185050 519742
rect 185211 519710 185245 519748
rect 185947 519714 185981 519752
rect 186315 519710 186349 519748
rect 187053 519719 187085 519743
rect 187419 519710 187453 519752
rect 172211 519548 172485 519710
rect 172487 519548 173589 519710
rect 173591 519548 174693 519710
rect 174789 519536 174875 519693
rect 174879 519548 175981 519710
rect 175983 519548 177085 519710
rect 177087 519548 178189 519710
rect 178191 519548 179293 519710
rect 179295 519548 179845 519710
rect 179941 519536 180027 519693
rect 180031 519548 181133 519710
rect 181135 519548 182237 519710
rect 182239 519548 183341 519710
rect 183343 519548 184445 519710
rect 184447 519548 184997 519710
rect 185093 519536 185179 519693
rect 185183 519548 186285 519710
rect 186287 519548 187021 519710
rect 187207 519548 187481 519710
rect 172211 518664 172485 518826
rect 172487 518664 173589 518826
rect 173591 518664 174693 518826
rect 174695 518664 175797 518826
rect 175799 518664 176901 518826
rect 176903 518664 177269 518826
rect 177365 518681 177451 518838
rect 177455 518664 178557 518826
rect 178559 518664 179661 518826
rect 179663 518664 180765 518826
rect 180767 518664 181869 518826
rect 181871 518664 182421 518826
rect 182517 518681 182603 518838
rect 182607 518664 183709 518826
rect 183711 518664 184813 518826
rect 184815 518664 185917 518826
rect 185919 518664 187021 518826
rect 187207 518664 187481 518826
rect 172239 518622 172273 518664
rect 172515 518622 172549 518664
rect 173619 518622 173653 518664
rect 174723 518654 174757 518664
rect 174722 518632 174757 518654
rect 174723 518626 174757 518632
rect 174907 518622 174941 518660
rect 175827 518626 175861 518664
rect 176011 518622 176045 518660
rect 176931 518626 176965 518664
rect 177115 518622 177149 518660
rect 177298 518632 177322 518654
rect 177483 518626 177517 518664
rect 178219 518622 178253 518660
rect 178587 518626 178621 518664
rect 179323 518622 179357 518660
rect 179691 518626 179725 518664
rect 179874 518632 179898 518654
rect 180059 518622 180093 518660
rect 180795 518626 180829 518664
rect 181163 518622 181197 518660
rect 181899 518626 181933 518664
rect 182267 518622 182301 518660
rect 182450 518632 182474 518654
rect 182635 518626 182669 518664
rect 183371 518622 183405 518660
rect 183739 518626 183773 518664
rect 184475 518622 184509 518660
rect 184843 518626 184877 518664
rect 185026 518632 185050 518654
rect 185211 518622 185245 518660
rect 185947 518626 185981 518664
rect 186315 518622 186349 518660
rect 187053 518631 187085 518655
rect 187419 518622 187453 518664
rect 172211 518460 172485 518622
rect 172487 518460 173589 518622
rect 173591 518460 174693 518622
rect 174789 518448 174875 518605
rect 174879 518460 175981 518622
rect 175983 518460 177085 518622
rect 177087 518460 178189 518622
rect 178191 518460 179293 518622
rect 179295 518460 179845 518622
rect 179941 518448 180027 518605
rect 180031 518460 181133 518622
rect 181135 518460 182237 518622
rect 182239 518460 183341 518622
rect 183343 518460 184445 518622
rect 184447 518460 184997 518622
rect 185093 518448 185179 518605
rect 185183 518460 186285 518622
rect 186287 518460 187021 518622
rect 187207 518460 187481 518622
rect 172211 517576 172485 517738
rect 172487 517576 173589 517738
rect 173591 517576 174693 517738
rect 174695 517576 175797 517738
rect 175799 517576 176901 517738
rect 176903 517576 177269 517738
rect 177365 517593 177451 517750
rect 177455 517576 178557 517738
rect 178559 517576 179661 517738
rect 179663 517576 180765 517738
rect 180767 517576 181869 517738
rect 181871 517576 182421 517738
rect 182517 517593 182603 517750
rect 182607 517576 183709 517738
rect 183711 517576 184813 517738
rect 184815 517576 185917 517738
rect 185919 517576 187021 517738
rect 187207 517576 187481 517738
rect 172239 517534 172273 517576
rect 172515 517534 172549 517576
rect 173619 517534 173653 517576
rect 174723 517566 174757 517576
rect 174722 517544 174757 517566
rect 174723 517538 174757 517544
rect 174907 517534 174941 517572
rect 175827 517538 175861 517576
rect 176011 517534 176045 517572
rect 176931 517538 176965 517576
rect 177115 517534 177149 517572
rect 177298 517544 177322 517566
rect 177483 517538 177517 517576
rect 178219 517534 178253 517572
rect 178587 517538 178621 517576
rect 179323 517534 179357 517572
rect 179691 517538 179725 517576
rect 179874 517544 179898 517566
rect 180059 517534 180093 517572
rect 180795 517538 180829 517576
rect 181163 517534 181197 517572
rect 181899 517538 181933 517576
rect 182267 517534 182301 517572
rect 182450 517544 182474 517566
rect 182635 517538 182669 517576
rect 183371 517534 183405 517572
rect 183739 517538 183773 517576
rect 184475 517534 184509 517572
rect 184843 517538 184877 517576
rect 185026 517544 185050 517566
rect 185211 517534 185245 517572
rect 185947 517538 185981 517576
rect 186315 517534 186349 517572
rect 187053 517543 187085 517567
rect 187419 517534 187453 517576
rect 172211 517372 172485 517534
rect 172487 517372 173589 517534
rect 173591 517372 174693 517534
rect 174789 517360 174875 517517
rect 174879 517372 175981 517534
rect 175983 517372 177085 517534
rect 177087 517372 178189 517534
rect 178191 517372 179293 517534
rect 179295 517372 179845 517534
rect 179941 517360 180027 517517
rect 180031 517372 181133 517534
rect 181135 517372 182237 517534
rect 182239 517372 183341 517534
rect 183343 517372 184445 517534
rect 184447 517372 184997 517534
rect 185093 517360 185179 517517
rect 185183 517372 186285 517534
rect 186287 517372 187021 517534
rect 187207 517372 187481 517534
rect 172211 516488 172485 516650
rect 172487 516488 173589 516650
rect 173591 516488 174693 516650
rect 174695 516488 175797 516650
rect 175799 516488 176901 516650
rect 176903 516488 177269 516650
rect 177365 516505 177451 516662
rect 177455 516488 178557 516650
rect 178559 516488 179661 516650
rect 179663 516488 180765 516650
rect 180767 516488 181869 516650
rect 181871 516488 182421 516650
rect 182517 516505 182603 516662
rect 182607 516488 183709 516650
rect 183711 516488 184813 516650
rect 184815 516488 185917 516650
rect 185919 516488 187021 516650
rect 187207 516488 187481 516650
rect 172239 516446 172273 516488
rect 172515 516446 172549 516488
rect 173619 516446 173653 516488
rect 174723 516478 174757 516488
rect 174722 516456 174757 516478
rect 174723 516450 174757 516456
rect 174907 516446 174941 516484
rect 175827 516450 175861 516488
rect 176011 516446 176045 516484
rect 176931 516450 176965 516488
rect 177115 516446 177149 516484
rect 177298 516456 177322 516478
rect 177483 516450 177517 516488
rect 178219 516446 178253 516484
rect 178587 516450 178621 516488
rect 179323 516446 179357 516484
rect 179691 516450 179725 516488
rect 179874 516456 179898 516478
rect 180059 516446 180093 516484
rect 180795 516450 180829 516488
rect 181163 516446 181197 516484
rect 181899 516450 181933 516488
rect 182267 516446 182301 516484
rect 182450 516456 182474 516478
rect 182635 516450 182669 516488
rect 183371 516446 183405 516484
rect 183739 516450 183773 516488
rect 184475 516446 184509 516484
rect 184843 516450 184877 516488
rect 185026 516456 185050 516478
rect 185211 516446 185245 516484
rect 185947 516450 185981 516488
rect 186315 516446 186349 516484
rect 187053 516455 187085 516479
rect 187419 516446 187453 516488
rect 172211 516284 172485 516446
rect 172487 516284 173589 516446
rect 173591 516284 174693 516446
rect 174789 516272 174875 516429
rect 174879 516284 175981 516446
rect 175983 516284 177085 516446
rect 177087 516284 178189 516446
rect 178191 516284 179293 516446
rect 179295 516284 179845 516446
rect 179941 516272 180027 516429
rect 180031 516284 181133 516446
rect 181135 516284 182237 516446
rect 182239 516284 183341 516446
rect 183343 516284 184445 516446
rect 184447 516284 184997 516446
rect 185093 516272 185179 516429
rect 185183 516284 186285 516446
rect 186287 516284 187021 516446
rect 187207 516284 187481 516446
rect 172211 515400 172485 515562
rect 172487 515400 173221 515562
rect 173407 515400 173955 515536
rect 173959 515400 174693 515562
rect 174789 515417 174875 515574
rect 174879 515400 175981 515562
rect 175983 515400 177085 515562
rect 177087 515400 177361 515562
rect 177365 515417 177451 515574
rect 177455 515400 178557 515562
rect 178559 515400 179661 515562
rect 179663 515400 179937 515562
rect 179941 515417 180027 515574
rect 180031 515400 181133 515562
rect 181135 515400 181869 515562
rect 182055 515400 182329 515556
rect 182517 515417 182603 515574
rect 182607 515400 183709 515562
rect 183711 515400 184813 515562
rect 184815 515400 185089 515562
rect 185093 515417 185179 515574
rect 185183 515400 186285 515562
rect 186379 515400 186927 515536
rect 186931 515400 187205 515562
rect 187207 515400 187481 515562
rect 172239 515362 172273 515400
rect 172515 515362 172549 515400
rect 173253 515369 173285 515391
rect 173435 515362 173469 515400
rect 173987 515362 174021 515400
rect 174722 515368 174746 515390
rect 174907 515362 174941 515400
rect 176011 515362 176045 515400
rect 177115 515362 177149 515400
rect 177483 515362 177517 515400
rect 178587 515362 178621 515400
rect 179691 515362 179725 515400
rect 180059 515362 180093 515400
rect 181163 515362 181197 515400
rect 181901 515369 181933 515391
rect 182265 515362 182299 515400
rect 182361 515369 182393 515391
rect 182635 515362 182669 515400
rect 183739 515362 183773 515400
rect 184843 515362 184877 515400
rect 185211 515362 185245 515400
rect 186314 515368 186338 515390
rect 186407 515362 186441 515400
rect 186959 515362 186993 515400
rect 187419 515362 187453 515400
<< nmos >>
rect 164732 540079 164762 541079
rect 164939 540086 164969 541086
rect 165035 540086 165065 541086
rect 165131 540086 165161 541086
rect 165227 540086 165257 541086
rect 165323 540086 165353 541086
rect 165419 540086 165449 541086
rect 165515 540086 165545 541086
rect 165611 540086 165641 541086
rect 165707 540086 165737 541086
rect 165803 540086 165833 541086
rect 165899 540086 165929 541086
rect 165995 540086 166025 541086
rect 166212 540079 166242 540279
rect 166412 540079 166442 541079
rect 168532 540079 168562 541079
rect 168739 540086 168769 541086
rect 168835 540086 168865 541086
rect 168931 540086 168961 541086
rect 169027 540086 169057 541086
rect 169123 540086 169153 541086
rect 169219 540086 169249 541086
rect 169315 540086 169345 541086
rect 169411 540086 169441 541086
rect 169507 540086 169537 541086
rect 169603 540086 169633 541086
rect 169699 540086 169729 541086
rect 169795 540086 169825 541086
rect 170012 540079 170042 540279
rect 170212 540079 170242 541079
rect 172232 540079 172262 541079
rect 172439 540086 172469 541086
rect 172535 540086 172565 541086
rect 172631 540086 172661 541086
rect 172727 540086 172757 541086
rect 172823 540086 172853 541086
rect 172919 540086 172949 541086
rect 173015 540086 173045 541086
rect 173111 540086 173141 541086
rect 173207 540086 173237 541086
rect 173303 540086 173333 541086
rect 173399 540086 173429 541086
rect 173495 540086 173525 541086
rect 173712 540079 173742 540279
rect 173912 540079 173942 541079
rect 175732 540079 175762 541079
rect 175939 540086 175969 541086
rect 176035 540086 176065 541086
rect 176131 540086 176161 541086
rect 176227 540086 176257 541086
rect 176323 540086 176353 541086
rect 176419 540086 176449 541086
rect 176515 540086 176545 541086
rect 176611 540086 176641 541086
rect 176707 540086 176737 541086
rect 176803 540086 176833 541086
rect 176899 540086 176929 541086
rect 176995 540086 177025 541086
rect 177212 540079 177242 540279
rect 177412 540079 177442 541079
rect 179332 540079 179362 541079
rect 179539 540086 179569 541086
rect 179635 540086 179665 541086
rect 179731 540086 179761 541086
rect 179827 540086 179857 541086
rect 179923 540086 179953 541086
rect 180019 540086 180049 541086
rect 180115 540086 180145 541086
rect 180211 540086 180241 541086
rect 180307 540086 180337 541086
rect 180403 540086 180433 541086
rect 180499 540086 180529 541086
rect 180595 540086 180625 541086
rect 180812 540079 180842 540279
rect 181012 540079 181042 541079
rect 182632 540079 182662 541079
rect 182839 540086 182869 541086
rect 182935 540086 182965 541086
rect 183031 540086 183061 541086
rect 183127 540086 183157 541086
rect 183223 540086 183253 541086
rect 183319 540086 183349 541086
rect 183415 540086 183445 541086
rect 183511 540086 183541 541086
rect 183607 540086 183637 541086
rect 183703 540086 183733 541086
rect 183799 540086 183829 541086
rect 183895 540086 183925 541086
rect 184112 540079 184142 540279
rect 184312 540079 184342 541079
rect 185932 540079 185962 541079
rect 186139 540086 186169 541086
rect 186235 540086 186265 541086
rect 186331 540086 186361 541086
rect 186427 540086 186457 541086
rect 186523 540086 186553 541086
rect 186619 540086 186649 541086
rect 186715 540086 186745 541086
rect 186811 540086 186841 541086
rect 186907 540086 186937 541086
rect 187003 540086 187033 541086
rect 187099 540086 187129 541086
rect 187195 540086 187225 541086
rect 187412 540079 187442 540279
rect 187612 540079 187642 541079
rect 189232 540079 189262 541079
rect 189439 540086 189469 541086
rect 189535 540086 189565 541086
rect 189631 540086 189661 541086
rect 189727 540086 189757 541086
rect 189823 540086 189853 541086
rect 189919 540086 189949 541086
rect 190015 540086 190045 541086
rect 190111 540086 190141 541086
rect 190207 540086 190237 541086
rect 190303 540086 190333 541086
rect 190399 540086 190429 541086
rect 190495 540086 190525 541086
rect 190712 540079 190742 540279
rect 190912 540079 190942 541079
rect 158712 538229 158912 538429
rect 159088 538229 159288 538429
rect 159346 538229 159546 538429
rect 159604 538229 159804 538429
rect 159862 538229 160062 538429
rect 160120 538229 160320 538429
rect 160378 538229 160578 538429
rect 160636 538229 160836 538429
rect 160894 538229 161094 538429
rect 161152 538229 161352 538429
rect 161532 538229 161732 538429
rect 161932 538229 162132 538429
rect 162312 538229 162512 538429
<< scnmos >>
rect 172289 530454 172407 530564
rect 172573 530480 172603 530564
rect 172659 530480 172689 530564
rect 172745 530480 172775 530564
rect 172831 530480 172861 530564
rect 172928 530480 172958 530564
rect 173117 530454 174063 530564
rect 174221 530454 174615 530564
rect 174965 530480 174995 530564
rect 175051 530480 175081 530564
rect 175137 530480 175167 530564
rect 175223 530480 175253 530564
rect 175320 530480 175350 530564
rect 175601 530434 175631 530564
rect 175809 530480 175839 530564
rect 175900 530480 175930 530564
rect 176049 530480 176079 530564
rect 176145 530492 176175 530564
rect 176254 530492 176284 530564
rect 176353 530436 176383 530564
rect 176485 530480 176515 530564
rect 176557 530480 176587 530564
rect 176723 530492 176753 530564
rect 176819 530492 176849 530564
rect 176914 530480 176944 530564
rect 177169 530480 177199 530564
rect 177253 530480 177283 530564
rect 177736 530434 177766 530564
rect 177831 530480 177931 530564
rect 178089 530480 178189 530564
rect 178243 530480 178273 530564
rect 178453 530460 178483 530564
rect 178541 530460 178571 530564
rect 178737 530480 178767 530564
rect 178823 530480 178853 530564
rect 178909 530480 178939 530564
rect 178995 530480 179025 530564
rect 179092 530480 179122 530564
rect 179282 530480 179312 530564
rect 179379 530480 179409 530564
rect 179465 530480 179495 530564
rect 179551 530480 179581 530564
rect 179637 530480 179667 530564
rect 180293 530434 180323 530564
rect 180402 530480 180432 530564
rect 180498 530480 180528 530564
rect 180623 530480 180653 530564
rect 180719 530480 180749 530564
rect 180887 530480 180917 530564
rect 181259 530480 181289 530564
rect 181427 530480 181457 530564
rect 181523 530480 181553 530564
rect 181648 530480 181678 530564
rect 181744 530480 181774 530564
rect 181853 530434 181883 530564
rect 182042 530480 182072 530564
rect 182139 530480 182169 530564
rect 182225 530480 182255 530564
rect 182311 530480 182341 530564
rect 182397 530480 182427 530564
rect 182685 530454 182895 530564
rect 183146 530480 183176 530564
rect 183243 530480 183273 530564
rect 183329 530480 183359 530564
rect 183415 530480 183445 530564
rect 183501 530480 183531 530564
rect 183697 530454 184643 530564
rect 184801 530454 185011 530564
rect 185262 530480 185292 530564
rect 185359 530480 185389 530564
rect 185445 530480 185475 530564
rect 185531 530480 185561 530564
rect 185617 530480 185647 530564
rect 185813 530454 186759 530564
rect 187285 530454 187403 530564
rect 172289 529570 172407 529680
rect 172565 529570 173511 529680
rect 173669 529570 174615 529680
rect 174887 529570 174917 529654
rect 174971 529570 175071 529654
rect 175229 529570 175329 529654
rect 175394 529570 175424 529700
rect 175601 529570 175631 529654
rect 175685 529570 175715 529654
rect 175940 529570 175970 529654
rect 176035 529570 176065 529642
rect 176131 529570 176161 529642
rect 176297 529570 176327 529654
rect 176369 529570 176399 529654
rect 176501 529570 176531 529698
rect 176600 529570 176630 529642
rect 176709 529570 176739 529642
rect 176805 529570 176835 529654
rect 176954 529570 176984 529654
rect 177045 529570 177075 529654
rect 177253 529570 177283 529700
rect 177671 529570 177701 529654
rect 177839 529570 177869 529654
rect 177935 529570 177965 529654
rect 178060 529570 178090 529654
rect 178156 529570 178186 529654
rect 178265 529570 178295 529700
rect 178453 529570 178483 529700
rect 178661 529570 178691 529654
rect 178752 529570 178782 529654
rect 178901 529570 178931 529654
rect 178997 529570 179027 529642
rect 179106 529570 179136 529642
rect 179205 529570 179235 529698
rect 179337 529570 179367 529654
rect 179409 529570 179439 529654
rect 179575 529570 179605 529642
rect 179671 529570 179701 529642
rect 179766 529570 179796 529654
rect 180021 529570 180051 529654
rect 180105 529570 180135 529654
rect 180293 529570 180323 529654
rect 180377 529570 180407 529654
rect 180632 529570 180662 529654
rect 180727 529570 180757 529642
rect 180823 529570 180853 529642
rect 180989 529570 181019 529654
rect 181061 529570 181091 529654
rect 181193 529570 181223 529698
rect 181292 529570 181322 529642
rect 181401 529570 181431 529642
rect 181497 529570 181527 529654
rect 181646 529570 181676 529654
rect 181737 529570 181767 529654
rect 181945 529570 181975 529700
rect 182133 529570 182343 529680
rect 182704 529570 182734 529700
rect 182799 529570 182899 529654
rect 183057 529570 183157 529654
rect 183211 529570 183241 529654
rect 183421 529570 184367 529680
rect 184525 529570 185471 529680
rect 185629 529570 186575 529680
rect 186733 529570 187127 529680
rect 187285 529570 187403 529680
rect 172289 529366 172407 529476
rect 172565 529366 173511 529476
rect 173669 529366 174615 529476
rect 175187 529392 175217 529476
rect 175355 529392 175385 529476
rect 175451 529392 175481 529476
rect 175576 529392 175606 529476
rect 175672 529392 175702 529476
rect 175781 529346 175811 529476
rect 175987 529392 176017 529476
rect 176073 529392 176103 529476
rect 176159 529392 176189 529476
rect 176245 529392 176275 529476
rect 176331 529392 176361 529476
rect 176417 529392 176447 529476
rect 176503 529392 176533 529476
rect 176589 529392 176619 529476
rect 176674 529392 176704 529476
rect 176760 529392 176790 529476
rect 176846 529392 176876 529476
rect 176932 529392 176962 529476
rect 177018 529392 177048 529476
rect 177104 529392 177134 529476
rect 177190 529392 177220 529476
rect 177276 529392 177306 529476
rect 177362 529392 177392 529476
rect 177448 529392 177478 529476
rect 177534 529392 177564 529476
rect 177620 529392 177650 529476
rect 177809 529392 177839 529476
rect 177893 529392 177923 529476
rect 178148 529392 178178 529476
rect 178243 529404 178273 529476
rect 178339 529404 178369 529476
rect 178505 529392 178535 529476
rect 178577 529392 178607 529476
rect 178709 529348 178739 529476
rect 178808 529404 178838 529476
rect 178917 529404 178947 529476
rect 179013 529392 179043 529476
rect 179162 529392 179192 529476
rect 179253 529392 179283 529476
rect 179461 529346 179491 529476
rect 179741 529372 179771 529476
rect 179829 529372 179859 529476
rect 180109 529366 180503 529476
rect 180754 529392 180784 529476
rect 180840 529392 180870 529476
rect 180926 529392 180956 529476
rect 181012 529392 181042 529476
rect 181098 529392 181128 529476
rect 181184 529392 181214 529476
rect 181270 529392 181300 529476
rect 181356 529392 181386 529476
rect 181442 529392 181472 529476
rect 181528 529392 181558 529476
rect 181614 529392 181644 529476
rect 181700 529392 181730 529476
rect 181785 529392 181815 529476
rect 181871 529392 181901 529476
rect 181957 529392 181987 529476
rect 182043 529392 182073 529476
rect 182129 529392 182159 529476
rect 182215 529392 182245 529476
rect 182301 529392 182331 529476
rect 182387 529392 182417 529476
rect 182593 529372 182623 529476
rect 182681 529372 182711 529476
rect 182869 529366 183815 529476
rect 183973 529366 184919 529476
rect 185261 529366 186207 529476
rect 186365 529366 186943 529476
rect 187285 529366 187403 529476
rect 172289 528482 172407 528592
rect 172565 528482 173511 528592
rect 173669 528482 174615 528592
rect 174773 528482 175719 528592
rect 175969 528482 175999 528586
rect 176057 528482 176087 528586
rect 176245 528482 176275 528586
rect 176333 528482 176363 528586
rect 176567 528482 176597 528566
rect 176735 528482 176765 528566
rect 176831 528482 176861 528566
rect 176956 528482 176986 528566
rect 177052 528482 177082 528566
rect 177161 528482 177191 528612
rect 177552 528482 177582 528612
rect 177647 528482 177747 528566
rect 177905 528482 178005 528566
rect 178059 528482 178089 528566
rect 178454 528482 178484 528566
rect 178540 528482 178570 528566
rect 178626 528482 178656 528566
rect 178712 528482 178742 528566
rect 178798 528482 178828 528566
rect 178884 528482 178914 528566
rect 178970 528482 179000 528566
rect 179056 528482 179086 528566
rect 179142 528482 179172 528566
rect 179228 528482 179258 528566
rect 179314 528482 179344 528566
rect 179400 528482 179430 528566
rect 179485 528482 179515 528566
rect 179571 528482 179601 528566
rect 179657 528482 179687 528566
rect 179743 528482 179773 528566
rect 179829 528482 179859 528566
rect 179915 528482 179945 528566
rect 180001 528482 180031 528566
rect 180087 528482 180117 528566
rect 180293 528482 180323 528586
rect 180381 528482 180411 528586
rect 180569 528482 180599 528566
rect 180653 528482 180683 528566
rect 180908 528482 180938 528566
rect 181003 528482 181033 528554
rect 181099 528482 181129 528554
rect 181265 528482 181295 528566
rect 181337 528482 181367 528566
rect 181469 528482 181499 528610
rect 181568 528482 181598 528554
rect 181677 528482 181707 528554
rect 181773 528482 181803 528566
rect 181922 528482 181952 528566
rect 182013 528482 182043 528566
rect 182221 528482 182251 528612
rect 182685 528482 183631 528592
rect 183789 528482 184735 528592
rect 184893 528482 185839 528592
rect 185997 528482 186943 528592
rect 187285 528482 187403 528592
rect 172289 528278 172407 528388
rect 172565 528278 173511 528388
rect 173669 528278 174615 528388
rect 174957 528278 175903 528388
rect 176153 528304 176183 528388
rect 176237 528304 176267 528388
rect 176492 528304 176522 528388
rect 176587 528316 176617 528388
rect 176683 528316 176713 528388
rect 176849 528304 176879 528388
rect 176921 528304 176951 528388
rect 177053 528260 177083 528388
rect 177152 528316 177182 528388
rect 177261 528316 177291 528388
rect 177357 528304 177387 528388
rect 177506 528304 177536 528388
rect 177597 528304 177627 528388
rect 177805 528258 177835 528388
rect 177993 528284 178023 528388
rect 178081 528284 178111 528388
rect 178269 528278 178847 528388
rect 179005 528258 179035 528388
rect 179114 528304 179144 528388
rect 179210 528304 179240 528388
rect 179335 528304 179365 528388
rect 179431 528304 179461 528388
rect 179599 528304 179629 528388
rect 180109 528278 180687 528388
rect 181029 528258 181059 528388
rect 181138 528304 181168 528388
rect 181234 528304 181264 528388
rect 181359 528304 181389 528388
rect 181455 528304 181485 528388
rect 181623 528304 181653 528388
rect 181857 528278 182803 528388
rect 182961 528278 183907 528388
rect 184065 528278 185011 528388
rect 185261 528278 186207 528388
rect 186365 528278 186943 528388
rect 187285 528278 187403 528388
rect 172289 527394 172407 527504
rect 172565 527394 173511 527504
rect 173669 527394 174615 527504
rect 174773 527394 175719 527504
rect 175877 527394 176271 527504
rect 176448 527394 176478 527524
rect 176543 527394 176643 527478
rect 176801 527394 176901 527478
rect 176955 527394 176985 527478
rect 177165 527394 177283 527504
rect 177533 527394 178479 527504
rect 178637 527394 178847 527504
rect 179024 527394 179054 527524
rect 179119 527394 179219 527478
rect 179377 527394 179477 527478
rect 179531 527394 179561 527478
rect 179741 527394 180687 527504
rect 180845 527394 181791 527504
rect 181949 527394 182343 527504
rect 182685 527394 183631 527504
rect 183789 527394 184735 527504
rect 184893 527394 185839 527504
rect 185997 527394 186943 527504
rect 187285 527394 187403 527504
rect 172289 527190 172407 527300
rect 172565 527190 173511 527300
rect 173669 527190 174615 527300
rect 174957 527190 175903 527300
rect 176061 527190 177007 527300
rect 177165 527190 178111 527300
rect 178269 527190 179215 527300
rect 179373 527190 179767 527300
rect 180109 527190 181055 527300
rect 181213 527190 182159 527300
rect 182317 527190 183263 527300
rect 183421 527190 184367 527300
rect 184525 527190 184919 527300
rect 185261 527190 186207 527300
rect 186365 527190 186943 527300
rect 187285 527190 187403 527300
rect 172289 526306 172407 526416
rect 172565 526306 173511 526416
rect 173669 526306 174615 526416
rect 174773 526306 175719 526416
rect 175877 526306 176823 526416
rect 176981 526306 177191 526416
rect 177533 526306 178479 526416
rect 178637 526306 179583 526416
rect 179741 526306 180687 526416
rect 180845 526306 181791 526416
rect 181949 526306 182343 526416
rect 182685 526306 183631 526416
rect 183789 526306 184735 526416
rect 184893 526306 185839 526416
rect 185997 526306 186943 526416
rect 187285 526306 187403 526416
rect 172289 526102 172407 526212
rect 172565 526102 173511 526212
rect 173669 526102 174615 526212
rect 174957 526102 175903 526212
rect 176061 526102 177007 526212
rect 177165 526102 178111 526212
rect 178269 526102 179215 526212
rect 179373 526102 179767 526212
rect 180109 526102 181055 526212
rect 181213 526102 182159 526212
rect 182317 526102 183263 526212
rect 183421 526102 184367 526212
rect 184525 526102 184919 526212
rect 185261 526102 186207 526212
rect 186365 526102 186943 526212
rect 187285 526102 187403 526212
rect 172289 525218 172407 525328
rect 172565 525218 173511 525328
rect 173669 525218 174615 525328
rect 174773 525218 175719 525328
rect 175877 525218 176823 525328
rect 176981 525218 177191 525328
rect 177533 525218 178479 525328
rect 178637 525218 179583 525328
rect 179741 525218 180687 525328
rect 180845 525218 181791 525328
rect 181949 525218 182343 525328
rect 182685 525218 183631 525328
rect 183789 525218 184735 525328
rect 184893 525218 185839 525328
rect 185997 525218 186943 525328
rect 187285 525218 187403 525328
rect 172289 525014 172407 525124
rect 172565 525014 173511 525124
rect 173669 525014 174615 525124
rect 174957 525014 175903 525124
rect 176061 525014 177007 525124
rect 177165 525014 178111 525124
rect 178269 525014 179215 525124
rect 179373 525014 179767 525124
rect 180109 525014 181055 525124
rect 181213 525014 182159 525124
rect 182317 525014 183263 525124
rect 183421 525014 184367 525124
rect 184525 525014 184919 525124
rect 185261 525014 186207 525124
rect 186365 525014 186943 525124
rect 187285 525014 187403 525124
rect 172289 524130 172407 524240
rect 172565 524130 173511 524240
rect 173669 524130 174615 524240
rect 174773 524130 175719 524240
rect 175877 524130 176823 524240
rect 176981 524130 177191 524240
rect 177533 524130 178479 524240
rect 178637 524130 179583 524240
rect 179741 524130 180687 524240
rect 180845 524130 181791 524240
rect 181949 524130 182343 524240
rect 182685 524130 183631 524240
rect 183789 524130 184735 524240
rect 184893 524130 185839 524240
rect 185997 524130 186943 524240
rect 187285 524130 187403 524240
rect 172289 523926 172407 524036
rect 172565 523926 173511 524036
rect 173669 523926 174615 524036
rect 174957 523926 175903 524036
rect 176061 523926 177007 524036
rect 177165 523926 178111 524036
rect 178269 523926 179215 524036
rect 179373 523926 179767 524036
rect 180109 523926 181055 524036
rect 181213 523926 182159 524036
rect 182317 523926 183263 524036
rect 183421 523926 184367 524036
rect 184525 523926 184919 524036
rect 185261 523926 186207 524036
rect 186365 523926 186943 524036
rect 187285 523926 187403 524036
rect 172289 523042 172407 523152
rect 172565 523042 173511 523152
rect 173669 523042 174615 523152
rect 174773 523042 175719 523152
rect 175877 523042 176823 523152
rect 176981 523042 177191 523152
rect 177533 523042 178479 523152
rect 178637 523042 179583 523152
rect 179741 523042 180687 523152
rect 180845 523042 181791 523152
rect 181949 523042 182343 523152
rect 182685 523042 183631 523152
rect 183789 523042 184735 523152
rect 184893 523042 185839 523152
rect 185997 523042 186943 523152
rect 187285 523042 187403 523152
rect 172289 522838 172407 522948
rect 172565 522838 173511 522948
rect 173669 522838 174615 522948
rect 174957 522838 175903 522948
rect 176061 522838 177007 522948
rect 177165 522838 178111 522948
rect 178269 522838 179215 522948
rect 179373 522838 179767 522948
rect 180109 522838 181055 522948
rect 181213 522838 182159 522948
rect 182317 522838 183263 522948
rect 183421 522838 184367 522948
rect 184525 522838 184919 522948
rect 185261 522838 186207 522948
rect 186365 522838 186943 522948
rect 187285 522838 187403 522948
rect 172289 521954 172407 522064
rect 172565 521954 173511 522064
rect 173669 521954 174615 522064
rect 174773 521954 175719 522064
rect 175877 521954 176823 522064
rect 176981 521954 177191 522064
rect 177533 521954 178479 522064
rect 178637 521954 179583 522064
rect 179741 521954 180687 522064
rect 180845 521954 181791 522064
rect 181949 521954 182343 522064
rect 182685 521954 183631 522064
rect 183789 521954 184735 522064
rect 184893 521954 185839 522064
rect 185997 521954 186943 522064
rect 187285 521954 187403 522064
rect 172289 521750 172407 521860
rect 172565 521750 173511 521860
rect 173669 521750 174615 521860
rect 174957 521750 175903 521860
rect 176061 521750 177007 521860
rect 177165 521750 178111 521860
rect 178269 521750 179215 521860
rect 179373 521750 179767 521860
rect 180109 521750 181055 521860
rect 181213 521750 182159 521860
rect 182317 521750 183263 521860
rect 183421 521750 184367 521860
rect 184525 521750 184919 521860
rect 185261 521750 186207 521860
rect 186365 521750 186943 521860
rect 187285 521750 187403 521860
rect 172289 520866 172407 520976
rect 172565 520866 173511 520976
rect 173669 520866 174615 520976
rect 174773 520866 175719 520976
rect 175877 520866 176823 520976
rect 176981 520866 177191 520976
rect 177533 520866 178479 520976
rect 178637 520866 179583 520976
rect 179741 520866 180687 520976
rect 180845 520866 181791 520976
rect 181949 520866 182343 520976
rect 182685 520866 183631 520976
rect 183789 520866 184735 520976
rect 184893 520866 185839 520976
rect 185997 520866 186943 520976
rect 187285 520866 187403 520976
rect 172289 520662 172407 520772
rect 172565 520662 173511 520772
rect 173669 520662 174615 520772
rect 174957 520662 175903 520772
rect 176061 520662 177007 520772
rect 177165 520662 178111 520772
rect 178269 520662 179215 520772
rect 179373 520662 179767 520772
rect 180109 520662 181055 520772
rect 181213 520662 182159 520772
rect 182317 520662 183263 520772
rect 183421 520662 184367 520772
rect 184525 520662 184919 520772
rect 185261 520662 186207 520772
rect 186365 520662 186943 520772
rect 187285 520662 187403 520772
rect 172289 519778 172407 519888
rect 172565 519778 173511 519888
rect 173669 519778 174615 519888
rect 174773 519778 175719 519888
rect 175877 519778 176823 519888
rect 176981 519778 177191 519888
rect 177533 519778 178479 519888
rect 178637 519778 179583 519888
rect 179741 519778 180687 519888
rect 180845 519778 181791 519888
rect 181949 519778 182343 519888
rect 182685 519778 183631 519888
rect 183789 519778 184735 519888
rect 184893 519778 185839 519888
rect 185997 519778 186943 519888
rect 187285 519778 187403 519888
rect 172289 519574 172407 519684
rect 172565 519574 173511 519684
rect 173669 519574 174615 519684
rect 174957 519574 175903 519684
rect 176061 519574 177007 519684
rect 177165 519574 178111 519684
rect 178269 519574 179215 519684
rect 179373 519574 179767 519684
rect 180109 519574 181055 519684
rect 181213 519574 182159 519684
rect 182317 519574 183263 519684
rect 183421 519574 184367 519684
rect 184525 519574 184919 519684
rect 185261 519574 186207 519684
rect 186365 519574 186943 519684
rect 187285 519574 187403 519684
rect 172289 518690 172407 518800
rect 172565 518690 173511 518800
rect 173669 518690 174615 518800
rect 174773 518690 175719 518800
rect 175877 518690 176823 518800
rect 176981 518690 177191 518800
rect 177533 518690 178479 518800
rect 178637 518690 179583 518800
rect 179741 518690 180687 518800
rect 180845 518690 181791 518800
rect 181949 518690 182343 518800
rect 182685 518690 183631 518800
rect 183789 518690 184735 518800
rect 184893 518690 185839 518800
rect 185997 518690 186943 518800
rect 187285 518690 187403 518800
rect 172289 518486 172407 518596
rect 172565 518486 173511 518596
rect 173669 518486 174615 518596
rect 174957 518486 175903 518596
rect 176061 518486 177007 518596
rect 177165 518486 178111 518596
rect 178269 518486 179215 518596
rect 179373 518486 179767 518596
rect 180109 518486 181055 518596
rect 181213 518486 182159 518596
rect 182317 518486 183263 518596
rect 183421 518486 184367 518596
rect 184525 518486 184919 518596
rect 185261 518486 186207 518596
rect 186365 518486 186943 518596
rect 187285 518486 187403 518596
rect 172289 517602 172407 517712
rect 172565 517602 173511 517712
rect 173669 517602 174615 517712
rect 174773 517602 175719 517712
rect 175877 517602 176823 517712
rect 176981 517602 177191 517712
rect 177533 517602 178479 517712
rect 178637 517602 179583 517712
rect 179741 517602 180687 517712
rect 180845 517602 181791 517712
rect 181949 517602 182343 517712
rect 182685 517602 183631 517712
rect 183789 517602 184735 517712
rect 184893 517602 185839 517712
rect 185997 517602 186943 517712
rect 187285 517602 187403 517712
rect 172289 517398 172407 517508
rect 172565 517398 173511 517508
rect 173669 517398 174615 517508
rect 174957 517398 175903 517508
rect 176061 517398 177007 517508
rect 177165 517398 178111 517508
rect 178269 517398 179215 517508
rect 179373 517398 179767 517508
rect 180109 517398 181055 517508
rect 181213 517398 182159 517508
rect 182317 517398 183263 517508
rect 183421 517398 184367 517508
rect 184525 517398 184919 517508
rect 185261 517398 186207 517508
rect 186365 517398 186943 517508
rect 187285 517398 187403 517508
rect 172289 516514 172407 516624
rect 172565 516514 173511 516624
rect 173669 516514 174615 516624
rect 174773 516514 175719 516624
rect 175877 516514 176823 516624
rect 176981 516514 177191 516624
rect 177533 516514 178479 516624
rect 178637 516514 179583 516624
rect 179741 516514 180687 516624
rect 180845 516514 181791 516624
rect 181949 516514 182343 516624
rect 182685 516514 183631 516624
rect 183789 516514 184735 516624
rect 184893 516514 185839 516624
rect 185997 516514 186943 516624
rect 187285 516514 187403 516624
rect 172289 516310 172407 516420
rect 172565 516310 173511 516420
rect 173669 516310 174615 516420
rect 174957 516310 175903 516420
rect 176061 516310 177007 516420
rect 177165 516310 178111 516420
rect 178269 516310 179215 516420
rect 179373 516310 179767 516420
rect 180109 516310 181055 516420
rect 181213 516310 182159 516420
rect 182317 516310 183263 516420
rect 183421 516310 184367 516420
rect 184525 516310 184919 516420
rect 185261 516310 186207 516420
rect 186365 516310 186943 516420
rect 187285 516310 187403 516420
rect 172289 515426 172407 515536
rect 172565 515426 173143 515536
rect 173486 515426 173516 515510
rect 173583 515426 173613 515510
rect 173669 515426 173699 515510
rect 173755 515426 173785 515510
rect 173841 515426 173871 515510
rect 174037 515426 174615 515536
rect 174957 515426 175903 515536
rect 176061 515426 177007 515536
rect 177165 515426 177283 515536
rect 177533 515426 178479 515536
rect 178637 515426 179583 515536
rect 179741 515426 179859 515536
rect 180109 515426 181055 515536
rect 181213 515426 181791 515536
rect 182133 515426 182163 515530
rect 182221 515426 182251 515530
rect 182685 515426 183631 515536
rect 183789 515426 184735 515536
rect 184893 515426 185011 515536
rect 185261 515426 186207 515536
rect 186458 515426 186488 515510
rect 186555 515426 186585 515510
rect 186641 515426 186671 515510
rect 186727 515426 186757 515510
rect 186813 515426 186843 515510
rect 187009 515426 187127 515536
rect 187285 515426 187403 515536
<< pmos >>
rect 164716 538557 164746 539557
rect 164943 538564 164973 539564
rect 165039 538564 165069 539564
rect 165135 538564 165165 539564
rect 165231 538564 165261 539564
rect 165327 538564 165357 539564
rect 165423 538564 165453 539564
rect 165519 538564 165549 539564
rect 165615 538564 165645 539564
rect 165711 538564 165741 539564
rect 165807 538564 165837 539564
rect 165903 538564 165933 539564
rect 165999 538564 166029 539564
rect 166216 538957 166246 539557
rect 166416 538557 166446 539557
rect 168516 538557 168546 539557
rect 168743 538564 168773 539564
rect 168839 538564 168869 539564
rect 168935 538564 168965 539564
rect 169031 538564 169061 539564
rect 169127 538564 169157 539564
rect 169223 538564 169253 539564
rect 169319 538564 169349 539564
rect 169415 538564 169445 539564
rect 169511 538564 169541 539564
rect 169607 538564 169637 539564
rect 169703 538564 169733 539564
rect 169799 538564 169829 539564
rect 170016 538957 170046 539557
rect 170216 538557 170246 539557
rect 172216 538557 172246 539557
rect 172443 538564 172473 539564
rect 172539 538564 172569 539564
rect 172635 538564 172665 539564
rect 172731 538564 172761 539564
rect 172827 538564 172857 539564
rect 172923 538564 172953 539564
rect 173019 538564 173049 539564
rect 173115 538564 173145 539564
rect 173211 538564 173241 539564
rect 173307 538564 173337 539564
rect 173403 538564 173433 539564
rect 173499 538564 173529 539564
rect 173716 538957 173746 539557
rect 173916 538557 173946 539557
rect 175716 538557 175746 539557
rect 175943 538564 175973 539564
rect 176039 538564 176069 539564
rect 176135 538564 176165 539564
rect 176231 538564 176261 539564
rect 176327 538564 176357 539564
rect 176423 538564 176453 539564
rect 176519 538564 176549 539564
rect 176615 538564 176645 539564
rect 176711 538564 176741 539564
rect 176807 538564 176837 539564
rect 176903 538564 176933 539564
rect 176999 538564 177029 539564
rect 177216 538957 177246 539557
rect 177416 538557 177446 539557
rect 179316 538557 179346 539557
rect 179543 538564 179573 539564
rect 179639 538564 179669 539564
rect 179735 538564 179765 539564
rect 179831 538564 179861 539564
rect 179927 538564 179957 539564
rect 180023 538564 180053 539564
rect 180119 538564 180149 539564
rect 180215 538564 180245 539564
rect 180311 538564 180341 539564
rect 180407 538564 180437 539564
rect 180503 538564 180533 539564
rect 180599 538564 180629 539564
rect 180816 538957 180846 539557
rect 181016 538557 181046 539557
rect 182616 538557 182646 539557
rect 182843 538564 182873 539564
rect 182939 538564 182969 539564
rect 183035 538564 183065 539564
rect 183131 538564 183161 539564
rect 183227 538564 183257 539564
rect 183323 538564 183353 539564
rect 183419 538564 183449 539564
rect 183515 538564 183545 539564
rect 183611 538564 183641 539564
rect 183707 538564 183737 539564
rect 183803 538564 183833 539564
rect 183899 538564 183929 539564
rect 184116 538957 184146 539557
rect 184316 538557 184346 539557
rect 185916 538557 185946 539557
rect 186143 538564 186173 539564
rect 186239 538564 186269 539564
rect 186335 538564 186365 539564
rect 186431 538564 186461 539564
rect 186527 538564 186557 539564
rect 186623 538564 186653 539564
rect 186719 538564 186749 539564
rect 186815 538564 186845 539564
rect 186911 538564 186941 539564
rect 187007 538564 187037 539564
rect 187103 538564 187133 539564
rect 187199 538564 187229 539564
rect 187416 538957 187446 539557
rect 187616 538557 187646 539557
rect 189216 538557 189246 539557
rect 189443 538564 189473 539564
rect 189539 538564 189569 539564
rect 189635 538564 189665 539564
rect 189731 538564 189761 539564
rect 189827 538564 189857 539564
rect 189923 538564 189953 539564
rect 190019 538564 190049 539564
rect 190115 538564 190145 539564
rect 190211 538564 190241 539564
rect 190307 538564 190337 539564
rect 190403 538564 190433 539564
rect 190499 538564 190529 539564
rect 190716 538957 190746 539557
rect 190916 538557 190946 539557
rect 161306 537057 161336 537657
rect 161510 537057 161540 537657
rect 161606 537057 161636 537657
rect 161702 537057 161732 537657
rect 161910 537057 161940 537657
rect 162006 537057 162036 537657
rect 162102 537057 162132 537657
rect 162326 537057 162356 537657
rect 157796 536037 157996 536637
rect 158174 536037 158374 536637
rect 158432 536037 158632 536637
rect 158690 536037 158890 536637
rect 158948 536037 159148 536637
rect 159206 536037 159406 536637
rect 159464 536037 159664 536637
rect 159722 536037 159922 536637
rect 159980 536037 160180 536637
rect 160238 536037 160438 536637
rect 160496 536037 160696 536637
rect 160880 536037 161080 536637
rect 161138 536037 161338 536637
rect 161396 536037 161596 536637
rect 161778 536037 161978 536637
rect 162036 536037 162236 536637
rect 162416 536037 162616 536637
<< scpmoshvt >>
rect 172289 530114 172407 530288
rect 172574 530114 172604 530314
rect 172660 530114 172690 530314
rect 172746 530114 172776 530314
rect 172832 530114 172862 530314
rect 172928 530114 172958 530314
rect 173117 530114 174063 530288
rect 174221 530114 174615 530288
rect 174966 530114 174996 530314
rect 175052 530114 175082 530314
rect 175138 530114 175168 530314
rect 175224 530114 175254 530314
rect 175320 530114 175350 530314
rect 175601 530114 175631 530314
rect 175816 530114 175846 530198
rect 175900 530114 175930 530198
rect 176008 530114 176038 530198
rect 176092 530114 176122 530198
rect 176178 530114 176208 530198
rect 176277 530114 176307 530282
rect 176474 530114 176504 530198
rect 176571 530114 176601 530198
rect 176711 530114 176741 530198
rect 176810 530114 176840 530198
rect 176902 530114 176932 530198
rect 177169 530120 177199 530248
rect 177253 530120 177283 530248
rect 177736 530114 177766 530314
rect 177831 530114 177931 530198
rect 178089 530114 178189 530198
rect 178243 530114 178273 530198
rect 178453 530114 178483 530272
rect 178541 530114 178571 530272
rect 178738 530114 178768 530314
rect 178824 530114 178854 530314
rect 178910 530114 178940 530314
rect 178996 530114 179026 530314
rect 179092 530114 179122 530314
rect 179282 530114 179312 530314
rect 179378 530114 179408 530314
rect 179464 530114 179494 530314
rect 179550 530114 179580 530314
rect 179636 530114 179666 530314
rect 180293 530114 180323 530314
rect 180402 530153 180432 530237
rect 180505 530153 180535 530237
rect 180719 530153 180749 530237
rect 180791 530153 180821 530237
rect 180887 530153 180917 530237
rect 181259 530153 181289 530237
rect 181355 530153 181385 530237
rect 181427 530153 181457 530237
rect 181641 530153 181671 530237
rect 181744 530153 181774 530237
rect 181853 530114 181883 530314
rect 182042 530114 182072 530314
rect 182138 530114 182168 530314
rect 182224 530114 182254 530314
rect 182310 530114 182340 530314
rect 182396 530114 182426 530314
rect 182685 530114 182895 530288
rect 183146 530114 183176 530314
rect 183242 530114 183272 530314
rect 183328 530114 183358 530314
rect 183414 530114 183444 530314
rect 183500 530114 183530 530314
rect 183697 530114 184643 530288
rect 184801 530114 185011 530288
rect 185262 530114 185292 530314
rect 185358 530114 185388 530314
rect 185444 530114 185474 530314
rect 185530 530114 185560 530314
rect 185616 530114 185646 530314
rect 185813 530114 186759 530288
rect 187285 530114 187403 530288
rect 172289 529846 172407 530020
rect 172565 529846 173511 530020
rect 173669 529846 174615 530020
rect 174887 529936 174917 530020
rect 174971 529936 175071 530020
rect 175229 529936 175329 530020
rect 175394 529820 175424 530020
rect 175601 529886 175631 530014
rect 175685 529886 175715 530014
rect 175952 529936 175982 530020
rect 176044 529936 176074 530020
rect 176143 529936 176173 530020
rect 176283 529936 176313 530020
rect 176380 529936 176410 530020
rect 176577 529852 176607 530020
rect 176676 529936 176706 530020
rect 176762 529936 176792 530020
rect 176846 529936 176876 530020
rect 176954 529936 176984 530020
rect 177038 529936 177068 530020
rect 177253 529820 177283 530020
rect 177671 529897 177701 529981
rect 177767 529897 177797 529981
rect 177839 529897 177869 529981
rect 178053 529897 178083 529981
rect 178156 529897 178186 529981
rect 178265 529820 178295 530020
rect 178453 529820 178483 530020
rect 178668 529936 178698 530020
rect 178752 529936 178782 530020
rect 178860 529936 178890 530020
rect 178944 529936 178974 530020
rect 179030 529936 179060 530020
rect 179129 529852 179159 530020
rect 179326 529936 179356 530020
rect 179423 529936 179453 530020
rect 179563 529936 179593 530020
rect 179662 529936 179692 530020
rect 179754 529936 179784 530020
rect 180021 529886 180051 530014
rect 180105 529886 180135 530014
rect 180293 529886 180323 530014
rect 180377 529886 180407 530014
rect 180644 529936 180674 530020
rect 180736 529936 180766 530020
rect 180835 529936 180865 530020
rect 180975 529936 181005 530020
rect 181072 529936 181102 530020
rect 181269 529852 181299 530020
rect 181368 529936 181398 530020
rect 181454 529936 181484 530020
rect 181538 529936 181568 530020
rect 181646 529936 181676 530020
rect 181730 529936 181760 530020
rect 181945 529820 181975 530020
rect 182133 529846 182343 530020
rect 182704 529820 182734 530020
rect 182799 529936 182899 530020
rect 183057 529936 183157 530020
rect 183211 529936 183241 530020
rect 183421 529846 184367 530020
rect 184525 529846 185471 530020
rect 185629 529846 186575 530020
rect 186733 529846 187127 530020
rect 187285 529846 187403 530020
rect 172289 529026 172407 529200
rect 172565 529026 173511 529200
rect 173669 529026 174615 529200
rect 175187 529065 175217 529149
rect 175283 529065 175313 529149
rect 175355 529065 175385 529149
rect 175569 529065 175599 529149
rect 175672 529065 175702 529149
rect 175781 529026 175811 529226
rect 175987 529026 176017 529226
rect 176073 529026 176103 529226
rect 176159 529026 176189 529226
rect 176245 529026 176275 529226
rect 176331 529026 176361 529226
rect 176417 529026 176447 529226
rect 176503 529026 176533 529226
rect 176589 529026 176619 529226
rect 176674 529026 176704 529226
rect 176760 529026 176790 529226
rect 176846 529026 176876 529226
rect 176932 529026 176962 529226
rect 177018 529026 177048 529226
rect 177104 529026 177134 529226
rect 177190 529026 177220 529226
rect 177276 529026 177306 529226
rect 177362 529026 177392 529226
rect 177448 529026 177478 529226
rect 177534 529026 177564 529226
rect 177620 529026 177650 529226
rect 177809 529032 177839 529160
rect 177893 529032 177923 529160
rect 178160 529026 178190 529110
rect 178252 529026 178282 529110
rect 178351 529026 178381 529110
rect 178491 529026 178521 529110
rect 178588 529026 178618 529110
rect 178785 529026 178815 529194
rect 178884 529026 178914 529110
rect 178970 529026 179000 529110
rect 179054 529026 179084 529110
rect 179162 529026 179192 529110
rect 179246 529026 179276 529110
rect 179461 529026 179491 529226
rect 179741 529026 179771 529184
rect 179829 529026 179859 529184
rect 180109 529026 180503 529200
rect 180754 529026 180784 529226
rect 180840 529026 180870 529226
rect 180926 529026 180956 529226
rect 181012 529026 181042 529226
rect 181098 529026 181128 529226
rect 181184 529026 181214 529226
rect 181270 529026 181300 529226
rect 181356 529026 181386 529226
rect 181442 529026 181472 529226
rect 181528 529026 181558 529226
rect 181614 529026 181644 529226
rect 181700 529026 181730 529226
rect 181785 529026 181815 529226
rect 181871 529026 181901 529226
rect 181957 529026 181987 529226
rect 182043 529026 182073 529226
rect 182129 529026 182159 529226
rect 182215 529026 182245 529226
rect 182301 529026 182331 529226
rect 182387 529026 182417 529226
rect 182593 529026 182623 529184
rect 182681 529026 182711 529184
rect 182869 529026 183815 529200
rect 183973 529026 184919 529200
rect 185261 529026 186207 529200
rect 186365 529026 186943 529200
rect 187285 529026 187403 529200
rect 172289 528758 172407 528932
rect 172565 528758 173511 528932
rect 173669 528758 174615 528932
rect 174773 528758 175719 528932
rect 175969 528774 175999 528932
rect 176057 528774 176087 528932
rect 176245 528774 176275 528932
rect 176333 528774 176363 528932
rect 176567 528809 176597 528893
rect 176663 528809 176693 528893
rect 176735 528809 176765 528893
rect 176949 528809 176979 528893
rect 177052 528809 177082 528893
rect 177161 528732 177191 528932
rect 177552 528732 177582 528932
rect 177647 528848 177747 528932
rect 177905 528848 178005 528932
rect 178059 528848 178089 528932
rect 178454 528732 178484 528932
rect 178540 528732 178570 528932
rect 178626 528732 178656 528932
rect 178712 528732 178742 528932
rect 178798 528732 178828 528932
rect 178884 528732 178914 528932
rect 178970 528732 179000 528932
rect 179056 528732 179086 528932
rect 179142 528732 179172 528932
rect 179228 528732 179258 528932
rect 179314 528732 179344 528932
rect 179400 528732 179430 528932
rect 179485 528732 179515 528932
rect 179571 528732 179601 528932
rect 179657 528732 179687 528932
rect 179743 528732 179773 528932
rect 179829 528732 179859 528932
rect 179915 528732 179945 528932
rect 180001 528732 180031 528932
rect 180087 528732 180117 528932
rect 180293 528774 180323 528932
rect 180381 528774 180411 528932
rect 180569 528798 180599 528926
rect 180653 528798 180683 528926
rect 180920 528848 180950 528932
rect 181012 528848 181042 528932
rect 181111 528848 181141 528932
rect 181251 528848 181281 528932
rect 181348 528848 181378 528932
rect 181545 528764 181575 528932
rect 181644 528848 181674 528932
rect 181730 528848 181760 528932
rect 181814 528848 181844 528932
rect 181922 528848 181952 528932
rect 182006 528848 182036 528932
rect 182221 528732 182251 528932
rect 182685 528758 183631 528932
rect 183789 528758 184735 528932
rect 184893 528758 185839 528932
rect 185997 528758 186943 528932
rect 187285 528758 187403 528932
rect 172289 527938 172407 528112
rect 172565 527938 173511 528112
rect 173669 527938 174615 528112
rect 174957 527938 175903 528112
rect 176153 527944 176183 528072
rect 176237 527944 176267 528072
rect 176504 527938 176534 528022
rect 176596 527938 176626 528022
rect 176695 527938 176725 528022
rect 176835 527938 176865 528022
rect 176932 527938 176962 528022
rect 177129 527938 177159 528106
rect 177228 527938 177258 528022
rect 177314 527938 177344 528022
rect 177398 527938 177428 528022
rect 177506 527938 177536 528022
rect 177590 527938 177620 528022
rect 177805 527938 177835 528138
rect 177993 527938 178023 528096
rect 178081 527938 178111 528096
rect 178269 527938 178847 528112
rect 179005 527938 179035 528138
rect 179114 527977 179144 528061
rect 179217 527977 179247 528061
rect 179431 527977 179461 528061
rect 179503 527977 179533 528061
rect 179599 527977 179629 528061
rect 180109 527938 180687 528112
rect 181029 527938 181059 528138
rect 181138 527977 181168 528061
rect 181241 527977 181271 528061
rect 181455 527977 181485 528061
rect 181527 527977 181557 528061
rect 181623 527977 181653 528061
rect 181857 527938 182803 528112
rect 182961 527938 183907 528112
rect 184065 527938 185011 528112
rect 185261 527938 186207 528112
rect 186365 527938 186943 528112
rect 187285 527938 187403 528112
rect 172289 527670 172407 527844
rect 172565 527670 173511 527844
rect 173669 527670 174615 527844
rect 174773 527670 175719 527844
rect 175877 527670 176271 527844
rect 176448 527644 176478 527844
rect 176543 527760 176643 527844
rect 176801 527760 176901 527844
rect 176955 527760 176985 527844
rect 177165 527670 177283 527844
rect 177533 527670 178479 527844
rect 178637 527670 178847 527844
rect 179024 527644 179054 527844
rect 179119 527760 179219 527844
rect 179377 527760 179477 527844
rect 179531 527760 179561 527844
rect 179741 527670 180687 527844
rect 180845 527670 181791 527844
rect 181949 527670 182343 527844
rect 182685 527670 183631 527844
rect 183789 527670 184735 527844
rect 184893 527670 185839 527844
rect 185997 527670 186943 527844
rect 187285 527670 187403 527844
rect 172289 526850 172407 527024
rect 172565 526850 173511 527024
rect 173669 526850 174615 527024
rect 174957 526850 175903 527024
rect 176061 526850 177007 527024
rect 177165 526850 178111 527024
rect 178269 526850 179215 527024
rect 179373 526850 179767 527024
rect 180109 526850 181055 527024
rect 181213 526850 182159 527024
rect 182317 526850 183263 527024
rect 183421 526850 184367 527024
rect 184525 526850 184919 527024
rect 185261 526850 186207 527024
rect 186365 526850 186943 527024
rect 187285 526850 187403 527024
rect 172289 526582 172407 526756
rect 172565 526582 173511 526756
rect 173669 526582 174615 526756
rect 174773 526582 175719 526756
rect 175877 526582 176823 526756
rect 176981 526582 177191 526756
rect 177533 526582 178479 526756
rect 178637 526582 179583 526756
rect 179741 526582 180687 526756
rect 180845 526582 181791 526756
rect 181949 526582 182343 526756
rect 182685 526582 183631 526756
rect 183789 526582 184735 526756
rect 184893 526582 185839 526756
rect 185997 526582 186943 526756
rect 187285 526582 187403 526756
rect 172289 525762 172407 525936
rect 172565 525762 173511 525936
rect 173669 525762 174615 525936
rect 174957 525762 175903 525936
rect 176061 525762 177007 525936
rect 177165 525762 178111 525936
rect 178269 525762 179215 525936
rect 179373 525762 179767 525936
rect 180109 525762 181055 525936
rect 181213 525762 182159 525936
rect 182317 525762 183263 525936
rect 183421 525762 184367 525936
rect 184525 525762 184919 525936
rect 185261 525762 186207 525936
rect 186365 525762 186943 525936
rect 187285 525762 187403 525936
rect 172289 525494 172407 525668
rect 172565 525494 173511 525668
rect 173669 525494 174615 525668
rect 174773 525494 175719 525668
rect 175877 525494 176823 525668
rect 176981 525494 177191 525668
rect 177533 525494 178479 525668
rect 178637 525494 179583 525668
rect 179741 525494 180687 525668
rect 180845 525494 181791 525668
rect 181949 525494 182343 525668
rect 182685 525494 183631 525668
rect 183789 525494 184735 525668
rect 184893 525494 185839 525668
rect 185997 525494 186943 525668
rect 187285 525494 187403 525668
rect 172289 524674 172407 524848
rect 172565 524674 173511 524848
rect 173669 524674 174615 524848
rect 174957 524674 175903 524848
rect 176061 524674 177007 524848
rect 177165 524674 178111 524848
rect 178269 524674 179215 524848
rect 179373 524674 179767 524848
rect 180109 524674 181055 524848
rect 181213 524674 182159 524848
rect 182317 524674 183263 524848
rect 183421 524674 184367 524848
rect 184525 524674 184919 524848
rect 185261 524674 186207 524848
rect 186365 524674 186943 524848
rect 187285 524674 187403 524848
rect 172289 524406 172407 524580
rect 172565 524406 173511 524580
rect 173669 524406 174615 524580
rect 174773 524406 175719 524580
rect 175877 524406 176823 524580
rect 176981 524406 177191 524580
rect 177533 524406 178479 524580
rect 178637 524406 179583 524580
rect 179741 524406 180687 524580
rect 180845 524406 181791 524580
rect 181949 524406 182343 524580
rect 182685 524406 183631 524580
rect 183789 524406 184735 524580
rect 184893 524406 185839 524580
rect 185997 524406 186943 524580
rect 187285 524406 187403 524580
rect 172289 523586 172407 523760
rect 172565 523586 173511 523760
rect 173669 523586 174615 523760
rect 174957 523586 175903 523760
rect 176061 523586 177007 523760
rect 177165 523586 178111 523760
rect 178269 523586 179215 523760
rect 179373 523586 179767 523760
rect 180109 523586 181055 523760
rect 181213 523586 182159 523760
rect 182317 523586 183263 523760
rect 183421 523586 184367 523760
rect 184525 523586 184919 523760
rect 185261 523586 186207 523760
rect 186365 523586 186943 523760
rect 187285 523586 187403 523760
rect 172289 523318 172407 523492
rect 172565 523318 173511 523492
rect 173669 523318 174615 523492
rect 174773 523318 175719 523492
rect 175877 523318 176823 523492
rect 176981 523318 177191 523492
rect 177533 523318 178479 523492
rect 178637 523318 179583 523492
rect 179741 523318 180687 523492
rect 180845 523318 181791 523492
rect 181949 523318 182343 523492
rect 182685 523318 183631 523492
rect 183789 523318 184735 523492
rect 184893 523318 185839 523492
rect 185997 523318 186943 523492
rect 187285 523318 187403 523492
rect 172289 522498 172407 522672
rect 172565 522498 173511 522672
rect 173669 522498 174615 522672
rect 174957 522498 175903 522672
rect 176061 522498 177007 522672
rect 177165 522498 178111 522672
rect 178269 522498 179215 522672
rect 179373 522498 179767 522672
rect 180109 522498 181055 522672
rect 181213 522498 182159 522672
rect 182317 522498 183263 522672
rect 183421 522498 184367 522672
rect 184525 522498 184919 522672
rect 185261 522498 186207 522672
rect 186365 522498 186943 522672
rect 187285 522498 187403 522672
rect 172289 522230 172407 522404
rect 172565 522230 173511 522404
rect 173669 522230 174615 522404
rect 174773 522230 175719 522404
rect 175877 522230 176823 522404
rect 176981 522230 177191 522404
rect 177533 522230 178479 522404
rect 178637 522230 179583 522404
rect 179741 522230 180687 522404
rect 180845 522230 181791 522404
rect 181949 522230 182343 522404
rect 182685 522230 183631 522404
rect 183789 522230 184735 522404
rect 184893 522230 185839 522404
rect 185997 522230 186943 522404
rect 187285 522230 187403 522404
rect 172289 521410 172407 521584
rect 172565 521410 173511 521584
rect 173669 521410 174615 521584
rect 174957 521410 175903 521584
rect 176061 521410 177007 521584
rect 177165 521410 178111 521584
rect 178269 521410 179215 521584
rect 179373 521410 179767 521584
rect 180109 521410 181055 521584
rect 181213 521410 182159 521584
rect 182317 521410 183263 521584
rect 183421 521410 184367 521584
rect 184525 521410 184919 521584
rect 185261 521410 186207 521584
rect 186365 521410 186943 521584
rect 187285 521410 187403 521584
rect 172289 521142 172407 521316
rect 172565 521142 173511 521316
rect 173669 521142 174615 521316
rect 174773 521142 175719 521316
rect 175877 521142 176823 521316
rect 176981 521142 177191 521316
rect 177533 521142 178479 521316
rect 178637 521142 179583 521316
rect 179741 521142 180687 521316
rect 180845 521142 181791 521316
rect 181949 521142 182343 521316
rect 182685 521142 183631 521316
rect 183789 521142 184735 521316
rect 184893 521142 185839 521316
rect 185997 521142 186943 521316
rect 187285 521142 187403 521316
rect 172289 520322 172407 520496
rect 172565 520322 173511 520496
rect 173669 520322 174615 520496
rect 174957 520322 175903 520496
rect 176061 520322 177007 520496
rect 177165 520322 178111 520496
rect 178269 520322 179215 520496
rect 179373 520322 179767 520496
rect 180109 520322 181055 520496
rect 181213 520322 182159 520496
rect 182317 520322 183263 520496
rect 183421 520322 184367 520496
rect 184525 520322 184919 520496
rect 185261 520322 186207 520496
rect 186365 520322 186943 520496
rect 187285 520322 187403 520496
rect 172289 520054 172407 520228
rect 172565 520054 173511 520228
rect 173669 520054 174615 520228
rect 174773 520054 175719 520228
rect 175877 520054 176823 520228
rect 176981 520054 177191 520228
rect 177533 520054 178479 520228
rect 178637 520054 179583 520228
rect 179741 520054 180687 520228
rect 180845 520054 181791 520228
rect 181949 520054 182343 520228
rect 182685 520054 183631 520228
rect 183789 520054 184735 520228
rect 184893 520054 185839 520228
rect 185997 520054 186943 520228
rect 187285 520054 187403 520228
rect 172289 519234 172407 519408
rect 172565 519234 173511 519408
rect 173669 519234 174615 519408
rect 174957 519234 175903 519408
rect 176061 519234 177007 519408
rect 177165 519234 178111 519408
rect 178269 519234 179215 519408
rect 179373 519234 179767 519408
rect 180109 519234 181055 519408
rect 181213 519234 182159 519408
rect 182317 519234 183263 519408
rect 183421 519234 184367 519408
rect 184525 519234 184919 519408
rect 185261 519234 186207 519408
rect 186365 519234 186943 519408
rect 187285 519234 187403 519408
rect 172289 518966 172407 519140
rect 172565 518966 173511 519140
rect 173669 518966 174615 519140
rect 174773 518966 175719 519140
rect 175877 518966 176823 519140
rect 176981 518966 177191 519140
rect 177533 518966 178479 519140
rect 178637 518966 179583 519140
rect 179741 518966 180687 519140
rect 180845 518966 181791 519140
rect 181949 518966 182343 519140
rect 182685 518966 183631 519140
rect 183789 518966 184735 519140
rect 184893 518966 185839 519140
rect 185997 518966 186943 519140
rect 187285 518966 187403 519140
rect 172289 518146 172407 518320
rect 172565 518146 173511 518320
rect 173669 518146 174615 518320
rect 174957 518146 175903 518320
rect 176061 518146 177007 518320
rect 177165 518146 178111 518320
rect 178269 518146 179215 518320
rect 179373 518146 179767 518320
rect 180109 518146 181055 518320
rect 181213 518146 182159 518320
rect 182317 518146 183263 518320
rect 183421 518146 184367 518320
rect 184525 518146 184919 518320
rect 185261 518146 186207 518320
rect 186365 518146 186943 518320
rect 187285 518146 187403 518320
rect 172289 517878 172407 518052
rect 172565 517878 173511 518052
rect 173669 517878 174615 518052
rect 174773 517878 175719 518052
rect 175877 517878 176823 518052
rect 176981 517878 177191 518052
rect 177533 517878 178479 518052
rect 178637 517878 179583 518052
rect 179741 517878 180687 518052
rect 180845 517878 181791 518052
rect 181949 517878 182343 518052
rect 182685 517878 183631 518052
rect 183789 517878 184735 518052
rect 184893 517878 185839 518052
rect 185997 517878 186943 518052
rect 187285 517878 187403 518052
rect 172289 517058 172407 517232
rect 172565 517058 173511 517232
rect 173669 517058 174615 517232
rect 174957 517058 175903 517232
rect 176061 517058 177007 517232
rect 177165 517058 178111 517232
rect 178269 517058 179215 517232
rect 179373 517058 179767 517232
rect 180109 517058 181055 517232
rect 181213 517058 182159 517232
rect 182317 517058 183263 517232
rect 183421 517058 184367 517232
rect 184525 517058 184919 517232
rect 185261 517058 186207 517232
rect 186365 517058 186943 517232
rect 187285 517058 187403 517232
rect 172289 516790 172407 516964
rect 172565 516790 173511 516964
rect 173669 516790 174615 516964
rect 174773 516790 175719 516964
rect 175877 516790 176823 516964
rect 176981 516790 177191 516964
rect 177533 516790 178479 516964
rect 178637 516790 179583 516964
rect 179741 516790 180687 516964
rect 180845 516790 181791 516964
rect 181949 516790 182343 516964
rect 182685 516790 183631 516964
rect 183789 516790 184735 516964
rect 184893 516790 185839 516964
rect 185997 516790 186943 516964
rect 187285 516790 187403 516964
rect 172289 515970 172407 516144
rect 172565 515970 173511 516144
rect 173669 515970 174615 516144
rect 174957 515970 175903 516144
rect 176061 515970 177007 516144
rect 177165 515970 178111 516144
rect 178269 515970 179215 516144
rect 179373 515970 179767 516144
rect 180109 515970 181055 516144
rect 181213 515970 182159 516144
rect 182317 515970 183263 516144
rect 183421 515970 184367 516144
rect 184525 515970 184919 516144
rect 185261 515970 186207 516144
rect 186365 515970 186943 516144
rect 187285 515970 187403 516144
rect 172289 515702 172407 515876
rect 172565 515702 173143 515876
rect 173486 515676 173516 515876
rect 173582 515676 173612 515876
rect 173668 515676 173698 515876
rect 173754 515676 173784 515876
rect 173840 515676 173870 515876
rect 174037 515702 174615 515876
rect 174957 515702 175903 515876
rect 176061 515702 177007 515876
rect 177165 515702 177283 515876
rect 177533 515702 178479 515876
rect 178637 515702 179583 515876
rect 179741 515702 179859 515876
rect 180109 515702 181055 515876
rect 181213 515702 181791 515876
rect 182133 515718 182163 515876
rect 182221 515718 182251 515876
rect 182685 515702 183631 515876
rect 183789 515702 184735 515876
rect 184893 515702 185011 515876
rect 185261 515702 186207 515876
rect 186458 515676 186488 515876
rect 186554 515676 186584 515876
rect 186640 515676 186670 515876
rect 186726 515676 186756 515876
rect 186812 515676 186842 515876
rect 187009 515702 187127 515876
rect 187285 515702 187403 515876
<< ndiff >>
rect 164674 541067 164732 541079
rect 164674 540091 164686 541067
rect 164720 540091 164732 541067
rect 164674 540079 164732 540091
rect 164762 541067 164820 541079
rect 164762 540091 164774 541067
rect 164808 540091 164820 541067
rect 164762 540079 164820 540091
rect 164877 541074 164939 541086
rect 164877 540098 164889 541074
rect 164923 540098 164939 541074
rect 164877 540086 164939 540098
rect 164969 541074 165035 541086
rect 164969 540098 164985 541074
rect 165019 540098 165035 541074
rect 164969 540086 165035 540098
rect 165065 541074 165131 541086
rect 165065 540098 165081 541074
rect 165115 540098 165131 541074
rect 165065 540086 165131 540098
rect 165161 541074 165227 541086
rect 165161 540098 165177 541074
rect 165211 540098 165227 541074
rect 165161 540086 165227 540098
rect 165257 541074 165323 541086
rect 165257 540098 165273 541074
rect 165307 540098 165323 541074
rect 165257 540086 165323 540098
rect 165353 541074 165419 541086
rect 165353 540098 165369 541074
rect 165403 540098 165419 541074
rect 165353 540086 165419 540098
rect 165449 541074 165515 541086
rect 165449 540098 165465 541074
rect 165499 540098 165515 541074
rect 165449 540086 165515 540098
rect 165545 541074 165611 541086
rect 165545 540098 165561 541074
rect 165595 540098 165611 541074
rect 165545 540086 165611 540098
rect 165641 541074 165707 541086
rect 165641 540098 165657 541074
rect 165691 540098 165707 541074
rect 165641 540086 165707 540098
rect 165737 541074 165803 541086
rect 165737 540098 165753 541074
rect 165787 540098 165803 541074
rect 165737 540086 165803 540098
rect 165833 541074 165899 541086
rect 165833 540098 165849 541074
rect 165883 540098 165899 541074
rect 165833 540086 165899 540098
rect 165929 541074 165995 541086
rect 165929 540098 165945 541074
rect 165979 540098 165995 541074
rect 165929 540086 165995 540098
rect 166025 541074 166087 541086
rect 166025 540098 166041 541074
rect 166075 540098 166087 541074
rect 166354 541067 166412 541079
rect 166025 540086 166087 540098
rect 166154 540267 166212 540279
rect 166154 540091 166166 540267
rect 166200 540091 166212 540267
rect 166154 540079 166212 540091
rect 166242 540267 166300 540279
rect 166242 540091 166254 540267
rect 166288 540091 166300 540267
rect 166242 540079 166300 540091
rect 166354 540091 166366 541067
rect 166400 540091 166412 541067
rect 166354 540079 166412 540091
rect 166442 541067 166500 541079
rect 166442 540091 166454 541067
rect 166488 540091 166500 541067
rect 166442 540079 166500 540091
rect 168474 541067 168532 541079
rect 168474 540091 168486 541067
rect 168520 540091 168532 541067
rect 168474 540079 168532 540091
rect 168562 541067 168620 541079
rect 168562 540091 168574 541067
rect 168608 540091 168620 541067
rect 168562 540079 168620 540091
rect 168677 541074 168739 541086
rect 168677 540098 168689 541074
rect 168723 540098 168739 541074
rect 168677 540086 168739 540098
rect 168769 541074 168835 541086
rect 168769 540098 168785 541074
rect 168819 540098 168835 541074
rect 168769 540086 168835 540098
rect 168865 541074 168931 541086
rect 168865 540098 168881 541074
rect 168915 540098 168931 541074
rect 168865 540086 168931 540098
rect 168961 541074 169027 541086
rect 168961 540098 168977 541074
rect 169011 540098 169027 541074
rect 168961 540086 169027 540098
rect 169057 541074 169123 541086
rect 169057 540098 169073 541074
rect 169107 540098 169123 541074
rect 169057 540086 169123 540098
rect 169153 541074 169219 541086
rect 169153 540098 169169 541074
rect 169203 540098 169219 541074
rect 169153 540086 169219 540098
rect 169249 541074 169315 541086
rect 169249 540098 169265 541074
rect 169299 540098 169315 541074
rect 169249 540086 169315 540098
rect 169345 541074 169411 541086
rect 169345 540098 169361 541074
rect 169395 540098 169411 541074
rect 169345 540086 169411 540098
rect 169441 541074 169507 541086
rect 169441 540098 169457 541074
rect 169491 540098 169507 541074
rect 169441 540086 169507 540098
rect 169537 541074 169603 541086
rect 169537 540098 169553 541074
rect 169587 540098 169603 541074
rect 169537 540086 169603 540098
rect 169633 541074 169699 541086
rect 169633 540098 169649 541074
rect 169683 540098 169699 541074
rect 169633 540086 169699 540098
rect 169729 541074 169795 541086
rect 169729 540098 169745 541074
rect 169779 540098 169795 541074
rect 169729 540086 169795 540098
rect 169825 541074 169887 541086
rect 169825 540098 169841 541074
rect 169875 540098 169887 541074
rect 170154 541067 170212 541079
rect 169825 540086 169887 540098
rect 169954 540267 170012 540279
rect 169954 540091 169966 540267
rect 170000 540091 170012 540267
rect 169954 540079 170012 540091
rect 170042 540267 170100 540279
rect 170042 540091 170054 540267
rect 170088 540091 170100 540267
rect 170042 540079 170100 540091
rect 170154 540091 170166 541067
rect 170200 540091 170212 541067
rect 170154 540079 170212 540091
rect 170242 541067 170300 541079
rect 170242 540091 170254 541067
rect 170288 540091 170300 541067
rect 170242 540079 170300 540091
rect 172174 541067 172232 541079
rect 172174 540091 172186 541067
rect 172220 540091 172232 541067
rect 172174 540079 172232 540091
rect 172262 541067 172320 541079
rect 172262 540091 172274 541067
rect 172308 540091 172320 541067
rect 172262 540079 172320 540091
rect 172377 541074 172439 541086
rect 172377 540098 172389 541074
rect 172423 540098 172439 541074
rect 172377 540086 172439 540098
rect 172469 541074 172535 541086
rect 172469 540098 172485 541074
rect 172519 540098 172535 541074
rect 172469 540086 172535 540098
rect 172565 541074 172631 541086
rect 172565 540098 172581 541074
rect 172615 540098 172631 541074
rect 172565 540086 172631 540098
rect 172661 541074 172727 541086
rect 172661 540098 172677 541074
rect 172711 540098 172727 541074
rect 172661 540086 172727 540098
rect 172757 541074 172823 541086
rect 172757 540098 172773 541074
rect 172807 540098 172823 541074
rect 172757 540086 172823 540098
rect 172853 541074 172919 541086
rect 172853 540098 172869 541074
rect 172903 540098 172919 541074
rect 172853 540086 172919 540098
rect 172949 541074 173015 541086
rect 172949 540098 172965 541074
rect 172999 540098 173015 541074
rect 172949 540086 173015 540098
rect 173045 541074 173111 541086
rect 173045 540098 173061 541074
rect 173095 540098 173111 541074
rect 173045 540086 173111 540098
rect 173141 541074 173207 541086
rect 173141 540098 173157 541074
rect 173191 540098 173207 541074
rect 173141 540086 173207 540098
rect 173237 541074 173303 541086
rect 173237 540098 173253 541074
rect 173287 540098 173303 541074
rect 173237 540086 173303 540098
rect 173333 541074 173399 541086
rect 173333 540098 173349 541074
rect 173383 540098 173399 541074
rect 173333 540086 173399 540098
rect 173429 541074 173495 541086
rect 173429 540098 173445 541074
rect 173479 540098 173495 541074
rect 173429 540086 173495 540098
rect 173525 541074 173587 541086
rect 173525 540098 173541 541074
rect 173575 540098 173587 541074
rect 173854 541067 173912 541079
rect 173525 540086 173587 540098
rect 173654 540267 173712 540279
rect 173654 540091 173666 540267
rect 173700 540091 173712 540267
rect 173654 540079 173712 540091
rect 173742 540267 173800 540279
rect 173742 540091 173754 540267
rect 173788 540091 173800 540267
rect 173742 540079 173800 540091
rect 173854 540091 173866 541067
rect 173900 540091 173912 541067
rect 173854 540079 173912 540091
rect 173942 541067 174000 541079
rect 173942 540091 173954 541067
rect 173988 540091 174000 541067
rect 173942 540079 174000 540091
rect 175674 541067 175732 541079
rect 175674 540091 175686 541067
rect 175720 540091 175732 541067
rect 175674 540079 175732 540091
rect 175762 541067 175820 541079
rect 175762 540091 175774 541067
rect 175808 540091 175820 541067
rect 175762 540079 175820 540091
rect 175877 541074 175939 541086
rect 175877 540098 175889 541074
rect 175923 540098 175939 541074
rect 175877 540086 175939 540098
rect 175969 541074 176035 541086
rect 175969 540098 175985 541074
rect 176019 540098 176035 541074
rect 175969 540086 176035 540098
rect 176065 541074 176131 541086
rect 176065 540098 176081 541074
rect 176115 540098 176131 541074
rect 176065 540086 176131 540098
rect 176161 541074 176227 541086
rect 176161 540098 176177 541074
rect 176211 540098 176227 541074
rect 176161 540086 176227 540098
rect 176257 541074 176323 541086
rect 176257 540098 176273 541074
rect 176307 540098 176323 541074
rect 176257 540086 176323 540098
rect 176353 541074 176419 541086
rect 176353 540098 176369 541074
rect 176403 540098 176419 541074
rect 176353 540086 176419 540098
rect 176449 541074 176515 541086
rect 176449 540098 176465 541074
rect 176499 540098 176515 541074
rect 176449 540086 176515 540098
rect 176545 541074 176611 541086
rect 176545 540098 176561 541074
rect 176595 540098 176611 541074
rect 176545 540086 176611 540098
rect 176641 541074 176707 541086
rect 176641 540098 176657 541074
rect 176691 540098 176707 541074
rect 176641 540086 176707 540098
rect 176737 541074 176803 541086
rect 176737 540098 176753 541074
rect 176787 540098 176803 541074
rect 176737 540086 176803 540098
rect 176833 541074 176899 541086
rect 176833 540098 176849 541074
rect 176883 540098 176899 541074
rect 176833 540086 176899 540098
rect 176929 541074 176995 541086
rect 176929 540098 176945 541074
rect 176979 540098 176995 541074
rect 176929 540086 176995 540098
rect 177025 541074 177087 541086
rect 177025 540098 177041 541074
rect 177075 540098 177087 541074
rect 177354 541067 177412 541079
rect 177025 540086 177087 540098
rect 177154 540267 177212 540279
rect 177154 540091 177166 540267
rect 177200 540091 177212 540267
rect 177154 540079 177212 540091
rect 177242 540267 177300 540279
rect 177242 540091 177254 540267
rect 177288 540091 177300 540267
rect 177242 540079 177300 540091
rect 177354 540091 177366 541067
rect 177400 540091 177412 541067
rect 177354 540079 177412 540091
rect 177442 541067 177500 541079
rect 177442 540091 177454 541067
rect 177488 540091 177500 541067
rect 177442 540079 177500 540091
rect 179274 541067 179332 541079
rect 179274 540091 179286 541067
rect 179320 540091 179332 541067
rect 179274 540079 179332 540091
rect 179362 541067 179420 541079
rect 179362 540091 179374 541067
rect 179408 540091 179420 541067
rect 179362 540079 179420 540091
rect 179477 541074 179539 541086
rect 179477 540098 179489 541074
rect 179523 540098 179539 541074
rect 179477 540086 179539 540098
rect 179569 541074 179635 541086
rect 179569 540098 179585 541074
rect 179619 540098 179635 541074
rect 179569 540086 179635 540098
rect 179665 541074 179731 541086
rect 179665 540098 179681 541074
rect 179715 540098 179731 541074
rect 179665 540086 179731 540098
rect 179761 541074 179827 541086
rect 179761 540098 179777 541074
rect 179811 540098 179827 541074
rect 179761 540086 179827 540098
rect 179857 541074 179923 541086
rect 179857 540098 179873 541074
rect 179907 540098 179923 541074
rect 179857 540086 179923 540098
rect 179953 541074 180019 541086
rect 179953 540098 179969 541074
rect 180003 540098 180019 541074
rect 179953 540086 180019 540098
rect 180049 541074 180115 541086
rect 180049 540098 180065 541074
rect 180099 540098 180115 541074
rect 180049 540086 180115 540098
rect 180145 541074 180211 541086
rect 180145 540098 180161 541074
rect 180195 540098 180211 541074
rect 180145 540086 180211 540098
rect 180241 541074 180307 541086
rect 180241 540098 180257 541074
rect 180291 540098 180307 541074
rect 180241 540086 180307 540098
rect 180337 541074 180403 541086
rect 180337 540098 180353 541074
rect 180387 540098 180403 541074
rect 180337 540086 180403 540098
rect 180433 541074 180499 541086
rect 180433 540098 180449 541074
rect 180483 540098 180499 541074
rect 180433 540086 180499 540098
rect 180529 541074 180595 541086
rect 180529 540098 180545 541074
rect 180579 540098 180595 541074
rect 180529 540086 180595 540098
rect 180625 541074 180687 541086
rect 180625 540098 180641 541074
rect 180675 540098 180687 541074
rect 180954 541067 181012 541079
rect 180625 540086 180687 540098
rect 180754 540267 180812 540279
rect 180754 540091 180766 540267
rect 180800 540091 180812 540267
rect 180754 540079 180812 540091
rect 180842 540267 180900 540279
rect 180842 540091 180854 540267
rect 180888 540091 180900 540267
rect 180842 540079 180900 540091
rect 180954 540091 180966 541067
rect 181000 540091 181012 541067
rect 180954 540079 181012 540091
rect 181042 541067 181100 541079
rect 181042 540091 181054 541067
rect 181088 540091 181100 541067
rect 181042 540079 181100 540091
rect 182574 541067 182632 541079
rect 182574 540091 182586 541067
rect 182620 540091 182632 541067
rect 182574 540079 182632 540091
rect 182662 541067 182720 541079
rect 182662 540091 182674 541067
rect 182708 540091 182720 541067
rect 182662 540079 182720 540091
rect 182777 541074 182839 541086
rect 182777 540098 182789 541074
rect 182823 540098 182839 541074
rect 182777 540086 182839 540098
rect 182869 541074 182935 541086
rect 182869 540098 182885 541074
rect 182919 540098 182935 541074
rect 182869 540086 182935 540098
rect 182965 541074 183031 541086
rect 182965 540098 182981 541074
rect 183015 540098 183031 541074
rect 182965 540086 183031 540098
rect 183061 541074 183127 541086
rect 183061 540098 183077 541074
rect 183111 540098 183127 541074
rect 183061 540086 183127 540098
rect 183157 541074 183223 541086
rect 183157 540098 183173 541074
rect 183207 540098 183223 541074
rect 183157 540086 183223 540098
rect 183253 541074 183319 541086
rect 183253 540098 183269 541074
rect 183303 540098 183319 541074
rect 183253 540086 183319 540098
rect 183349 541074 183415 541086
rect 183349 540098 183365 541074
rect 183399 540098 183415 541074
rect 183349 540086 183415 540098
rect 183445 541074 183511 541086
rect 183445 540098 183461 541074
rect 183495 540098 183511 541074
rect 183445 540086 183511 540098
rect 183541 541074 183607 541086
rect 183541 540098 183557 541074
rect 183591 540098 183607 541074
rect 183541 540086 183607 540098
rect 183637 541074 183703 541086
rect 183637 540098 183653 541074
rect 183687 540098 183703 541074
rect 183637 540086 183703 540098
rect 183733 541074 183799 541086
rect 183733 540098 183749 541074
rect 183783 540098 183799 541074
rect 183733 540086 183799 540098
rect 183829 541074 183895 541086
rect 183829 540098 183845 541074
rect 183879 540098 183895 541074
rect 183829 540086 183895 540098
rect 183925 541074 183987 541086
rect 183925 540098 183941 541074
rect 183975 540098 183987 541074
rect 184254 541067 184312 541079
rect 183925 540086 183987 540098
rect 184054 540267 184112 540279
rect 184054 540091 184066 540267
rect 184100 540091 184112 540267
rect 184054 540079 184112 540091
rect 184142 540267 184200 540279
rect 184142 540091 184154 540267
rect 184188 540091 184200 540267
rect 184142 540079 184200 540091
rect 184254 540091 184266 541067
rect 184300 540091 184312 541067
rect 184254 540079 184312 540091
rect 184342 541067 184400 541079
rect 184342 540091 184354 541067
rect 184388 540091 184400 541067
rect 184342 540079 184400 540091
rect 185874 541067 185932 541079
rect 185874 540091 185886 541067
rect 185920 540091 185932 541067
rect 185874 540079 185932 540091
rect 185962 541067 186020 541079
rect 185962 540091 185974 541067
rect 186008 540091 186020 541067
rect 185962 540079 186020 540091
rect 186077 541074 186139 541086
rect 186077 540098 186089 541074
rect 186123 540098 186139 541074
rect 186077 540086 186139 540098
rect 186169 541074 186235 541086
rect 186169 540098 186185 541074
rect 186219 540098 186235 541074
rect 186169 540086 186235 540098
rect 186265 541074 186331 541086
rect 186265 540098 186281 541074
rect 186315 540098 186331 541074
rect 186265 540086 186331 540098
rect 186361 541074 186427 541086
rect 186361 540098 186377 541074
rect 186411 540098 186427 541074
rect 186361 540086 186427 540098
rect 186457 541074 186523 541086
rect 186457 540098 186473 541074
rect 186507 540098 186523 541074
rect 186457 540086 186523 540098
rect 186553 541074 186619 541086
rect 186553 540098 186569 541074
rect 186603 540098 186619 541074
rect 186553 540086 186619 540098
rect 186649 541074 186715 541086
rect 186649 540098 186665 541074
rect 186699 540098 186715 541074
rect 186649 540086 186715 540098
rect 186745 541074 186811 541086
rect 186745 540098 186761 541074
rect 186795 540098 186811 541074
rect 186745 540086 186811 540098
rect 186841 541074 186907 541086
rect 186841 540098 186857 541074
rect 186891 540098 186907 541074
rect 186841 540086 186907 540098
rect 186937 541074 187003 541086
rect 186937 540098 186953 541074
rect 186987 540098 187003 541074
rect 186937 540086 187003 540098
rect 187033 541074 187099 541086
rect 187033 540098 187049 541074
rect 187083 540098 187099 541074
rect 187033 540086 187099 540098
rect 187129 541074 187195 541086
rect 187129 540098 187145 541074
rect 187179 540098 187195 541074
rect 187129 540086 187195 540098
rect 187225 541074 187287 541086
rect 187225 540098 187241 541074
rect 187275 540098 187287 541074
rect 187554 541067 187612 541079
rect 187225 540086 187287 540098
rect 187354 540267 187412 540279
rect 187354 540091 187366 540267
rect 187400 540091 187412 540267
rect 187354 540079 187412 540091
rect 187442 540267 187500 540279
rect 187442 540091 187454 540267
rect 187488 540091 187500 540267
rect 187442 540079 187500 540091
rect 187554 540091 187566 541067
rect 187600 540091 187612 541067
rect 187554 540079 187612 540091
rect 187642 541067 187700 541079
rect 187642 540091 187654 541067
rect 187688 540091 187700 541067
rect 187642 540079 187700 540091
rect 189174 541067 189232 541079
rect 189174 540091 189186 541067
rect 189220 540091 189232 541067
rect 189174 540079 189232 540091
rect 189262 541067 189320 541079
rect 189262 540091 189274 541067
rect 189308 540091 189320 541067
rect 189262 540079 189320 540091
rect 189377 541074 189439 541086
rect 189377 540098 189389 541074
rect 189423 540098 189439 541074
rect 189377 540086 189439 540098
rect 189469 541074 189535 541086
rect 189469 540098 189485 541074
rect 189519 540098 189535 541074
rect 189469 540086 189535 540098
rect 189565 541074 189631 541086
rect 189565 540098 189581 541074
rect 189615 540098 189631 541074
rect 189565 540086 189631 540098
rect 189661 541074 189727 541086
rect 189661 540098 189677 541074
rect 189711 540098 189727 541074
rect 189661 540086 189727 540098
rect 189757 541074 189823 541086
rect 189757 540098 189773 541074
rect 189807 540098 189823 541074
rect 189757 540086 189823 540098
rect 189853 541074 189919 541086
rect 189853 540098 189869 541074
rect 189903 540098 189919 541074
rect 189853 540086 189919 540098
rect 189949 541074 190015 541086
rect 189949 540098 189965 541074
rect 189999 540098 190015 541074
rect 189949 540086 190015 540098
rect 190045 541074 190111 541086
rect 190045 540098 190061 541074
rect 190095 540098 190111 541074
rect 190045 540086 190111 540098
rect 190141 541074 190207 541086
rect 190141 540098 190157 541074
rect 190191 540098 190207 541074
rect 190141 540086 190207 540098
rect 190237 541074 190303 541086
rect 190237 540098 190253 541074
rect 190287 540098 190303 541074
rect 190237 540086 190303 540098
rect 190333 541074 190399 541086
rect 190333 540098 190349 541074
rect 190383 540098 190399 541074
rect 190333 540086 190399 540098
rect 190429 541074 190495 541086
rect 190429 540098 190445 541074
rect 190479 540098 190495 541074
rect 190429 540086 190495 540098
rect 190525 541074 190587 541086
rect 190525 540098 190541 541074
rect 190575 540098 190587 541074
rect 190854 541067 190912 541079
rect 190525 540086 190587 540098
rect 190654 540267 190712 540279
rect 190654 540091 190666 540267
rect 190700 540091 190712 540267
rect 190654 540079 190712 540091
rect 190742 540267 190800 540279
rect 190742 540091 190754 540267
rect 190788 540091 190800 540267
rect 190742 540079 190800 540091
rect 190854 540091 190866 541067
rect 190900 540091 190912 541067
rect 190854 540079 190912 540091
rect 190942 541067 191000 541079
rect 190942 540091 190954 541067
rect 190988 540091 191000 541067
rect 190942 540079 191000 540091
rect 158654 538417 158712 538429
rect 158654 538241 158666 538417
rect 158700 538241 158712 538417
rect 158654 538229 158712 538241
rect 158912 538417 158970 538429
rect 158912 538241 158924 538417
rect 158958 538241 158970 538417
rect 158912 538229 158970 538241
rect 159030 538417 159088 538429
rect 159030 538241 159042 538417
rect 159076 538241 159088 538417
rect 159030 538229 159088 538241
rect 159288 538417 159346 538429
rect 159288 538241 159300 538417
rect 159334 538241 159346 538417
rect 159288 538229 159346 538241
rect 159546 538417 159604 538429
rect 159546 538241 159558 538417
rect 159592 538241 159604 538417
rect 159546 538229 159604 538241
rect 159804 538417 159862 538429
rect 159804 538241 159816 538417
rect 159850 538241 159862 538417
rect 159804 538229 159862 538241
rect 160062 538417 160120 538429
rect 160062 538241 160074 538417
rect 160108 538241 160120 538417
rect 160062 538229 160120 538241
rect 160320 538417 160378 538429
rect 160320 538241 160332 538417
rect 160366 538241 160378 538417
rect 160320 538229 160378 538241
rect 160578 538417 160636 538429
rect 160578 538241 160590 538417
rect 160624 538241 160636 538417
rect 160578 538229 160636 538241
rect 160836 538417 160894 538429
rect 160836 538241 160848 538417
rect 160882 538241 160894 538417
rect 160836 538229 160894 538241
rect 161094 538417 161152 538429
rect 161094 538241 161106 538417
rect 161140 538241 161152 538417
rect 161094 538229 161152 538241
rect 161352 538417 161410 538429
rect 161352 538241 161364 538417
rect 161398 538241 161410 538417
rect 161352 538229 161410 538241
rect 161474 538417 161532 538429
rect 161474 538241 161486 538417
rect 161520 538241 161532 538417
rect 161474 538229 161532 538241
rect 161732 538417 161790 538429
rect 161732 538241 161744 538417
rect 161778 538241 161790 538417
rect 161732 538229 161790 538241
rect 161874 538417 161932 538429
rect 161874 538241 161886 538417
rect 161920 538241 161932 538417
rect 161874 538229 161932 538241
rect 162132 538417 162190 538429
rect 162132 538241 162144 538417
rect 162178 538241 162190 538417
rect 162132 538229 162190 538241
rect 162254 538417 162312 538429
rect 162254 538241 162266 538417
rect 162300 538241 162312 538417
rect 162254 538229 162312 538241
rect 162512 538417 162570 538429
rect 162512 538241 162524 538417
rect 162558 538241 162570 538417
rect 162512 538229 162570 538241
rect 172237 530531 172289 530564
rect 172237 530497 172245 530531
rect 172279 530497 172289 530531
rect 172237 530454 172289 530497
rect 172407 530531 172459 530564
rect 172407 530497 172417 530531
rect 172451 530497 172459 530531
rect 172407 530454 172459 530497
rect 172515 530548 172573 530564
rect 172515 530514 172528 530548
rect 172562 530514 172573 530548
rect 172515 530480 172573 530514
rect 172603 530526 172659 530564
rect 172603 530492 172614 530526
rect 172648 530492 172659 530526
rect 172603 530480 172659 530492
rect 172689 530548 172745 530564
rect 172689 530514 172700 530548
rect 172734 530514 172745 530548
rect 172689 530480 172745 530514
rect 172775 530526 172831 530564
rect 172775 530492 172786 530526
rect 172820 530492 172831 530526
rect 172775 530480 172831 530492
rect 172861 530548 172928 530564
rect 172861 530514 172883 530548
rect 172917 530514 172928 530548
rect 172861 530480 172928 530514
rect 172958 530544 173011 530564
rect 172958 530510 172969 530544
rect 173003 530510 173011 530544
rect 172958 530480 173011 530510
rect 173065 530533 173117 530564
rect 173065 530499 173073 530533
rect 173107 530499 173117 530533
rect 173065 530454 173117 530499
rect 174063 530533 174115 530564
rect 174063 530499 174073 530533
rect 174107 530499 174115 530533
rect 174063 530454 174115 530499
rect 174169 530533 174221 530564
rect 174169 530499 174177 530533
rect 174211 530499 174221 530533
rect 174169 530454 174221 530499
rect 174615 530533 174667 530564
rect 174907 530548 174965 530564
rect 174615 530499 174625 530533
rect 174659 530499 174667 530533
rect 174615 530454 174667 530499
rect 174907 530514 174920 530548
rect 174954 530514 174965 530548
rect 174907 530480 174965 530514
rect 174995 530526 175051 530564
rect 174995 530492 175006 530526
rect 175040 530492 175051 530526
rect 174995 530480 175051 530492
rect 175081 530548 175137 530564
rect 175081 530514 175092 530548
rect 175126 530514 175137 530548
rect 175081 530480 175137 530514
rect 175167 530526 175223 530564
rect 175167 530492 175178 530526
rect 175212 530492 175223 530526
rect 175167 530480 175223 530492
rect 175253 530548 175320 530564
rect 175253 530514 175275 530548
rect 175309 530514 175320 530548
rect 175253 530480 175320 530514
rect 175350 530544 175403 530564
rect 175350 530510 175361 530544
rect 175395 530510 175403 530544
rect 175350 530480 175403 530510
rect 175549 530502 175601 530564
rect 175549 530468 175557 530502
rect 175591 530468 175601 530502
rect 175549 530434 175601 530468
rect 175631 530552 175703 530564
rect 175631 530518 175641 530552
rect 175675 530518 175703 530552
rect 175631 530480 175703 530518
rect 175757 530536 175809 530564
rect 175757 530502 175765 530536
rect 175799 530502 175809 530536
rect 175757 530480 175809 530502
rect 175839 530480 175900 530564
rect 175930 530556 176049 530564
rect 175930 530522 175983 530556
rect 176017 530522 176049 530556
rect 175930 530480 176049 530522
rect 176079 530492 176145 530564
rect 176175 530552 176254 530564
rect 176175 530518 176195 530552
rect 176229 530518 176254 530552
rect 176175 530492 176254 530518
rect 176284 530556 176353 530564
rect 176284 530522 176305 530556
rect 176339 530522 176353 530556
rect 176284 530492 176353 530522
rect 176079 530480 176129 530492
rect 175631 530434 175681 530480
rect 176299 530436 176353 530492
rect 176383 530552 176485 530564
rect 176383 530518 176417 530552
rect 176451 530518 176485 530552
rect 176383 530480 176485 530518
rect 176515 530480 176557 530564
rect 176587 530492 176723 530564
rect 176753 530550 176819 530564
rect 176753 530516 176763 530550
rect 176797 530516 176819 530550
rect 176753 530492 176819 530516
rect 176849 530550 176914 530564
rect 176849 530516 176870 530550
rect 176904 530516 176914 530550
rect 176849 530492 176914 530516
rect 176587 530480 176705 530492
rect 176383 530436 176433 530480
rect 176864 530480 176914 530492
rect 176944 530556 177049 530564
rect 176944 530522 177003 530556
rect 177037 530522 177049 530556
rect 176944 530480 177049 530522
rect 177117 530526 177169 530564
rect 177117 530492 177125 530526
rect 177159 530492 177169 530526
rect 177117 530480 177169 530492
rect 177199 530552 177253 530564
rect 177199 530518 177209 530552
rect 177243 530518 177253 530552
rect 177199 530480 177253 530518
rect 177283 530526 177335 530564
rect 177283 530492 177293 530526
rect 177327 530492 177335 530526
rect 177283 530480 177335 530492
rect 177684 530526 177736 530564
rect 177684 530492 177692 530526
rect 177726 530492 177736 530526
rect 177684 530434 177736 530492
rect 177766 530552 177831 530564
rect 177766 530518 177782 530552
rect 177816 530518 177831 530552
rect 177766 530480 177831 530518
rect 177931 530526 177983 530564
rect 177931 530492 177941 530526
rect 177975 530492 177983 530526
rect 177931 530480 177983 530492
rect 178037 530526 178089 530564
rect 178037 530492 178045 530526
rect 178079 530492 178089 530526
rect 178037 530480 178089 530492
rect 178189 530552 178243 530564
rect 178189 530518 178199 530552
rect 178233 530518 178243 530552
rect 178189 530480 178243 530518
rect 178273 530526 178325 530564
rect 178273 530492 178283 530526
rect 178317 530492 178325 530526
rect 178273 530480 178325 530492
rect 178401 530522 178453 530564
rect 178401 530488 178409 530522
rect 178443 530488 178453 530522
rect 177766 530434 177816 530480
rect 178401 530460 178453 530488
rect 178483 530552 178541 530564
rect 178483 530518 178495 530552
rect 178529 530518 178541 530552
rect 178483 530460 178541 530518
rect 178571 530539 178623 530564
rect 178571 530505 178581 530539
rect 178615 530505 178623 530539
rect 178571 530460 178623 530505
rect 178679 530548 178737 530564
rect 178679 530514 178692 530548
rect 178726 530514 178737 530548
rect 178679 530480 178737 530514
rect 178767 530526 178823 530564
rect 178767 530492 178778 530526
rect 178812 530492 178823 530526
rect 178767 530480 178823 530492
rect 178853 530548 178909 530564
rect 178853 530514 178864 530548
rect 178898 530514 178909 530548
rect 178853 530480 178909 530514
rect 178939 530526 178995 530564
rect 178939 530492 178950 530526
rect 178984 530492 178995 530526
rect 178939 530480 178995 530492
rect 179025 530548 179092 530564
rect 179025 530514 179047 530548
rect 179081 530514 179092 530548
rect 179025 530480 179092 530514
rect 179122 530544 179175 530564
rect 179122 530510 179133 530544
rect 179167 530510 179175 530544
rect 179122 530480 179175 530510
rect 179229 530544 179282 530564
rect 179229 530510 179237 530544
rect 179271 530510 179282 530544
rect 179229 530480 179282 530510
rect 179312 530548 179379 530564
rect 179312 530514 179323 530548
rect 179357 530514 179379 530548
rect 179312 530480 179379 530514
rect 179409 530526 179465 530564
rect 179409 530492 179420 530526
rect 179454 530492 179465 530526
rect 179409 530480 179465 530492
rect 179495 530548 179551 530564
rect 179495 530514 179506 530548
rect 179540 530514 179551 530548
rect 179495 530480 179551 530514
rect 179581 530526 179637 530564
rect 179581 530492 179592 530526
rect 179626 530492 179637 530526
rect 179581 530480 179637 530492
rect 179667 530548 179725 530564
rect 179667 530514 179678 530548
rect 179712 530514 179725 530548
rect 179667 530480 179725 530514
rect 180241 530533 180293 530564
rect 180241 530499 180249 530533
rect 180283 530499 180293 530533
rect 180241 530434 180293 530499
rect 180323 530552 180402 530564
rect 180323 530518 180333 530552
rect 180367 530518 180402 530552
rect 180323 530480 180402 530518
rect 180432 530480 180498 530564
rect 180528 530537 180623 530564
rect 180528 530503 180540 530537
rect 180574 530503 180623 530537
rect 180528 530480 180623 530503
rect 180653 530480 180719 530564
rect 180749 530537 180887 530564
rect 180749 530503 180775 530537
rect 180809 530503 180843 530537
rect 180877 530503 180887 530537
rect 180749 530480 180887 530503
rect 180917 530537 180969 530564
rect 180917 530503 180927 530537
rect 180961 530503 180969 530537
rect 180917 530480 180969 530503
rect 181207 530537 181259 530564
rect 181207 530503 181215 530537
rect 181249 530503 181259 530537
rect 181207 530480 181259 530503
rect 181289 530537 181427 530564
rect 181289 530503 181299 530537
rect 181333 530503 181367 530537
rect 181401 530503 181427 530537
rect 181289 530480 181427 530503
rect 181457 530480 181523 530564
rect 181553 530537 181648 530564
rect 181553 530503 181602 530537
rect 181636 530503 181648 530537
rect 181553 530480 181648 530503
rect 181678 530480 181744 530564
rect 181774 530552 181853 530564
rect 181774 530518 181809 530552
rect 181843 530518 181853 530552
rect 181774 530480 181853 530518
rect 180323 530434 180375 530480
rect 181801 530434 181853 530480
rect 181883 530533 181935 530564
rect 181883 530499 181893 530533
rect 181927 530499 181935 530533
rect 181883 530434 181935 530499
rect 181989 530544 182042 530564
rect 181989 530510 181997 530544
rect 182031 530510 182042 530544
rect 181989 530480 182042 530510
rect 182072 530548 182139 530564
rect 182072 530514 182083 530548
rect 182117 530514 182139 530548
rect 182072 530480 182139 530514
rect 182169 530526 182225 530564
rect 182169 530492 182180 530526
rect 182214 530492 182225 530526
rect 182169 530480 182225 530492
rect 182255 530548 182311 530564
rect 182255 530514 182266 530548
rect 182300 530514 182311 530548
rect 182255 530480 182311 530514
rect 182341 530526 182397 530564
rect 182341 530492 182352 530526
rect 182386 530492 182397 530526
rect 182341 530480 182397 530492
rect 182427 530548 182485 530564
rect 182427 530514 182438 530548
rect 182472 530514 182485 530548
rect 182427 530480 182485 530514
rect 182633 530526 182685 530564
rect 182633 530492 182641 530526
rect 182675 530492 182685 530526
rect 182633 530454 182685 530492
rect 182895 530526 182947 530564
rect 182895 530492 182905 530526
rect 182939 530492 182947 530526
rect 182895 530454 182947 530492
rect 183093 530544 183146 530564
rect 183093 530510 183101 530544
rect 183135 530510 183146 530544
rect 183093 530480 183146 530510
rect 183176 530548 183243 530564
rect 183176 530514 183187 530548
rect 183221 530514 183243 530548
rect 183176 530480 183243 530514
rect 183273 530526 183329 530564
rect 183273 530492 183284 530526
rect 183318 530492 183329 530526
rect 183273 530480 183329 530492
rect 183359 530548 183415 530564
rect 183359 530514 183370 530548
rect 183404 530514 183415 530548
rect 183359 530480 183415 530514
rect 183445 530526 183501 530564
rect 183445 530492 183456 530526
rect 183490 530492 183501 530526
rect 183445 530480 183501 530492
rect 183531 530548 183589 530564
rect 183531 530514 183542 530548
rect 183576 530514 183589 530548
rect 183531 530480 183589 530514
rect 183645 530533 183697 530564
rect 183645 530499 183653 530533
rect 183687 530499 183697 530533
rect 183645 530454 183697 530499
rect 184643 530533 184695 530564
rect 184643 530499 184653 530533
rect 184687 530499 184695 530533
rect 184643 530454 184695 530499
rect 184749 530526 184801 530564
rect 184749 530492 184757 530526
rect 184791 530492 184801 530526
rect 184749 530454 184801 530492
rect 185011 530526 185063 530564
rect 185011 530492 185021 530526
rect 185055 530492 185063 530526
rect 185011 530454 185063 530492
rect 185209 530544 185262 530564
rect 185209 530510 185217 530544
rect 185251 530510 185262 530544
rect 185209 530480 185262 530510
rect 185292 530548 185359 530564
rect 185292 530514 185303 530548
rect 185337 530514 185359 530548
rect 185292 530480 185359 530514
rect 185389 530526 185445 530564
rect 185389 530492 185400 530526
rect 185434 530492 185445 530526
rect 185389 530480 185445 530492
rect 185475 530548 185531 530564
rect 185475 530514 185486 530548
rect 185520 530514 185531 530548
rect 185475 530480 185531 530514
rect 185561 530526 185617 530564
rect 185561 530492 185572 530526
rect 185606 530492 185617 530526
rect 185561 530480 185617 530492
rect 185647 530548 185705 530564
rect 185647 530514 185658 530548
rect 185692 530514 185705 530548
rect 185647 530480 185705 530514
rect 185761 530533 185813 530564
rect 185761 530499 185769 530533
rect 185803 530499 185813 530533
rect 185761 530454 185813 530499
rect 186759 530533 186811 530564
rect 186759 530499 186769 530533
rect 186803 530499 186811 530533
rect 186759 530454 186811 530499
rect 187233 530531 187285 530564
rect 187233 530497 187241 530531
rect 187275 530497 187285 530531
rect 187233 530454 187285 530497
rect 187403 530531 187455 530564
rect 187403 530497 187413 530531
rect 187447 530497 187455 530531
rect 187403 530454 187455 530497
rect 172237 529637 172289 529680
rect 172237 529603 172245 529637
rect 172279 529603 172289 529637
rect 172237 529570 172289 529603
rect 172407 529637 172459 529680
rect 172407 529603 172417 529637
rect 172451 529603 172459 529637
rect 172407 529570 172459 529603
rect 172513 529635 172565 529680
rect 172513 529601 172521 529635
rect 172555 529601 172565 529635
rect 172513 529570 172565 529601
rect 173511 529635 173563 529680
rect 173511 529601 173521 529635
rect 173555 529601 173563 529635
rect 173511 529570 173563 529601
rect 173617 529635 173669 529680
rect 173617 529601 173625 529635
rect 173659 529601 173669 529635
rect 173617 529570 173669 529601
rect 174615 529635 174667 529680
rect 175344 529654 175394 529700
rect 174615 529601 174625 529635
rect 174659 529601 174667 529635
rect 174615 529570 174667 529601
rect 174835 529642 174887 529654
rect 174835 529608 174843 529642
rect 174877 529608 174887 529642
rect 174835 529570 174887 529608
rect 174917 529616 174971 529654
rect 174917 529582 174927 529616
rect 174961 529582 174971 529616
rect 174917 529570 174971 529582
rect 175071 529642 175123 529654
rect 175071 529608 175081 529642
rect 175115 529608 175123 529642
rect 175071 529570 175123 529608
rect 175177 529642 175229 529654
rect 175177 529608 175185 529642
rect 175219 529608 175229 529642
rect 175177 529570 175229 529608
rect 175329 529616 175394 529654
rect 175329 529582 175344 529616
rect 175378 529582 175394 529616
rect 175329 529570 175394 529582
rect 175424 529642 175476 529700
rect 175424 529608 175434 529642
rect 175468 529608 175476 529642
rect 175424 529570 175476 529608
rect 175549 529642 175601 529654
rect 175549 529608 175557 529642
rect 175591 529608 175601 529642
rect 175549 529570 175601 529608
rect 175631 529616 175685 529654
rect 175631 529582 175641 529616
rect 175675 529582 175685 529616
rect 175631 529570 175685 529582
rect 175715 529642 175767 529654
rect 175715 529608 175725 529642
rect 175759 529608 175767 529642
rect 175715 529570 175767 529608
rect 175835 529612 175940 529654
rect 175835 529578 175847 529612
rect 175881 529578 175940 529612
rect 175835 529570 175940 529578
rect 175970 529642 176020 529654
rect 176451 529654 176501 529698
rect 176179 529642 176297 529654
rect 175970 529618 176035 529642
rect 175970 529584 175980 529618
rect 176014 529584 176035 529618
rect 175970 529570 176035 529584
rect 176065 529618 176131 529642
rect 176065 529584 176087 529618
rect 176121 529584 176131 529618
rect 176065 529570 176131 529584
rect 176161 529570 176297 529642
rect 176327 529570 176369 529654
rect 176399 529616 176501 529654
rect 176399 529582 176433 529616
rect 176467 529582 176501 529616
rect 176399 529570 176501 529582
rect 176531 529642 176585 529698
rect 177203 529654 177253 529700
rect 176755 529642 176805 529654
rect 176531 529612 176600 529642
rect 176531 529578 176545 529612
rect 176579 529578 176600 529612
rect 176531 529570 176600 529578
rect 176630 529616 176709 529642
rect 176630 529582 176655 529616
rect 176689 529582 176709 529616
rect 176630 529570 176709 529582
rect 176739 529570 176805 529642
rect 176835 529612 176954 529654
rect 176835 529578 176867 529612
rect 176901 529578 176954 529612
rect 176835 529570 176954 529578
rect 176984 529570 177045 529654
rect 177075 529632 177127 529654
rect 177075 529598 177085 529632
rect 177119 529598 177127 529632
rect 177075 529570 177127 529598
rect 177181 529616 177253 529654
rect 177181 529582 177209 529616
rect 177243 529582 177253 529616
rect 177181 529570 177253 529582
rect 177283 529666 177335 529700
rect 177283 529632 177293 529666
rect 177327 529632 177335 529666
rect 177283 529570 177335 529632
rect 178213 529654 178265 529700
rect 177619 529631 177671 529654
rect 177619 529597 177627 529631
rect 177661 529597 177671 529631
rect 177619 529570 177671 529597
rect 177701 529631 177839 529654
rect 177701 529597 177711 529631
rect 177745 529597 177779 529631
rect 177813 529597 177839 529631
rect 177701 529570 177839 529597
rect 177869 529570 177935 529654
rect 177965 529631 178060 529654
rect 177965 529597 178014 529631
rect 178048 529597 178060 529631
rect 177965 529570 178060 529597
rect 178090 529570 178156 529654
rect 178186 529616 178265 529654
rect 178186 529582 178221 529616
rect 178255 529582 178265 529616
rect 178186 529570 178265 529582
rect 178295 529635 178347 529700
rect 178295 529601 178305 529635
rect 178339 529601 178347 529635
rect 178295 529570 178347 529601
rect 178401 529666 178453 529700
rect 178401 529632 178409 529666
rect 178443 529632 178453 529666
rect 178401 529570 178453 529632
rect 178483 529654 178533 529700
rect 178483 529616 178555 529654
rect 178483 529582 178493 529616
rect 178527 529582 178555 529616
rect 178483 529570 178555 529582
rect 178609 529632 178661 529654
rect 178609 529598 178617 529632
rect 178651 529598 178661 529632
rect 178609 529570 178661 529598
rect 178691 529570 178752 529654
rect 178782 529612 178901 529654
rect 178782 529578 178835 529612
rect 178869 529578 178901 529612
rect 178782 529570 178901 529578
rect 178931 529642 178981 529654
rect 179151 529642 179205 529698
rect 178931 529570 178997 529642
rect 179027 529616 179106 529642
rect 179027 529582 179047 529616
rect 179081 529582 179106 529616
rect 179027 529570 179106 529582
rect 179136 529612 179205 529642
rect 179136 529578 179157 529612
rect 179191 529578 179205 529612
rect 179136 529570 179205 529578
rect 179235 529654 179285 529698
rect 179235 529616 179337 529654
rect 179235 529582 179269 529616
rect 179303 529582 179337 529616
rect 179235 529570 179337 529582
rect 179367 529570 179409 529654
rect 179439 529642 179557 529654
rect 179716 529642 179766 529654
rect 179439 529570 179575 529642
rect 179605 529618 179671 529642
rect 179605 529584 179615 529618
rect 179649 529584 179671 529618
rect 179605 529570 179671 529584
rect 179701 529618 179766 529642
rect 179701 529584 179722 529618
rect 179756 529584 179766 529618
rect 179701 529570 179766 529584
rect 179796 529612 179901 529654
rect 179796 529578 179855 529612
rect 179889 529578 179901 529612
rect 179796 529570 179901 529578
rect 179969 529642 180021 529654
rect 179969 529608 179977 529642
rect 180011 529608 180021 529642
rect 179969 529570 180021 529608
rect 180051 529616 180105 529654
rect 180051 529582 180061 529616
rect 180095 529582 180105 529616
rect 180051 529570 180105 529582
rect 180135 529642 180187 529654
rect 180135 529608 180145 529642
rect 180179 529608 180187 529642
rect 180135 529570 180187 529608
rect 180241 529642 180293 529654
rect 180241 529608 180249 529642
rect 180283 529608 180293 529642
rect 180241 529570 180293 529608
rect 180323 529616 180377 529654
rect 180323 529582 180333 529616
rect 180367 529582 180377 529616
rect 180323 529570 180377 529582
rect 180407 529642 180459 529654
rect 180407 529608 180417 529642
rect 180451 529608 180459 529642
rect 180407 529570 180459 529608
rect 180527 529612 180632 529654
rect 180527 529578 180539 529612
rect 180573 529578 180632 529612
rect 180527 529570 180632 529578
rect 180662 529642 180712 529654
rect 181143 529654 181193 529698
rect 180871 529642 180989 529654
rect 180662 529618 180727 529642
rect 180662 529584 180672 529618
rect 180706 529584 180727 529618
rect 180662 529570 180727 529584
rect 180757 529618 180823 529642
rect 180757 529584 180779 529618
rect 180813 529584 180823 529618
rect 180757 529570 180823 529584
rect 180853 529570 180989 529642
rect 181019 529570 181061 529654
rect 181091 529616 181193 529654
rect 181091 529582 181125 529616
rect 181159 529582 181193 529616
rect 181091 529570 181193 529582
rect 181223 529642 181277 529698
rect 181895 529654 181945 529700
rect 181447 529642 181497 529654
rect 181223 529612 181292 529642
rect 181223 529578 181237 529612
rect 181271 529578 181292 529612
rect 181223 529570 181292 529578
rect 181322 529616 181401 529642
rect 181322 529582 181347 529616
rect 181381 529582 181401 529616
rect 181322 529570 181401 529582
rect 181431 529570 181497 529642
rect 181527 529612 181646 529654
rect 181527 529578 181559 529612
rect 181593 529578 181646 529612
rect 181527 529570 181646 529578
rect 181676 529570 181737 529654
rect 181767 529632 181819 529654
rect 181767 529598 181777 529632
rect 181811 529598 181819 529632
rect 181767 529570 181819 529598
rect 181873 529616 181945 529654
rect 181873 529582 181901 529616
rect 181935 529582 181945 529616
rect 181873 529570 181945 529582
rect 181975 529666 182027 529700
rect 181975 529632 181985 529666
rect 182019 529632 182027 529666
rect 181975 529570 182027 529632
rect 182081 529642 182133 529680
rect 182081 529608 182089 529642
rect 182123 529608 182133 529642
rect 182081 529570 182133 529608
rect 182343 529642 182395 529680
rect 182343 529608 182353 529642
rect 182387 529608 182395 529642
rect 182343 529570 182395 529608
rect 182652 529642 182704 529700
rect 182652 529608 182660 529642
rect 182694 529608 182704 529642
rect 182652 529570 182704 529608
rect 182734 529654 182784 529700
rect 182734 529616 182799 529654
rect 182734 529582 182750 529616
rect 182784 529582 182799 529616
rect 182734 529570 182799 529582
rect 182899 529642 182951 529654
rect 182899 529608 182909 529642
rect 182943 529608 182951 529642
rect 182899 529570 182951 529608
rect 183005 529642 183057 529654
rect 183005 529608 183013 529642
rect 183047 529608 183057 529642
rect 183005 529570 183057 529608
rect 183157 529616 183211 529654
rect 183157 529582 183167 529616
rect 183201 529582 183211 529616
rect 183157 529570 183211 529582
rect 183241 529642 183293 529654
rect 183241 529608 183251 529642
rect 183285 529608 183293 529642
rect 183241 529570 183293 529608
rect 183369 529635 183421 529680
rect 183369 529601 183377 529635
rect 183411 529601 183421 529635
rect 183369 529570 183421 529601
rect 184367 529635 184419 529680
rect 184367 529601 184377 529635
rect 184411 529601 184419 529635
rect 184367 529570 184419 529601
rect 184473 529635 184525 529680
rect 184473 529601 184481 529635
rect 184515 529601 184525 529635
rect 184473 529570 184525 529601
rect 185471 529635 185523 529680
rect 185471 529601 185481 529635
rect 185515 529601 185523 529635
rect 185471 529570 185523 529601
rect 185577 529635 185629 529680
rect 185577 529601 185585 529635
rect 185619 529601 185629 529635
rect 185577 529570 185629 529601
rect 186575 529635 186627 529680
rect 186575 529601 186585 529635
rect 186619 529601 186627 529635
rect 186575 529570 186627 529601
rect 186681 529635 186733 529680
rect 186681 529601 186689 529635
rect 186723 529601 186733 529635
rect 186681 529570 186733 529601
rect 187127 529635 187179 529680
rect 187127 529601 187137 529635
rect 187171 529601 187179 529635
rect 187127 529570 187179 529601
rect 187233 529637 187285 529680
rect 187233 529603 187241 529637
rect 187275 529603 187285 529637
rect 187233 529570 187285 529603
rect 187403 529637 187455 529680
rect 187403 529603 187413 529637
rect 187447 529603 187455 529637
rect 187403 529570 187455 529603
rect 172237 529443 172289 529476
rect 172237 529409 172245 529443
rect 172279 529409 172289 529443
rect 172237 529366 172289 529409
rect 172407 529443 172459 529476
rect 172407 529409 172417 529443
rect 172451 529409 172459 529443
rect 172407 529366 172459 529409
rect 172513 529445 172565 529476
rect 172513 529411 172521 529445
rect 172555 529411 172565 529445
rect 172513 529366 172565 529411
rect 173511 529445 173563 529476
rect 173511 529411 173521 529445
rect 173555 529411 173563 529445
rect 173511 529366 173563 529411
rect 173617 529445 173669 529476
rect 173617 529411 173625 529445
rect 173659 529411 173669 529445
rect 173617 529366 173669 529411
rect 174615 529445 174667 529476
rect 174615 529411 174625 529445
rect 174659 529411 174667 529445
rect 174615 529366 174667 529411
rect 175135 529449 175187 529476
rect 175135 529415 175143 529449
rect 175177 529415 175187 529449
rect 175135 529392 175187 529415
rect 175217 529449 175355 529476
rect 175217 529415 175227 529449
rect 175261 529415 175295 529449
rect 175329 529415 175355 529449
rect 175217 529392 175355 529415
rect 175385 529392 175451 529476
rect 175481 529449 175576 529476
rect 175481 529415 175530 529449
rect 175564 529415 175576 529449
rect 175481 529392 175576 529415
rect 175606 529392 175672 529476
rect 175702 529464 175781 529476
rect 175702 529430 175737 529464
rect 175771 529430 175781 529464
rect 175702 529392 175781 529430
rect 175729 529346 175781 529392
rect 175811 529445 175863 529476
rect 175811 529411 175821 529445
rect 175855 529411 175863 529445
rect 175811 529346 175863 529411
rect 175934 529460 175987 529476
rect 175934 529426 175942 529460
rect 175976 529426 175987 529460
rect 175934 529392 175987 529426
rect 176017 529451 176073 529476
rect 176017 529417 176028 529451
rect 176062 529417 176073 529451
rect 176017 529392 176073 529417
rect 176103 529460 176159 529476
rect 176103 529426 176114 529460
rect 176148 529426 176159 529460
rect 176103 529392 176159 529426
rect 176189 529451 176245 529476
rect 176189 529417 176200 529451
rect 176234 529417 176245 529451
rect 176189 529392 176245 529417
rect 176275 529460 176331 529476
rect 176275 529426 176286 529460
rect 176320 529426 176331 529460
rect 176275 529392 176331 529426
rect 176361 529451 176417 529476
rect 176361 529417 176372 529451
rect 176406 529417 176417 529451
rect 176361 529392 176417 529417
rect 176447 529460 176503 529476
rect 176447 529426 176458 529460
rect 176492 529426 176503 529460
rect 176447 529392 176503 529426
rect 176533 529451 176589 529476
rect 176533 529417 176544 529451
rect 176578 529417 176589 529451
rect 176533 529392 176589 529417
rect 176619 529460 176674 529476
rect 176619 529426 176629 529460
rect 176663 529426 176674 529460
rect 176619 529392 176674 529426
rect 176704 529451 176760 529476
rect 176704 529417 176715 529451
rect 176749 529417 176760 529451
rect 176704 529392 176760 529417
rect 176790 529460 176846 529476
rect 176790 529426 176801 529460
rect 176835 529426 176846 529460
rect 176790 529392 176846 529426
rect 176876 529451 176932 529476
rect 176876 529417 176887 529451
rect 176921 529417 176932 529451
rect 176876 529392 176932 529417
rect 176962 529460 177018 529476
rect 176962 529426 176973 529460
rect 177007 529426 177018 529460
rect 176962 529392 177018 529426
rect 177048 529451 177104 529476
rect 177048 529417 177059 529451
rect 177093 529417 177104 529451
rect 177048 529392 177104 529417
rect 177134 529460 177190 529476
rect 177134 529426 177145 529460
rect 177179 529426 177190 529460
rect 177134 529392 177190 529426
rect 177220 529451 177276 529476
rect 177220 529417 177231 529451
rect 177265 529417 177276 529451
rect 177220 529392 177276 529417
rect 177306 529451 177362 529476
rect 177306 529417 177317 529451
rect 177351 529417 177362 529451
rect 177306 529392 177362 529417
rect 177392 529451 177448 529476
rect 177392 529417 177403 529451
rect 177437 529417 177448 529451
rect 177392 529392 177448 529417
rect 177478 529451 177534 529476
rect 177478 529417 177489 529451
rect 177523 529417 177534 529451
rect 177478 529392 177534 529417
rect 177564 529451 177620 529476
rect 177564 529417 177575 529451
rect 177609 529417 177620 529451
rect 177564 529392 177620 529417
rect 177650 529464 177703 529476
rect 177650 529430 177661 529464
rect 177695 529430 177703 529464
rect 177650 529392 177703 529430
rect 177757 529438 177809 529476
rect 177757 529404 177765 529438
rect 177799 529404 177809 529438
rect 177757 529392 177809 529404
rect 177839 529464 177893 529476
rect 177839 529430 177849 529464
rect 177883 529430 177893 529464
rect 177839 529392 177893 529430
rect 177923 529438 177975 529476
rect 177923 529404 177933 529438
rect 177967 529404 177975 529438
rect 177923 529392 177975 529404
rect 178043 529468 178148 529476
rect 178043 529434 178055 529468
rect 178089 529434 178148 529468
rect 178043 529392 178148 529434
rect 178178 529462 178243 529476
rect 178178 529428 178188 529462
rect 178222 529428 178243 529462
rect 178178 529404 178243 529428
rect 178273 529462 178339 529476
rect 178273 529428 178295 529462
rect 178329 529428 178339 529462
rect 178273 529404 178339 529428
rect 178369 529404 178505 529476
rect 178178 529392 178228 529404
rect 178387 529392 178505 529404
rect 178535 529392 178577 529476
rect 178607 529464 178709 529476
rect 178607 529430 178641 529464
rect 178675 529430 178709 529464
rect 178607 529392 178709 529430
rect 178659 529348 178709 529392
rect 178739 529468 178808 529476
rect 178739 529434 178753 529468
rect 178787 529434 178808 529468
rect 178739 529404 178808 529434
rect 178838 529464 178917 529476
rect 178838 529430 178863 529464
rect 178897 529430 178917 529464
rect 178838 529404 178917 529430
rect 178947 529404 179013 529476
rect 178739 529348 178793 529404
rect 178963 529392 179013 529404
rect 179043 529468 179162 529476
rect 179043 529434 179075 529468
rect 179109 529434 179162 529468
rect 179043 529392 179162 529434
rect 179192 529392 179253 529476
rect 179283 529448 179335 529476
rect 179283 529414 179293 529448
rect 179327 529414 179335 529448
rect 179283 529392 179335 529414
rect 179389 529464 179461 529476
rect 179389 529430 179417 529464
rect 179451 529430 179461 529464
rect 179389 529392 179461 529430
rect 179411 529346 179461 529392
rect 179491 529414 179543 529476
rect 179491 529380 179501 529414
rect 179535 529380 179543 529414
rect 179491 529346 179543 529380
rect 179689 529451 179741 529476
rect 179689 529417 179697 529451
rect 179731 529417 179741 529451
rect 179689 529372 179741 529417
rect 179771 529464 179829 529476
rect 179771 529430 179783 529464
rect 179817 529430 179829 529464
rect 179771 529372 179829 529430
rect 179859 529434 179911 529476
rect 179859 529400 179869 529434
rect 179903 529400 179911 529434
rect 179859 529372 179911 529400
rect 180057 529445 180109 529476
rect 180057 529411 180065 529445
rect 180099 529411 180109 529445
rect 180057 529366 180109 529411
rect 180503 529445 180555 529476
rect 180503 529411 180513 529445
rect 180547 529411 180555 529445
rect 180503 529366 180555 529411
rect 180701 529464 180754 529476
rect 180701 529430 180709 529464
rect 180743 529430 180754 529464
rect 180701 529392 180754 529430
rect 180784 529451 180840 529476
rect 180784 529417 180795 529451
rect 180829 529417 180840 529451
rect 180784 529392 180840 529417
rect 180870 529451 180926 529476
rect 180870 529417 180881 529451
rect 180915 529417 180926 529451
rect 180870 529392 180926 529417
rect 180956 529451 181012 529476
rect 180956 529417 180967 529451
rect 181001 529417 181012 529451
rect 180956 529392 181012 529417
rect 181042 529451 181098 529476
rect 181042 529417 181053 529451
rect 181087 529417 181098 529451
rect 181042 529392 181098 529417
rect 181128 529451 181184 529476
rect 181128 529417 181139 529451
rect 181173 529417 181184 529451
rect 181128 529392 181184 529417
rect 181214 529460 181270 529476
rect 181214 529426 181225 529460
rect 181259 529426 181270 529460
rect 181214 529392 181270 529426
rect 181300 529451 181356 529476
rect 181300 529417 181311 529451
rect 181345 529417 181356 529451
rect 181300 529392 181356 529417
rect 181386 529460 181442 529476
rect 181386 529426 181397 529460
rect 181431 529426 181442 529460
rect 181386 529392 181442 529426
rect 181472 529451 181528 529476
rect 181472 529417 181483 529451
rect 181517 529417 181528 529451
rect 181472 529392 181528 529417
rect 181558 529460 181614 529476
rect 181558 529426 181569 529460
rect 181603 529426 181614 529460
rect 181558 529392 181614 529426
rect 181644 529451 181700 529476
rect 181644 529417 181655 529451
rect 181689 529417 181700 529451
rect 181644 529392 181700 529417
rect 181730 529460 181785 529476
rect 181730 529426 181741 529460
rect 181775 529426 181785 529460
rect 181730 529392 181785 529426
rect 181815 529451 181871 529476
rect 181815 529417 181826 529451
rect 181860 529417 181871 529451
rect 181815 529392 181871 529417
rect 181901 529460 181957 529476
rect 181901 529426 181912 529460
rect 181946 529426 181957 529460
rect 181901 529392 181957 529426
rect 181987 529451 182043 529476
rect 181987 529417 181998 529451
rect 182032 529417 182043 529451
rect 181987 529392 182043 529417
rect 182073 529460 182129 529476
rect 182073 529426 182084 529460
rect 182118 529426 182129 529460
rect 182073 529392 182129 529426
rect 182159 529451 182215 529476
rect 182159 529417 182170 529451
rect 182204 529417 182215 529451
rect 182159 529392 182215 529417
rect 182245 529460 182301 529476
rect 182245 529426 182256 529460
rect 182290 529426 182301 529460
rect 182245 529392 182301 529426
rect 182331 529451 182387 529476
rect 182331 529417 182342 529451
rect 182376 529417 182387 529451
rect 182331 529392 182387 529417
rect 182417 529460 182470 529476
rect 182417 529426 182428 529460
rect 182462 529426 182470 529460
rect 182417 529392 182470 529426
rect 182541 529434 182593 529476
rect 182541 529400 182549 529434
rect 182583 529400 182593 529434
rect 182541 529372 182593 529400
rect 182623 529464 182681 529476
rect 182623 529430 182635 529464
rect 182669 529430 182681 529464
rect 182623 529372 182681 529430
rect 182711 529451 182763 529476
rect 182711 529417 182721 529451
rect 182755 529417 182763 529451
rect 182711 529372 182763 529417
rect 182817 529445 182869 529476
rect 182817 529411 182825 529445
rect 182859 529411 182869 529445
rect 182817 529366 182869 529411
rect 183815 529445 183867 529476
rect 183815 529411 183825 529445
rect 183859 529411 183867 529445
rect 183815 529366 183867 529411
rect 183921 529445 183973 529476
rect 183921 529411 183929 529445
rect 183963 529411 183973 529445
rect 183921 529366 183973 529411
rect 184919 529445 184971 529476
rect 184919 529411 184929 529445
rect 184963 529411 184971 529445
rect 184919 529366 184971 529411
rect 185209 529445 185261 529476
rect 185209 529411 185217 529445
rect 185251 529411 185261 529445
rect 185209 529366 185261 529411
rect 186207 529445 186259 529476
rect 186207 529411 186217 529445
rect 186251 529411 186259 529445
rect 186207 529366 186259 529411
rect 186313 529445 186365 529476
rect 186313 529411 186321 529445
rect 186355 529411 186365 529445
rect 186313 529366 186365 529411
rect 186943 529445 186995 529476
rect 186943 529411 186953 529445
rect 186987 529411 186995 529445
rect 186943 529366 186995 529411
rect 187233 529443 187285 529476
rect 187233 529409 187241 529443
rect 187275 529409 187285 529443
rect 187233 529366 187285 529409
rect 187403 529443 187455 529476
rect 187403 529409 187413 529443
rect 187447 529409 187455 529443
rect 187403 529366 187455 529409
rect 172237 528549 172289 528592
rect 172237 528515 172245 528549
rect 172279 528515 172289 528549
rect 172237 528482 172289 528515
rect 172407 528549 172459 528592
rect 172407 528515 172417 528549
rect 172451 528515 172459 528549
rect 172407 528482 172459 528515
rect 172513 528547 172565 528592
rect 172513 528513 172521 528547
rect 172555 528513 172565 528547
rect 172513 528482 172565 528513
rect 173511 528547 173563 528592
rect 173511 528513 173521 528547
rect 173555 528513 173563 528547
rect 173511 528482 173563 528513
rect 173617 528547 173669 528592
rect 173617 528513 173625 528547
rect 173659 528513 173669 528547
rect 173617 528482 173669 528513
rect 174615 528547 174667 528592
rect 174615 528513 174625 528547
rect 174659 528513 174667 528547
rect 174615 528482 174667 528513
rect 174721 528547 174773 528592
rect 174721 528513 174729 528547
rect 174763 528513 174773 528547
rect 174721 528482 174773 528513
rect 175719 528547 175771 528592
rect 175719 528513 175729 528547
rect 175763 528513 175771 528547
rect 175719 528482 175771 528513
rect 175917 528541 175969 528586
rect 175917 528507 175925 528541
rect 175959 528507 175969 528541
rect 175917 528482 175969 528507
rect 175999 528528 176057 528586
rect 175999 528494 176011 528528
rect 176045 528494 176057 528528
rect 175999 528482 176057 528494
rect 176087 528558 176139 528586
rect 176087 528524 176097 528558
rect 176131 528524 176139 528558
rect 176087 528482 176139 528524
rect 176193 528541 176245 528586
rect 176193 528507 176201 528541
rect 176235 528507 176245 528541
rect 176193 528482 176245 528507
rect 176275 528528 176333 528586
rect 176275 528494 176287 528528
rect 176321 528494 176333 528528
rect 176275 528482 176333 528494
rect 176363 528558 176415 528586
rect 177109 528566 177161 528612
rect 176363 528524 176373 528558
rect 176407 528524 176415 528558
rect 176363 528482 176415 528524
rect 176515 528543 176567 528566
rect 176515 528509 176523 528543
rect 176557 528509 176567 528543
rect 176515 528482 176567 528509
rect 176597 528543 176735 528566
rect 176597 528509 176607 528543
rect 176641 528509 176675 528543
rect 176709 528509 176735 528543
rect 176597 528482 176735 528509
rect 176765 528482 176831 528566
rect 176861 528543 176956 528566
rect 176861 528509 176910 528543
rect 176944 528509 176956 528543
rect 176861 528482 176956 528509
rect 176986 528482 177052 528566
rect 177082 528528 177161 528566
rect 177082 528494 177117 528528
rect 177151 528494 177161 528528
rect 177082 528482 177161 528494
rect 177191 528547 177243 528612
rect 177191 528513 177201 528547
rect 177235 528513 177243 528547
rect 177191 528482 177243 528513
rect 177500 528554 177552 528612
rect 177500 528520 177508 528554
rect 177542 528520 177552 528554
rect 177500 528482 177552 528520
rect 177582 528566 177632 528612
rect 177582 528528 177647 528566
rect 177582 528494 177598 528528
rect 177632 528494 177647 528528
rect 177582 528482 177647 528494
rect 177747 528554 177799 528566
rect 177747 528520 177757 528554
rect 177791 528520 177799 528554
rect 177747 528482 177799 528520
rect 177853 528554 177905 528566
rect 177853 528520 177861 528554
rect 177895 528520 177905 528554
rect 177853 528482 177905 528520
rect 178005 528528 178059 528566
rect 178005 528494 178015 528528
rect 178049 528494 178059 528528
rect 178005 528482 178059 528494
rect 178089 528554 178141 528566
rect 178089 528520 178099 528554
rect 178133 528520 178141 528554
rect 178089 528482 178141 528520
rect 178401 528528 178454 528566
rect 178401 528494 178409 528528
rect 178443 528494 178454 528528
rect 178401 528482 178454 528494
rect 178484 528541 178540 528566
rect 178484 528507 178495 528541
rect 178529 528507 178540 528541
rect 178484 528482 178540 528507
rect 178570 528541 178626 528566
rect 178570 528507 178581 528541
rect 178615 528507 178626 528541
rect 178570 528482 178626 528507
rect 178656 528541 178712 528566
rect 178656 528507 178667 528541
rect 178701 528507 178712 528541
rect 178656 528482 178712 528507
rect 178742 528541 178798 528566
rect 178742 528507 178753 528541
rect 178787 528507 178798 528541
rect 178742 528482 178798 528507
rect 178828 528541 178884 528566
rect 178828 528507 178839 528541
rect 178873 528507 178884 528541
rect 178828 528482 178884 528507
rect 178914 528532 178970 528566
rect 178914 528498 178925 528532
rect 178959 528498 178970 528532
rect 178914 528482 178970 528498
rect 179000 528541 179056 528566
rect 179000 528507 179011 528541
rect 179045 528507 179056 528541
rect 179000 528482 179056 528507
rect 179086 528532 179142 528566
rect 179086 528498 179097 528532
rect 179131 528498 179142 528532
rect 179086 528482 179142 528498
rect 179172 528541 179228 528566
rect 179172 528507 179183 528541
rect 179217 528507 179228 528541
rect 179172 528482 179228 528507
rect 179258 528532 179314 528566
rect 179258 528498 179269 528532
rect 179303 528498 179314 528532
rect 179258 528482 179314 528498
rect 179344 528541 179400 528566
rect 179344 528507 179355 528541
rect 179389 528507 179400 528541
rect 179344 528482 179400 528507
rect 179430 528532 179485 528566
rect 179430 528498 179441 528532
rect 179475 528498 179485 528532
rect 179430 528482 179485 528498
rect 179515 528541 179571 528566
rect 179515 528507 179526 528541
rect 179560 528507 179571 528541
rect 179515 528482 179571 528507
rect 179601 528532 179657 528566
rect 179601 528498 179612 528532
rect 179646 528498 179657 528532
rect 179601 528482 179657 528498
rect 179687 528541 179743 528566
rect 179687 528507 179698 528541
rect 179732 528507 179743 528541
rect 179687 528482 179743 528507
rect 179773 528532 179829 528566
rect 179773 528498 179784 528532
rect 179818 528498 179829 528532
rect 179773 528482 179829 528498
rect 179859 528541 179915 528566
rect 179859 528507 179870 528541
rect 179904 528507 179915 528541
rect 179859 528482 179915 528507
rect 179945 528532 180001 528566
rect 179945 528498 179956 528532
rect 179990 528498 180001 528532
rect 179945 528482 180001 528498
rect 180031 528541 180087 528566
rect 180031 528507 180042 528541
rect 180076 528507 180087 528541
rect 180031 528482 180087 528507
rect 180117 528532 180170 528566
rect 180117 528498 180128 528532
rect 180162 528498 180170 528532
rect 180117 528482 180170 528498
rect 180241 528541 180293 528586
rect 180241 528507 180249 528541
rect 180283 528507 180293 528541
rect 180241 528482 180293 528507
rect 180323 528528 180381 528586
rect 180323 528494 180335 528528
rect 180369 528494 180381 528528
rect 180323 528482 180381 528494
rect 180411 528558 180463 528586
rect 180411 528524 180421 528558
rect 180455 528524 180463 528558
rect 180411 528482 180463 528524
rect 180517 528554 180569 528566
rect 180517 528520 180525 528554
rect 180559 528520 180569 528554
rect 180517 528482 180569 528520
rect 180599 528528 180653 528566
rect 180599 528494 180609 528528
rect 180643 528494 180653 528528
rect 180599 528482 180653 528494
rect 180683 528554 180735 528566
rect 180683 528520 180693 528554
rect 180727 528520 180735 528554
rect 180683 528482 180735 528520
rect 180803 528524 180908 528566
rect 180803 528490 180815 528524
rect 180849 528490 180908 528524
rect 180803 528482 180908 528490
rect 180938 528554 180988 528566
rect 181419 528566 181469 528610
rect 181147 528554 181265 528566
rect 180938 528530 181003 528554
rect 180938 528496 180948 528530
rect 180982 528496 181003 528530
rect 180938 528482 181003 528496
rect 181033 528530 181099 528554
rect 181033 528496 181055 528530
rect 181089 528496 181099 528530
rect 181033 528482 181099 528496
rect 181129 528482 181265 528554
rect 181295 528482 181337 528566
rect 181367 528528 181469 528566
rect 181367 528494 181401 528528
rect 181435 528494 181469 528528
rect 181367 528482 181469 528494
rect 181499 528554 181553 528610
rect 182171 528566 182221 528612
rect 181723 528554 181773 528566
rect 181499 528524 181568 528554
rect 181499 528490 181513 528524
rect 181547 528490 181568 528524
rect 181499 528482 181568 528490
rect 181598 528528 181677 528554
rect 181598 528494 181623 528528
rect 181657 528494 181677 528528
rect 181598 528482 181677 528494
rect 181707 528482 181773 528554
rect 181803 528524 181922 528566
rect 181803 528490 181835 528524
rect 181869 528490 181922 528524
rect 181803 528482 181922 528490
rect 181952 528482 182013 528566
rect 182043 528544 182095 528566
rect 182043 528510 182053 528544
rect 182087 528510 182095 528544
rect 182043 528482 182095 528510
rect 182149 528528 182221 528566
rect 182149 528494 182177 528528
rect 182211 528494 182221 528528
rect 182149 528482 182221 528494
rect 182251 528578 182303 528612
rect 182251 528544 182261 528578
rect 182295 528544 182303 528578
rect 182251 528482 182303 528544
rect 182633 528547 182685 528592
rect 182633 528513 182641 528547
rect 182675 528513 182685 528547
rect 182633 528482 182685 528513
rect 183631 528547 183683 528592
rect 183631 528513 183641 528547
rect 183675 528513 183683 528547
rect 183631 528482 183683 528513
rect 183737 528547 183789 528592
rect 183737 528513 183745 528547
rect 183779 528513 183789 528547
rect 183737 528482 183789 528513
rect 184735 528547 184787 528592
rect 184735 528513 184745 528547
rect 184779 528513 184787 528547
rect 184735 528482 184787 528513
rect 184841 528547 184893 528592
rect 184841 528513 184849 528547
rect 184883 528513 184893 528547
rect 184841 528482 184893 528513
rect 185839 528547 185891 528592
rect 185839 528513 185849 528547
rect 185883 528513 185891 528547
rect 185839 528482 185891 528513
rect 185945 528547 185997 528592
rect 185945 528513 185953 528547
rect 185987 528513 185997 528547
rect 185945 528482 185997 528513
rect 186943 528547 186995 528592
rect 186943 528513 186953 528547
rect 186987 528513 186995 528547
rect 186943 528482 186995 528513
rect 187233 528549 187285 528592
rect 187233 528515 187241 528549
rect 187275 528515 187285 528549
rect 187233 528482 187285 528515
rect 187403 528549 187455 528592
rect 187403 528515 187413 528549
rect 187447 528515 187455 528549
rect 187403 528482 187455 528515
rect 172237 528355 172289 528388
rect 172237 528321 172245 528355
rect 172279 528321 172289 528355
rect 172237 528278 172289 528321
rect 172407 528355 172459 528388
rect 172407 528321 172417 528355
rect 172451 528321 172459 528355
rect 172407 528278 172459 528321
rect 172513 528357 172565 528388
rect 172513 528323 172521 528357
rect 172555 528323 172565 528357
rect 172513 528278 172565 528323
rect 173511 528357 173563 528388
rect 173511 528323 173521 528357
rect 173555 528323 173563 528357
rect 173511 528278 173563 528323
rect 173617 528357 173669 528388
rect 173617 528323 173625 528357
rect 173659 528323 173669 528357
rect 173617 528278 173669 528323
rect 174615 528357 174667 528388
rect 174615 528323 174625 528357
rect 174659 528323 174667 528357
rect 174615 528278 174667 528323
rect 174905 528357 174957 528388
rect 174905 528323 174913 528357
rect 174947 528323 174957 528357
rect 174905 528278 174957 528323
rect 175903 528357 175955 528388
rect 175903 528323 175913 528357
rect 175947 528323 175955 528357
rect 175903 528278 175955 528323
rect 176101 528350 176153 528388
rect 176101 528316 176109 528350
rect 176143 528316 176153 528350
rect 176101 528304 176153 528316
rect 176183 528376 176237 528388
rect 176183 528342 176193 528376
rect 176227 528342 176237 528376
rect 176183 528304 176237 528342
rect 176267 528350 176319 528388
rect 176267 528316 176277 528350
rect 176311 528316 176319 528350
rect 176267 528304 176319 528316
rect 176387 528380 176492 528388
rect 176387 528346 176399 528380
rect 176433 528346 176492 528380
rect 176387 528304 176492 528346
rect 176522 528374 176587 528388
rect 176522 528340 176532 528374
rect 176566 528340 176587 528374
rect 176522 528316 176587 528340
rect 176617 528374 176683 528388
rect 176617 528340 176639 528374
rect 176673 528340 176683 528374
rect 176617 528316 176683 528340
rect 176713 528316 176849 528388
rect 176522 528304 176572 528316
rect 176731 528304 176849 528316
rect 176879 528304 176921 528388
rect 176951 528376 177053 528388
rect 176951 528342 176985 528376
rect 177019 528342 177053 528376
rect 176951 528304 177053 528342
rect 177003 528260 177053 528304
rect 177083 528380 177152 528388
rect 177083 528346 177097 528380
rect 177131 528346 177152 528380
rect 177083 528316 177152 528346
rect 177182 528376 177261 528388
rect 177182 528342 177207 528376
rect 177241 528342 177261 528376
rect 177182 528316 177261 528342
rect 177291 528316 177357 528388
rect 177083 528260 177137 528316
rect 177307 528304 177357 528316
rect 177387 528380 177506 528388
rect 177387 528346 177419 528380
rect 177453 528346 177506 528380
rect 177387 528304 177506 528346
rect 177536 528304 177597 528388
rect 177627 528360 177679 528388
rect 177627 528326 177637 528360
rect 177671 528326 177679 528360
rect 177627 528304 177679 528326
rect 177733 528376 177805 528388
rect 177733 528342 177761 528376
rect 177795 528342 177805 528376
rect 177733 528304 177805 528342
rect 177755 528258 177805 528304
rect 177835 528326 177887 528388
rect 177835 528292 177845 528326
rect 177879 528292 177887 528326
rect 177835 528258 177887 528292
rect 177941 528346 177993 528388
rect 177941 528312 177949 528346
rect 177983 528312 177993 528346
rect 177941 528284 177993 528312
rect 178023 528376 178081 528388
rect 178023 528342 178035 528376
rect 178069 528342 178081 528376
rect 178023 528284 178081 528342
rect 178111 528363 178163 528388
rect 178111 528329 178121 528363
rect 178155 528329 178163 528363
rect 178111 528284 178163 528329
rect 178217 528357 178269 528388
rect 178217 528323 178225 528357
rect 178259 528323 178269 528357
rect 178217 528278 178269 528323
rect 178847 528357 178899 528388
rect 178847 528323 178857 528357
rect 178891 528323 178899 528357
rect 178847 528278 178899 528323
rect 178953 528357 179005 528388
rect 178953 528323 178961 528357
rect 178995 528323 179005 528357
rect 178953 528258 179005 528323
rect 179035 528376 179114 528388
rect 179035 528342 179045 528376
rect 179079 528342 179114 528376
rect 179035 528304 179114 528342
rect 179144 528304 179210 528388
rect 179240 528361 179335 528388
rect 179240 528327 179252 528361
rect 179286 528327 179335 528361
rect 179240 528304 179335 528327
rect 179365 528304 179431 528388
rect 179461 528361 179599 528388
rect 179461 528327 179487 528361
rect 179521 528327 179555 528361
rect 179589 528327 179599 528361
rect 179461 528304 179599 528327
rect 179629 528361 179681 528388
rect 179629 528327 179639 528361
rect 179673 528327 179681 528361
rect 179629 528304 179681 528327
rect 179035 528258 179087 528304
rect 180057 528357 180109 528388
rect 180057 528323 180065 528357
rect 180099 528323 180109 528357
rect 180057 528278 180109 528323
rect 180687 528357 180739 528388
rect 180687 528323 180697 528357
rect 180731 528323 180739 528357
rect 180687 528278 180739 528323
rect 180977 528357 181029 528388
rect 180977 528323 180985 528357
rect 181019 528323 181029 528357
rect 180977 528258 181029 528323
rect 181059 528376 181138 528388
rect 181059 528342 181069 528376
rect 181103 528342 181138 528376
rect 181059 528304 181138 528342
rect 181168 528304 181234 528388
rect 181264 528361 181359 528388
rect 181264 528327 181276 528361
rect 181310 528327 181359 528361
rect 181264 528304 181359 528327
rect 181389 528304 181455 528388
rect 181485 528361 181623 528388
rect 181485 528327 181511 528361
rect 181545 528327 181579 528361
rect 181613 528327 181623 528361
rect 181485 528304 181623 528327
rect 181653 528361 181705 528388
rect 181653 528327 181663 528361
rect 181697 528327 181705 528361
rect 181653 528304 181705 528327
rect 181805 528357 181857 528388
rect 181805 528323 181813 528357
rect 181847 528323 181857 528357
rect 181059 528258 181111 528304
rect 181805 528278 181857 528323
rect 182803 528357 182855 528388
rect 182803 528323 182813 528357
rect 182847 528323 182855 528357
rect 182803 528278 182855 528323
rect 182909 528357 182961 528388
rect 182909 528323 182917 528357
rect 182951 528323 182961 528357
rect 182909 528278 182961 528323
rect 183907 528357 183959 528388
rect 183907 528323 183917 528357
rect 183951 528323 183959 528357
rect 183907 528278 183959 528323
rect 184013 528357 184065 528388
rect 184013 528323 184021 528357
rect 184055 528323 184065 528357
rect 184013 528278 184065 528323
rect 185011 528357 185063 528388
rect 185011 528323 185021 528357
rect 185055 528323 185063 528357
rect 185011 528278 185063 528323
rect 185209 528357 185261 528388
rect 185209 528323 185217 528357
rect 185251 528323 185261 528357
rect 185209 528278 185261 528323
rect 186207 528357 186259 528388
rect 186207 528323 186217 528357
rect 186251 528323 186259 528357
rect 186207 528278 186259 528323
rect 186313 528357 186365 528388
rect 186313 528323 186321 528357
rect 186355 528323 186365 528357
rect 186313 528278 186365 528323
rect 186943 528357 186995 528388
rect 186943 528323 186953 528357
rect 186987 528323 186995 528357
rect 186943 528278 186995 528323
rect 187233 528355 187285 528388
rect 187233 528321 187241 528355
rect 187275 528321 187285 528355
rect 187233 528278 187285 528321
rect 187403 528355 187455 528388
rect 187403 528321 187413 528355
rect 187447 528321 187455 528355
rect 187403 528278 187455 528321
rect 172237 527461 172289 527504
rect 172237 527427 172245 527461
rect 172279 527427 172289 527461
rect 172237 527394 172289 527427
rect 172407 527461 172459 527504
rect 172407 527427 172417 527461
rect 172451 527427 172459 527461
rect 172407 527394 172459 527427
rect 172513 527459 172565 527504
rect 172513 527425 172521 527459
rect 172555 527425 172565 527459
rect 172513 527394 172565 527425
rect 173511 527459 173563 527504
rect 173511 527425 173521 527459
rect 173555 527425 173563 527459
rect 173511 527394 173563 527425
rect 173617 527459 173669 527504
rect 173617 527425 173625 527459
rect 173659 527425 173669 527459
rect 173617 527394 173669 527425
rect 174615 527459 174667 527504
rect 174615 527425 174625 527459
rect 174659 527425 174667 527459
rect 174615 527394 174667 527425
rect 174721 527459 174773 527504
rect 174721 527425 174729 527459
rect 174763 527425 174773 527459
rect 174721 527394 174773 527425
rect 175719 527459 175771 527504
rect 175719 527425 175729 527459
rect 175763 527425 175771 527459
rect 175719 527394 175771 527425
rect 175825 527459 175877 527504
rect 175825 527425 175833 527459
rect 175867 527425 175877 527459
rect 175825 527394 175877 527425
rect 176271 527459 176323 527504
rect 176271 527425 176281 527459
rect 176315 527425 176323 527459
rect 176271 527394 176323 527425
rect 176396 527466 176448 527524
rect 176396 527432 176404 527466
rect 176438 527432 176448 527466
rect 176396 527394 176448 527432
rect 176478 527478 176528 527524
rect 176478 527440 176543 527478
rect 176478 527406 176494 527440
rect 176528 527406 176543 527440
rect 176478 527394 176543 527406
rect 176643 527466 176695 527478
rect 176643 527432 176653 527466
rect 176687 527432 176695 527466
rect 176643 527394 176695 527432
rect 176749 527466 176801 527478
rect 176749 527432 176757 527466
rect 176791 527432 176801 527466
rect 176749 527394 176801 527432
rect 176901 527440 176955 527478
rect 176901 527406 176911 527440
rect 176945 527406 176955 527440
rect 176901 527394 176955 527406
rect 176985 527466 177037 527478
rect 176985 527432 176995 527466
rect 177029 527432 177037 527466
rect 176985 527394 177037 527432
rect 177113 527461 177165 527504
rect 177113 527427 177121 527461
rect 177155 527427 177165 527461
rect 177113 527394 177165 527427
rect 177283 527461 177335 527504
rect 177283 527427 177293 527461
rect 177327 527427 177335 527461
rect 177283 527394 177335 527427
rect 177481 527459 177533 527504
rect 177481 527425 177489 527459
rect 177523 527425 177533 527459
rect 177481 527394 177533 527425
rect 178479 527459 178531 527504
rect 178479 527425 178489 527459
rect 178523 527425 178531 527459
rect 178479 527394 178531 527425
rect 178585 527466 178637 527504
rect 178585 527432 178593 527466
rect 178627 527432 178637 527466
rect 178585 527394 178637 527432
rect 178847 527466 178899 527504
rect 178847 527432 178857 527466
rect 178891 527432 178899 527466
rect 178847 527394 178899 527432
rect 178972 527466 179024 527524
rect 178972 527432 178980 527466
rect 179014 527432 179024 527466
rect 178972 527394 179024 527432
rect 179054 527478 179104 527524
rect 179054 527440 179119 527478
rect 179054 527406 179070 527440
rect 179104 527406 179119 527440
rect 179054 527394 179119 527406
rect 179219 527466 179271 527478
rect 179219 527432 179229 527466
rect 179263 527432 179271 527466
rect 179219 527394 179271 527432
rect 179325 527466 179377 527478
rect 179325 527432 179333 527466
rect 179367 527432 179377 527466
rect 179325 527394 179377 527432
rect 179477 527440 179531 527478
rect 179477 527406 179487 527440
rect 179521 527406 179531 527440
rect 179477 527394 179531 527406
rect 179561 527466 179613 527478
rect 179561 527432 179571 527466
rect 179605 527432 179613 527466
rect 179561 527394 179613 527432
rect 179689 527459 179741 527504
rect 179689 527425 179697 527459
rect 179731 527425 179741 527459
rect 179689 527394 179741 527425
rect 180687 527459 180739 527504
rect 180687 527425 180697 527459
rect 180731 527425 180739 527459
rect 180687 527394 180739 527425
rect 180793 527459 180845 527504
rect 180793 527425 180801 527459
rect 180835 527425 180845 527459
rect 180793 527394 180845 527425
rect 181791 527459 181843 527504
rect 181791 527425 181801 527459
rect 181835 527425 181843 527459
rect 181791 527394 181843 527425
rect 181897 527459 181949 527504
rect 181897 527425 181905 527459
rect 181939 527425 181949 527459
rect 181897 527394 181949 527425
rect 182343 527459 182395 527504
rect 182343 527425 182353 527459
rect 182387 527425 182395 527459
rect 182343 527394 182395 527425
rect 182633 527459 182685 527504
rect 182633 527425 182641 527459
rect 182675 527425 182685 527459
rect 182633 527394 182685 527425
rect 183631 527459 183683 527504
rect 183631 527425 183641 527459
rect 183675 527425 183683 527459
rect 183631 527394 183683 527425
rect 183737 527459 183789 527504
rect 183737 527425 183745 527459
rect 183779 527425 183789 527459
rect 183737 527394 183789 527425
rect 184735 527459 184787 527504
rect 184735 527425 184745 527459
rect 184779 527425 184787 527459
rect 184735 527394 184787 527425
rect 184841 527459 184893 527504
rect 184841 527425 184849 527459
rect 184883 527425 184893 527459
rect 184841 527394 184893 527425
rect 185839 527459 185891 527504
rect 185839 527425 185849 527459
rect 185883 527425 185891 527459
rect 185839 527394 185891 527425
rect 185945 527459 185997 527504
rect 185945 527425 185953 527459
rect 185987 527425 185997 527459
rect 185945 527394 185997 527425
rect 186943 527459 186995 527504
rect 186943 527425 186953 527459
rect 186987 527425 186995 527459
rect 186943 527394 186995 527425
rect 187233 527461 187285 527504
rect 187233 527427 187241 527461
rect 187275 527427 187285 527461
rect 187233 527394 187285 527427
rect 187403 527461 187455 527504
rect 187403 527427 187413 527461
rect 187447 527427 187455 527461
rect 187403 527394 187455 527427
rect 172237 527267 172289 527300
rect 172237 527233 172245 527267
rect 172279 527233 172289 527267
rect 172237 527190 172289 527233
rect 172407 527267 172459 527300
rect 172407 527233 172417 527267
rect 172451 527233 172459 527267
rect 172407 527190 172459 527233
rect 172513 527269 172565 527300
rect 172513 527235 172521 527269
rect 172555 527235 172565 527269
rect 172513 527190 172565 527235
rect 173511 527269 173563 527300
rect 173511 527235 173521 527269
rect 173555 527235 173563 527269
rect 173511 527190 173563 527235
rect 173617 527269 173669 527300
rect 173617 527235 173625 527269
rect 173659 527235 173669 527269
rect 173617 527190 173669 527235
rect 174615 527269 174667 527300
rect 174615 527235 174625 527269
rect 174659 527235 174667 527269
rect 174615 527190 174667 527235
rect 174905 527269 174957 527300
rect 174905 527235 174913 527269
rect 174947 527235 174957 527269
rect 174905 527190 174957 527235
rect 175903 527269 175955 527300
rect 175903 527235 175913 527269
rect 175947 527235 175955 527269
rect 175903 527190 175955 527235
rect 176009 527269 176061 527300
rect 176009 527235 176017 527269
rect 176051 527235 176061 527269
rect 176009 527190 176061 527235
rect 177007 527269 177059 527300
rect 177007 527235 177017 527269
rect 177051 527235 177059 527269
rect 177007 527190 177059 527235
rect 177113 527269 177165 527300
rect 177113 527235 177121 527269
rect 177155 527235 177165 527269
rect 177113 527190 177165 527235
rect 178111 527269 178163 527300
rect 178111 527235 178121 527269
rect 178155 527235 178163 527269
rect 178111 527190 178163 527235
rect 178217 527269 178269 527300
rect 178217 527235 178225 527269
rect 178259 527235 178269 527269
rect 178217 527190 178269 527235
rect 179215 527269 179267 527300
rect 179215 527235 179225 527269
rect 179259 527235 179267 527269
rect 179215 527190 179267 527235
rect 179321 527269 179373 527300
rect 179321 527235 179329 527269
rect 179363 527235 179373 527269
rect 179321 527190 179373 527235
rect 179767 527269 179819 527300
rect 179767 527235 179777 527269
rect 179811 527235 179819 527269
rect 179767 527190 179819 527235
rect 180057 527269 180109 527300
rect 180057 527235 180065 527269
rect 180099 527235 180109 527269
rect 180057 527190 180109 527235
rect 181055 527269 181107 527300
rect 181055 527235 181065 527269
rect 181099 527235 181107 527269
rect 181055 527190 181107 527235
rect 181161 527269 181213 527300
rect 181161 527235 181169 527269
rect 181203 527235 181213 527269
rect 181161 527190 181213 527235
rect 182159 527269 182211 527300
rect 182159 527235 182169 527269
rect 182203 527235 182211 527269
rect 182159 527190 182211 527235
rect 182265 527269 182317 527300
rect 182265 527235 182273 527269
rect 182307 527235 182317 527269
rect 182265 527190 182317 527235
rect 183263 527269 183315 527300
rect 183263 527235 183273 527269
rect 183307 527235 183315 527269
rect 183263 527190 183315 527235
rect 183369 527269 183421 527300
rect 183369 527235 183377 527269
rect 183411 527235 183421 527269
rect 183369 527190 183421 527235
rect 184367 527269 184419 527300
rect 184367 527235 184377 527269
rect 184411 527235 184419 527269
rect 184367 527190 184419 527235
rect 184473 527269 184525 527300
rect 184473 527235 184481 527269
rect 184515 527235 184525 527269
rect 184473 527190 184525 527235
rect 184919 527269 184971 527300
rect 184919 527235 184929 527269
rect 184963 527235 184971 527269
rect 184919 527190 184971 527235
rect 185209 527269 185261 527300
rect 185209 527235 185217 527269
rect 185251 527235 185261 527269
rect 185209 527190 185261 527235
rect 186207 527269 186259 527300
rect 186207 527235 186217 527269
rect 186251 527235 186259 527269
rect 186207 527190 186259 527235
rect 186313 527269 186365 527300
rect 186313 527235 186321 527269
rect 186355 527235 186365 527269
rect 186313 527190 186365 527235
rect 186943 527269 186995 527300
rect 186943 527235 186953 527269
rect 186987 527235 186995 527269
rect 186943 527190 186995 527235
rect 187233 527267 187285 527300
rect 187233 527233 187241 527267
rect 187275 527233 187285 527267
rect 187233 527190 187285 527233
rect 187403 527267 187455 527300
rect 187403 527233 187413 527267
rect 187447 527233 187455 527267
rect 187403 527190 187455 527233
rect 172237 526373 172289 526416
rect 172237 526339 172245 526373
rect 172279 526339 172289 526373
rect 172237 526306 172289 526339
rect 172407 526373 172459 526416
rect 172407 526339 172417 526373
rect 172451 526339 172459 526373
rect 172407 526306 172459 526339
rect 172513 526371 172565 526416
rect 172513 526337 172521 526371
rect 172555 526337 172565 526371
rect 172513 526306 172565 526337
rect 173511 526371 173563 526416
rect 173511 526337 173521 526371
rect 173555 526337 173563 526371
rect 173511 526306 173563 526337
rect 173617 526371 173669 526416
rect 173617 526337 173625 526371
rect 173659 526337 173669 526371
rect 173617 526306 173669 526337
rect 174615 526371 174667 526416
rect 174615 526337 174625 526371
rect 174659 526337 174667 526371
rect 174615 526306 174667 526337
rect 174721 526371 174773 526416
rect 174721 526337 174729 526371
rect 174763 526337 174773 526371
rect 174721 526306 174773 526337
rect 175719 526371 175771 526416
rect 175719 526337 175729 526371
rect 175763 526337 175771 526371
rect 175719 526306 175771 526337
rect 175825 526371 175877 526416
rect 175825 526337 175833 526371
rect 175867 526337 175877 526371
rect 175825 526306 175877 526337
rect 176823 526371 176875 526416
rect 176823 526337 176833 526371
rect 176867 526337 176875 526371
rect 176823 526306 176875 526337
rect 176929 526378 176981 526416
rect 176929 526344 176937 526378
rect 176971 526344 176981 526378
rect 176929 526306 176981 526344
rect 177191 526378 177243 526416
rect 177191 526344 177201 526378
rect 177235 526344 177243 526378
rect 177191 526306 177243 526344
rect 177481 526371 177533 526416
rect 177481 526337 177489 526371
rect 177523 526337 177533 526371
rect 177481 526306 177533 526337
rect 178479 526371 178531 526416
rect 178479 526337 178489 526371
rect 178523 526337 178531 526371
rect 178479 526306 178531 526337
rect 178585 526371 178637 526416
rect 178585 526337 178593 526371
rect 178627 526337 178637 526371
rect 178585 526306 178637 526337
rect 179583 526371 179635 526416
rect 179583 526337 179593 526371
rect 179627 526337 179635 526371
rect 179583 526306 179635 526337
rect 179689 526371 179741 526416
rect 179689 526337 179697 526371
rect 179731 526337 179741 526371
rect 179689 526306 179741 526337
rect 180687 526371 180739 526416
rect 180687 526337 180697 526371
rect 180731 526337 180739 526371
rect 180687 526306 180739 526337
rect 180793 526371 180845 526416
rect 180793 526337 180801 526371
rect 180835 526337 180845 526371
rect 180793 526306 180845 526337
rect 181791 526371 181843 526416
rect 181791 526337 181801 526371
rect 181835 526337 181843 526371
rect 181791 526306 181843 526337
rect 181897 526371 181949 526416
rect 181897 526337 181905 526371
rect 181939 526337 181949 526371
rect 181897 526306 181949 526337
rect 182343 526371 182395 526416
rect 182343 526337 182353 526371
rect 182387 526337 182395 526371
rect 182343 526306 182395 526337
rect 182633 526371 182685 526416
rect 182633 526337 182641 526371
rect 182675 526337 182685 526371
rect 182633 526306 182685 526337
rect 183631 526371 183683 526416
rect 183631 526337 183641 526371
rect 183675 526337 183683 526371
rect 183631 526306 183683 526337
rect 183737 526371 183789 526416
rect 183737 526337 183745 526371
rect 183779 526337 183789 526371
rect 183737 526306 183789 526337
rect 184735 526371 184787 526416
rect 184735 526337 184745 526371
rect 184779 526337 184787 526371
rect 184735 526306 184787 526337
rect 184841 526371 184893 526416
rect 184841 526337 184849 526371
rect 184883 526337 184893 526371
rect 184841 526306 184893 526337
rect 185839 526371 185891 526416
rect 185839 526337 185849 526371
rect 185883 526337 185891 526371
rect 185839 526306 185891 526337
rect 185945 526371 185997 526416
rect 185945 526337 185953 526371
rect 185987 526337 185997 526371
rect 185945 526306 185997 526337
rect 186943 526371 186995 526416
rect 186943 526337 186953 526371
rect 186987 526337 186995 526371
rect 186943 526306 186995 526337
rect 187233 526373 187285 526416
rect 187233 526339 187241 526373
rect 187275 526339 187285 526373
rect 187233 526306 187285 526339
rect 187403 526373 187455 526416
rect 187403 526339 187413 526373
rect 187447 526339 187455 526373
rect 187403 526306 187455 526339
rect 172237 526179 172289 526212
rect 172237 526145 172245 526179
rect 172279 526145 172289 526179
rect 172237 526102 172289 526145
rect 172407 526179 172459 526212
rect 172407 526145 172417 526179
rect 172451 526145 172459 526179
rect 172407 526102 172459 526145
rect 172513 526181 172565 526212
rect 172513 526147 172521 526181
rect 172555 526147 172565 526181
rect 172513 526102 172565 526147
rect 173511 526181 173563 526212
rect 173511 526147 173521 526181
rect 173555 526147 173563 526181
rect 173511 526102 173563 526147
rect 173617 526181 173669 526212
rect 173617 526147 173625 526181
rect 173659 526147 173669 526181
rect 173617 526102 173669 526147
rect 174615 526181 174667 526212
rect 174615 526147 174625 526181
rect 174659 526147 174667 526181
rect 174615 526102 174667 526147
rect 174905 526181 174957 526212
rect 174905 526147 174913 526181
rect 174947 526147 174957 526181
rect 174905 526102 174957 526147
rect 175903 526181 175955 526212
rect 175903 526147 175913 526181
rect 175947 526147 175955 526181
rect 175903 526102 175955 526147
rect 176009 526181 176061 526212
rect 176009 526147 176017 526181
rect 176051 526147 176061 526181
rect 176009 526102 176061 526147
rect 177007 526181 177059 526212
rect 177007 526147 177017 526181
rect 177051 526147 177059 526181
rect 177007 526102 177059 526147
rect 177113 526181 177165 526212
rect 177113 526147 177121 526181
rect 177155 526147 177165 526181
rect 177113 526102 177165 526147
rect 178111 526181 178163 526212
rect 178111 526147 178121 526181
rect 178155 526147 178163 526181
rect 178111 526102 178163 526147
rect 178217 526181 178269 526212
rect 178217 526147 178225 526181
rect 178259 526147 178269 526181
rect 178217 526102 178269 526147
rect 179215 526181 179267 526212
rect 179215 526147 179225 526181
rect 179259 526147 179267 526181
rect 179215 526102 179267 526147
rect 179321 526181 179373 526212
rect 179321 526147 179329 526181
rect 179363 526147 179373 526181
rect 179321 526102 179373 526147
rect 179767 526181 179819 526212
rect 179767 526147 179777 526181
rect 179811 526147 179819 526181
rect 179767 526102 179819 526147
rect 180057 526181 180109 526212
rect 180057 526147 180065 526181
rect 180099 526147 180109 526181
rect 180057 526102 180109 526147
rect 181055 526181 181107 526212
rect 181055 526147 181065 526181
rect 181099 526147 181107 526181
rect 181055 526102 181107 526147
rect 181161 526181 181213 526212
rect 181161 526147 181169 526181
rect 181203 526147 181213 526181
rect 181161 526102 181213 526147
rect 182159 526181 182211 526212
rect 182159 526147 182169 526181
rect 182203 526147 182211 526181
rect 182159 526102 182211 526147
rect 182265 526181 182317 526212
rect 182265 526147 182273 526181
rect 182307 526147 182317 526181
rect 182265 526102 182317 526147
rect 183263 526181 183315 526212
rect 183263 526147 183273 526181
rect 183307 526147 183315 526181
rect 183263 526102 183315 526147
rect 183369 526181 183421 526212
rect 183369 526147 183377 526181
rect 183411 526147 183421 526181
rect 183369 526102 183421 526147
rect 184367 526181 184419 526212
rect 184367 526147 184377 526181
rect 184411 526147 184419 526181
rect 184367 526102 184419 526147
rect 184473 526181 184525 526212
rect 184473 526147 184481 526181
rect 184515 526147 184525 526181
rect 184473 526102 184525 526147
rect 184919 526181 184971 526212
rect 184919 526147 184929 526181
rect 184963 526147 184971 526181
rect 184919 526102 184971 526147
rect 185209 526181 185261 526212
rect 185209 526147 185217 526181
rect 185251 526147 185261 526181
rect 185209 526102 185261 526147
rect 186207 526181 186259 526212
rect 186207 526147 186217 526181
rect 186251 526147 186259 526181
rect 186207 526102 186259 526147
rect 186313 526181 186365 526212
rect 186313 526147 186321 526181
rect 186355 526147 186365 526181
rect 186313 526102 186365 526147
rect 186943 526181 186995 526212
rect 186943 526147 186953 526181
rect 186987 526147 186995 526181
rect 186943 526102 186995 526147
rect 187233 526179 187285 526212
rect 187233 526145 187241 526179
rect 187275 526145 187285 526179
rect 187233 526102 187285 526145
rect 187403 526179 187455 526212
rect 187403 526145 187413 526179
rect 187447 526145 187455 526179
rect 187403 526102 187455 526145
rect 172237 525285 172289 525328
rect 172237 525251 172245 525285
rect 172279 525251 172289 525285
rect 172237 525218 172289 525251
rect 172407 525285 172459 525328
rect 172407 525251 172417 525285
rect 172451 525251 172459 525285
rect 172407 525218 172459 525251
rect 172513 525283 172565 525328
rect 172513 525249 172521 525283
rect 172555 525249 172565 525283
rect 172513 525218 172565 525249
rect 173511 525283 173563 525328
rect 173511 525249 173521 525283
rect 173555 525249 173563 525283
rect 173511 525218 173563 525249
rect 173617 525283 173669 525328
rect 173617 525249 173625 525283
rect 173659 525249 173669 525283
rect 173617 525218 173669 525249
rect 174615 525283 174667 525328
rect 174615 525249 174625 525283
rect 174659 525249 174667 525283
rect 174615 525218 174667 525249
rect 174721 525283 174773 525328
rect 174721 525249 174729 525283
rect 174763 525249 174773 525283
rect 174721 525218 174773 525249
rect 175719 525283 175771 525328
rect 175719 525249 175729 525283
rect 175763 525249 175771 525283
rect 175719 525218 175771 525249
rect 175825 525283 175877 525328
rect 175825 525249 175833 525283
rect 175867 525249 175877 525283
rect 175825 525218 175877 525249
rect 176823 525283 176875 525328
rect 176823 525249 176833 525283
rect 176867 525249 176875 525283
rect 176823 525218 176875 525249
rect 176929 525290 176981 525328
rect 176929 525256 176937 525290
rect 176971 525256 176981 525290
rect 176929 525218 176981 525256
rect 177191 525290 177243 525328
rect 177191 525256 177201 525290
rect 177235 525256 177243 525290
rect 177191 525218 177243 525256
rect 177481 525283 177533 525328
rect 177481 525249 177489 525283
rect 177523 525249 177533 525283
rect 177481 525218 177533 525249
rect 178479 525283 178531 525328
rect 178479 525249 178489 525283
rect 178523 525249 178531 525283
rect 178479 525218 178531 525249
rect 178585 525283 178637 525328
rect 178585 525249 178593 525283
rect 178627 525249 178637 525283
rect 178585 525218 178637 525249
rect 179583 525283 179635 525328
rect 179583 525249 179593 525283
rect 179627 525249 179635 525283
rect 179583 525218 179635 525249
rect 179689 525283 179741 525328
rect 179689 525249 179697 525283
rect 179731 525249 179741 525283
rect 179689 525218 179741 525249
rect 180687 525283 180739 525328
rect 180687 525249 180697 525283
rect 180731 525249 180739 525283
rect 180687 525218 180739 525249
rect 180793 525283 180845 525328
rect 180793 525249 180801 525283
rect 180835 525249 180845 525283
rect 180793 525218 180845 525249
rect 181791 525283 181843 525328
rect 181791 525249 181801 525283
rect 181835 525249 181843 525283
rect 181791 525218 181843 525249
rect 181897 525283 181949 525328
rect 181897 525249 181905 525283
rect 181939 525249 181949 525283
rect 181897 525218 181949 525249
rect 182343 525283 182395 525328
rect 182343 525249 182353 525283
rect 182387 525249 182395 525283
rect 182343 525218 182395 525249
rect 182633 525283 182685 525328
rect 182633 525249 182641 525283
rect 182675 525249 182685 525283
rect 182633 525218 182685 525249
rect 183631 525283 183683 525328
rect 183631 525249 183641 525283
rect 183675 525249 183683 525283
rect 183631 525218 183683 525249
rect 183737 525283 183789 525328
rect 183737 525249 183745 525283
rect 183779 525249 183789 525283
rect 183737 525218 183789 525249
rect 184735 525283 184787 525328
rect 184735 525249 184745 525283
rect 184779 525249 184787 525283
rect 184735 525218 184787 525249
rect 184841 525283 184893 525328
rect 184841 525249 184849 525283
rect 184883 525249 184893 525283
rect 184841 525218 184893 525249
rect 185839 525283 185891 525328
rect 185839 525249 185849 525283
rect 185883 525249 185891 525283
rect 185839 525218 185891 525249
rect 185945 525283 185997 525328
rect 185945 525249 185953 525283
rect 185987 525249 185997 525283
rect 185945 525218 185997 525249
rect 186943 525283 186995 525328
rect 186943 525249 186953 525283
rect 186987 525249 186995 525283
rect 186943 525218 186995 525249
rect 187233 525285 187285 525328
rect 187233 525251 187241 525285
rect 187275 525251 187285 525285
rect 187233 525218 187285 525251
rect 187403 525285 187455 525328
rect 187403 525251 187413 525285
rect 187447 525251 187455 525285
rect 187403 525218 187455 525251
rect 172237 525091 172289 525124
rect 172237 525057 172245 525091
rect 172279 525057 172289 525091
rect 172237 525014 172289 525057
rect 172407 525091 172459 525124
rect 172407 525057 172417 525091
rect 172451 525057 172459 525091
rect 172407 525014 172459 525057
rect 172513 525093 172565 525124
rect 172513 525059 172521 525093
rect 172555 525059 172565 525093
rect 172513 525014 172565 525059
rect 173511 525093 173563 525124
rect 173511 525059 173521 525093
rect 173555 525059 173563 525093
rect 173511 525014 173563 525059
rect 173617 525093 173669 525124
rect 173617 525059 173625 525093
rect 173659 525059 173669 525093
rect 173617 525014 173669 525059
rect 174615 525093 174667 525124
rect 174615 525059 174625 525093
rect 174659 525059 174667 525093
rect 174615 525014 174667 525059
rect 174905 525093 174957 525124
rect 174905 525059 174913 525093
rect 174947 525059 174957 525093
rect 174905 525014 174957 525059
rect 175903 525093 175955 525124
rect 175903 525059 175913 525093
rect 175947 525059 175955 525093
rect 175903 525014 175955 525059
rect 176009 525093 176061 525124
rect 176009 525059 176017 525093
rect 176051 525059 176061 525093
rect 176009 525014 176061 525059
rect 177007 525093 177059 525124
rect 177007 525059 177017 525093
rect 177051 525059 177059 525093
rect 177007 525014 177059 525059
rect 177113 525093 177165 525124
rect 177113 525059 177121 525093
rect 177155 525059 177165 525093
rect 177113 525014 177165 525059
rect 178111 525093 178163 525124
rect 178111 525059 178121 525093
rect 178155 525059 178163 525093
rect 178111 525014 178163 525059
rect 178217 525093 178269 525124
rect 178217 525059 178225 525093
rect 178259 525059 178269 525093
rect 178217 525014 178269 525059
rect 179215 525093 179267 525124
rect 179215 525059 179225 525093
rect 179259 525059 179267 525093
rect 179215 525014 179267 525059
rect 179321 525093 179373 525124
rect 179321 525059 179329 525093
rect 179363 525059 179373 525093
rect 179321 525014 179373 525059
rect 179767 525093 179819 525124
rect 179767 525059 179777 525093
rect 179811 525059 179819 525093
rect 179767 525014 179819 525059
rect 180057 525093 180109 525124
rect 180057 525059 180065 525093
rect 180099 525059 180109 525093
rect 180057 525014 180109 525059
rect 181055 525093 181107 525124
rect 181055 525059 181065 525093
rect 181099 525059 181107 525093
rect 181055 525014 181107 525059
rect 181161 525093 181213 525124
rect 181161 525059 181169 525093
rect 181203 525059 181213 525093
rect 181161 525014 181213 525059
rect 182159 525093 182211 525124
rect 182159 525059 182169 525093
rect 182203 525059 182211 525093
rect 182159 525014 182211 525059
rect 182265 525093 182317 525124
rect 182265 525059 182273 525093
rect 182307 525059 182317 525093
rect 182265 525014 182317 525059
rect 183263 525093 183315 525124
rect 183263 525059 183273 525093
rect 183307 525059 183315 525093
rect 183263 525014 183315 525059
rect 183369 525093 183421 525124
rect 183369 525059 183377 525093
rect 183411 525059 183421 525093
rect 183369 525014 183421 525059
rect 184367 525093 184419 525124
rect 184367 525059 184377 525093
rect 184411 525059 184419 525093
rect 184367 525014 184419 525059
rect 184473 525093 184525 525124
rect 184473 525059 184481 525093
rect 184515 525059 184525 525093
rect 184473 525014 184525 525059
rect 184919 525093 184971 525124
rect 184919 525059 184929 525093
rect 184963 525059 184971 525093
rect 184919 525014 184971 525059
rect 185209 525093 185261 525124
rect 185209 525059 185217 525093
rect 185251 525059 185261 525093
rect 185209 525014 185261 525059
rect 186207 525093 186259 525124
rect 186207 525059 186217 525093
rect 186251 525059 186259 525093
rect 186207 525014 186259 525059
rect 186313 525093 186365 525124
rect 186313 525059 186321 525093
rect 186355 525059 186365 525093
rect 186313 525014 186365 525059
rect 186943 525093 186995 525124
rect 186943 525059 186953 525093
rect 186987 525059 186995 525093
rect 186943 525014 186995 525059
rect 187233 525091 187285 525124
rect 187233 525057 187241 525091
rect 187275 525057 187285 525091
rect 187233 525014 187285 525057
rect 187403 525091 187455 525124
rect 187403 525057 187413 525091
rect 187447 525057 187455 525091
rect 187403 525014 187455 525057
rect 172237 524197 172289 524240
rect 172237 524163 172245 524197
rect 172279 524163 172289 524197
rect 172237 524130 172289 524163
rect 172407 524197 172459 524240
rect 172407 524163 172417 524197
rect 172451 524163 172459 524197
rect 172407 524130 172459 524163
rect 172513 524195 172565 524240
rect 172513 524161 172521 524195
rect 172555 524161 172565 524195
rect 172513 524130 172565 524161
rect 173511 524195 173563 524240
rect 173511 524161 173521 524195
rect 173555 524161 173563 524195
rect 173511 524130 173563 524161
rect 173617 524195 173669 524240
rect 173617 524161 173625 524195
rect 173659 524161 173669 524195
rect 173617 524130 173669 524161
rect 174615 524195 174667 524240
rect 174615 524161 174625 524195
rect 174659 524161 174667 524195
rect 174615 524130 174667 524161
rect 174721 524195 174773 524240
rect 174721 524161 174729 524195
rect 174763 524161 174773 524195
rect 174721 524130 174773 524161
rect 175719 524195 175771 524240
rect 175719 524161 175729 524195
rect 175763 524161 175771 524195
rect 175719 524130 175771 524161
rect 175825 524195 175877 524240
rect 175825 524161 175833 524195
rect 175867 524161 175877 524195
rect 175825 524130 175877 524161
rect 176823 524195 176875 524240
rect 176823 524161 176833 524195
rect 176867 524161 176875 524195
rect 176823 524130 176875 524161
rect 176929 524202 176981 524240
rect 176929 524168 176937 524202
rect 176971 524168 176981 524202
rect 176929 524130 176981 524168
rect 177191 524202 177243 524240
rect 177191 524168 177201 524202
rect 177235 524168 177243 524202
rect 177191 524130 177243 524168
rect 177481 524195 177533 524240
rect 177481 524161 177489 524195
rect 177523 524161 177533 524195
rect 177481 524130 177533 524161
rect 178479 524195 178531 524240
rect 178479 524161 178489 524195
rect 178523 524161 178531 524195
rect 178479 524130 178531 524161
rect 178585 524195 178637 524240
rect 178585 524161 178593 524195
rect 178627 524161 178637 524195
rect 178585 524130 178637 524161
rect 179583 524195 179635 524240
rect 179583 524161 179593 524195
rect 179627 524161 179635 524195
rect 179583 524130 179635 524161
rect 179689 524195 179741 524240
rect 179689 524161 179697 524195
rect 179731 524161 179741 524195
rect 179689 524130 179741 524161
rect 180687 524195 180739 524240
rect 180687 524161 180697 524195
rect 180731 524161 180739 524195
rect 180687 524130 180739 524161
rect 180793 524195 180845 524240
rect 180793 524161 180801 524195
rect 180835 524161 180845 524195
rect 180793 524130 180845 524161
rect 181791 524195 181843 524240
rect 181791 524161 181801 524195
rect 181835 524161 181843 524195
rect 181791 524130 181843 524161
rect 181897 524195 181949 524240
rect 181897 524161 181905 524195
rect 181939 524161 181949 524195
rect 181897 524130 181949 524161
rect 182343 524195 182395 524240
rect 182343 524161 182353 524195
rect 182387 524161 182395 524195
rect 182343 524130 182395 524161
rect 182633 524195 182685 524240
rect 182633 524161 182641 524195
rect 182675 524161 182685 524195
rect 182633 524130 182685 524161
rect 183631 524195 183683 524240
rect 183631 524161 183641 524195
rect 183675 524161 183683 524195
rect 183631 524130 183683 524161
rect 183737 524195 183789 524240
rect 183737 524161 183745 524195
rect 183779 524161 183789 524195
rect 183737 524130 183789 524161
rect 184735 524195 184787 524240
rect 184735 524161 184745 524195
rect 184779 524161 184787 524195
rect 184735 524130 184787 524161
rect 184841 524195 184893 524240
rect 184841 524161 184849 524195
rect 184883 524161 184893 524195
rect 184841 524130 184893 524161
rect 185839 524195 185891 524240
rect 185839 524161 185849 524195
rect 185883 524161 185891 524195
rect 185839 524130 185891 524161
rect 185945 524195 185997 524240
rect 185945 524161 185953 524195
rect 185987 524161 185997 524195
rect 185945 524130 185997 524161
rect 186943 524195 186995 524240
rect 186943 524161 186953 524195
rect 186987 524161 186995 524195
rect 186943 524130 186995 524161
rect 187233 524197 187285 524240
rect 187233 524163 187241 524197
rect 187275 524163 187285 524197
rect 187233 524130 187285 524163
rect 187403 524197 187455 524240
rect 187403 524163 187413 524197
rect 187447 524163 187455 524197
rect 187403 524130 187455 524163
rect 172237 524003 172289 524036
rect 172237 523969 172245 524003
rect 172279 523969 172289 524003
rect 172237 523926 172289 523969
rect 172407 524003 172459 524036
rect 172407 523969 172417 524003
rect 172451 523969 172459 524003
rect 172407 523926 172459 523969
rect 172513 524005 172565 524036
rect 172513 523971 172521 524005
rect 172555 523971 172565 524005
rect 172513 523926 172565 523971
rect 173511 524005 173563 524036
rect 173511 523971 173521 524005
rect 173555 523971 173563 524005
rect 173511 523926 173563 523971
rect 173617 524005 173669 524036
rect 173617 523971 173625 524005
rect 173659 523971 173669 524005
rect 173617 523926 173669 523971
rect 174615 524005 174667 524036
rect 174615 523971 174625 524005
rect 174659 523971 174667 524005
rect 174615 523926 174667 523971
rect 174905 524005 174957 524036
rect 174905 523971 174913 524005
rect 174947 523971 174957 524005
rect 174905 523926 174957 523971
rect 175903 524005 175955 524036
rect 175903 523971 175913 524005
rect 175947 523971 175955 524005
rect 175903 523926 175955 523971
rect 176009 524005 176061 524036
rect 176009 523971 176017 524005
rect 176051 523971 176061 524005
rect 176009 523926 176061 523971
rect 177007 524005 177059 524036
rect 177007 523971 177017 524005
rect 177051 523971 177059 524005
rect 177007 523926 177059 523971
rect 177113 524005 177165 524036
rect 177113 523971 177121 524005
rect 177155 523971 177165 524005
rect 177113 523926 177165 523971
rect 178111 524005 178163 524036
rect 178111 523971 178121 524005
rect 178155 523971 178163 524005
rect 178111 523926 178163 523971
rect 178217 524005 178269 524036
rect 178217 523971 178225 524005
rect 178259 523971 178269 524005
rect 178217 523926 178269 523971
rect 179215 524005 179267 524036
rect 179215 523971 179225 524005
rect 179259 523971 179267 524005
rect 179215 523926 179267 523971
rect 179321 524005 179373 524036
rect 179321 523971 179329 524005
rect 179363 523971 179373 524005
rect 179321 523926 179373 523971
rect 179767 524005 179819 524036
rect 179767 523971 179777 524005
rect 179811 523971 179819 524005
rect 179767 523926 179819 523971
rect 180057 524005 180109 524036
rect 180057 523971 180065 524005
rect 180099 523971 180109 524005
rect 180057 523926 180109 523971
rect 181055 524005 181107 524036
rect 181055 523971 181065 524005
rect 181099 523971 181107 524005
rect 181055 523926 181107 523971
rect 181161 524005 181213 524036
rect 181161 523971 181169 524005
rect 181203 523971 181213 524005
rect 181161 523926 181213 523971
rect 182159 524005 182211 524036
rect 182159 523971 182169 524005
rect 182203 523971 182211 524005
rect 182159 523926 182211 523971
rect 182265 524005 182317 524036
rect 182265 523971 182273 524005
rect 182307 523971 182317 524005
rect 182265 523926 182317 523971
rect 183263 524005 183315 524036
rect 183263 523971 183273 524005
rect 183307 523971 183315 524005
rect 183263 523926 183315 523971
rect 183369 524005 183421 524036
rect 183369 523971 183377 524005
rect 183411 523971 183421 524005
rect 183369 523926 183421 523971
rect 184367 524005 184419 524036
rect 184367 523971 184377 524005
rect 184411 523971 184419 524005
rect 184367 523926 184419 523971
rect 184473 524005 184525 524036
rect 184473 523971 184481 524005
rect 184515 523971 184525 524005
rect 184473 523926 184525 523971
rect 184919 524005 184971 524036
rect 184919 523971 184929 524005
rect 184963 523971 184971 524005
rect 184919 523926 184971 523971
rect 185209 524005 185261 524036
rect 185209 523971 185217 524005
rect 185251 523971 185261 524005
rect 185209 523926 185261 523971
rect 186207 524005 186259 524036
rect 186207 523971 186217 524005
rect 186251 523971 186259 524005
rect 186207 523926 186259 523971
rect 186313 524005 186365 524036
rect 186313 523971 186321 524005
rect 186355 523971 186365 524005
rect 186313 523926 186365 523971
rect 186943 524005 186995 524036
rect 186943 523971 186953 524005
rect 186987 523971 186995 524005
rect 186943 523926 186995 523971
rect 187233 524003 187285 524036
rect 187233 523969 187241 524003
rect 187275 523969 187285 524003
rect 187233 523926 187285 523969
rect 187403 524003 187455 524036
rect 187403 523969 187413 524003
rect 187447 523969 187455 524003
rect 187403 523926 187455 523969
rect 172237 523109 172289 523152
rect 172237 523075 172245 523109
rect 172279 523075 172289 523109
rect 172237 523042 172289 523075
rect 172407 523109 172459 523152
rect 172407 523075 172417 523109
rect 172451 523075 172459 523109
rect 172407 523042 172459 523075
rect 172513 523107 172565 523152
rect 172513 523073 172521 523107
rect 172555 523073 172565 523107
rect 172513 523042 172565 523073
rect 173511 523107 173563 523152
rect 173511 523073 173521 523107
rect 173555 523073 173563 523107
rect 173511 523042 173563 523073
rect 173617 523107 173669 523152
rect 173617 523073 173625 523107
rect 173659 523073 173669 523107
rect 173617 523042 173669 523073
rect 174615 523107 174667 523152
rect 174615 523073 174625 523107
rect 174659 523073 174667 523107
rect 174615 523042 174667 523073
rect 174721 523107 174773 523152
rect 174721 523073 174729 523107
rect 174763 523073 174773 523107
rect 174721 523042 174773 523073
rect 175719 523107 175771 523152
rect 175719 523073 175729 523107
rect 175763 523073 175771 523107
rect 175719 523042 175771 523073
rect 175825 523107 175877 523152
rect 175825 523073 175833 523107
rect 175867 523073 175877 523107
rect 175825 523042 175877 523073
rect 176823 523107 176875 523152
rect 176823 523073 176833 523107
rect 176867 523073 176875 523107
rect 176823 523042 176875 523073
rect 176929 523114 176981 523152
rect 176929 523080 176937 523114
rect 176971 523080 176981 523114
rect 176929 523042 176981 523080
rect 177191 523114 177243 523152
rect 177191 523080 177201 523114
rect 177235 523080 177243 523114
rect 177191 523042 177243 523080
rect 177481 523107 177533 523152
rect 177481 523073 177489 523107
rect 177523 523073 177533 523107
rect 177481 523042 177533 523073
rect 178479 523107 178531 523152
rect 178479 523073 178489 523107
rect 178523 523073 178531 523107
rect 178479 523042 178531 523073
rect 178585 523107 178637 523152
rect 178585 523073 178593 523107
rect 178627 523073 178637 523107
rect 178585 523042 178637 523073
rect 179583 523107 179635 523152
rect 179583 523073 179593 523107
rect 179627 523073 179635 523107
rect 179583 523042 179635 523073
rect 179689 523107 179741 523152
rect 179689 523073 179697 523107
rect 179731 523073 179741 523107
rect 179689 523042 179741 523073
rect 180687 523107 180739 523152
rect 180687 523073 180697 523107
rect 180731 523073 180739 523107
rect 180687 523042 180739 523073
rect 180793 523107 180845 523152
rect 180793 523073 180801 523107
rect 180835 523073 180845 523107
rect 180793 523042 180845 523073
rect 181791 523107 181843 523152
rect 181791 523073 181801 523107
rect 181835 523073 181843 523107
rect 181791 523042 181843 523073
rect 181897 523107 181949 523152
rect 181897 523073 181905 523107
rect 181939 523073 181949 523107
rect 181897 523042 181949 523073
rect 182343 523107 182395 523152
rect 182343 523073 182353 523107
rect 182387 523073 182395 523107
rect 182343 523042 182395 523073
rect 182633 523107 182685 523152
rect 182633 523073 182641 523107
rect 182675 523073 182685 523107
rect 182633 523042 182685 523073
rect 183631 523107 183683 523152
rect 183631 523073 183641 523107
rect 183675 523073 183683 523107
rect 183631 523042 183683 523073
rect 183737 523107 183789 523152
rect 183737 523073 183745 523107
rect 183779 523073 183789 523107
rect 183737 523042 183789 523073
rect 184735 523107 184787 523152
rect 184735 523073 184745 523107
rect 184779 523073 184787 523107
rect 184735 523042 184787 523073
rect 184841 523107 184893 523152
rect 184841 523073 184849 523107
rect 184883 523073 184893 523107
rect 184841 523042 184893 523073
rect 185839 523107 185891 523152
rect 185839 523073 185849 523107
rect 185883 523073 185891 523107
rect 185839 523042 185891 523073
rect 185945 523107 185997 523152
rect 185945 523073 185953 523107
rect 185987 523073 185997 523107
rect 185945 523042 185997 523073
rect 186943 523107 186995 523152
rect 186943 523073 186953 523107
rect 186987 523073 186995 523107
rect 186943 523042 186995 523073
rect 187233 523109 187285 523152
rect 187233 523075 187241 523109
rect 187275 523075 187285 523109
rect 187233 523042 187285 523075
rect 187403 523109 187455 523152
rect 187403 523075 187413 523109
rect 187447 523075 187455 523109
rect 187403 523042 187455 523075
rect 172237 522915 172289 522948
rect 172237 522881 172245 522915
rect 172279 522881 172289 522915
rect 172237 522838 172289 522881
rect 172407 522915 172459 522948
rect 172407 522881 172417 522915
rect 172451 522881 172459 522915
rect 172407 522838 172459 522881
rect 172513 522917 172565 522948
rect 172513 522883 172521 522917
rect 172555 522883 172565 522917
rect 172513 522838 172565 522883
rect 173511 522917 173563 522948
rect 173511 522883 173521 522917
rect 173555 522883 173563 522917
rect 173511 522838 173563 522883
rect 173617 522917 173669 522948
rect 173617 522883 173625 522917
rect 173659 522883 173669 522917
rect 173617 522838 173669 522883
rect 174615 522917 174667 522948
rect 174615 522883 174625 522917
rect 174659 522883 174667 522917
rect 174615 522838 174667 522883
rect 174905 522917 174957 522948
rect 174905 522883 174913 522917
rect 174947 522883 174957 522917
rect 174905 522838 174957 522883
rect 175903 522917 175955 522948
rect 175903 522883 175913 522917
rect 175947 522883 175955 522917
rect 175903 522838 175955 522883
rect 176009 522917 176061 522948
rect 176009 522883 176017 522917
rect 176051 522883 176061 522917
rect 176009 522838 176061 522883
rect 177007 522917 177059 522948
rect 177007 522883 177017 522917
rect 177051 522883 177059 522917
rect 177007 522838 177059 522883
rect 177113 522917 177165 522948
rect 177113 522883 177121 522917
rect 177155 522883 177165 522917
rect 177113 522838 177165 522883
rect 178111 522917 178163 522948
rect 178111 522883 178121 522917
rect 178155 522883 178163 522917
rect 178111 522838 178163 522883
rect 178217 522917 178269 522948
rect 178217 522883 178225 522917
rect 178259 522883 178269 522917
rect 178217 522838 178269 522883
rect 179215 522917 179267 522948
rect 179215 522883 179225 522917
rect 179259 522883 179267 522917
rect 179215 522838 179267 522883
rect 179321 522917 179373 522948
rect 179321 522883 179329 522917
rect 179363 522883 179373 522917
rect 179321 522838 179373 522883
rect 179767 522917 179819 522948
rect 179767 522883 179777 522917
rect 179811 522883 179819 522917
rect 179767 522838 179819 522883
rect 180057 522917 180109 522948
rect 180057 522883 180065 522917
rect 180099 522883 180109 522917
rect 180057 522838 180109 522883
rect 181055 522917 181107 522948
rect 181055 522883 181065 522917
rect 181099 522883 181107 522917
rect 181055 522838 181107 522883
rect 181161 522917 181213 522948
rect 181161 522883 181169 522917
rect 181203 522883 181213 522917
rect 181161 522838 181213 522883
rect 182159 522917 182211 522948
rect 182159 522883 182169 522917
rect 182203 522883 182211 522917
rect 182159 522838 182211 522883
rect 182265 522917 182317 522948
rect 182265 522883 182273 522917
rect 182307 522883 182317 522917
rect 182265 522838 182317 522883
rect 183263 522917 183315 522948
rect 183263 522883 183273 522917
rect 183307 522883 183315 522917
rect 183263 522838 183315 522883
rect 183369 522917 183421 522948
rect 183369 522883 183377 522917
rect 183411 522883 183421 522917
rect 183369 522838 183421 522883
rect 184367 522917 184419 522948
rect 184367 522883 184377 522917
rect 184411 522883 184419 522917
rect 184367 522838 184419 522883
rect 184473 522917 184525 522948
rect 184473 522883 184481 522917
rect 184515 522883 184525 522917
rect 184473 522838 184525 522883
rect 184919 522917 184971 522948
rect 184919 522883 184929 522917
rect 184963 522883 184971 522917
rect 184919 522838 184971 522883
rect 185209 522917 185261 522948
rect 185209 522883 185217 522917
rect 185251 522883 185261 522917
rect 185209 522838 185261 522883
rect 186207 522917 186259 522948
rect 186207 522883 186217 522917
rect 186251 522883 186259 522917
rect 186207 522838 186259 522883
rect 186313 522917 186365 522948
rect 186313 522883 186321 522917
rect 186355 522883 186365 522917
rect 186313 522838 186365 522883
rect 186943 522917 186995 522948
rect 186943 522883 186953 522917
rect 186987 522883 186995 522917
rect 186943 522838 186995 522883
rect 187233 522915 187285 522948
rect 187233 522881 187241 522915
rect 187275 522881 187285 522915
rect 187233 522838 187285 522881
rect 187403 522915 187455 522948
rect 187403 522881 187413 522915
rect 187447 522881 187455 522915
rect 187403 522838 187455 522881
rect 172237 522021 172289 522064
rect 172237 521987 172245 522021
rect 172279 521987 172289 522021
rect 172237 521954 172289 521987
rect 172407 522021 172459 522064
rect 172407 521987 172417 522021
rect 172451 521987 172459 522021
rect 172407 521954 172459 521987
rect 172513 522019 172565 522064
rect 172513 521985 172521 522019
rect 172555 521985 172565 522019
rect 172513 521954 172565 521985
rect 173511 522019 173563 522064
rect 173511 521985 173521 522019
rect 173555 521985 173563 522019
rect 173511 521954 173563 521985
rect 173617 522019 173669 522064
rect 173617 521985 173625 522019
rect 173659 521985 173669 522019
rect 173617 521954 173669 521985
rect 174615 522019 174667 522064
rect 174615 521985 174625 522019
rect 174659 521985 174667 522019
rect 174615 521954 174667 521985
rect 174721 522019 174773 522064
rect 174721 521985 174729 522019
rect 174763 521985 174773 522019
rect 174721 521954 174773 521985
rect 175719 522019 175771 522064
rect 175719 521985 175729 522019
rect 175763 521985 175771 522019
rect 175719 521954 175771 521985
rect 175825 522019 175877 522064
rect 175825 521985 175833 522019
rect 175867 521985 175877 522019
rect 175825 521954 175877 521985
rect 176823 522019 176875 522064
rect 176823 521985 176833 522019
rect 176867 521985 176875 522019
rect 176823 521954 176875 521985
rect 176929 522026 176981 522064
rect 176929 521992 176937 522026
rect 176971 521992 176981 522026
rect 176929 521954 176981 521992
rect 177191 522026 177243 522064
rect 177191 521992 177201 522026
rect 177235 521992 177243 522026
rect 177191 521954 177243 521992
rect 177481 522019 177533 522064
rect 177481 521985 177489 522019
rect 177523 521985 177533 522019
rect 177481 521954 177533 521985
rect 178479 522019 178531 522064
rect 178479 521985 178489 522019
rect 178523 521985 178531 522019
rect 178479 521954 178531 521985
rect 178585 522019 178637 522064
rect 178585 521985 178593 522019
rect 178627 521985 178637 522019
rect 178585 521954 178637 521985
rect 179583 522019 179635 522064
rect 179583 521985 179593 522019
rect 179627 521985 179635 522019
rect 179583 521954 179635 521985
rect 179689 522019 179741 522064
rect 179689 521985 179697 522019
rect 179731 521985 179741 522019
rect 179689 521954 179741 521985
rect 180687 522019 180739 522064
rect 180687 521985 180697 522019
rect 180731 521985 180739 522019
rect 180687 521954 180739 521985
rect 180793 522019 180845 522064
rect 180793 521985 180801 522019
rect 180835 521985 180845 522019
rect 180793 521954 180845 521985
rect 181791 522019 181843 522064
rect 181791 521985 181801 522019
rect 181835 521985 181843 522019
rect 181791 521954 181843 521985
rect 181897 522019 181949 522064
rect 181897 521985 181905 522019
rect 181939 521985 181949 522019
rect 181897 521954 181949 521985
rect 182343 522019 182395 522064
rect 182343 521985 182353 522019
rect 182387 521985 182395 522019
rect 182343 521954 182395 521985
rect 182633 522019 182685 522064
rect 182633 521985 182641 522019
rect 182675 521985 182685 522019
rect 182633 521954 182685 521985
rect 183631 522019 183683 522064
rect 183631 521985 183641 522019
rect 183675 521985 183683 522019
rect 183631 521954 183683 521985
rect 183737 522019 183789 522064
rect 183737 521985 183745 522019
rect 183779 521985 183789 522019
rect 183737 521954 183789 521985
rect 184735 522019 184787 522064
rect 184735 521985 184745 522019
rect 184779 521985 184787 522019
rect 184735 521954 184787 521985
rect 184841 522019 184893 522064
rect 184841 521985 184849 522019
rect 184883 521985 184893 522019
rect 184841 521954 184893 521985
rect 185839 522019 185891 522064
rect 185839 521985 185849 522019
rect 185883 521985 185891 522019
rect 185839 521954 185891 521985
rect 185945 522019 185997 522064
rect 185945 521985 185953 522019
rect 185987 521985 185997 522019
rect 185945 521954 185997 521985
rect 186943 522019 186995 522064
rect 186943 521985 186953 522019
rect 186987 521985 186995 522019
rect 186943 521954 186995 521985
rect 187233 522021 187285 522064
rect 187233 521987 187241 522021
rect 187275 521987 187285 522021
rect 187233 521954 187285 521987
rect 187403 522021 187455 522064
rect 187403 521987 187413 522021
rect 187447 521987 187455 522021
rect 187403 521954 187455 521987
rect 172237 521827 172289 521860
rect 172237 521793 172245 521827
rect 172279 521793 172289 521827
rect 172237 521750 172289 521793
rect 172407 521827 172459 521860
rect 172407 521793 172417 521827
rect 172451 521793 172459 521827
rect 172407 521750 172459 521793
rect 172513 521829 172565 521860
rect 172513 521795 172521 521829
rect 172555 521795 172565 521829
rect 172513 521750 172565 521795
rect 173511 521829 173563 521860
rect 173511 521795 173521 521829
rect 173555 521795 173563 521829
rect 173511 521750 173563 521795
rect 173617 521829 173669 521860
rect 173617 521795 173625 521829
rect 173659 521795 173669 521829
rect 173617 521750 173669 521795
rect 174615 521829 174667 521860
rect 174615 521795 174625 521829
rect 174659 521795 174667 521829
rect 174615 521750 174667 521795
rect 174905 521829 174957 521860
rect 174905 521795 174913 521829
rect 174947 521795 174957 521829
rect 174905 521750 174957 521795
rect 175903 521829 175955 521860
rect 175903 521795 175913 521829
rect 175947 521795 175955 521829
rect 175903 521750 175955 521795
rect 176009 521829 176061 521860
rect 176009 521795 176017 521829
rect 176051 521795 176061 521829
rect 176009 521750 176061 521795
rect 177007 521829 177059 521860
rect 177007 521795 177017 521829
rect 177051 521795 177059 521829
rect 177007 521750 177059 521795
rect 177113 521829 177165 521860
rect 177113 521795 177121 521829
rect 177155 521795 177165 521829
rect 177113 521750 177165 521795
rect 178111 521829 178163 521860
rect 178111 521795 178121 521829
rect 178155 521795 178163 521829
rect 178111 521750 178163 521795
rect 178217 521829 178269 521860
rect 178217 521795 178225 521829
rect 178259 521795 178269 521829
rect 178217 521750 178269 521795
rect 179215 521829 179267 521860
rect 179215 521795 179225 521829
rect 179259 521795 179267 521829
rect 179215 521750 179267 521795
rect 179321 521829 179373 521860
rect 179321 521795 179329 521829
rect 179363 521795 179373 521829
rect 179321 521750 179373 521795
rect 179767 521829 179819 521860
rect 179767 521795 179777 521829
rect 179811 521795 179819 521829
rect 179767 521750 179819 521795
rect 180057 521829 180109 521860
rect 180057 521795 180065 521829
rect 180099 521795 180109 521829
rect 180057 521750 180109 521795
rect 181055 521829 181107 521860
rect 181055 521795 181065 521829
rect 181099 521795 181107 521829
rect 181055 521750 181107 521795
rect 181161 521829 181213 521860
rect 181161 521795 181169 521829
rect 181203 521795 181213 521829
rect 181161 521750 181213 521795
rect 182159 521829 182211 521860
rect 182159 521795 182169 521829
rect 182203 521795 182211 521829
rect 182159 521750 182211 521795
rect 182265 521829 182317 521860
rect 182265 521795 182273 521829
rect 182307 521795 182317 521829
rect 182265 521750 182317 521795
rect 183263 521829 183315 521860
rect 183263 521795 183273 521829
rect 183307 521795 183315 521829
rect 183263 521750 183315 521795
rect 183369 521829 183421 521860
rect 183369 521795 183377 521829
rect 183411 521795 183421 521829
rect 183369 521750 183421 521795
rect 184367 521829 184419 521860
rect 184367 521795 184377 521829
rect 184411 521795 184419 521829
rect 184367 521750 184419 521795
rect 184473 521829 184525 521860
rect 184473 521795 184481 521829
rect 184515 521795 184525 521829
rect 184473 521750 184525 521795
rect 184919 521829 184971 521860
rect 184919 521795 184929 521829
rect 184963 521795 184971 521829
rect 184919 521750 184971 521795
rect 185209 521829 185261 521860
rect 185209 521795 185217 521829
rect 185251 521795 185261 521829
rect 185209 521750 185261 521795
rect 186207 521829 186259 521860
rect 186207 521795 186217 521829
rect 186251 521795 186259 521829
rect 186207 521750 186259 521795
rect 186313 521829 186365 521860
rect 186313 521795 186321 521829
rect 186355 521795 186365 521829
rect 186313 521750 186365 521795
rect 186943 521829 186995 521860
rect 186943 521795 186953 521829
rect 186987 521795 186995 521829
rect 186943 521750 186995 521795
rect 187233 521827 187285 521860
rect 187233 521793 187241 521827
rect 187275 521793 187285 521827
rect 187233 521750 187285 521793
rect 187403 521827 187455 521860
rect 187403 521793 187413 521827
rect 187447 521793 187455 521827
rect 187403 521750 187455 521793
rect 172237 520933 172289 520976
rect 172237 520899 172245 520933
rect 172279 520899 172289 520933
rect 172237 520866 172289 520899
rect 172407 520933 172459 520976
rect 172407 520899 172417 520933
rect 172451 520899 172459 520933
rect 172407 520866 172459 520899
rect 172513 520931 172565 520976
rect 172513 520897 172521 520931
rect 172555 520897 172565 520931
rect 172513 520866 172565 520897
rect 173511 520931 173563 520976
rect 173511 520897 173521 520931
rect 173555 520897 173563 520931
rect 173511 520866 173563 520897
rect 173617 520931 173669 520976
rect 173617 520897 173625 520931
rect 173659 520897 173669 520931
rect 173617 520866 173669 520897
rect 174615 520931 174667 520976
rect 174615 520897 174625 520931
rect 174659 520897 174667 520931
rect 174615 520866 174667 520897
rect 174721 520931 174773 520976
rect 174721 520897 174729 520931
rect 174763 520897 174773 520931
rect 174721 520866 174773 520897
rect 175719 520931 175771 520976
rect 175719 520897 175729 520931
rect 175763 520897 175771 520931
rect 175719 520866 175771 520897
rect 175825 520931 175877 520976
rect 175825 520897 175833 520931
rect 175867 520897 175877 520931
rect 175825 520866 175877 520897
rect 176823 520931 176875 520976
rect 176823 520897 176833 520931
rect 176867 520897 176875 520931
rect 176823 520866 176875 520897
rect 176929 520938 176981 520976
rect 176929 520904 176937 520938
rect 176971 520904 176981 520938
rect 176929 520866 176981 520904
rect 177191 520938 177243 520976
rect 177191 520904 177201 520938
rect 177235 520904 177243 520938
rect 177191 520866 177243 520904
rect 177481 520931 177533 520976
rect 177481 520897 177489 520931
rect 177523 520897 177533 520931
rect 177481 520866 177533 520897
rect 178479 520931 178531 520976
rect 178479 520897 178489 520931
rect 178523 520897 178531 520931
rect 178479 520866 178531 520897
rect 178585 520931 178637 520976
rect 178585 520897 178593 520931
rect 178627 520897 178637 520931
rect 178585 520866 178637 520897
rect 179583 520931 179635 520976
rect 179583 520897 179593 520931
rect 179627 520897 179635 520931
rect 179583 520866 179635 520897
rect 179689 520931 179741 520976
rect 179689 520897 179697 520931
rect 179731 520897 179741 520931
rect 179689 520866 179741 520897
rect 180687 520931 180739 520976
rect 180687 520897 180697 520931
rect 180731 520897 180739 520931
rect 180687 520866 180739 520897
rect 180793 520931 180845 520976
rect 180793 520897 180801 520931
rect 180835 520897 180845 520931
rect 180793 520866 180845 520897
rect 181791 520931 181843 520976
rect 181791 520897 181801 520931
rect 181835 520897 181843 520931
rect 181791 520866 181843 520897
rect 181897 520931 181949 520976
rect 181897 520897 181905 520931
rect 181939 520897 181949 520931
rect 181897 520866 181949 520897
rect 182343 520931 182395 520976
rect 182343 520897 182353 520931
rect 182387 520897 182395 520931
rect 182343 520866 182395 520897
rect 182633 520931 182685 520976
rect 182633 520897 182641 520931
rect 182675 520897 182685 520931
rect 182633 520866 182685 520897
rect 183631 520931 183683 520976
rect 183631 520897 183641 520931
rect 183675 520897 183683 520931
rect 183631 520866 183683 520897
rect 183737 520931 183789 520976
rect 183737 520897 183745 520931
rect 183779 520897 183789 520931
rect 183737 520866 183789 520897
rect 184735 520931 184787 520976
rect 184735 520897 184745 520931
rect 184779 520897 184787 520931
rect 184735 520866 184787 520897
rect 184841 520931 184893 520976
rect 184841 520897 184849 520931
rect 184883 520897 184893 520931
rect 184841 520866 184893 520897
rect 185839 520931 185891 520976
rect 185839 520897 185849 520931
rect 185883 520897 185891 520931
rect 185839 520866 185891 520897
rect 185945 520931 185997 520976
rect 185945 520897 185953 520931
rect 185987 520897 185997 520931
rect 185945 520866 185997 520897
rect 186943 520931 186995 520976
rect 186943 520897 186953 520931
rect 186987 520897 186995 520931
rect 186943 520866 186995 520897
rect 187233 520933 187285 520976
rect 187233 520899 187241 520933
rect 187275 520899 187285 520933
rect 187233 520866 187285 520899
rect 187403 520933 187455 520976
rect 187403 520899 187413 520933
rect 187447 520899 187455 520933
rect 187403 520866 187455 520899
rect 172237 520739 172289 520772
rect 172237 520705 172245 520739
rect 172279 520705 172289 520739
rect 172237 520662 172289 520705
rect 172407 520739 172459 520772
rect 172407 520705 172417 520739
rect 172451 520705 172459 520739
rect 172407 520662 172459 520705
rect 172513 520741 172565 520772
rect 172513 520707 172521 520741
rect 172555 520707 172565 520741
rect 172513 520662 172565 520707
rect 173511 520741 173563 520772
rect 173511 520707 173521 520741
rect 173555 520707 173563 520741
rect 173511 520662 173563 520707
rect 173617 520741 173669 520772
rect 173617 520707 173625 520741
rect 173659 520707 173669 520741
rect 173617 520662 173669 520707
rect 174615 520741 174667 520772
rect 174615 520707 174625 520741
rect 174659 520707 174667 520741
rect 174615 520662 174667 520707
rect 174905 520741 174957 520772
rect 174905 520707 174913 520741
rect 174947 520707 174957 520741
rect 174905 520662 174957 520707
rect 175903 520741 175955 520772
rect 175903 520707 175913 520741
rect 175947 520707 175955 520741
rect 175903 520662 175955 520707
rect 176009 520741 176061 520772
rect 176009 520707 176017 520741
rect 176051 520707 176061 520741
rect 176009 520662 176061 520707
rect 177007 520741 177059 520772
rect 177007 520707 177017 520741
rect 177051 520707 177059 520741
rect 177007 520662 177059 520707
rect 177113 520741 177165 520772
rect 177113 520707 177121 520741
rect 177155 520707 177165 520741
rect 177113 520662 177165 520707
rect 178111 520741 178163 520772
rect 178111 520707 178121 520741
rect 178155 520707 178163 520741
rect 178111 520662 178163 520707
rect 178217 520741 178269 520772
rect 178217 520707 178225 520741
rect 178259 520707 178269 520741
rect 178217 520662 178269 520707
rect 179215 520741 179267 520772
rect 179215 520707 179225 520741
rect 179259 520707 179267 520741
rect 179215 520662 179267 520707
rect 179321 520741 179373 520772
rect 179321 520707 179329 520741
rect 179363 520707 179373 520741
rect 179321 520662 179373 520707
rect 179767 520741 179819 520772
rect 179767 520707 179777 520741
rect 179811 520707 179819 520741
rect 179767 520662 179819 520707
rect 180057 520741 180109 520772
rect 180057 520707 180065 520741
rect 180099 520707 180109 520741
rect 180057 520662 180109 520707
rect 181055 520741 181107 520772
rect 181055 520707 181065 520741
rect 181099 520707 181107 520741
rect 181055 520662 181107 520707
rect 181161 520741 181213 520772
rect 181161 520707 181169 520741
rect 181203 520707 181213 520741
rect 181161 520662 181213 520707
rect 182159 520741 182211 520772
rect 182159 520707 182169 520741
rect 182203 520707 182211 520741
rect 182159 520662 182211 520707
rect 182265 520741 182317 520772
rect 182265 520707 182273 520741
rect 182307 520707 182317 520741
rect 182265 520662 182317 520707
rect 183263 520741 183315 520772
rect 183263 520707 183273 520741
rect 183307 520707 183315 520741
rect 183263 520662 183315 520707
rect 183369 520741 183421 520772
rect 183369 520707 183377 520741
rect 183411 520707 183421 520741
rect 183369 520662 183421 520707
rect 184367 520741 184419 520772
rect 184367 520707 184377 520741
rect 184411 520707 184419 520741
rect 184367 520662 184419 520707
rect 184473 520741 184525 520772
rect 184473 520707 184481 520741
rect 184515 520707 184525 520741
rect 184473 520662 184525 520707
rect 184919 520741 184971 520772
rect 184919 520707 184929 520741
rect 184963 520707 184971 520741
rect 184919 520662 184971 520707
rect 185209 520741 185261 520772
rect 185209 520707 185217 520741
rect 185251 520707 185261 520741
rect 185209 520662 185261 520707
rect 186207 520741 186259 520772
rect 186207 520707 186217 520741
rect 186251 520707 186259 520741
rect 186207 520662 186259 520707
rect 186313 520741 186365 520772
rect 186313 520707 186321 520741
rect 186355 520707 186365 520741
rect 186313 520662 186365 520707
rect 186943 520741 186995 520772
rect 186943 520707 186953 520741
rect 186987 520707 186995 520741
rect 186943 520662 186995 520707
rect 187233 520739 187285 520772
rect 187233 520705 187241 520739
rect 187275 520705 187285 520739
rect 187233 520662 187285 520705
rect 187403 520739 187455 520772
rect 187403 520705 187413 520739
rect 187447 520705 187455 520739
rect 187403 520662 187455 520705
rect 172237 519845 172289 519888
rect 172237 519811 172245 519845
rect 172279 519811 172289 519845
rect 172237 519778 172289 519811
rect 172407 519845 172459 519888
rect 172407 519811 172417 519845
rect 172451 519811 172459 519845
rect 172407 519778 172459 519811
rect 172513 519843 172565 519888
rect 172513 519809 172521 519843
rect 172555 519809 172565 519843
rect 172513 519778 172565 519809
rect 173511 519843 173563 519888
rect 173511 519809 173521 519843
rect 173555 519809 173563 519843
rect 173511 519778 173563 519809
rect 173617 519843 173669 519888
rect 173617 519809 173625 519843
rect 173659 519809 173669 519843
rect 173617 519778 173669 519809
rect 174615 519843 174667 519888
rect 174615 519809 174625 519843
rect 174659 519809 174667 519843
rect 174615 519778 174667 519809
rect 174721 519843 174773 519888
rect 174721 519809 174729 519843
rect 174763 519809 174773 519843
rect 174721 519778 174773 519809
rect 175719 519843 175771 519888
rect 175719 519809 175729 519843
rect 175763 519809 175771 519843
rect 175719 519778 175771 519809
rect 175825 519843 175877 519888
rect 175825 519809 175833 519843
rect 175867 519809 175877 519843
rect 175825 519778 175877 519809
rect 176823 519843 176875 519888
rect 176823 519809 176833 519843
rect 176867 519809 176875 519843
rect 176823 519778 176875 519809
rect 176929 519850 176981 519888
rect 176929 519816 176937 519850
rect 176971 519816 176981 519850
rect 176929 519778 176981 519816
rect 177191 519850 177243 519888
rect 177191 519816 177201 519850
rect 177235 519816 177243 519850
rect 177191 519778 177243 519816
rect 177481 519843 177533 519888
rect 177481 519809 177489 519843
rect 177523 519809 177533 519843
rect 177481 519778 177533 519809
rect 178479 519843 178531 519888
rect 178479 519809 178489 519843
rect 178523 519809 178531 519843
rect 178479 519778 178531 519809
rect 178585 519843 178637 519888
rect 178585 519809 178593 519843
rect 178627 519809 178637 519843
rect 178585 519778 178637 519809
rect 179583 519843 179635 519888
rect 179583 519809 179593 519843
rect 179627 519809 179635 519843
rect 179583 519778 179635 519809
rect 179689 519843 179741 519888
rect 179689 519809 179697 519843
rect 179731 519809 179741 519843
rect 179689 519778 179741 519809
rect 180687 519843 180739 519888
rect 180687 519809 180697 519843
rect 180731 519809 180739 519843
rect 180687 519778 180739 519809
rect 180793 519843 180845 519888
rect 180793 519809 180801 519843
rect 180835 519809 180845 519843
rect 180793 519778 180845 519809
rect 181791 519843 181843 519888
rect 181791 519809 181801 519843
rect 181835 519809 181843 519843
rect 181791 519778 181843 519809
rect 181897 519843 181949 519888
rect 181897 519809 181905 519843
rect 181939 519809 181949 519843
rect 181897 519778 181949 519809
rect 182343 519843 182395 519888
rect 182343 519809 182353 519843
rect 182387 519809 182395 519843
rect 182343 519778 182395 519809
rect 182633 519843 182685 519888
rect 182633 519809 182641 519843
rect 182675 519809 182685 519843
rect 182633 519778 182685 519809
rect 183631 519843 183683 519888
rect 183631 519809 183641 519843
rect 183675 519809 183683 519843
rect 183631 519778 183683 519809
rect 183737 519843 183789 519888
rect 183737 519809 183745 519843
rect 183779 519809 183789 519843
rect 183737 519778 183789 519809
rect 184735 519843 184787 519888
rect 184735 519809 184745 519843
rect 184779 519809 184787 519843
rect 184735 519778 184787 519809
rect 184841 519843 184893 519888
rect 184841 519809 184849 519843
rect 184883 519809 184893 519843
rect 184841 519778 184893 519809
rect 185839 519843 185891 519888
rect 185839 519809 185849 519843
rect 185883 519809 185891 519843
rect 185839 519778 185891 519809
rect 185945 519843 185997 519888
rect 185945 519809 185953 519843
rect 185987 519809 185997 519843
rect 185945 519778 185997 519809
rect 186943 519843 186995 519888
rect 186943 519809 186953 519843
rect 186987 519809 186995 519843
rect 186943 519778 186995 519809
rect 187233 519845 187285 519888
rect 187233 519811 187241 519845
rect 187275 519811 187285 519845
rect 187233 519778 187285 519811
rect 187403 519845 187455 519888
rect 187403 519811 187413 519845
rect 187447 519811 187455 519845
rect 187403 519778 187455 519811
rect 172237 519651 172289 519684
rect 172237 519617 172245 519651
rect 172279 519617 172289 519651
rect 172237 519574 172289 519617
rect 172407 519651 172459 519684
rect 172407 519617 172417 519651
rect 172451 519617 172459 519651
rect 172407 519574 172459 519617
rect 172513 519653 172565 519684
rect 172513 519619 172521 519653
rect 172555 519619 172565 519653
rect 172513 519574 172565 519619
rect 173511 519653 173563 519684
rect 173511 519619 173521 519653
rect 173555 519619 173563 519653
rect 173511 519574 173563 519619
rect 173617 519653 173669 519684
rect 173617 519619 173625 519653
rect 173659 519619 173669 519653
rect 173617 519574 173669 519619
rect 174615 519653 174667 519684
rect 174615 519619 174625 519653
rect 174659 519619 174667 519653
rect 174615 519574 174667 519619
rect 174905 519653 174957 519684
rect 174905 519619 174913 519653
rect 174947 519619 174957 519653
rect 174905 519574 174957 519619
rect 175903 519653 175955 519684
rect 175903 519619 175913 519653
rect 175947 519619 175955 519653
rect 175903 519574 175955 519619
rect 176009 519653 176061 519684
rect 176009 519619 176017 519653
rect 176051 519619 176061 519653
rect 176009 519574 176061 519619
rect 177007 519653 177059 519684
rect 177007 519619 177017 519653
rect 177051 519619 177059 519653
rect 177007 519574 177059 519619
rect 177113 519653 177165 519684
rect 177113 519619 177121 519653
rect 177155 519619 177165 519653
rect 177113 519574 177165 519619
rect 178111 519653 178163 519684
rect 178111 519619 178121 519653
rect 178155 519619 178163 519653
rect 178111 519574 178163 519619
rect 178217 519653 178269 519684
rect 178217 519619 178225 519653
rect 178259 519619 178269 519653
rect 178217 519574 178269 519619
rect 179215 519653 179267 519684
rect 179215 519619 179225 519653
rect 179259 519619 179267 519653
rect 179215 519574 179267 519619
rect 179321 519653 179373 519684
rect 179321 519619 179329 519653
rect 179363 519619 179373 519653
rect 179321 519574 179373 519619
rect 179767 519653 179819 519684
rect 179767 519619 179777 519653
rect 179811 519619 179819 519653
rect 179767 519574 179819 519619
rect 180057 519653 180109 519684
rect 180057 519619 180065 519653
rect 180099 519619 180109 519653
rect 180057 519574 180109 519619
rect 181055 519653 181107 519684
rect 181055 519619 181065 519653
rect 181099 519619 181107 519653
rect 181055 519574 181107 519619
rect 181161 519653 181213 519684
rect 181161 519619 181169 519653
rect 181203 519619 181213 519653
rect 181161 519574 181213 519619
rect 182159 519653 182211 519684
rect 182159 519619 182169 519653
rect 182203 519619 182211 519653
rect 182159 519574 182211 519619
rect 182265 519653 182317 519684
rect 182265 519619 182273 519653
rect 182307 519619 182317 519653
rect 182265 519574 182317 519619
rect 183263 519653 183315 519684
rect 183263 519619 183273 519653
rect 183307 519619 183315 519653
rect 183263 519574 183315 519619
rect 183369 519653 183421 519684
rect 183369 519619 183377 519653
rect 183411 519619 183421 519653
rect 183369 519574 183421 519619
rect 184367 519653 184419 519684
rect 184367 519619 184377 519653
rect 184411 519619 184419 519653
rect 184367 519574 184419 519619
rect 184473 519653 184525 519684
rect 184473 519619 184481 519653
rect 184515 519619 184525 519653
rect 184473 519574 184525 519619
rect 184919 519653 184971 519684
rect 184919 519619 184929 519653
rect 184963 519619 184971 519653
rect 184919 519574 184971 519619
rect 185209 519653 185261 519684
rect 185209 519619 185217 519653
rect 185251 519619 185261 519653
rect 185209 519574 185261 519619
rect 186207 519653 186259 519684
rect 186207 519619 186217 519653
rect 186251 519619 186259 519653
rect 186207 519574 186259 519619
rect 186313 519653 186365 519684
rect 186313 519619 186321 519653
rect 186355 519619 186365 519653
rect 186313 519574 186365 519619
rect 186943 519653 186995 519684
rect 186943 519619 186953 519653
rect 186987 519619 186995 519653
rect 186943 519574 186995 519619
rect 187233 519651 187285 519684
rect 187233 519617 187241 519651
rect 187275 519617 187285 519651
rect 187233 519574 187285 519617
rect 187403 519651 187455 519684
rect 187403 519617 187413 519651
rect 187447 519617 187455 519651
rect 187403 519574 187455 519617
rect 172237 518757 172289 518800
rect 172237 518723 172245 518757
rect 172279 518723 172289 518757
rect 172237 518690 172289 518723
rect 172407 518757 172459 518800
rect 172407 518723 172417 518757
rect 172451 518723 172459 518757
rect 172407 518690 172459 518723
rect 172513 518755 172565 518800
rect 172513 518721 172521 518755
rect 172555 518721 172565 518755
rect 172513 518690 172565 518721
rect 173511 518755 173563 518800
rect 173511 518721 173521 518755
rect 173555 518721 173563 518755
rect 173511 518690 173563 518721
rect 173617 518755 173669 518800
rect 173617 518721 173625 518755
rect 173659 518721 173669 518755
rect 173617 518690 173669 518721
rect 174615 518755 174667 518800
rect 174615 518721 174625 518755
rect 174659 518721 174667 518755
rect 174615 518690 174667 518721
rect 174721 518755 174773 518800
rect 174721 518721 174729 518755
rect 174763 518721 174773 518755
rect 174721 518690 174773 518721
rect 175719 518755 175771 518800
rect 175719 518721 175729 518755
rect 175763 518721 175771 518755
rect 175719 518690 175771 518721
rect 175825 518755 175877 518800
rect 175825 518721 175833 518755
rect 175867 518721 175877 518755
rect 175825 518690 175877 518721
rect 176823 518755 176875 518800
rect 176823 518721 176833 518755
rect 176867 518721 176875 518755
rect 176823 518690 176875 518721
rect 176929 518762 176981 518800
rect 176929 518728 176937 518762
rect 176971 518728 176981 518762
rect 176929 518690 176981 518728
rect 177191 518762 177243 518800
rect 177191 518728 177201 518762
rect 177235 518728 177243 518762
rect 177191 518690 177243 518728
rect 177481 518755 177533 518800
rect 177481 518721 177489 518755
rect 177523 518721 177533 518755
rect 177481 518690 177533 518721
rect 178479 518755 178531 518800
rect 178479 518721 178489 518755
rect 178523 518721 178531 518755
rect 178479 518690 178531 518721
rect 178585 518755 178637 518800
rect 178585 518721 178593 518755
rect 178627 518721 178637 518755
rect 178585 518690 178637 518721
rect 179583 518755 179635 518800
rect 179583 518721 179593 518755
rect 179627 518721 179635 518755
rect 179583 518690 179635 518721
rect 179689 518755 179741 518800
rect 179689 518721 179697 518755
rect 179731 518721 179741 518755
rect 179689 518690 179741 518721
rect 180687 518755 180739 518800
rect 180687 518721 180697 518755
rect 180731 518721 180739 518755
rect 180687 518690 180739 518721
rect 180793 518755 180845 518800
rect 180793 518721 180801 518755
rect 180835 518721 180845 518755
rect 180793 518690 180845 518721
rect 181791 518755 181843 518800
rect 181791 518721 181801 518755
rect 181835 518721 181843 518755
rect 181791 518690 181843 518721
rect 181897 518755 181949 518800
rect 181897 518721 181905 518755
rect 181939 518721 181949 518755
rect 181897 518690 181949 518721
rect 182343 518755 182395 518800
rect 182343 518721 182353 518755
rect 182387 518721 182395 518755
rect 182343 518690 182395 518721
rect 182633 518755 182685 518800
rect 182633 518721 182641 518755
rect 182675 518721 182685 518755
rect 182633 518690 182685 518721
rect 183631 518755 183683 518800
rect 183631 518721 183641 518755
rect 183675 518721 183683 518755
rect 183631 518690 183683 518721
rect 183737 518755 183789 518800
rect 183737 518721 183745 518755
rect 183779 518721 183789 518755
rect 183737 518690 183789 518721
rect 184735 518755 184787 518800
rect 184735 518721 184745 518755
rect 184779 518721 184787 518755
rect 184735 518690 184787 518721
rect 184841 518755 184893 518800
rect 184841 518721 184849 518755
rect 184883 518721 184893 518755
rect 184841 518690 184893 518721
rect 185839 518755 185891 518800
rect 185839 518721 185849 518755
rect 185883 518721 185891 518755
rect 185839 518690 185891 518721
rect 185945 518755 185997 518800
rect 185945 518721 185953 518755
rect 185987 518721 185997 518755
rect 185945 518690 185997 518721
rect 186943 518755 186995 518800
rect 186943 518721 186953 518755
rect 186987 518721 186995 518755
rect 186943 518690 186995 518721
rect 187233 518757 187285 518800
rect 187233 518723 187241 518757
rect 187275 518723 187285 518757
rect 187233 518690 187285 518723
rect 187403 518757 187455 518800
rect 187403 518723 187413 518757
rect 187447 518723 187455 518757
rect 187403 518690 187455 518723
rect 172237 518563 172289 518596
rect 172237 518529 172245 518563
rect 172279 518529 172289 518563
rect 172237 518486 172289 518529
rect 172407 518563 172459 518596
rect 172407 518529 172417 518563
rect 172451 518529 172459 518563
rect 172407 518486 172459 518529
rect 172513 518565 172565 518596
rect 172513 518531 172521 518565
rect 172555 518531 172565 518565
rect 172513 518486 172565 518531
rect 173511 518565 173563 518596
rect 173511 518531 173521 518565
rect 173555 518531 173563 518565
rect 173511 518486 173563 518531
rect 173617 518565 173669 518596
rect 173617 518531 173625 518565
rect 173659 518531 173669 518565
rect 173617 518486 173669 518531
rect 174615 518565 174667 518596
rect 174615 518531 174625 518565
rect 174659 518531 174667 518565
rect 174615 518486 174667 518531
rect 174905 518565 174957 518596
rect 174905 518531 174913 518565
rect 174947 518531 174957 518565
rect 174905 518486 174957 518531
rect 175903 518565 175955 518596
rect 175903 518531 175913 518565
rect 175947 518531 175955 518565
rect 175903 518486 175955 518531
rect 176009 518565 176061 518596
rect 176009 518531 176017 518565
rect 176051 518531 176061 518565
rect 176009 518486 176061 518531
rect 177007 518565 177059 518596
rect 177007 518531 177017 518565
rect 177051 518531 177059 518565
rect 177007 518486 177059 518531
rect 177113 518565 177165 518596
rect 177113 518531 177121 518565
rect 177155 518531 177165 518565
rect 177113 518486 177165 518531
rect 178111 518565 178163 518596
rect 178111 518531 178121 518565
rect 178155 518531 178163 518565
rect 178111 518486 178163 518531
rect 178217 518565 178269 518596
rect 178217 518531 178225 518565
rect 178259 518531 178269 518565
rect 178217 518486 178269 518531
rect 179215 518565 179267 518596
rect 179215 518531 179225 518565
rect 179259 518531 179267 518565
rect 179215 518486 179267 518531
rect 179321 518565 179373 518596
rect 179321 518531 179329 518565
rect 179363 518531 179373 518565
rect 179321 518486 179373 518531
rect 179767 518565 179819 518596
rect 179767 518531 179777 518565
rect 179811 518531 179819 518565
rect 179767 518486 179819 518531
rect 180057 518565 180109 518596
rect 180057 518531 180065 518565
rect 180099 518531 180109 518565
rect 180057 518486 180109 518531
rect 181055 518565 181107 518596
rect 181055 518531 181065 518565
rect 181099 518531 181107 518565
rect 181055 518486 181107 518531
rect 181161 518565 181213 518596
rect 181161 518531 181169 518565
rect 181203 518531 181213 518565
rect 181161 518486 181213 518531
rect 182159 518565 182211 518596
rect 182159 518531 182169 518565
rect 182203 518531 182211 518565
rect 182159 518486 182211 518531
rect 182265 518565 182317 518596
rect 182265 518531 182273 518565
rect 182307 518531 182317 518565
rect 182265 518486 182317 518531
rect 183263 518565 183315 518596
rect 183263 518531 183273 518565
rect 183307 518531 183315 518565
rect 183263 518486 183315 518531
rect 183369 518565 183421 518596
rect 183369 518531 183377 518565
rect 183411 518531 183421 518565
rect 183369 518486 183421 518531
rect 184367 518565 184419 518596
rect 184367 518531 184377 518565
rect 184411 518531 184419 518565
rect 184367 518486 184419 518531
rect 184473 518565 184525 518596
rect 184473 518531 184481 518565
rect 184515 518531 184525 518565
rect 184473 518486 184525 518531
rect 184919 518565 184971 518596
rect 184919 518531 184929 518565
rect 184963 518531 184971 518565
rect 184919 518486 184971 518531
rect 185209 518565 185261 518596
rect 185209 518531 185217 518565
rect 185251 518531 185261 518565
rect 185209 518486 185261 518531
rect 186207 518565 186259 518596
rect 186207 518531 186217 518565
rect 186251 518531 186259 518565
rect 186207 518486 186259 518531
rect 186313 518565 186365 518596
rect 186313 518531 186321 518565
rect 186355 518531 186365 518565
rect 186313 518486 186365 518531
rect 186943 518565 186995 518596
rect 186943 518531 186953 518565
rect 186987 518531 186995 518565
rect 186943 518486 186995 518531
rect 187233 518563 187285 518596
rect 187233 518529 187241 518563
rect 187275 518529 187285 518563
rect 187233 518486 187285 518529
rect 187403 518563 187455 518596
rect 187403 518529 187413 518563
rect 187447 518529 187455 518563
rect 187403 518486 187455 518529
rect 172237 517669 172289 517712
rect 172237 517635 172245 517669
rect 172279 517635 172289 517669
rect 172237 517602 172289 517635
rect 172407 517669 172459 517712
rect 172407 517635 172417 517669
rect 172451 517635 172459 517669
rect 172407 517602 172459 517635
rect 172513 517667 172565 517712
rect 172513 517633 172521 517667
rect 172555 517633 172565 517667
rect 172513 517602 172565 517633
rect 173511 517667 173563 517712
rect 173511 517633 173521 517667
rect 173555 517633 173563 517667
rect 173511 517602 173563 517633
rect 173617 517667 173669 517712
rect 173617 517633 173625 517667
rect 173659 517633 173669 517667
rect 173617 517602 173669 517633
rect 174615 517667 174667 517712
rect 174615 517633 174625 517667
rect 174659 517633 174667 517667
rect 174615 517602 174667 517633
rect 174721 517667 174773 517712
rect 174721 517633 174729 517667
rect 174763 517633 174773 517667
rect 174721 517602 174773 517633
rect 175719 517667 175771 517712
rect 175719 517633 175729 517667
rect 175763 517633 175771 517667
rect 175719 517602 175771 517633
rect 175825 517667 175877 517712
rect 175825 517633 175833 517667
rect 175867 517633 175877 517667
rect 175825 517602 175877 517633
rect 176823 517667 176875 517712
rect 176823 517633 176833 517667
rect 176867 517633 176875 517667
rect 176823 517602 176875 517633
rect 176929 517674 176981 517712
rect 176929 517640 176937 517674
rect 176971 517640 176981 517674
rect 176929 517602 176981 517640
rect 177191 517674 177243 517712
rect 177191 517640 177201 517674
rect 177235 517640 177243 517674
rect 177191 517602 177243 517640
rect 177481 517667 177533 517712
rect 177481 517633 177489 517667
rect 177523 517633 177533 517667
rect 177481 517602 177533 517633
rect 178479 517667 178531 517712
rect 178479 517633 178489 517667
rect 178523 517633 178531 517667
rect 178479 517602 178531 517633
rect 178585 517667 178637 517712
rect 178585 517633 178593 517667
rect 178627 517633 178637 517667
rect 178585 517602 178637 517633
rect 179583 517667 179635 517712
rect 179583 517633 179593 517667
rect 179627 517633 179635 517667
rect 179583 517602 179635 517633
rect 179689 517667 179741 517712
rect 179689 517633 179697 517667
rect 179731 517633 179741 517667
rect 179689 517602 179741 517633
rect 180687 517667 180739 517712
rect 180687 517633 180697 517667
rect 180731 517633 180739 517667
rect 180687 517602 180739 517633
rect 180793 517667 180845 517712
rect 180793 517633 180801 517667
rect 180835 517633 180845 517667
rect 180793 517602 180845 517633
rect 181791 517667 181843 517712
rect 181791 517633 181801 517667
rect 181835 517633 181843 517667
rect 181791 517602 181843 517633
rect 181897 517667 181949 517712
rect 181897 517633 181905 517667
rect 181939 517633 181949 517667
rect 181897 517602 181949 517633
rect 182343 517667 182395 517712
rect 182343 517633 182353 517667
rect 182387 517633 182395 517667
rect 182343 517602 182395 517633
rect 182633 517667 182685 517712
rect 182633 517633 182641 517667
rect 182675 517633 182685 517667
rect 182633 517602 182685 517633
rect 183631 517667 183683 517712
rect 183631 517633 183641 517667
rect 183675 517633 183683 517667
rect 183631 517602 183683 517633
rect 183737 517667 183789 517712
rect 183737 517633 183745 517667
rect 183779 517633 183789 517667
rect 183737 517602 183789 517633
rect 184735 517667 184787 517712
rect 184735 517633 184745 517667
rect 184779 517633 184787 517667
rect 184735 517602 184787 517633
rect 184841 517667 184893 517712
rect 184841 517633 184849 517667
rect 184883 517633 184893 517667
rect 184841 517602 184893 517633
rect 185839 517667 185891 517712
rect 185839 517633 185849 517667
rect 185883 517633 185891 517667
rect 185839 517602 185891 517633
rect 185945 517667 185997 517712
rect 185945 517633 185953 517667
rect 185987 517633 185997 517667
rect 185945 517602 185997 517633
rect 186943 517667 186995 517712
rect 186943 517633 186953 517667
rect 186987 517633 186995 517667
rect 186943 517602 186995 517633
rect 187233 517669 187285 517712
rect 187233 517635 187241 517669
rect 187275 517635 187285 517669
rect 187233 517602 187285 517635
rect 187403 517669 187455 517712
rect 187403 517635 187413 517669
rect 187447 517635 187455 517669
rect 187403 517602 187455 517635
rect 172237 517475 172289 517508
rect 172237 517441 172245 517475
rect 172279 517441 172289 517475
rect 172237 517398 172289 517441
rect 172407 517475 172459 517508
rect 172407 517441 172417 517475
rect 172451 517441 172459 517475
rect 172407 517398 172459 517441
rect 172513 517477 172565 517508
rect 172513 517443 172521 517477
rect 172555 517443 172565 517477
rect 172513 517398 172565 517443
rect 173511 517477 173563 517508
rect 173511 517443 173521 517477
rect 173555 517443 173563 517477
rect 173511 517398 173563 517443
rect 173617 517477 173669 517508
rect 173617 517443 173625 517477
rect 173659 517443 173669 517477
rect 173617 517398 173669 517443
rect 174615 517477 174667 517508
rect 174615 517443 174625 517477
rect 174659 517443 174667 517477
rect 174615 517398 174667 517443
rect 174905 517477 174957 517508
rect 174905 517443 174913 517477
rect 174947 517443 174957 517477
rect 174905 517398 174957 517443
rect 175903 517477 175955 517508
rect 175903 517443 175913 517477
rect 175947 517443 175955 517477
rect 175903 517398 175955 517443
rect 176009 517477 176061 517508
rect 176009 517443 176017 517477
rect 176051 517443 176061 517477
rect 176009 517398 176061 517443
rect 177007 517477 177059 517508
rect 177007 517443 177017 517477
rect 177051 517443 177059 517477
rect 177007 517398 177059 517443
rect 177113 517477 177165 517508
rect 177113 517443 177121 517477
rect 177155 517443 177165 517477
rect 177113 517398 177165 517443
rect 178111 517477 178163 517508
rect 178111 517443 178121 517477
rect 178155 517443 178163 517477
rect 178111 517398 178163 517443
rect 178217 517477 178269 517508
rect 178217 517443 178225 517477
rect 178259 517443 178269 517477
rect 178217 517398 178269 517443
rect 179215 517477 179267 517508
rect 179215 517443 179225 517477
rect 179259 517443 179267 517477
rect 179215 517398 179267 517443
rect 179321 517477 179373 517508
rect 179321 517443 179329 517477
rect 179363 517443 179373 517477
rect 179321 517398 179373 517443
rect 179767 517477 179819 517508
rect 179767 517443 179777 517477
rect 179811 517443 179819 517477
rect 179767 517398 179819 517443
rect 180057 517477 180109 517508
rect 180057 517443 180065 517477
rect 180099 517443 180109 517477
rect 180057 517398 180109 517443
rect 181055 517477 181107 517508
rect 181055 517443 181065 517477
rect 181099 517443 181107 517477
rect 181055 517398 181107 517443
rect 181161 517477 181213 517508
rect 181161 517443 181169 517477
rect 181203 517443 181213 517477
rect 181161 517398 181213 517443
rect 182159 517477 182211 517508
rect 182159 517443 182169 517477
rect 182203 517443 182211 517477
rect 182159 517398 182211 517443
rect 182265 517477 182317 517508
rect 182265 517443 182273 517477
rect 182307 517443 182317 517477
rect 182265 517398 182317 517443
rect 183263 517477 183315 517508
rect 183263 517443 183273 517477
rect 183307 517443 183315 517477
rect 183263 517398 183315 517443
rect 183369 517477 183421 517508
rect 183369 517443 183377 517477
rect 183411 517443 183421 517477
rect 183369 517398 183421 517443
rect 184367 517477 184419 517508
rect 184367 517443 184377 517477
rect 184411 517443 184419 517477
rect 184367 517398 184419 517443
rect 184473 517477 184525 517508
rect 184473 517443 184481 517477
rect 184515 517443 184525 517477
rect 184473 517398 184525 517443
rect 184919 517477 184971 517508
rect 184919 517443 184929 517477
rect 184963 517443 184971 517477
rect 184919 517398 184971 517443
rect 185209 517477 185261 517508
rect 185209 517443 185217 517477
rect 185251 517443 185261 517477
rect 185209 517398 185261 517443
rect 186207 517477 186259 517508
rect 186207 517443 186217 517477
rect 186251 517443 186259 517477
rect 186207 517398 186259 517443
rect 186313 517477 186365 517508
rect 186313 517443 186321 517477
rect 186355 517443 186365 517477
rect 186313 517398 186365 517443
rect 186943 517477 186995 517508
rect 186943 517443 186953 517477
rect 186987 517443 186995 517477
rect 186943 517398 186995 517443
rect 187233 517475 187285 517508
rect 187233 517441 187241 517475
rect 187275 517441 187285 517475
rect 187233 517398 187285 517441
rect 187403 517475 187455 517508
rect 187403 517441 187413 517475
rect 187447 517441 187455 517475
rect 187403 517398 187455 517441
rect 172237 516581 172289 516624
rect 172237 516547 172245 516581
rect 172279 516547 172289 516581
rect 172237 516514 172289 516547
rect 172407 516581 172459 516624
rect 172407 516547 172417 516581
rect 172451 516547 172459 516581
rect 172407 516514 172459 516547
rect 172513 516579 172565 516624
rect 172513 516545 172521 516579
rect 172555 516545 172565 516579
rect 172513 516514 172565 516545
rect 173511 516579 173563 516624
rect 173511 516545 173521 516579
rect 173555 516545 173563 516579
rect 173511 516514 173563 516545
rect 173617 516579 173669 516624
rect 173617 516545 173625 516579
rect 173659 516545 173669 516579
rect 173617 516514 173669 516545
rect 174615 516579 174667 516624
rect 174615 516545 174625 516579
rect 174659 516545 174667 516579
rect 174615 516514 174667 516545
rect 174721 516579 174773 516624
rect 174721 516545 174729 516579
rect 174763 516545 174773 516579
rect 174721 516514 174773 516545
rect 175719 516579 175771 516624
rect 175719 516545 175729 516579
rect 175763 516545 175771 516579
rect 175719 516514 175771 516545
rect 175825 516579 175877 516624
rect 175825 516545 175833 516579
rect 175867 516545 175877 516579
rect 175825 516514 175877 516545
rect 176823 516579 176875 516624
rect 176823 516545 176833 516579
rect 176867 516545 176875 516579
rect 176823 516514 176875 516545
rect 176929 516586 176981 516624
rect 176929 516552 176937 516586
rect 176971 516552 176981 516586
rect 176929 516514 176981 516552
rect 177191 516586 177243 516624
rect 177191 516552 177201 516586
rect 177235 516552 177243 516586
rect 177191 516514 177243 516552
rect 177481 516579 177533 516624
rect 177481 516545 177489 516579
rect 177523 516545 177533 516579
rect 177481 516514 177533 516545
rect 178479 516579 178531 516624
rect 178479 516545 178489 516579
rect 178523 516545 178531 516579
rect 178479 516514 178531 516545
rect 178585 516579 178637 516624
rect 178585 516545 178593 516579
rect 178627 516545 178637 516579
rect 178585 516514 178637 516545
rect 179583 516579 179635 516624
rect 179583 516545 179593 516579
rect 179627 516545 179635 516579
rect 179583 516514 179635 516545
rect 179689 516579 179741 516624
rect 179689 516545 179697 516579
rect 179731 516545 179741 516579
rect 179689 516514 179741 516545
rect 180687 516579 180739 516624
rect 180687 516545 180697 516579
rect 180731 516545 180739 516579
rect 180687 516514 180739 516545
rect 180793 516579 180845 516624
rect 180793 516545 180801 516579
rect 180835 516545 180845 516579
rect 180793 516514 180845 516545
rect 181791 516579 181843 516624
rect 181791 516545 181801 516579
rect 181835 516545 181843 516579
rect 181791 516514 181843 516545
rect 181897 516579 181949 516624
rect 181897 516545 181905 516579
rect 181939 516545 181949 516579
rect 181897 516514 181949 516545
rect 182343 516579 182395 516624
rect 182343 516545 182353 516579
rect 182387 516545 182395 516579
rect 182343 516514 182395 516545
rect 182633 516579 182685 516624
rect 182633 516545 182641 516579
rect 182675 516545 182685 516579
rect 182633 516514 182685 516545
rect 183631 516579 183683 516624
rect 183631 516545 183641 516579
rect 183675 516545 183683 516579
rect 183631 516514 183683 516545
rect 183737 516579 183789 516624
rect 183737 516545 183745 516579
rect 183779 516545 183789 516579
rect 183737 516514 183789 516545
rect 184735 516579 184787 516624
rect 184735 516545 184745 516579
rect 184779 516545 184787 516579
rect 184735 516514 184787 516545
rect 184841 516579 184893 516624
rect 184841 516545 184849 516579
rect 184883 516545 184893 516579
rect 184841 516514 184893 516545
rect 185839 516579 185891 516624
rect 185839 516545 185849 516579
rect 185883 516545 185891 516579
rect 185839 516514 185891 516545
rect 185945 516579 185997 516624
rect 185945 516545 185953 516579
rect 185987 516545 185997 516579
rect 185945 516514 185997 516545
rect 186943 516579 186995 516624
rect 186943 516545 186953 516579
rect 186987 516545 186995 516579
rect 186943 516514 186995 516545
rect 187233 516581 187285 516624
rect 187233 516547 187241 516581
rect 187275 516547 187285 516581
rect 187233 516514 187285 516547
rect 187403 516581 187455 516624
rect 187403 516547 187413 516581
rect 187447 516547 187455 516581
rect 187403 516514 187455 516547
rect 172237 516387 172289 516420
rect 172237 516353 172245 516387
rect 172279 516353 172289 516387
rect 172237 516310 172289 516353
rect 172407 516387 172459 516420
rect 172407 516353 172417 516387
rect 172451 516353 172459 516387
rect 172407 516310 172459 516353
rect 172513 516389 172565 516420
rect 172513 516355 172521 516389
rect 172555 516355 172565 516389
rect 172513 516310 172565 516355
rect 173511 516389 173563 516420
rect 173511 516355 173521 516389
rect 173555 516355 173563 516389
rect 173511 516310 173563 516355
rect 173617 516389 173669 516420
rect 173617 516355 173625 516389
rect 173659 516355 173669 516389
rect 173617 516310 173669 516355
rect 174615 516389 174667 516420
rect 174615 516355 174625 516389
rect 174659 516355 174667 516389
rect 174615 516310 174667 516355
rect 174905 516389 174957 516420
rect 174905 516355 174913 516389
rect 174947 516355 174957 516389
rect 174905 516310 174957 516355
rect 175903 516389 175955 516420
rect 175903 516355 175913 516389
rect 175947 516355 175955 516389
rect 175903 516310 175955 516355
rect 176009 516389 176061 516420
rect 176009 516355 176017 516389
rect 176051 516355 176061 516389
rect 176009 516310 176061 516355
rect 177007 516389 177059 516420
rect 177007 516355 177017 516389
rect 177051 516355 177059 516389
rect 177007 516310 177059 516355
rect 177113 516389 177165 516420
rect 177113 516355 177121 516389
rect 177155 516355 177165 516389
rect 177113 516310 177165 516355
rect 178111 516389 178163 516420
rect 178111 516355 178121 516389
rect 178155 516355 178163 516389
rect 178111 516310 178163 516355
rect 178217 516389 178269 516420
rect 178217 516355 178225 516389
rect 178259 516355 178269 516389
rect 178217 516310 178269 516355
rect 179215 516389 179267 516420
rect 179215 516355 179225 516389
rect 179259 516355 179267 516389
rect 179215 516310 179267 516355
rect 179321 516389 179373 516420
rect 179321 516355 179329 516389
rect 179363 516355 179373 516389
rect 179321 516310 179373 516355
rect 179767 516389 179819 516420
rect 179767 516355 179777 516389
rect 179811 516355 179819 516389
rect 179767 516310 179819 516355
rect 180057 516389 180109 516420
rect 180057 516355 180065 516389
rect 180099 516355 180109 516389
rect 180057 516310 180109 516355
rect 181055 516389 181107 516420
rect 181055 516355 181065 516389
rect 181099 516355 181107 516389
rect 181055 516310 181107 516355
rect 181161 516389 181213 516420
rect 181161 516355 181169 516389
rect 181203 516355 181213 516389
rect 181161 516310 181213 516355
rect 182159 516389 182211 516420
rect 182159 516355 182169 516389
rect 182203 516355 182211 516389
rect 182159 516310 182211 516355
rect 182265 516389 182317 516420
rect 182265 516355 182273 516389
rect 182307 516355 182317 516389
rect 182265 516310 182317 516355
rect 183263 516389 183315 516420
rect 183263 516355 183273 516389
rect 183307 516355 183315 516389
rect 183263 516310 183315 516355
rect 183369 516389 183421 516420
rect 183369 516355 183377 516389
rect 183411 516355 183421 516389
rect 183369 516310 183421 516355
rect 184367 516389 184419 516420
rect 184367 516355 184377 516389
rect 184411 516355 184419 516389
rect 184367 516310 184419 516355
rect 184473 516389 184525 516420
rect 184473 516355 184481 516389
rect 184515 516355 184525 516389
rect 184473 516310 184525 516355
rect 184919 516389 184971 516420
rect 184919 516355 184929 516389
rect 184963 516355 184971 516389
rect 184919 516310 184971 516355
rect 185209 516389 185261 516420
rect 185209 516355 185217 516389
rect 185251 516355 185261 516389
rect 185209 516310 185261 516355
rect 186207 516389 186259 516420
rect 186207 516355 186217 516389
rect 186251 516355 186259 516389
rect 186207 516310 186259 516355
rect 186313 516389 186365 516420
rect 186313 516355 186321 516389
rect 186355 516355 186365 516389
rect 186313 516310 186365 516355
rect 186943 516389 186995 516420
rect 186943 516355 186953 516389
rect 186987 516355 186995 516389
rect 186943 516310 186995 516355
rect 187233 516387 187285 516420
rect 187233 516353 187241 516387
rect 187275 516353 187285 516387
rect 187233 516310 187285 516353
rect 187403 516387 187455 516420
rect 187403 516353 187413 516387
rect 187447 516353 187455 516387
rect 187403 516310 187455 516353
rect 172237 515493 172289 515536
rect 172237 515459 172245 515493
rect 172279 515459 172289 515493
rect 172237 515426 172289 515459
rect 172407 515493 172459 515536
rect 172407 515459 172417 515493
rect 172451 515459 172459 515493
rect 172407 515426 172459 515459
rect 172513 515491 172565 515536
rect 172513 515457 172521 515491
rect 172555 515457 172565 515491
rect 172513 515426 172565 515457
rect 173143 515491 173195 515536
rect 173143 515457 173153 515491
rect 173187 515457 173195 515491
rect 173143 515426 173195 515457
rect 173433 515480 173486 515510
rect 173433 515446 173441 515480
rect 173475 515446 173486 515480
rect 173433 515426 173486 515446
rect 173516 515476 173583 515510
rect 173516 515442 173527 515476
rect 173561 515442 173583 515476
rect 173516 515426 173583 515442
rect 173613 515498 173669 515510
rect 173613 515464 173624 515498
rect 173658 515464 173669 515498
rect 173613 515426 173669 515464
rect 173699 515476 173755 515510
rect 173699 515442 173710 515476
rect 173744 515442 173755 515476
rect 173699 515426 173755 515442
rect 173785 515498 173841 515510
rect 173785 515464 173796 515498
rect 173830 515464 173841 515498
rect 173785 515426 173841 515464
rect 173871 515476 173929 515510
rect 173871 515442 173882 515476
rect 173916 515442 173929 515476
rect 173871 515426 173929 515442
rect 173985 515491 174037 515536
rect 173985 515457 173993 515491
rect 174027 515457 174037 515491
rect 173985 515426 174037 515457
rect 174615 515491 174667 515536
rect 174615 515457 174625 515491
rect 174659 515457 174667 515491
rect 174615 515426 174667 515457
rect 174905 515491 174957 515536
rect 174905 515457 174913 515491
rect 174947 515457 174957 515491
rect 174905 515426 174957 515457
rect 175903 515491 175955 515536
rect 175903 515457 175913 515491
rect 175947 515457 175955 515491
rect 175903 515426 175955 515457
rect 176009 515491 176061 515536
rect 176009 515457 176017 515491
rect 176051 515457 176061 515491
rect 176009 515426 176061 515457
rect 177007 515491 177059 515536
rect 177007 515457 177017 515491
rect 177051 515457 177059 515491
rect 177007 515426 177059 515457
rect 177113 515493 177165 515536
rect 177113 515459 177121 515493
rect 177155 515459 177165 515493
rect 177113 515426 177165 515459
rect 177283 515493 177335 515536
rect 177283 515459 177293 515493
rect 177327 515459 177335 515493
rect 177283 515426 177335 515459
rect 177481 515491 177533 515536
rect 177481 515457 177489 515491
rect 177523 515457 177533 515491
rect 177481 515426 177533 515457
rect 178479 515491 178531 515536
rect 178479 515457 178489 515491
rect 178523 515457 178531 515491
rect 178479 515426 178531 515457
rect 178585 515491 178637 515536
rect 178585 515457 178593 515491
rect 178627 515457 178637 515491
rect 178585 515426 178637 515457
rect 179583 515491 179635 515536
rect 179583 515457 179593 515491
rect 179627 515457 179635 515491
rect 179583 515426 179635 515457
rect 179689 515493 179741 515536
rect 179689 515459 179697 515493
rect 179731 515459 179741 515493
rect 179689 515426 179741 515459
rect 179859 515493 179911 515536
rect 179859 515459 179869 515493
rect 179903 515459 179911 515493
rect 179859 515426 179911 515459
rect 180057 515491 180109 515536
rect 180057 515457 180065 515491
rect 180099 515457 180109 515491
rect 180057 515426 180109 515457
rect 181055 515491 181107 515536
rect 181055 515457 181065 515491
rect 181099 515457 181107 515491
rect 181055 515426 181107 515457
rect 181161 515491 181213 515536
rect 181161 515457 181169 515491
rect 181203 515457 181213 515491
rect 181161 515426 181213 515457
rect 181791 515491 181843 515536
rect 181791 515457 181801 515491
rect 181835 515457 181843 515491
rect 181791 515426 181843 515457
rect 182081 515502 182133 515530
rect 182081 515468 182089 515502
rect 182123 515468 182133 515502
rect 182081 515426 182133 515468
rect 182163 515472 182221 515530
rect 182163 515438 182175 515472
rect 182209 515438 182221 515472
rect 182163 515426 182221 515438
rect 182251 515485 182303 515530
rect 182251 515451 182261 515485
rect 182295 515451 182303 515485
rect 182251 515426 182303 515451
rect 182633 515491 182685 515536
rect 182633 515457 182641 515491
rect 182675 515457 182685 515491
rect 182633 515426 182685 515457
rect 183631 515491 183683 515536
rect 183631 515457 183641 515491
rect 183675 515457 183683 515491
rect 183631 515426 183683 515457
rect 183737 515491 183789 515536
rect 183737 515457 183745 515491
rect 183779 515457 183789 515491
rect 183737 515426 183789 515457
rect 184735 515491 184787 515536
rect 184735 515457 184745 515491
rect 184779 515457 184787 515491
rect 184735 515426 184787 515457
rect 184841 515493 184893 515536
rect 184841 515459 184849 515493
rect 184883 515459 184893 515493
rect 184841 515426 184893 515459
rect 185011 515493 185063 515536
rect 185011 515459 185021 515493
rect 185055 515459 185063 515493
rect 185011 515426 185063 515459
rect 185209 515491 185261 515536
rect 185209 515457 185217 515491
rect 185251 515457 185261 515491
rect 185209 515426 185261 515457
rect 186207 515491 186259 515536
rect 186207 515457 186217 515491
rect 186251 515457 186259 515491
rect 186207 515426 186259 515457
rect 186405 515480 186458 515510
rect 186405 515446 186413 515480
rect 186447 515446 186458 515480
rect 186405 515426 186458 515446
rect 186488 515476 186555 515510
rect 186488 515442 186499 515476
rect 186533 515442 186555 515476
rect 186488 515426 186555 515442
rect 186585 515498 186641 515510
rect 186585 515464 186596 515498
rect 186630 515464 186641 515498
rect 186585 515426 186641 515464
rect 186671 515476 186727 515510
rect 186671 515442 186682 515476
rect 186716 515442 186727 515476
rect 186671 515426 186727 515442
rect 186757 515498 186813 515510
rect 186757 515464 186768 515498
rect 186802 515464 186813 515498
rect 186757 515426 186813 515464
rect 186843 515476 186901 515510
rect 186843 515442 186854 515476
rect 186888 515442 186901 515476
rect 186843 515426 186901 515442
rect 186957 515493 187009 515536
rect 186957 515459 186965 515493
rect 186999 515459 187009 515493
rect 186957 515426 187009 515459
rect 187127 515493 187179 515536
rect 187127 515459 187137 515493
rect 187171 515459 187179 515493
rect 187127 515426 187179 515459
rect 187233 515493 187285 515536
rect 187233 515459 187241 515493
rect 187275 515459 187285 515493
rect 187233 515426 187285 515459
rect 187403 515493 187455 515536
rect 187403 515459 187413 515493
rect 187447 515459 187455 515493
rect 187403 515426 187455 515459
<< pdiff >>
rect 164658 539545 164716 539557
rect 164658 538569 164670 539545
rect 164704 538569 164716 539545
rect 164658 538557 164716 538569
rect 164746 539545 164804 539557
rect 164746 538569 164758 539545
rect 164792 538569 164804 539545
rect 164746 538557 164804 538569
rect 164881 539552 164943 539564
rect 164881 538576 164893 539552
rect 164927 538576 164943 539552
rect 164881 538564 164943 538576
rect 164973 539552 165039 539564
rect 164973 538576 164989 539552
rect 165023 538576 165039 539552
rect 164973 538564 165039 538576
rect 165069 539552 165135 539564
rect 165069 538576 165085 539552
rect 165119 538576 165135 539552
rect 165069 538564 165135 538576
rect 165165 539552 165231 539564
rect 165165 538576 165181 539552
rect 165215 538576 165231 539552
rect 165165 538564 165231 538576
rect 165261 539552 165327 539564
rect 165261 538576 165277 539552
rect 165311 538576 165327 539552
rect 165261 538564 165327 538576
rect 165357 539552 165423 539564
rect 165357 538576 165373 539552
rect 165407 538576 165423 539552
rect 165357 538564 165423 538576
rect 165453 539552 165519 539564
rect 165453 538576 165469 539552
rect 165503 538576 165519 539552
rect 165453 538564 165519 538576
rect 165549 539552 165615 539564
rect 165549 538576 165565 539552
rect 165599 538576 165615 539552
rect 165549 538564 165615 538576
rect 165645 539552 165711 539564
rect 165645 538576 165661 539552
rect 165695 538576 165711 539552
rect 165645 538564 165711 538576
rect 165741 539552 165807 539564
rect 165741 538576 165757 539552
rect 165791 538576 165807 539552
rect 165741 538564 165807 538576
rect 165837 539552 165903 539564
rect 165837 538576 165853 539552
rect 165887 538576 165903 539552
rect 165837 538564 165903 538576
rect 165933 539552 165999 539564
rect 165933 538576 165949 539552
rect 165983 538576 165999 539552
rect 165933 538564 165999 538576
rect 166029 539552 166091 539564
rect 166029 538576 166045 539552
rect 166079 538576 166091 539552
rect 166158 539545 166216 539557
rect 166158 538969 166170 539545
rect 166204 538969 166216 539545
rect 166158 538957 166216 538969
rect 166246 539545 166304 539557
rect 166246 538969 166258 539545
rect 166292 538969 166304 539545
rect 166246 538957 166304 538969
rect 166358 539545 166416 539557
rect 166029 538564 166091 538576
rect 166358 538569 166370 539545
rect 166404 538569 166416 539545
rect 166358 538557 166416 538569
rect 166446 539545 166504 539557
rect 166446 538569 166458 539545
rect 166492 538569 166504 539545
rect 166446 538557 166504 538569
rect 168458 539545 168516 539557
rect 168458 538569 168470 539545
rect 168504 538569 168516 539545
rect 168458 538557 168516 538569
rect 168546 539545 168604 539557
rect 168546 538569 168558 539545
rect 168592 538569 168604 539545
rect 168546 538557 168604 538569
rect 168681 539552 168743 539564
rect 168681 538576 168693 539552
rect 168727 538576 168743 539552
rect 168681 538564 168743 538576
rect 168773 539552 168839 539564
rect 168773 538576 168789 539552
rect 168823 538576 168839 539552
rect 168773 538564 168839 538576
rect 168869 539552 168935 539564
rect 168869 538576 168885 539552
rect 168919 538576 168935 539552
rect 168869 538564 168935 538576
rect 168965 539552 169031 539564
rect 168965 538576 168981 539552
rect 169015 538576 169031 539552
rect 168965 538564 169031 538576
rect 169061 539552 169127 539564
rect 169061 538576 169077 539552
rect 169111 538576 169127 539552
rect 169061 538564 169127 538576
rect 169157 539552 169223 539564
rect 169157 538576 169173 539552
rect 169207 538576 169223 539552
rect 169157 538564 169223 538576
rect 169253 539552 169319 539564
rect 169253 538576 169269 539552
rect 169303 538576 169319 539552
rect 169253 538564 169319 538576
rect 169349 539552 169415 539564
rect 169349 538576 169365 539552
rect 169399 538576 169415 539552
rect 169349 538564 169415 538576
rect 169445 539552 169511 539564
rect 169445 538576 169461 539552
rect 169495 538576 169511 539552
rect 169445 538564 169511 538576
rect 169541 539552 169607 539564
rect 169541 538576 169557 539552
rect 169591 538576 169607 539552
rect 169541 538564 169607 538576
rect 169637 539552 169703 539564
rect 169637 538576 169653 539552
rect 169687 538576 169703 539552
rect 169637 538564 169703 538576
rect 169733 539552 169799 539564
rect 169733 538576 169749 539552
rect 169783 538576 169799 539552
rect 169733 538564 169799 538576
rect 169829 539552 169891 539564
rect 169829 538576 169845 539552
rect 169879 538576 169891 539552
rect 169958 539545 170016 539557
rect 169958 538969 169970 539545
rect 170004 538969 170016 539545
rect 169958 538957 170016 538969
rect 170046 539545 170104 539557
rect 170046 538969 170058 539545
rect 170092 538969 170104 539545
rect 170046 538957 170104 538969
rect 170158 539545 170216 539557
rect 169829 538564 169891 538576
rect 170158 538569 170170 539545
rect 170204 538569 170216 539545
rect 170158 538557 170216 538569
rect 170246 539545 170304 539557
rect 170246 538569 170258 539545
rect 170292 538569 170304 539545
rect 170246 538557 170304 538569
rect 172158 539545 172216 539557
rect 172158 538569 172170 539545
rect 172204 538569 172216 539545
rect 172158 538557 172216 538569
rect 172246 539545 172304 539557
rect 172246 538569 172258 539545
rect 172292 538569 172304 539545
rect 172246 538557 172304 538569
rect 172381 539552 172443 539564
rect 172381 538576 172393 539552
rect 172427 538576 172443 539552
rect 172381 538564 172443 538576
rect 172473 539552 172539 539564
rect 172473 538576 172489 539552
rect 172523 538576 172539 539552
rect 172473 538564 172539 538576
rect 172569 539552 172635 539564
rect 172569 538576 172585 539552
rect 172619 538576 172635 539552
rect 172569 538564 172635 538576
rect 172665 539552 172731 539564
rect 172665 538576 172681 539552
rect 172715 538576 172731 539552
rect 172665 538564 172731 538576
rect 172761 539552 172827 539564
rect 172761 538576 172777 539552
rect 172811 538576 172827 539552
rect 172761 538564 172827 538576
rect 172857 539552 172923 539564
rect 172857 538576 172873 539552
rect 172907 538576 172923 539552
rect 172857 538564 172923 538576
rect 172953 539552 173019 539564
rect 172953 538576 172969 539552
rect 173003 538576 173019 539552
rect 172953 538564 173019 538576
rect 173049 539552 173115 539564
rect 173049 538576 173065 539552
rect 173099 538576 173115 539552
rect 173049 538564 173115 538576
rect 173145 539552 173211 539564
rect 173145 538576 173161 539552
rect 173195 538576 173211 539552
rect 173145 538564 173211 538576
rect 173241 539552 173307 539564
rect 173241 538576 173257 539552
rect 173291 538576 173307 539552
rect 173241 538564 173307 538576
rect 173337 539552 173403 539564
rect 173337 538576 173353 539552
rect 173387 538576 173403 539552
rect 173337 538564 173403 538576
rect 173433 539552 173499 539564
rect 173433 538576 173449 539552
rect 173483 538576 173499 539552
rect 173433 538564 173499 538576
rect 173529 539552 173591 539564
rect 173529 538576 173545 539552
rect 173579 538576 173591 539552
rect 173658 539545 173716 539557
rect 173658 538969 173670 539545
rect 173704 538969 173716 539545
rect 173658 538957 173716 538969
rect 173746 539545 173804 539557
rect 173746 538969 173758 539545
rect 173792 538969 173804 539545
rect 173746 538957 173804 538969
rect 173858 539545 173916 539557
rect 173529 538564 173591 538576
rect 173858 538569 173870 539545
rect 173904 538569 173916 539545
rect 173858 538557 173916 538569
rect 173946 539545 174004 539557
rect 173946 538569 173958 539545
rect 173992 538569 174004 539545
rect 173946 538557 174004 538569
rect 175658 539545 175716 539557
rect 175658 538569 175670 539545
rect 175704 538569 175716 539545
rect 175658 538557 175716 538569
rect 175746 539545 175804 539557
rect 175746 538569 175758 539545
rect 175792 538569 175804 539545
rect 175746 538557 175804 538569
rect 175881 539552 175943 539564
rect 175881 538576 175893 539552
rect 175927 538576 175943 539552
rect 175881 538564 175943 538576
rect 175973 539552 176039 539564
rect 175973 538576 175989 539552
rect 176023 538576 176039 539552
rect 175973 538564 176039 538576
rect 176069 539552 176135 539564
rect 176069 538576 176085 539552
rect 176119 538576 176135 539552
rect 176069 538564 176135 538576
rect 176165 539552 176231 539564
rect 176165 538576 176181 539552
rect 176215 538576 176231 539552
rect 176165 538564 176231 538576
rect 176261 539552 176327 539564
rect 176261 538576 176277 539552
rect 176311 538576 176327 539552
rect 176261 538564 176327 538576
rect 176357 539552 176423 539564
rect 176357 538576 176373 539552
rect 176407 538576 176423 539552
rect 176357 538564 176423 538576
rect 176453 539552 176519 539564
rect 176453 538576 176469 539552
rect 176503 538576 176519 539552
rect 176453 538564 176519 538576
rect 176549 539552 176615 539564
rect 176549 538576 176565 539552
rect 176599 538576 176615 539552
rect 176549 538564 176615 538576
rect 176645 539552 176711 539564
rect 176645 538576 176661 539552
rect 176695 538576 176711 539552
rect 176645 538564 176711 538576
rect 176741 539552 176807 539564
rect 176741 538576 176757 539552
rect 176791 538576 176807 539552
rect 176741 538564 176807 538576
rect 176837 539552 176903 539564
rect 176837 538576 176853 539552
rect 176887 538576 176903 539552
rect 176837 538564 176903 538576
rect 176933 539552 176999 539564
rect 176933 538576 176949 539552
rect 176983 538576 176999 539552
rect 176933 538564 176999 538576
rect 177029 539552 177091 539564
rect 177029 538576 177045 539552
rect 177079 538576 177091 539552
rect 177158 539545 177216 539557
rect 177158 538969 177170 539545
rect 177204 538969 177216 539545
rect 177158 538957 177216 538969
rect 177246 539545 177304 539557
rect 177246 538969 177258 539545
rect 177292 538969 177304 539545
rect 177246 538957 177304 538969
rect 177358 539545 177416 539557
rect 177029 538564 177091 538576
rect 177358 538569 177370 539545
rect 177404 538569 177416 539545
rect 177358 538557 177416 538569
rect 177446 539545 177504 539557
rect 177446 538569 177458 539545
rect 177492 538569 177504 539545
rect 177446 538557 177504 538569
rect 179258 539545 179316 539557
rect 179258 538569 179270 539545
rect 179304 538569 179316 539545
rect 179258 538557 179316 538569
rect 179346 539545 179404 539557
rect 179346 538569 179358 539545
rect 179392 538569 179404 539545
rect 179346 538557 179404 538569
rect 179481 539552 179543 539564
rect 179481 538576 179493 539552
rect 179527 538576 179543 539552
rect 179481 538564 179543 538576
rect 179573 539552 179639 539564
rect 179573 538576 179589 539552
rect 179623 538576 179639 539552
rect 179573 538564 179639 538576
rect 179669 539552 179735 539564
rect 179669 538576 179685 539552
rect 179719 538576 179735 539552
rect 179669 538564 179735 538576
rect 179765 539552 179831 539564
rect 179765 538576 179781 539552
rect 179815 538576 179831 539552
rect 179765 538564 179831 538576
rect 179861 539552 179927 539564
rect 179861 538576 179877 539552
rect 179911 538576 179927 539552
rect 179861 538564 179927 538576
rect 179957 539552 180023 539564
rect 179957 538576 179973 539552
rect 180007 538576 180023 539552
rect 179957 538564 180023 538576
rect 180053 539552 180119 539564
rect 180053 538576 180069 539552
rect 180103 538576 180119 539552
rect 180053 538564 180119 538576
rect 180149 539552 180215 539564
rect 180149 538576 180165 539552
rect 180199 538576 180215 539552
rect 180149 538564 180215 538576
rect 180245 539552 180311 539564
rect 180245 538576 180261 539552
rect 180295 538576 180311 539552
rect 180245 538564 180311 538576
rect 180341 539552 180407 539564
rect 180341 538576 180357 539552
rect 180391 538576 180407 539552
rect 180341 538564 180407 538576
rect 180437 539552 180503 539564
rect 180437 538576 180453 539552
rect 180487 538576 180503 539552
rect 180437 538564 180503 538576
rect 180533 539552 180599 539564
rect 180533 538576 180549 539552
rect 180583 538576 180599 539552
rect 180533 538564 180599 538576
rect 180629 539552 180691 539564
rect 180629 538576 180645 539552
rect 180679 538576 180691 539552
rect 180758 539545 180816 539557
rect 180758 538969 180770 539545
rect 180804 538969 180816 539545
rect 180758 538957 180816 538969
rect 180846 539545 180904 539557
rect 180846 538969 180858 539545
rect 180892 538969 180904 539545
rect 180846 538957 180904 538969
rect 180958 539545 181016 539557
rect 180629 538564 180691 538576
rect 180958 538569 180970 539545
rect 181004 538569 181016 539545
rect 180958 538557 181016 538569
rect 181046 539545 181104 539557
rect 181046 538569 181058 539545
rect 181092 538569 181104 539545
rect 181046 538557 181104 538569
rect 182558 539545 182616 539557
rect 182558 538569 182570 539545
rect 182604 538569 182616 539545
rect 182558 538557 182616 538569
rect 182646 539545 182704 539557
rect 182646 538569 182658 539545
rect 182692 538569 182704 539545
rect 182646 538557 182704 538569
rect 182781 539552 182843 539564
rect 182781 538576 182793 539552
rect 182827 538576 182843 539552
rect 182781 538564 182843 538576
rect 182873 539552 182939 539564
rect 182873 538576 182889 539552
rect 182923 538576 182939 539552
rect 182873 538564 182939 538576
rect 182969 539552 183035 539564
rect 182969 538576 182985 539552
rect 183019 538576 183035 539552
rect 182969 538564 183035 538576
rect 183065 539552 183131 539564
rect 183065 538576 183081 539552
rect 183115 538576 183131 539552
rect 183065 538564 183131 538576
rect 183161 539552 183227 539564
rect 183161 538576 183177 539552
rect 183211 538576 183227 539552
rect 183161 538564 183227 538576
rect 183257 539552 183323 539564
rect 183257 538576 183273 539552
rect 183307 538576 183323 539552
rect 183257 538564 183323 538576
rect 183353 539552 183419 539564
rect 183353 538576 183369 539552
rect 183403 538576 183419 539552
rect 183353 538564 183419 538576
rect 183449 539552 183515 539564
rect 183449 538576 183465 539552
rect 183499 538576 183515 539552
rect 183449 538564 183515 538576
rect 183545 539552 183611 539564
rect 183545 538576 183561 539552
rect 183595 538576 183611 539552
rect 183545 538564 183611 538576
rect 183641 539552 183707 539564
rect 183641 538576 183657 539552
rect 183691 538576 183707 539552
rect 183641 538564 183707 538576
rect 183737 539552 183803 539564
rect 183737 538576 183753 539552
rect 183787 538576 183803 539552
rect 183737 538564 183803 538576
rect 183833 539552 183899 539564
rect 183833 538576 183849 539552
rect 183883 538576 183899 539552
rect 183833 538564 183899 538576
rect 183929 539552 183991 539564
rect 183929 538576 183945 539552
rect 183979 538576 183991 539552
rect 184058 539545 184116 539557
rect 184058 538969 184070 539545
rect 184104 538969 184116 539545
rect 184058 538957 184116 538969
rect 184146 539545 184204 539557
rect 184146 538969 184158 539545
rect 184192 538969 184204 539545
rect 184146 538957 184204 538969
rect 184258 539545 184316 539557
rect 183929 538564 183991 538576
rect 184258 538569 184270 539545
rect 184304 538569 184316 539545
rect 184258 538557 184316 538569
rect 184346 539545 184404 539557
rect 184346 538569 184358 539545
rect 184392 538569 184404 539545
rect 184346 538557 184404 538569
rect 185858 539545 185916 539557
rect 185858 538569 185870 539545
rect 185904 538569 185916 539545
rect 185858 538557 185916 538569
rect 185946 539545 186004 539557
rect 185946 538569 185958 539545
rect 185992 538569 186004 539545
rect 185946 538557 186004 538569
rect 186081 539552 186143 539564
rect 186081 538576 186093 539552
rect 186127 538576 186143 539552
rect 186081 538564 186143 538576
rect 186173 539552 186239 539564
rect 186173 538576 186189 539552
rect 186223 538576 186239 539552
rect 186173 538564 186239 538576
rect 186269 539552 186335 539564
rect 186269 538576 186285 539552
rect 186319 538576 186335 539552
rect 186269 538564 186335 538576
rect 186365 539552 186431 539564
rect 186365 538576 186381 539552
rect 186415 538576 186431 539552
rect 186365 538564 186431 538576
rect 186461 539552 186527 539564
rect 186461 538576 186477 539552
rect 186511 538576 186527 539552
rect 186461 538564 186527 538576
rect 186557 539552 186623 539564
rect 186557 538576 186573 539552
rect 186607 538576 186623 539552
rect 186557 538564 186623 538576
rect 186653 539552 186719 539564
rect 186653 538576 186669 539552
rect 186703 538576 186719 539552
rect 186653 538564 186719 538576
rect 186749 539552 186815 539564
rect 186749 538576 186765 539552
rect 186799 538576 186815 539552
rect 186749 538564 186815 538576
rect 186845 539552 186911 539564
rect 186845 538576 186861 539552
rect 186895 538576 186911 539552
rect 186845 538564 186911 538576
rect 186941 539552 187007 539564
rect 186941 538576 186957 539552
rect 186991 538576 187007 539552
rect 186941 538564 187007 538576
rect 187037 539552 187103 539564
rect 187037 538576 187053 539552
rect 187087 538576 187103 539552
rect 187037 538564 187103 538576
rect 187133 539552 187199 539564
rect 187133 538576 187149 539552
rect 187183 538576 187199 539552
rect 187133 538564 187199 538576
rect 187229 539552 187291 539564
rect 187229 538576 187245 539552
rect 187279 538576 187291 539552
rect 187358 539545 187416 539557
rect 187358 538969 187370 539545
rect 187404 538969 187416 539545
rect 187358 538957 187416 538969
rect 187446 539545 187504 539557
rect 187446 538969 187458 539545
rect 187492 538969 187504 539545
rect 187446 538957 187504 538969
rect 187558 539545 187616 539557
rect 187229 538564 187291 538576
rect 187558 538569 187570 539545
rect 187604 538569 187616 539545
rect 187558 538557 187616 538569
rect 187646 539545 187704 539557
rect 187646 538569 187658 539545
rect 187692 538569 187704 539545
rect 187646 538557 187704 538569
rect 189158 539545 189216 539557
rect 189158 538569 189170 539545
rect 189204 538569 189216 539545
rect 189158 538557 189216 538569
rect 189246 539545 189304 539557
rect 189246 538569 189258 539545
rect 189292 538569 189304 539545
rect 189246 538557 189304 538569
rect 189381 539552 189443 539564
rect 189381 538576 189393 539552
rect 189427 538576 189443 539552
rect 189381 538564 189443 538576
rect 189473 539552 189539 539564
rect 189473 538576 189489 539552
rect 189523 538576 189539 539552
rect 189473 538564 189539 538576
rect 189569 539552 189635 539564
rect 189569 538576 189585 539552
rect 189619 538576 189635 539552
rect 189569 538564 189635 538576
rect 189665 539552 189731 539564
rect 189665 538576 189681 539552
rect 189715 538576 189731 539552
rect 189665 538564 189731 538576
rect 189761 539552 189827 539564
rect 189761 538576 189777 539552
rect 189811 538576 189827 539552
rect 189761 538564 189827 538576
rect 189857 539552 189923 539564
rect 189857 538576 189873 539552
rect 189907 538576 189923 539552
rect 189857 538564 189923 538576
rect 189953 539552 190019 539564
rect 189953 538576 189969 539552
rect 190003 538576 190019 539552
rect 189953 538564 190019 538576
rect 190049 539552 190115 539564
rect 190049 538576 190065 539552
rect 190099 538576 190115 539552
rect 190049 538564 190115 538576
rect 190145 539552 190211 539564
rect 190145 538576 190161 539552
rect 190195 538576 190211 539552
rect 190145 538564 190211 538576
rect 190241 539552 190307 539564
rect 190241 538576 190257 539552
rect 190291 538576 190307 539552
rect 190241 538564 190307 538576
rect 190337 539552 190403 539564
rect 190337 538576 190353 539552
rect 190387 538576 190403 539552
rect 190337 538564 190403 538576
rect 190433 539552 190499 539564
rect 190433 538576 190449 539552
rect 190483 538576 190499 539552
rect 190433 538564 190499 538576
rect 190529 539552 190591 539564
rect 190529 538576 190545 539552
rect 190579 538576 190591 539552
rect 190658 539545 190716 539557
rect 190658 538969 190670 539545
rect 190704 538969 190716 539545
rect 190658 538957 190716 538969
rect 190746 539545 190804 539557
rect 190746 538969 190758 539545
rect 190792 538969 190804 539545
rect 190746 538957 190804 538969
rect 190858 539545 190916 539557
rect 190529 538564 190591 538576
rect 190858 538569 190870 539545
rect 190904 538569 190916 539545
rect 190858 538557 190916 538569
rect 190946 539545 191004 539557
rect 190946 538569 190958 539545
rect 190992 538569 191004 539545
rect 190946 538557 191004 538569
rect 161248 537645 161306 537657
rect 161248 537069 161260 537645
rect 161294 537069 161306 537645
rect 161248 537057 161306 537069
rect 161336 537645 161394 537657
rect 161336 537069 161348 537645
rect 161382 537069 161394 537645
rect 161336 537057 161394 537069
rect 161448 537645 161510 537657
rect 161448 537069 161460 537645
rect 161494 537069 161510 537645
rect 161448 537057 161510 537069
rect 161540 537645 161606 537657
rect 161540 537069 161556 537645
rect 161590 537069 161606 537645
rect 161540 537057 161606 537069
rect 161636 537645 161702 537657
rect 161636 537069 161652 537645
rect 161686 537069 161702 537645
rect 161636 537057 161702 537069
rect 161732 537645 161794 537657
rect 161732 537069 161748 537645
rect 161782 537069 161794 537645
rect 161732 537057 161794 537069
rect 161848 537645 161910 537657
rect 161848 537069 161860 537645
rect 161894 537069 161910 537645
rect 161848 537057 161910 537069
rect 161940 537645 162006 537657
rect 161940 537069 161956 537645
rect 161990 537069 162006 537645
rect 161940 537057 162006 537069
rect 162036 537645 162102 537657
rect 162036 537069 162052 537645
rect 162086 537069 162102 537645
rect 162036 537057 162102 537069
rect 162132 537645 162194 537657
rect 162132 537069 162148 537645
rect 162182 537069 162194 537645
rect 162132 537057 162194 537069
rect 162268 537645 162326 537657
rect 162268 537069 162280 537645
rect 162314 537069 162326 537645
rect 162268 537057 162326 537069
rect 162356 537645 162414 537657
rect 162356 537069 162368 537645
rect 162402 537069 162414 537645
rect 162356 537057 162414 537069
rect 157738 536625 157796 536637
rect 157738 536049 157750 536625
rect 157784 536049 157796 536625
rect 157738 536037 157796 536049
rect 157996 536625 158054 536637
rect 157996 536049 158008 536625
rect 158042 536049 158054 536625
rect 157996 536037 158054 536049
rect 158116 536625 158174 536637
rect 158116 536049 158128 536625
rect 158162 536049 158174 536625
rect 158116 536037 158174 536049
rect 158374 536625 158432 536637
rect 158374 536049 158386 536625
rect 158420 536049 158432 536625
rect 158374 536037 158432 536049
rect 158632 536625 158690 536637
rect 158632 536049 158644 536625
rect 158678 536049 158690 536625
rect 158632 536037 158690 536049
rect 158890 536625 158948 536637
rect 158890 536049 158902 536625
rect 158936 536049 158948 536625
rect 158890 536037 158948 536049
rect 159148 536625 159206 536637
rect 159148 536049 159160 536625
rect 159194 536049 159206 536625
rect 159148 536037 159206 536049
rect 159406 536625 159464 536637
rect 159406 536049 159418 536625
rect 159452 536049 159464 536625
rect 159406 536037 159464 536049
rect 159664 536625 159722 536637
rect 159664 536049 159676 536625
rect 159710 536049 159722 536625
rect 159664 536037 159722 536049
rect 159922 536625 159980 536637
rect 159922 536049 159934 536625
rect 159968 536049 159980 536625
rect 159922 536037 159980 536049
rect 160180 536625 160238 536637
rect 160180 536049 160192 536625
rect 160226 536049 160238 536625
rect 160180 536037 160238 536049
rect 160438 536625 160496 536637
rect 160438 536049 160450 536625
rect 160484 536049 160496 536625
rect 160438 536037 160496 536049
rect 160696 536625 160754 536637
rect 160696 536049 160708 536625
rect 160742 536049 160754 536625
rect 160696 536037 160754 536049
rect 160822 536625 160880 536637
rect 160822 536049 160834 536625
rect 160868 536049 160880 536625
rect 160822 536037 160880 536049
rect 161080 536625 161138 536637
rect 161080 536049 161092 536625
rect 161126 536049 161138 536625
rect 161080 536037 161138 536049
rect 161338 536625 161396 536637
rect 161338 536049 161350 536625
rect 161384 536049 161396 536625
rect 161338 536037 161396 536049
rect 161596 536625 161654 536637
rect 161596 536049 161608 536625
rect 161642 536049 161654 536625
rect 161596 536037 161654 536049
rect 161720 536625 161778 536637
rect 161720 536049 161732 536625
rect 161766 536049 161778 536625
rect 161720 536037 161778 536049
rect 161978 536625 162036 536637
rect 161978 536049 161990 536625
rect 162024 536049 162036 536625
rect 161978 536037 162036 536049
rect 162236 536625 162294 536637
rect 162236 536049 162248 536625
rect 162282 536049 162294 536625
rect 162236 536037 162294 536049
rect 162358 536625 162416 536637
rect 162358 536049 162370 536625
rect 162404 536049 162416 536625
rect 162358 536037 162416 536049
rect 162616 536625 162674 536637
rect 162616 536049 162628 536625
rect 162662 536049 162674 536625
rect 162616 536037 162674 536049
rect 172237 530255 172289 530288
rect 172237 530221 172245 530255
rect 172279 530221 172289 530255
rect 172237 530160 172289 530221
rect 172237 530126 172245 530160
rect 172279 530126 172289 530160
rect 172237 530114 172289 530126
rect 172407 530255 172459 530288
rect 172407 530221 172417 530255
rect 172451 530221 172459 530255
rect 172407 530160 172459 530221
rect 172407 530126 172417 530160
rect 172451 530126 172459 530160
rect 172407 530114 172459 530126
rect 172514 530242 172574 530314
rect 172514 530208 172529 530242
rect 172563 530208 172574 530242
rect 172514 530174 172574 530208
rect 172514 530140 172529 530174
rect 172563 530140 172574 530174
rect 172514 530114 172574 530140
rect 172604 530304 172660 530314
rect 172604 530270 172615 530304
rect 172649 530270 172660 530304
rect 172604 530236 172660 530270
rect 172604 530202 172615 530236
rect 172649 530202 172660 530236
rect 172604 530168 172660 530202
rect 172604 530134 172615 530168
rect 172649 530134 172660 530168
rect 172604 530114 172660 530134
rect 172690 530160 172746 530314
rect 172690 530126 172701 530160
rect 172735 530126 172746 530160
rect 172690 530114 172746 530126
rect 172776 530195 172832 530314
rect 172776 530161 172787 530195
rect 172821 530161 172832 530195
rect 172776 530114 172832 530161
rect 172862 530228 172928 530314
rect 172862 530194 172883 530228
rect 172917 530194 172928 530228
rect 172862 530160 172928 530194
rect 172862 530126 172883 530160
rect 172917 530126 172928 530160
rect 172862 530114 172928 530126
rect 172958 530290 173011 530314
rect 172958 530256 172969 530290
rect 173003 530256 173011 530290
rect 172958 530168 173011 530256
rect 172958 530134 172969 530168
rect 173003 530134 173011 530168
rect 172958 530114 173011 530134
rect 173065 530160 173117 530288
rect 173065 530126 173073 530160
rect 173107 530126 173117 530160
rect 173065 530114 173117 530126
rect 174063 530160 174115 530288
rect 174063 530126 174073 530160
rect 174107 530126 174115 530160
rect 174063 530114 174115 530126
rect 174169 530262 174221 530288
rect 174169 530228 174177 530262
rect 174211 530228 174221 530262
rect 174169 530160 174221 530228
rect 174169 530126 174177 530160
rect 174211 530126 174221 530160
rect 174169 530114 174221 530126
rect 174615 530262 174667 530288
rect 174615 530228 174625 530262
rect 174659 530228 174667 530262
rect 174615 530160 174667 530228
rect 174615 530126 174625 530160
rect 174659 530126 174667 530160
rect 174906 530242 174966 530314
rect 174906 530208 174921 530242
rect 174955 530208 174966 530242
rect 174906 530174 174966 530208
rect 174906 530140 174921 530174
rect 174955 530140 174966 530174
rect 174615 530114 174667 530126
rect 174906 530114 174966 530140
rect 174996 530304 175052 530314
rect 174996 530270 175007 530304
rect 175041 530270 175052 530304
rect 174996 530236 175052 530270
rect 174996 530202 175007 530236
rect 175041 530202 175052 530236
rect 174996 530168 175052 530202
rect 174996 530134 175007 530168
rect 175041 530134 175052 530168
rect 174996 530114 175052 530134
rect 175082 530160 175138 530314
rect 175082 530126 175093 530160
rect 175127 530126 175138 530160
rect 175082 530114 175138 530126
rect 175168 530195 175224 530314
rect 175168 530161 175179 530195
rect 175213 530161 175224 530195
rect 175168 530114 175224 530161
rect 175254 530228 175320 530314
rect 175254 530194 175275 530228
rect 175309 530194 175320 530228
rect 175254 530160 175320 530194
rect 175254 530126 175275 530160
rect 175309 530126 175320 530160
rect 175254 530114 175320 530126
rect 175350 530290 175403 530314
rect 175350 530256 175361 530290
rect 175395 530256 175403 530290
rect 175350 530168 175403 530256
rect 175350 530134 175361 530168
rect 175395 530134 175403 530168
rect 175350 530114 175403 530134
rect 175549 530264 175601 530314
rect 175549 530230 175557 530264
rect 175591 530230 175601 530264
rect 175549 530196 175601 530230
rect 175549 530162 175557 530196
rect 175591 530162 175601 530196
rect 175549 530114 175601 530162
rect 175631 530242 175681 530314
rect 175631 530228 175697 530242
rect 175631 530194 175641 530228
rect 175675 530194 175697 530228
rect 176223 530198 176277 530282
rect 175631 530160 175697 530194
rect 175631 530126 175641 530160
rect 175675 530126 175697 530160
rect 175631 530114 175697 530126
rect 175762 530160 175816 530198
rect 175762 530126 175770 530160
rect 175804 530126 175816 530160
rect 175762 530114 175816 530126
rect 175846 530186 175900 530198
rect 175846 530152 175856 530186
rect 175890 530152 175900 530186
rect 175846 530114 175900 530152
rect 175930 530160 176008 530198
rect 175930 530126 175940 530160
rect 175974 530126 176008 530160
rect 175930 530114 176008 530126
rect 176038 530114 176092 530198
rect 176122 530161 176178 530198
rect 176122 530127 176132 530161
rect 176166 530127 176178 530161
rect 176122 530114 176178 530127
rect 176208 530168 176277 530198
rect 176208 530134 176229 530168
rect 176263 530134 176277 530168
rect 176208 530114 176277 530134
rect 176307 530160 176359 530282
rect 177117 530236 177169 530248
rect 177117 530202 177125 530236
rect 177159 530202 177169 530236
rect 176307 530126 176317 530160
rect 176351 530126 176359 530160
rect 176307 530114 176359 530126
rect 176422 530186 176474 530198
rect 176422 530152 176430 530186
rect 176464 530152 176474 530186
rect 176422 530114 176474 530152
rect 176504 530170 176571 530198
rect 176504 530136 176514 530170
rect 176548 530136 176571 530170
rect 176504 530114 176571 530136
rect 176601 530186 176711 530198
rect 176601 530152 176611 530186
rect 176645 530152 176711 530186
rect 176601 530114 176711 530152
rect 176741 530162 176810 530198
rect 176741 530128 176765 530162
rect 176799 530128 176810 530162
rect 176741 530114 176810 530128
rect 176840 530168 176902 530198
rect 176840 530134 176858 530168
rect 176892 530134 176902 530168
rect 176840 530114 176902 530134
rect 176932 530160 176984 530198
rect 176932 530126 176942 530160
rect 176976 530126 176984 530160
rect 176932 530114 176984 530126
rect 177117 530168 177169 530202
rect 177117 530134 177125 530168
rect 177159 530134 177169 530168
rect 177117 530120 177169 530134
rect 177199 530184 177253 530248
rect 177199 530150 177209 530184
rect 177243 530150 177253 530184
rect 177199 530120 177253 530150
rect 177283 530236 177335 530248
rect 177283 530202 177293 530236
rect 177327 530202 177335 530236
rect 177283 530168 177335 530202
rect 177283 530134 177293 530168
rect 177327 530134 177335 530168
rect 177283 530120 177335 530134
rect 177684 530186 177736 530314
rect 177684 530152 177692 530186
rect 177726 530152 177736 530186
rect 177684 530114 177736 530152
rect 177766 530198 177816 530314
rect 178401 530249 178453 530272
rect 178401 530215 178409 530249
rect 178443 530215 178453 530249
rect 177766 530160 177831 530198
rect 177766 530126 177782 530160
rect 177816 530126 177831 530160
rect 177766 530114 177831 530126
rect 177931 530186 177983 530198
rect 177931 530152 177941 530186
rect 177975 530152 177983 530186
rect 177931 530114 177983 530152
rect 178037 530186 178089 530198
rect 178037 530152 178045 530186
rect 178079 530152 178089 530186
rect 178037 530114 178089 530152
rect 178189 530160 178243 530198
rect 178189 530126 178199 530160
rect 178233 530126 178243 530160
rect 178189 530114 178243 530126
rect 178273 530186 178325 530198
rect 178273 530152 178283 530186
rect 178317 530152 178325 530186
rect 178273 530114 178325 530152
rect 178401 530168 178453 530215
rect 178401 530134 178409 530168
rect 178443 530134 178453 530168
rect 178401 530114 178453 530134
rect 178483 530236 178541 530272
rect 178483 530202 178495 530236
rect 178529 530202 178541 530236
rect 178483 530168 178541 530202
rect 178483 530134 178495 530168
rect 178529 530134 178541 530168
rect 178483 530114 178541 530134
rect 178571 530236 178623 530272
rect 178571 530202 178581 530236
rect 178615 530202 178623 530236
rect 178571 530168 178623 530202
rect 178571 530134 178581 530168
rect 178615 530134 178623 530168
rect 178571 530114 178623 530134
rect 178678 530242 178738 530314
rect 178678 530208 178693 530242
rect 178727 530208 178738 530242
rect 178678 530174 178738 530208
rect 178678 530140 178693 530174
rect 178727 530140 178738 530174
rect 178678 530114 178738 530140
rect 178768 530304 178824 530314
rect 178768 530270 178779 530304
rect 178813 530270 178824 530304
rect 178768 530236 178824 530270
rect 178768 530202 178779 530236
rect 178813 530202 178824 530236
rect 178768 530168 178824 530202
rect 178768 530134 178779 530168
rect 178813 530134 178824 530168
rect 178768 530114 178824 530134
rect 178854 530160 178910 530314
rect 178854 530126 178865 530160
rect 178899 530126 178910 530160
rect 178854 530114 178910 530126
rect 178940 530195 178996 530314
rect 178940 530161 178951 530195
rect 178985 530161 178996 530195
rect 178940 530114 178996 530161
rect 179026 530228 179092 530314
rect 179026 530194 179047 530228
rect 179081 530194 179092 530228
rect 179026 530160 179092 530194
rect 179026 530126 179047 530160
rect 179081 530126 179092 530160
rect 179026 530114 179092 530126
rect 179122 530290 179175 530314
rect 179122 530256 179133 530290
rect 179167 530256 179175 530290
rect 179122 530168 179175 530256
rect 179122 530134 179133 530168
rect 179167 530134 179175 530168
rect 179122 530114 179175 530134
rect 179229 530290 179282 530314
rect 179229 530256 179237 530290
rect 179271 530256 179282 530290
rect 179229 530168 179282 530256
rect 179229 530134 179237 530168
rect 179271 530134 179282 530168
rect 179229 530114 179282 530134
rect 179312 530228 179378 530314
rect 179312 530194 179323 530228
rect 179357 530194 179378 530228
rect 179312 530160 179378 530194
rect 179312 530126 179323 530160
rect 179357 530126 179378 530160
rect 179312 530114 179378 530126
rect 179408 530195 179464 530314
rect 179408 530161 179419 530195
rect 179453 530161 179464 530195
rect 179408 530114 179464 530161
rect 179494 530160 179550 530314
rect 179494 530126 179505 530160
rect 179539 530126 179550 530160
rect 179494 530114 179550 530126
rect 179580 530304 179636 530314
rect 179580 530270 179591 530304
rect 179625 530270 179636 530304
rect 179580 530236 179636 530270
rect 179580 530202 179591 530236
rect 179625 530202 179636 530236
rect 179580 530168 179636 530202
rect 179580 530134 179591 530168
rect 179625 530134 179636 530168
rect 179580 530114 179636 530134
rect 179666 530242 179726 530314
rect 179666 530208 179677 530242
rect 179711 530208 179726 530242
rect 179666 530174 179726 530208
rect 179666 530140 179677 530174
rect 179711 530140 179726 530174
rect 179666 530114 179726 530140
rect 180241 530296 180293 530314
rect 180241 530262 180249 530296
rect 180283 530262 180293 530296
rect 180241 530228 180293 530262
rect 180241 530194 180249 530228
rect 180283 530194 180293 530228
rect 180241 530160 180293 530194
rect 180241 530126 180249 530160
rect 180283 530126 180293 530160
rect 180241 530114 180293 530126
rect 180323 530296 180375 530314
rect 180323 530262 180333 530296
rect 180367 530262 180375 530296
rect 180323 530237 180375 530262
rect 181801 530296 181853 530314
rect 181801 530262 181809 530296
rect 181843 530262 181853 530296
rect 181801 530237 181853 530262
rect 180323 530228 180402 530237
rect 180323 530194 180333 530228
rect 180367 530194 180402 530228
rect 180323 530160 180402 530194
rect 180323 530126 180333 530160
rect 180367 530153 180402 530160
rect 180432 530153 180505 530237
rect 180535 530220 180719 530237
rect 180535 530186 180569 530220
rect 180603 530186 180644 530220
rect 180678 530186 180719 530220
rect 180535 530153 180719 530186
rect 180749 530153 180791 530237
rect 180821 530220 180887 530237
rect 180821 530186 180841 530220
rect 180875 530186 180887 530220
rect 180821 530153 180887 530186
rect 180917 530220 180973 530237
rect 180917 530186 180927 530220
rect 180961 530186 180973 530220
rect 180917 530153 180973 530186
rect 181203 530220 181259 530237
rect 181203 530186 181215 530220
rect 181249 530186 181259 530220
rect 181203 530153 181259 530186
rect 181289 530220 181355 530237
rect 181289 530186 181301 530220
rect 181335 530186 181355 530220
rect 181289 530153 181355 530186
rect 181385 530153 181427 530237
rect 181457 530220 181641 530237
rect 181457 530186 181498 530220
rect 181532 530186 181573 530220
rect 181607 530186 181641 530220
rect 181457 530153 181641 530186
rect 181671 530153 181744 530237
rect 181774 530228 181853 530237
rect 181774 530194 181809 530228
rect 181843 530194 181853 530228
rect 181774 530160 181853 530194
rect 181774 530153 181809 530160
rect 180367 530126 180375 530153
rect 180323 530114 180375 530126
rect 181801 530126 181809 530153
rect 181843 530126 181853 530160
rect 181801 530114 181853 530126
rect 181883 530296 181935 530314
rect 181883 530262 181893 530296
rect 181927 530262 181935 530296
rect 181883 530228 181935 530262
rect 181883 530194 181893 530228
rect 181927 530194 181935 530228
rect 181883 530160 181935 530194
rect 181883 530126 181893 530160
rect 181927 530126 181935 530160
rect 181883 530114 181935 530126
rect 181989 530290 182042 530314
rect 181989 530256 181997 530290
rect 182031 530256 182042 530290
rect 181989 530168 182042 530256
rect 181989 530134 181997 530168
rect 182031 530134 182042 530168
rect 181989 530114 182042 530134
rect 182072 530228 182138 530314
rect 182072 530194 182083 530228
rect 182117 530194 182138 530228
rect 182072 530160 182138 530194
rect 182072 530126 182083 530160
rect 182117 530126 182138 530160
rect 182072 530114 182138 530126
rect 182168 530195 182224 530314
rect 182168 530161 182179 530195
rect 182213 530161 182224 530195
rect 182168 530114 182224 530161
rect 182254 530160 182310 530314
rect 182254 530126 182265 530160
rect 182299 530126 182310 530160
rect 182254 530114 182310 530126
rect 182340 530304 182396 530314
rect 182340 530270 182351 530304
rect 182385 530270 182396 530304
rect 182340 530236 182396 530270
rect 182340 530202 182351 530236
rect 182385 530202 182396 530236
rect 182340 530168 182396 530202
rect 182340 530134 182351 530168
rect 182385 530134 182396 530168
rect 182340 530114 182396 530134
rect 182426 530242 182486 530314
rect 182426 530208 182437 530242
rect 182471 530208 182486 530242
rect 182426 530174 182486 530208
rect 182426 530140 182437 530174
rect 182471 530140 182486 530174
rect 182426 530114 182486 530140
rect 183093 530290 183146 530314
rect 182633 530262 182685 530288
rect 182633 530228 182641 530262
rect 182675 530228 182685 530262
rect 182633 530160 182685 530228
rect 182633 530126 182641 530160
rect 182675 530126 182685 530160
rect 182633 530114 182685 530126
rect 182895 530262 182947 530288
rect 182895 530228 182905 530262
rect 182939 530228 182947 530262
rect 182895 530160 182947 530228
rect 182895 530126 182905 530160
rect 182939 530126 182947 530160
rect 182895 530114 182947 530126
rect 183093 530256 183101 530290
rect 183135 530256 183146 530290
rect 183093 530168 183146 530256
rect 183093 530134 183101 530168
rect 183135 530134 183146 530168
rect 183093 530114 183146 530134
rect 183176 530228 183242 530314
rect 183176 530194 183187 530228
rect 183221 530194 183242 530228
rect 183176 530160 183242 530194
rect 183176 530126 183187 530160
rect 183221 530126 183242 530160
rect 183176 530114 183242 530126
rect 183272 530195 183328 530314
rect 183272 530161 183283 530195
rect 183317 530161 183328 530195
rect 183272 530114 183328 530161
rect 183358 530160 183414 530314
rect 183358 530126 183369 530160
rect 183403 530126 183414 530160
rect 183358 530114 183414 530126
rect 183444 530304 183500 530314
rect 183444 530270 183455 530304
rect 183489 530270 183500 530304
rect 183444 530236 183500 530270
rect 183444 530202 183455 530236
rect 183489 530202 183500 530236
rect 183444 530168 183500 530202
rect 183444 530134 183455 530168
rect 183489 530134 183500 530168
rect 183444 530114 183500 530134
rect 183530 530242 183590 530314
rect 183530 530208 183541 530242
rect 183575 530208 183590 530242
rect 183530 530174 183590 530208
rect 183530 530140 183541 530174
rect 183575 530140 183590 530174
rect 183530 530114 183590 530140
rect 183645 530160 183697 530288
rect 183645 530126 183653 530160
rect 183687 530126 183697 530160
rect 183645 530114 183697 530126
rect 184643 530160 184695 530288
rect 184643 530126 184653 530160
rect 184687 530126 184695 530160
rect 184643 530114 184695 530126
rect 184749 530262 184801 530288
rect 184749 530228 184757 530262
rect 184791 530228 184801 530262
rect 184749 530160 184801 530228
rect 184749 530126 184757 530160
rect 184791 530126 184801 530160
rect 184749 530114 184801 530126
rect 185011 530262 185063 530288
rect 185011 530228 185021 530262
rect 185055 530228 185063 530262
rect 185011 530160 185063 530228
rect 185011 530126 185021 530160
rect 185055 530126 185063 530160
rect 185209 530290 185262 530314
rect 185209 530256 185217 530290
rect 185251 530256 185262 530290
rect 185209 530168 185262 530256
rect 185209 530134 185217 530168
rect 185251 530134 185262 530168
rect 185011 530114 185063 530126
rect 185209 530114 185262 530134
rect 185292 530228 185358 530314
rect 185292 530194 185303 530228
rect 185337 530194 185358 530228
rect 185292 530160 185358 530194
rect 185292 530126 185303 530160
rect 185337 530126 185358 530160
rect 185292 530114 185358 530126
rect 185388 530195 185444 530314
rect 185388 530161 185399 530195
rect 185433 530161 185444 530195
rect 185388 530114 185444 530161
rect 185474 530160 185530 530314
rect 185474 530126 185485 530160
rect 185519 530126 185530 530160
rect 185474 530114 185530 530126
rect 185560 530304 185616 530314
rect 185560 530270 185571 530304
rect 185605 530270 185616 530304
rect 185560 530236 185616 530270
rect 185560 530202 185571 530236
rect 185605 530202 185616 530236
rect 185560 530168 185616 530202
rect 185560 530134 185571 530168
rect 185605 530134 185616 530168
rect 185560 530114 185616 530134
rect 185646 530242 185706 530314
rect 185646 530208 185657 530242
rect 185691 530208 185706 530242
rect 185646 530174 185706 530208
rect 185646 530140 185657 530174
rect 185691 530140 185706 530174
rect 185646 530114 185706 530140
rect 185761 530160 185813 530288
rect 185761 530126 185769 530160
rect 185803 530126 185813 530160
rect 185761 530114 185813 530126
rect 186759 530160 186811 530288
rect 186759 530126 186769 530160
rect 186803 530126 186811 530160
rect 186759 530114 186811 530126
rect 187233 530255 187285 530288
rect 187233 530221 187241 530255
rect 187275 530221 187285 530255
rect 187233 530160 187285 530221
rect 187233 530126 187241 530160
rect 187275 530126 187285 530160
rect 187233 530114 187285 530126
rect 187403 530255 187455 530288
rect 187403 530221 187413 530255
rect 187447 530221 187455 530255
rect 187403 530160 187455 530221
rect 187403 530126 187413 530160
rect 187447 530126 187455 530160
rect 187403 530114 187455 530126
rect 172237 530008 172289 530020
rect 172237 529974 172245 530008
rect 172279 529974 172289 530008
rect 172237 529913 172289 529974
rect 172237 529879 172245 529913
rect 172279 529879 172289 529913
rect 172237 529846 172289 529879
rect 172407 530008 172459 530020
rect 172407 529974 172417 530008
rect 172451 529974 172459 530008
rect 172407 529913 172459 529974
rect 172407 529879 172417 529913
rect 172451 529879 172459 529913
rect 172407 529846 172459 529879
rect 172513 530008 172565 530020
rect 172513 529974 172521 530008
rect 172555 529974 172565 530008
rect 172513 529846 172565 529974
rect 173511 530008 173563 530020
rect 173511 529974 173521 530008
rect 173555 529974 173563 530008
rect 173511 529846 173563 529974
rect 173617 530008 173669 530020
rect 173617 529974 173625 530008
rect 173659 529974 173669 530008
rect 173617 529846 173669 529974
rect 174615 530008 174667 530020
rect 174615 529974 174625 530008
rect 174659 529974 174667 530008
rect 174615 529846 174667 529974
rect 174835 529982 174887 530020
rect 174835 529948 174843 529982
rect 174877 529948 174887 529982
rect 174835 529936 174887 529948
rect 174917 530008 174971 530020
rect 174917 529974 174927 530008
rect 174961 529974 174971 530008
rect 174917 529936 174971 529974
rect 175071 529982 175123 530020
rect 175071 529948 175081 529982
rect 175115 529948 175123 529982
rect 175071 529936 175123 529948
rect 175177 529982 175229 530020
rect 175177 529948 175185 529982
rect 175219 529948 175229 529982
rect 175177 529936 175229 529948
rect 175329 530008 175394 530020
rect 175329 529974 175344 530008
rect 175378 529974 175394 530008
rect 175329 529936 175394 529974
rect 175344 529820 175394 529936
rect 175424 529982 175476 530020
rect 175424 529948 175434 529982
rect 175468 529948 175476 529982
rect 175424 529820 175476 529948
rect 175549 530000 175601 530014
rect 175549 529966 175557 530000
rect 175591 529966 175601 530000
rect 175549 529932 175601 529966
rect 175549 529898 175557 529932
rect 175591 529898 175601 529932
rect 175549 529886 175601 529898
rect 175631 529984 175685 530014
rect 175631 529950 175641 529984
rect 175675 529950 175685 529984
rect 175631 529886 175685 529950
rect 175715 530000 175767 530014
rect 175715 529966 175725 530000
rect 175759 529966 175767 530000
rect 175715 529932 175767 529966
rect 175900 530008 175952 530020
rect 175900 529974 175908 530008
rect 175942 529974 175952 530008
rect 175900 529936 175952 529974
rect 175982 530000 176044 530020
rect 175982 529966 175992 530000
rect 176026 529966 176044 530000
rect 175982 529936 176044 529966
rect 176074 530006 176143 530020
rect 176074 529972 176085 530006
rect 176119 529972 176143 530006
rect 176074 529936 176143 529972
rect 176173 529982 176283 530020
rect 176173 529948 176239 529982
rect 176273 529948 176283 529982
rect 176173 529936 176283 529948
rect 176313 529998 176380 530020
rect 176313 529964 176336 529998
rect 176370 529964 176380 529998
rect 176313 529936 176380 529964
rect 176410 529982 176462 530020
rect 176410 529948 176420 529982
rect 176454 529948 176462 529982
rect 176410 529936 176462 529948
rect 176525 530008 176577 530020
rect 176525 529974 176533 530008
rect 176567 529974 176577 530008
rect 175715 529898 175725 529932
rect 175759 529898 175767 529932
rect 175715 529886 175767 529898
rect 176525 529852 176577 529974
rect 176607 530000 176676 530020
rect 176607 529966 176621 530000
rect 176655 529966 176676 530000
rect 176607 529936 176676 529966
rect 176706 530007 176762 530020
rect 176706 529973 176718 530007
rect 176752 529973 176762 530007
rect 176706 529936 176762 529973
rect 176792 529936 176846 530020
rect 176876 530008 176954 530020
rect 176876 529974 176910 530008
rect 176944 529974 176954 530008
rect 176876 529936 176954 529974
rect 176984 529982 177038 530020
rect 176984 529948 176994 529982
rect 177028 529948 177038 529982
rect 176984 529936 177038 529948
rect 177068 530008 177122 530020
rect 177068 529974 177080 530008
rect 177114 529974 177122 530008
rect 177068 529936 177122 529974
rect 177187 530008 177253 530020
rect 177187 529974 177209 530008
rect 177243 529974 177253 530008
rect 177187 529940 177253 529974
rect 176607 529852 176661 529936
rect 177187 529906 177209 529940
rect 177243 529906 177253 529940
rect 177187 529892 177253 529906
rect 177203 529820 177253 529892
rect 177283 529972 177335 530020
rect 178213 530008 178265 530020
rect 177283 529938 177293 529972
rect 177327 529938 177335 529972
rect 177283 529904 177335 529938
rect 177283 529870 177293 529904
rect 177327 529870 177335 529904
rect 177283 529820 177335 529870
rect 178213 529981 178221 530008
rect 177615 529948 177671 529981
rect 177615 529914 177627 529948
rect 177661 529914 177671 529948
rect 177615 529897 177671 529914
rect 177701 529948 177767 529981
rect 177701 529914 177713 529948
rect 177747 529914 177767 529948
rect 177701 529897 177767 529914
rect 177797 529897 177839 529981
rect 177869 529948 178053 529981
rect 177869 529914 177910 529948
rect 177944 529914 177985 529948
rect 178019 529914 178053 529948
rect 177869 529897 178053 529914
rect 178083 529897 178156 529981
rect 178186 529974 178221 529981
rect 178255 529974 178265 530008
rect 178186 529940 178265 529974
rect 178186 529906 178221 529940
rect 178255 529906 178265 529940
rect 178186 529897 178265 529906
rect 178213 529872 178265 529897
rect 178213 529838 178221 529872
rect 178255 529838 178265 529872
rect 178213 529820 178265 529838
rect 178295 530008 178347 530020
rect 178295 529974 178305 530008
rect 178339 529974 178347 530008
rect 178295 529940 178347 529974
rect 178295 529906 178305 529940
rect 178339 529906 178347 529940
rect 178295 529872 178347 529906
rect 178295 529838 178305 529872
rect 178339 529838 178347 529872
rect 178295 529820 178347 529838
rect 178401 529972 178453 530020
rect 178401 529938 178409 529972
rect 178443 529938 178453 529972
rect 178401 529904 178453 529938
rect 178401 529870 178409 529904
rect 178443 529870 178453 529904
rect 178401 529820 178453 529870
rect 178483 530008 178549 530020
rect 178483 529974 178493 530008
rect 178527 529974 178549 530008
rect 178483 529940 178549 529974
rect 178483 529906 178493 529940
rect 178527 529906 178549 529940
rect 178614 530008 178668 530020
rect 178614 529974 178622 530008
rect 178656 529974 178668 530008
rect 178614 529936 178668 529974
rect 178698 529982 178752 530020
rect 178698 529948 178708 529982
rect 178742 529948 178752 529982
rect 178698 529936 178752 529948
rect 178782 530008 178860 530020
rect 178782 529974 178792 530008
rect 178826 529974 178860 530008
rect 178782 529936 178860 529974
rect 178890 529936 178944 530020
rect 178974 530007 179030 530020
rect 178974 529973 178984 530007
rect 179018 529973 179030 530007
rect 178974 529936 179030 529973
rect 179060 530000 179129 530020
rect 179060 529966 179081 530000
rect 179115 529966 179129 530000
rect 179060 529936 179129 529966
rect 178483 529892 178549 529906
rect 178483 529820 178533 529892
rect 179075 529852 179129 529936
rect 179159 530008 179211 530020
rect 179159 529974 179169 530008
rect 179203 529974 179211 530008
rect 179159 529852 179211 529974
rect 179274 529982 179326 530020
rect 179274 529948 179282 529982
rect 179316 529948 179326 529982
rect 179274 529936 179326 529948
rect 179356 529998 179423 530020
rect 179356 529964 179366 529998
rect 179400 529964 179423 529998
rect 179356 529936 179423 529964
rect 179453 529982 179563 530020
rect 179453 529948 179463 529982
rect 179497 529948 179563 529982
rect 179453 529936 179563 529948
rect 179593 530006 179662 530020
rect 179593 529972 179617 530006
rect 179651 529972 179662 530006
rect 179593 529936 179662 529972
rect 179692 530000 179754 530020
rect 179692 529966 179710 530000
rect 179744 529966 179754 530000
rect 179692 529936 179754 529966
rect 179784 530008 179836 530020
rect 179784 529974 179794 530008
rect 179828 529974 179836 530008
rect 179784 529936 179836 529974
rect 179969 530000 180021 530014
rect 179969 529966 179977 530000
rect 180011 529966 180021 530000
rect 179969 529932 180021 529966
rect 179969 529898 179977 529932
rect 180011 529898 180021 529932
rect 179969 529886 180021 529898
rect 180051 529984 180105 530014
rect 180051 529950 180061 529984
rect 180095 529950 180105 529984
rect 180051 529886 180105 529950
rect 180135 530000 180187 530014
rect 180135 529966 180145 530000
rect 180179 529966 180187 530000
rect 180135 529932 180187 529966
rect 180135 529898 180145 529932
rect 180179 529898 180187 529932
rect 180135 529886 180187 529898
rect 180241 530000 180293 530014
rect 180241 529966 180249 530000
rect 180283 529966 180293 530000
rect 180241 529932 180293 529966
rect 180241 529898 180249 529932
rect 180283 529898 180293 529932
rect 180241 529886 180293 529898
rect 180323 529984 180377 530014
rect 180323 529950 180333 529984
rect 180367 529950 180377 529984
rect 180323 529886 180377 529950
rect 180407 530000 180459 530014
rect 180407 529966 180417 530000
rect 180451 529966 180459 530000
rect 180407 529932 180459 529966
rect 180592 530008 180644 530020
rect 180592 529974 180600 530008
rect 180634 529974 180644 530008
rect 180592 529936 180644 529974
rect 180674 530000 180736 530020
rect 180674 529966 180684 530000
rect 180718 529966 180736 530000
rect 180674 529936 180736 529966
rect 180766 530006 180835 530020
rect 180766 529972 180777 530006
rect 180811 529972 180835 530006
rect 180766 529936 180835 529972
rect 180865 529982 180975 530020
rect 180865 529948 180931 529982
rect 180965 529948 180975 529982
rect 180865 529936 180975 529948
rect 181005 529998 181072 530020
rect 181005 529964 181028 529998
rect 181062 529964 181072 529998
rect 181005 529936 181072 529964
rect 181102 529982 181154 530020
rect 181102 529948 181112 529982
rect 181146 529948 181154 529982
rect 181102 529936 181154 529948
rect 181217 530008 181269 530020
rect 181217 529974 181225 530008
rect 181259 529974 181269 530008
rect 180407 529898 180417 529932
rect 180451 529898 180459 529932
rect 180407 529886 180459 529898
rect 181217 529852 181269 529974
rect 181299 530000 181368 530020
rect 181299 529966 181313 530000
rect 181347 529966 181368 530000
rect 181299 529936 181368 529966
rect 181398 530007 181454 530020
rect 181398 529973 181410 530007
rect 181444 529973 181454 530007
rect 181398 529936 181454 529973
rect 181484 529936 181538 530020
rect 181568 530008 181646 530020
rect 181568 529974 181602 530008
rect 181636 529974 181646 530008
rect 181568 529936 181646 529974
rect 181676 529982 181730 530020
rect 181676 529948 181686 529982
rect 181720 529948 181730 529982
rect 181676 529936 181730 529948
rect 181760 530008 181814 530020
rect 181760 529974 181772 530008
rect 181806 529974 181814 530008
rect 181760 529936 181814 529974
rect 181879 530008 181945 530020
rect 181879 529974 181901 530008
rect 181935 529974 181945 530008
rect 181879 529940 181945 529974
rect 181299 529852 181353 529936
rect 181879 529906 181901 529940
rect 181935 529906 181945 529940
rect 181879 529892 181945 529906
rect 181895 529820 181945 529892
rect 181975 529972 182027 530020
rect 181975 529938 181985 529972
rect 182019 529938 182027 529972
rect 181975 529904 182027 529938
rect 181975 529870 181985 529904
rect 182019 529870 182027 529904
rect 181975 529820 182027 529870
rect 182081 530008 182133 530020
rect 182081 529974 182089 530008
rect 182123 529974 182133 530008
rect 182081 529906 182133 529974
rect 182081 529872 182089 529906
rect 182123 529872 182133 529906
rect 182081 529846 182133 529872
rect 182343 530008 182395 530020
rect 182343 529974 182353 530008
rect 182387 529974 182395 530008
rect 182343 529906 182395 529974
rect 182343 529872 182353 529906
rect 182387 529872 182395 529906
rect 182343 529846 182395 529872
rect 182652 529982 182704 530020
rect 182652 529948 182660 529982
rect 182694 529948 182704 529982
rect 182652 529820 182704 529948
rect 182734 530008 182799 530020
rect 182734 529974 182750 530008
rect 182784 529974 182799 530008
rect 182734 529936 182799 529974
rect 182899 529982 182951 530020
rect 182899 529948 182909 529982
rect 182943 529948 182951 529982
rect 182899 529936 182951 529948
rect 183005 529982 183057 530020
rect 183005 529948 183013 529982
rect 183047 529948 183057 529982
rect 183005 529936 183057 529948
rect 183157 530008 183211 530020
rect 183157 529974 183167 530008
rect 183201 529974 183211 530008
rect 183157 529936 183211 529974
rect 183241 529982 183293 530020
rect 183241 529948 183251 529982
rect 183285 529948 183293 529982
rect 183241 529936 183293 529948
rect 183369 530008 183421 530020
rect 183369 529974 183377 530008
rect 183411 529974 183421 530008
rect 182734 529820 182784 529936
rect 183369 529846 183421 529974
rect 184367 530008 184419 530020
rect 184367 529974 184377 530008
rect 184411 529974 184419 530008
rect 184367 529846 184419 529974
rect 184473 530008 184525 530020
rect 184473 529974 184481 530008
rect 184515 529974 184525 530008
rect 184473 529846 184525 529974
rect 185471 530008 185523 530020
rect 185471 529974 185481 530008
rect 185515 529974 185523 530008
rect 185471 529846 185523 529974
rect 185577 530008 185629 530020
rect 185577 529974 185585 530008
rect 185619 529974 185629 530008
rect 185577 529846 185629 529974
rect 186575 530008 186627 530020
rect 186575 529974 186585 530008
rect 186619 529974 186627 530008
rect 186575 529846 186627 529974
rect 186681 530008 186733 530020
rect 186681 529974 186689 530008
rect 186723 529974 186733 530008
rect 186681 529906 186733 529974
rect 186681 529872 186689 529906
rect 186723 529872 186733 529906
rect 186681 529846 186733 529872
rect 187127 530008 187179 530020
rect 187127 529974 187137 530008
rect 187171 529974 187179 530008
rect 187127 529906 187179 529974
rect 187127 529872 187137 529906
rect 187171 529872 187179 529906
rect 187127 529846 187179 529872
rect 187233 530008 187285 530020
rect 187233 529974 187241 530008
rect 187275 529974 187285 530008
rect 187233 529913 187285 529974
rect 187233 529879 187241 529913
rect 187275 529879 187285 529913
rect 187233 529846 187285 529879
rect 187403 530008 187455 530020
rect 187403 529974 187413 530008
rect 187447 529974 187455 530008
rect 187403 529913 187455 529974
rect 187403 529879 187413 529913
rect 187447 529879 187455 529913
rect 187403 529846 187455 529879
rect 172237 529167 172289 529200
rect 172237 529133 172245 529167
rect 172279 529133 172289 529167
rect 172237 529072 172289 529133
rect 172237 529038 172245 529072
rect 172279 529038 172289 529072
rect 172237 529026 172289 529038
rect 172407 529167 172459 529200
rect 172407 529133 172417 529167
rect 172451 529133 172459 529167
rect 172407 529072 172459 529133
rect 172407 529038 172417 529072
rect 172451 529038 172459 529072
rect 172407 529026 172459 529038
rect 172513 529072 172565 529200
rect 172513 529038 172521 529072
rect 172555 529038 172565 529072
rect 172513 529026 172565 529038
rect 173511 529072 173563 529200
rect 173511 529038 173521 529072
rect 173555 529038 173563 529072
rect 173511 529026 173563 529038
rect 173617 529072 173669 529200
rect 173617 529038 173625 529072
rect 173659 529038 173669 529072
rect 173617 529026 173669 529038
rect 174615 529072 174667 529200
rect 174615 529038 174625 529072
rect 174659 529038 174667 529072
rect 175729 529208 175781 529226
rect 175729 529174 175737 529208
rect 175771 529174 175781 529208
rect 175729 529149 175781 529174
rect 175131 529132 175187 529149
rect 175131 529098 175143 529132
rect 175177 529098 175187 529132
rect 175131 529065 175187 529098
rect 175217 529132 175283 529149
rect 175217 529098 175229 529132
rect 175263 529098 175283 529132
rect 175217 529065 175283 529098
rect 175313 529065 175355 529149
rect 175385 529132 175569 529149
rect 175385 529098 175426 529132
rect 175460 529098 175501 529132
rect 175535 529098 175569 529132
rect 175385 529065 175569 529098
rect 175599 529065 175672 529149
rect 175702 529140 175781 529149
rect 175702 529106 175737 529140
rect 175771 529106 175781 529140
rect 175702 529072 175781 529106
rect 175702 529065 175737 529072
rect 174615 529026 174667 529038
rect 175729 529038 175737 529065
rect 175771 529038 175781 529072
rect 175729 529026 175781 529038
rect 175811 529208 175863 529226
rect 175811 529174 175821 529208
rect 175855 529174 175863 529208
rect 175811 529140 175863 529174
rect 175811 529106 175821 529140
rect 175855 529106 175863 529140
rect 175811 529072 175863 529106
rect 175811 529038 175821 529072
rect 175855 529038 175863 529072
rect 175811 529026 175863 529038
rect 175934 529096 175987 529226
rect 175934 529062 175942 529096
rect 175976 529062 175987 529096
rect 175934 529026 175987 529062
rect 176017 529202 176073 529226
rect 176017 529168 176028 529202
rect 176062 529168 176073 529202
rect 176017 529116 176073 529168
rect 176017 529082 176028 529116
rect 176062 529082 176073 529116
rect 176017 529026 176073 529082
rect 176103 529096 176159 529226
rect 176103 529062 176114 529096
rect 176148 529062 176159 529096
rect 176103 529026 176159 529062
rect 176189 529202 176245 529226
rect 176189 529168 176200 529202
rect 176234 529168 176245 529202
rect 176189 529116 176245 529168
rect 176189 529082 176200 529116
rect 176234 529082 176245 529116
rect 176189 529026 176245 529082
rect 176275 529096 176331 529226
rect 176275 529062 176286 529096
rect 176320 529062 176331 529096
rect 176275 529026 176331 529062
rect 176361 529202 176417 529226
rect 176361 529168 176372 529202
rect 176406 529168 176417 529202
rect 176361 529116 176417 529168
rect 176361 529082 176372 529116
rect 176406 529082 176417 529116
rect 176361 529026 176417 529082
rect 176447 529096 176503 529226
rect 176447 529062 176458 529096
rect 176492 529062 176503 529096
rect 176447 529026 176503 529062
rect 176533 529202 176589 529226
rect 176533 529168 176544 529202
rect 176578 529168 176589 529202
rect 176533 529116 176589 529168
rect 176533 529082 176544 529116
rect 176578 529082 176589 529116
rect 176533 529026 176589 529082
rect 176619 529096 176674 529226
rect 176619 529062 176629 529096
rect 176663 529062 176674 529096
rect 176619 529026 176674 529062
rect 176704 529202 176760 529226
rect 176704 529168 176715 529202
rect 176749 529168 176760 529202
rect 176704 529116 176760 529168
rect 176704 529082 176715 529116
rect 176749 529082 176760 529116
rect 176704 529026 176760 529082
rect 176790 529096 176846 529226
rect 176790 529062 176801 529096
rect 176835 529062 176846 529096
rect 176790 529026 176846 529062
rect 176876 529202 176932 529226
rect 176876 529168 176887 529202
rect 176921 529168 176932 529202
rect 176876 529116 176932 529168
rect 176876 529082 176887 529116
rect 176921 529082 176932 529116
rect 176876 529026 176932 529082
rect 176962 529096 177018 529226
rect 176962 529062 176973 529096
rect 177007 529062 177018 529096
rect 176962 529026 177018 529062
rect 177048 529202 177104 529226
rect 177048 529168 177059 529202
rect 177093 529168 177104 529202
rect 177048 529116 177104 529168
rect 177048 529082 177059 529116
rect 177093 529082 177104 529116
rect 177048 529026 177104 529082
rect 177134 529096 177190 529226
rect 177134 529062 177145 529096
rect 177179 529062 177190 529096
rect 177134 529026 177190 529062
rect 177220 529202 177276 529226
rect 177220 529168 177231 529202
rect 177265 529168 177276 529202
rect 177220 529116 177276 529168
rect 177220 529082 177231 529116
rect 177265 529082 177276 529116
rect 177220 529026 177276 529082
rect 177306 529140 177362 529226
rect 177306 529106 177317 529140
rect 177351 529106 177362 529140
rect 177306 529072 177362 529106
rect 177306 529038 177317 529072
rect 177351 529038 177362 529072
rect 177306 529026 177362 529038
rect 177392 529156 177448 529226
rect 177392 529122 177403 529156
rect 177437 529122 177448 529156
rect 177392 529088 177448 529122
rect 177392 529054 177403 529088
rect 177437 529054 177448 529088
rect 177392 529026 177448 529054
rect 177478 529140 177534 529226
rect 177478 529106 177489 529140
rect 177523 529106 177534 529140
rect 177478 529072 177534 529106
rect 177478 529038 177489 529072
rect 177523 529038 177534 529072
rect 177478 529026 177534 529038
rect 177564 529148 177620 529226
rect 177564 529114 177575 529148
rect 177609 529114 177620 529148
rect 177564 529080 177620 529114
rect 177564 529046 177575 529080
rect 177609 529046 177620 529080
rect 177564 529026 177620 529046
rect 177650 529140 177703 529226
rect 177650 529106 177661 529140
rect 177695 529106 177703 529140
rect 177650 529072 177703 529106
rect 177650 529038 177661 529072
rect 177695 529038 177703 529072
rect 177650 529026 177703 529038
rect 177757 529148 177809 529160
rect 177757 529114 177765 529148
rect 177799 529114 177809 529148
rect 177757 529080 177809 529114
rect 177757 529046 177765 529080
rect 177799 529046 177809 529080
rect 177757 529032 177809 529046
rect 177839 529096 177893 529160
rect 177839 529062 177849 529096
rect 177883 529062 177893 529096
rect 177839 529032 177893 529062
rect 177923 529148 177975 529160
rect 177923 529114 177933 529148
rect 177967 529114 177975 529148
rect 177923 529080 177975 529114
rect 177923 529046 177933 529080
rect 177967 529046 177975 529080
rect 177923 529032 177975 529046
rect 178108 529072 178160 529110
rect 178108 529038 178116 529072
rect 178150 529038 178160 529072
rect 178108 529026 178160 529038
rect 178190 529080 178252 529110
rect 178190 529046 178200 529080
rect 178234 529046 178252 529080
rect 178190 529026 178252 529046
rect 178282 529074 178351 529110
rect 178282 529040 178293 529074
rect 178327 529040 178351 529074
rect 178282 529026 178351 529040
rect 178381 529098 178491 529110
rect 178381 529064 178447 529098
rect 178481 529064 178491 529098
rect 178381 529026 178491 529064
rect 178521 529082 178588 529110
rect 178521 529048 178544 529082
rect 178578 529048 178588 529082
rect 178521 529026 178588 529048
rect 178618 529098 178670 529110
rect 178618 529064 178628 529098
rect 178662 529064 178670 529098
rect 178618 529026 178670 529064
rect 178733 529072 178785 529194
rect 178733 529038 178741 529072
rect 178775 529038 178785 529072
rect 178733 529026 178785 529038
rect 178815 529110 178869 529194
rect 179411 529154 179461 529226
rect 179395 529140 179461 529154
rect 178815 529080 178884 529110
rect 178815 529046 178829 529080
rect 178863 529046 178884 529080
rect 178815 529026 178884 529046
rect 178914 529073 178970 529110
rect 178914 529039 178926 529073
rect 178960 529039 178970 529073
rect 178914 529026 178970 529039
rect 179000 529026 179054 529110
rect 179084 529072 179162 529110
rect 179084 529038 179118 529072
rect 179152 529038 179162 529072
rect 179084 529026 179162 529038
rect 179192 529098 179246 529110
rect 179192 529064 179202 529098
rect 179236 529064 179246 529098
rect 179192 529026 179246 529064
rect 179276 529072 179330 529110
rect 179276 529038 179288 529072
rect 179322 529038 179330 529072
rect 179276 529026 179330 529038
rect 179395 529106 179417 529140
rect 179451 529106 179461 529140
rect 179395 529072 179461 529106
rect 179395 529038 179417 529072
rect 179451 529038 179461 529072
rect 179395 529026 179461 529038
rect 179491 529176 179543 529226
rect 179491 529142 179501 529176
rect 179535 529142 179543 529176
rect 179491 529108 179543 529142
rect 179491 529074 179501 529108
rect 179535 529074 179543 529108
rect 179491 529026 179543 529074
rect 179689 529148 179741 529184
rect 179689 529114 179697 529148
rect 179731 529114 179741 529148
rect 179689 529080 179741 529114
rect 179689 529046 179697 529080
rect 179731 529046 179741 529080
rect 179689 529026 179741 529046
rect 179771 529148 179829 529184
rect 179771 529114 179783 529148
rect 179817 529114 179829 529148
rect 179771 529080 179829 529114
rect 179771 529046 179783 529080
rect 179817 529046 179829 529080
rect 179771 529026 179829 529046
rect 179859 529161 179911 529184
rect 179859 529127 179869 529161
rect 179903 529127 179911 529161
rect 179859 529080 179911 529127
rect 179859 529046 179869 529080
rect 179903 529046 179911 529080
rect 179859 529026 179911 529046
rect 180057 529174 180109 529200
rect 180057 529140 180065 529174
rect 180099 529140 180109 529174
rect 180057 529072 180109 529140
rect 180057 529038 180065 529072
rect 180099 529038 180109 529072
rect 180057 529026 180109 529038
rect 180503 529174 180555 529200
rect 180503 529140 180513 529174
rect 180547 529140 180555 529174
rect 180503 529072 180555 529140
rect 180503 529038 180513 529072
rect 180547 529038 180555 529072
rect 180503 529026 180555 529038
rect 180701 529140 180754 529226
rect 180701 529106 180709 529140
rect 180743 529106 180754 529140
rect 180701 529072 180754 529106
rect 180701 529038 180709 529072
rect 180743 529038 180754 529072
rect 180701 529026 180754 529038
rect 180784 529148 180840 529226
rect 180784 529114 180795 529148
rect 180829 529114 180840 529148
rect 180784 529080 180840 529114
rect 180784 529046 180795 529080
rect 180829 529046 180840 529080
rect 180784 529026 180840 529046
rect 180870 529140 180926 529226
rect 180870 529106 180881 529140
rect 180915 529106 180926 529140
rect 180870 529072 180926 529106
rect 180870 529038 180881 529072
rect 180915 529038 180926 529072
rect 180870 529026 180926 529038
rect 180956 529156 181012 529226
rect 180956 529122 180967 529156
rect 181001 529122 181012 529156
rect 180956 529088 181012 529122
rect 180956 529054 180967 529088
rect 181001 529054 181012 529088
rect 180956 529026 181012 529054
rect 181042 529140 181098 529226
rect 181042 529106 181053 529140
rect 181087 529106 181098 529140
rect 181042 529072 181098 529106
rect 181042 529038 181053 529072
rect 181087 529038 181098 529072
rect 181042 529026 181098 529038
rect 181128 529202 181184 529226
rect 181128 529168 181139 529202
rect 181173 529168 181184 529202
rect 181128 529116 181184 529168
rect 181128 529082 181139 529116
rect 181173 529082 181184 529116
rect 181128 529026 181184 529082
rect 181214 529096 181270 529226
rect 181214 529062 181225 529096
rect 181259 529062 181270 529096
rect 181214 529026 181270 529062
rect 181300 529202 181356 529226
rect 181300 529168 181311 529202
rect 181345 529168 181356 529202
rect 181300 529116 181356 529168
rect 181300 529082 181311 529116
rect 181345 529082 181356 529116
rect 181300 529026 181356 529082
rect 181386 529096 181442 529226
rect 181386 529062 181397 529096
rect 181431 529062 181442 529096
rect 181386 529026 181442 529062
rect 181472 529202 181528 529226
rect 181472 529168 181483 529202
rect 181517 529168 181528 529202
rect 181472 529116 181528 529168
rect 181472 529082 181483 529116
rect 181517 529082 181528 529116
rect 181472 529026 181528 529082
rect 181558 529096 181614 529226
rect 181558 529062 181569 529096
rect 181603 529062 181614 529096
rect 181558 529026 181614 529062
rect 181644 529202 181700 529226
rect 181644 529168 181655 529202
rect 181689 529168 181700 529202
rect 181644 529116 181700 529168
rect 181644 529082 181655 529116
rect 181689 529082 181700 529116
rect 181644 529026 181700 529082
rect 181730 529096 181785 529226
rect 181730 529062 181741 529096
rect 181775 529062 181785 529096
rect 181730 529026 181785 529062
rect 181815 529202 181871 529226
rect 181815 529168 181826 529202
rect 181860 529168 181871 529202
rect 181815 529116 181871 529168
rect 181815 529082 181826 529116
rect 181860 529082 181871 529116
rect 181815 529026 181871 529082
rect 181901 529096 181957 529226
rect 181901 529062 181912 529096
rect 181946 529062 181957 529096
rect 181901 529026 181957 529062
rect 181987 529202 182043 529226
rect 181987 529168 181998 529202
rect 182032 529168 182043 529202
rect 181987 529116 182043 529168
rect 181987 529082 181998 529116
rect 182032 529082 182043 529116
rect 181987 529026 182043 529082
rect 182073 529096 182129 529226
rect 182073 529062 182084 529096
rect 182118 529062 182129 529096
rect 182073 529026 182129 529062
rect 182159 529202 182215 529226
rect 182159 529168 182170 529202
rect 182204 529168 182215 529202
rect 182159 529116 182215 529168
rect 182159 529082 182170 529116
rect 182204 529082 182215 529116
rect 182159 529026 182215 529082
rect 182245 529096 182301 529226
rect 182245 529062 182256 529096
rect 182290 529062 182301 529096
rect 182245 529026 182301 529062
rect 182331 529202 182387 529226
rect 182331 529168 182342 529202
rect 182376 529168 182387 529202
rect 182331 529116 182387 529168
rect 182331 529082 182342 529116
rect 182376 529082 182387 529116
rect 182331 529026 182387 529082
rect 182417 529096 182470 529226
rect 182417 529062 182428 529096
rect 182462 529062 182470 529096
rect 182417 529026 182470 529062
rect 182541 529161 182593 529184
rect 182541 529127 182549 529161
rect 182583 529127 182593 529161
rect 182541 529080 182593 529127
rect 182541 529046 182549 529080
rect 182583 529046 182593 529080
rect 182541 529026 182593 529046
rect 182623 529148 182681 529184
rect 182623 529114 182635 529148
rect 182669 529114 182681 529148
rect 182623 529080 182681 529114
rect 182623 529046 182635 529080
rect 182669 529046 182681 529080
rect 182623 529026 182681 529046
rect 182711 529148 182763 529184
rect 182711 529114 182721 529148
rect 182755 529114 182763 529148
rect 182711 529080 182763 529114
rect 182711 529046 182721 529080
rect 182755 529046 182763 529080
rect 182711 529026 182763 529046
rect 182817 529072 182869 529200
rect 182817 529038 182825 529072
rect 182859 529038 182869 529072
rect 182817 529026 182869 529038
rect 183815 529072 183867 529200
rect 183815 529038 183825 529072
rect 183859 529038 183867 529072
rect 183815 529026 183867 529038
rect 183921 529072 183973 529200
rect 183921 529038 183929 529072
rect 183963 529038 183973 529072
rect 183921 529026 183973 529038
rect 184919 529072 184971 529200
rect 184919 529038 184929 529072
rect 184963 529038 184971 529072
rect 185209 529072 185261 529200
rect 184919 529026 184971 529038
rect 185209 529038 185217 529072
rect 185251 529038 185261 529072
rect 185209 529026 185261 529038
rect 186207 529072 186259 529200
rect 186207 529038 186217 529072
rect 186251 529038 186259 529072
rect 186207 529026 186259 529038
rect 186313 529174 186365 529200
rect 186313 529140 186321 529174
rect 186355 529140 186365 529174
rect 186313 529072 186365 529140
rect 186313 529038 186321 529072
rect 186355 529038 186365 529072
rect 186313 529026 186365 529038
rect 186943 529174 186995 529200
rect 186943 529140 186953 529174
rect 186987 529140 186995 529174
rect 186943 529072 186995 529140
rect 186943 529038 186953 529072
rect 186987 529038 186995 529072
rect 186943 529026 186995 529038
rect 187233 529167 187285 529200
rect 187233 529133 187241 529167
rect 187275 529133 187285 529167
rect 187233 529072 187285 529133
rect 187233 529038 187241 529072
rect 187275 529038 187285 529072
rect 187233 529026 187285 529038
rect 187403 529167 187455 529200
rect 187403 529133 187413 529167
rect 187447 529133 187455 529167
rect 187403 529072 187455 529133
rect 187403 529038 187413 529072
rect 187447 529038 187455 529072
rect 187403 529026 187455 529038
rect 172237 528920 172289 528932
rect 172237 528886 172245 528920
rect 172279 528886 172289 528920
rect 172237 528825 172289 528886
rect 172237 528791 172245 528825
rect 172279 528791 172289 528825
rect 172237 528758 172289 528791
rect 172407 528920 172459 528932
rect 172407 528886 172417 528920
rect 172451 528886 172459 528920
rect 172407 528825 172459 528886
rect 172407 528791 172417 528825
rect 172451 528791 172459 528825
rect 172407 528758 172459 528791
rect 172513 528920 172565 528932
rect 172513 528886 172521 528920
rect 172555 528886 172565 528920
rect 172513 528758 172565 528886
rect 173511 528920 173563 528932
rect 173511 528886 173521 528920
rect 173555 528886 173563 528920
rect 173511 528758 173563 528886
rect 173617 528920 173669 528932
rect 173617 528886 173625 528920
rect 173659 528886 173669 528920
rect 173617 528758 173669 528886
rect 174615 528920 174667 528932
rect 174615 528886 174625 528920
rect 174659 528886 174667 528920
rect 174615 528758 174667 528886
rect 174721 528920 174773 528932
rect 174721 528886 174729 528920
rect 174763 528886 174773 528920
rect 174721 528758 174773 528886
rect 175719 528920 175771 528932
rect 175719 528886 175729 528920
rect 175763 528886 175771 528920
rect 175719 528758 175771 528886
rect 175917 528912 175969 528932
rect 175917 528878 175925 528912
rect 175959 528878 175969 528912
rect 175917 528844 175969 528878
rect 175917 528810 175925 528844
rect 175959 528810 175969 528844
rect 175917 528774 175969 528810
rect 175999 528912 176057 528932
rect 175999 528878 176011 528912
rect 176045 528878 176057 528912
rect 175999 528844 176057 528878
rect 175999 528810 176011 528844
rect 176045 528810 176057 528844
rect 175999 528774 176057 528810
rect 176087 528912 176139 528932
rect 176087 528878 176097 528912
rect 176131 528878 176139 528912
rect 176087 528831 176139 528878
rect 176087 528797 176097 528831
rect 176131 528797 176139 528831
rect 176087 528774 176139 528797
rect 176193 528912 176245 528932
rect 176193 528878 176201 528912
rect 176235 528878 176245 528912
rect 176193 528844 176245 528878
rect 176193 528810 176201 528844
rect 176235 528810 176245 528844
rect 176193 528774 176245 528810
rect 176275 528912 176333 528932
rect 176275 528878 176287 528912
rect 176321 528878 176333 528912
rect 176275 528844 176333 528878
rect 176275 528810 176287 528844
rect 176321 528810 176333 528844
rect 176275 528774 176333 528810
rect 176363 528912 176415 528932
rect 177109 528920 177161 528932
rect 176363 528878 176373 528912
rect 176407 528878 176415 528912
rect 177109 528893 177117 528920
rect 176363 528831 176415 528878
rect 176363 528797 176373 528831
rect 176407 528797 176415 528831
rect 176511 528860 176567 528893
rect 176511 528826 176523 528860
rect 176557 528826 176567 528860
rect 176511 528809 176567 528826
rect 176597 528860 176663 528893
rect 176597 528826 176609 528860
rect 176643 528826 176663 528860
rect 176597 528809 176663 528826
rect 176693 528809 176735 528893
rect 176765 528860 176949 528893
rect 176765 528826 176806 528860
rect 176840 528826 176881 528860
rect 176915 528826 176949 528860
rect 176765 528809 176949 528826
rect 176979 528809 177052 528893
rect 177082 528886 177117 528893
rect 177151 528886 177161 528920
rect 177082 528852 177161 528886
rect 177082 528818 177117 528852
rect 177151 528818 177161 528852
rect 177082 528809 177161 528818
rect 176363 528774 176415 528797
rect 177109 528784 177161 528809
rect 177109 528750 177117 528784
rect 177151 528750 177161 528784
rect 177109 528732 177161 528750
rect 177191 528920 177243 528932
rect 177191 528886 177201 528920
rect 177235 528886 177243 528920
rect 177191 528852 177243 528886
rect 177191 528818 177201 528852
rect 177235 528818 177243 528852
rect 177191 528784 177243 528818
rect 177191 528750 177201 528784
rect 177235 528750 177243 528784
rect 177191 528732 177243 528750
rect 177500 528894 177552 528932
rect 177500 528860 177508 528894
rect 177542 528860 177552 528894
rect 177500 528732 177552 528860
rect 177582 528920 177647 528932
rect 177582 528886 177598 528920
rect 177632 528886 177647 528920
rect 177582 528848 177647 528886
rect 177747 528894 177799 528932
rect 177747 528860 177757 528894
rect 177791 528860 177799 528894
rect 177747 528848 177799 528860
rect 177853 528894 177905 528932
rect 177853 528860 177861 528894
rect 177895 528860 177905 528894
rect 177853 528848 177905 528860
rect 178005 528920 178059 528932
rect 178005 528886 178015 528920
rect 178049 528886 178059 528920
rect 178005 528848 178059 528886
rect 178089 528894 178141 528932
rect 178089 528860 178099 528894
rect 178133 528860 178141 528894
rect 178089 528848 178141 528860
rect 178401 528920 178454 528932
rect 178401 528886 178409 528920
rect 178443 528886 178454 528920
rect 178401 528852 178454 528886
rect 177582 528732 177632 528848
rect 178401 528818 178409 528852
rect 178443 528818 178454 528852
rect 178401 528732 178454 528818
rect 178484 528912 178540 528932
rect 178484 528878 178495 528912
rect 178529 528878 178540 528912
rect 178484 528844 178540 528878
rect 178484 528810 178495 528844
rect 178529 528810 178540 528844
rect 178484 528732 178540 528810
rect 178570 528920 178626 528932
rect 178570 528886 178581 528920
rect 178615 528886 178626 528920
rect 178570 528852 178626 528886
rect 178570 528818 178581 528852
rect 178615 528818 178626 528852
rect 178570 528732 178626 528818
rect 178656 528904 178712 528932
rect 178656 528870 178667 528904
rect 178701 528870 178712 528904
rect 178656 528836 178712 528870
rect 178656 528802 178667 528836
rect 178701 528802 178712 528836
rect 178656 528732 178712 528802
rect 178742 528920 178798 528932
rect 178742 528886 178753 528920
rect 178787 528886 178798 528920
rect 178742 528852 178798 528886
rect 178742 528818 178753 528852
rect 178787 528818 178798 528852
rect 178742 528732 178798 528818
rect 178828 528876 178884 528932
rect 178828 528842 178839 528876
rect 178873 528842 178884 528876
rect 178828 528790 178884 528842
rect 178828 528756 178839 528790
rect 178873 528756 178884 528790
rect 178828 528732 178884 528756
rect 178914 528896 178970 528932
rect 178914 528862 178925 528896
rect 178959 528862 178970 528896
rect 178914 528732 178970 528862
rect 179000 528876 179056 528932
rect 179000 528842 179011 528876
rect 179045 528842 179056 528876
rect 179000 528790 179056 528842
rect 179000 528756 179011 528790
rect 179045 528756 179056 528790
rect 179000 528732 179056 528756
rect 179086 528896 179142 528932
rect 179086 528862 179097 528896
rect 179131 528862 179142 528896
rect 179086 528732 179142 528862
rect 179172 528876 179228 528932
rect 179172 528842 179183 528876
rect 179217 528842 179228 528876
rect 179172 528790 179228 528842
rect 179172 528756 179183 528790
rect 179217 528756 179228 528790
rect 179172 528732 179228 528756
rect 179258 528896 179314 528932
rect 179258 528862 179269 528896
rect 179303 528862 179314 528896
rect 179258 528732 179314 528862
rect 179344 528876 179400 528932
rect 179344 528842 179355 528876
rect 179389 528842 179400 528876
rect 179344 528790 179400 528842
rect 179344 528756 179355 528790
rect 179389 528756 179400 528790
rect 179344 528732 179400 528756
rect 179430 528896 179485 528932
rect 179430 528862 179441 528896
rect 179475 528862 179485 528896
rect 179430 528732 179485 528862
rect 179515 528876 179571 528932
rect 179515 528842 179526 528876
rect 179560 528842 179571 528876
rect 179515 528790 179571 528842
rect 179515 528756 179526 528790
rect 179560 528756 179571 528790
rect 179515 528732 179571 528756
rect 179601 528896 179657 528932
rect 179601 528862 179612 528896
rect 179646 528862 179657 528896
rect 179601 528732 179657 528862
rect 179687 528876 179743 528932
rect 179687 528842 179698 528876
rect 179732 528842 179743 528876
rect 179687 528790 179743 528842
rect 179687 528756 179698 528790
rect 179732 528756 179743 528790
rect 179687 528732 179743 528756
rect 179773 528896 179829 528932
rect 179773 528862 179784 528896
rect 179818 528862 179829 528896
rect 179773 528732 179829 528862
rect 179859 528876 179915 528932
rect 179859 528842 179870 528876
rect 179904 528842 179915 528876
rect 179859 528790 179915 528842
rect 179859 528756 179870 528790
rect 179904 528756 179915 528790
rect 179859 528732 179915 528756
rect 179945 528896 180001 528932
rect 179945 528862 179956 528896
rect 179990 528862 180001 528896
rect 179945 528732 180001 528862
rect 180031 528876 180087 528932
rect 180031 528842 180042 528876
rect 180076 528842 180087 528876
rect 180031 528790 180087 528842
rect 180031 528756 180042 528790
rect 180076 528756 180087 528790
rect 180031 528732 180087 528756
rect 180117 528896 180170 528932
rect 180117 528862 180128 528896
rect 180162 528862 180170 528896
rect 180117 528732 180170 528862
rect 180241 528912 180293 528932
rect 180241 528878 180249 528912
rect 180283 528878 180293 528912
rect 180241 528844 180293 528878
rect 180241 528810 180249 528844
rect 180283 528810 180293 528844
rect 180241 528774 180293 528810
rect 180323 528912 180381 528932
rect 180323 528878 180335 528912
rect 180369 528878 180381 528912
rect 180323 528844 180381 528878
rect 180323 528810 180335 528844
rect 180369 528810 180381 528844
rect 180323 528774 180381 528810
rect 180411 528912 180463 528932
rect 180411 528878 180421 528912
rect 180455 528878 180463 528912
rect 180411 528831 180463 528878
rect 180411 528797 180421 528831
rect 180455 528797 180463 528831
rect 180517 528912 180569 528926
rect 180517 528878 180525 528912
rect 180559 528878 180569 528912
rect 180517 528844 180569 528878
rect 180517 528810 180525 528844
rect 180559 528810 180569 528844
rect 180517 528798 180569 528810
rect 180599 528896 180653 528926
rect 180599 528862 180609 528896
rect 180643 528862 180653 528896
rect 180599 528798 180653 528862
rect 180683 528912 180735 528926
rect 180683 528878 180693 528912
rect 180727 528878 180735 528912
rect 180683 528844 180735 528878
rect 180868 528920 180920 528932
rect 180868 528886 180876 528920
rect 180910 528886 180920 528920
rect 180868 528848 180920 528886
rect 180950 528912 181012 528932
rect 180950 528878 180960 528912
rect 180994 528878 181012 528912
rect 180950 528848 181012 528878
rect 181042 528918 181111 528932
rect 181042 528884 181053 528918
rect 181087 528884 181111 528918
rect 181042 528848 181111 528884
rect 181141 528894 181251 528932
rect 181141 528860 181207 528894
rect 181241 528860 181251 528894
rect 181141 528848 181251 528860
rect 181281 528910 181348 528932
rect 181281 528876 181304 528910
rect 181338 528876 181348 528910
rect 181281 528848 181348 528876
rect 181378 528894 181430 528932
rect 181378 528860 181388 528894
rect 181422 528860 181430 528894
rect 181378 528848 181430 528860
rect 181493 528920 181545 528932
rect 181493 528886 181501 528920
rect 181535 528886 181545 528920
rect 180683 528810 180693 528844
rect 180727 528810 180735 528844
rect 180683 528798 180735 528810
rect 180411 528774 180463 528797
rect 181493 528764 181545 528886
rect 181575 528912 181644 528932
rect 181575 528878 181589 528912
rect 181623 528878 181644 528912
rect 181575 528848 181644 528878
rect 181674 528919 181730 528932
rect 181674 528885 181686 528919
rect 181720 528885 181730 528919
rect 181674 528848 181730 528885
rect 181760 528848 181814 528932
rect 181844 528920 181922 528932
rect 181844 528886 181878 528920
rect 181912 528886 181922 528920
rect 181844 528848 181922 528886
rect 181952 528894 182006 528932
rect 181952 528860 181962 528894
rect 181996 528860 182006 528894
rect 181952 528848 182006 528860
rect 182036 528920 182090 528932
rect 182036 528886 182048 528920
rect 182082 528886 182090 528920
rect 182036 528848 182090 528886
rect 182155 528920 182221 528932
rect 182155 528886 182177 528920
rect 182211 528886 182221 528920
rect 182155 528852 182221 528886
rect 181575 528764 181629 528848
rect 182155 528818 182177 528852
rect 182211 528818 182221 528852
rect 182155 528804 182221 528818
rect 182171 528732 182221 528804
rect 182251 528884 182303 528932
rect 182633 528920 182685 528932
rect 182251 528850 182261 528884
rect 182295 528850 182303 528884
rect 182251 528816 182303 528850
rect 182251 528782 182261 528816
rect 182295 528782 182303 528816
rect 182251 528732 182303 528782
rect 182633 528886 182641 528920
rect 182675 528886 182685 528920
rect 182633 528758 182685 528886
rect 183631 528920 183683 528932
rect 183631 528886 183641 528920
rect 183675 528886 183683 528920
rect 183631 528758 183683 528886
rect 183737 528920 183789 528932
rect 183737 528886 183745 528920
rect 183779 528886 183789 528920
rect 183737 528758 183789 528886
rect 184735 528920 184787 528932
rect 184735 528886 184745 528920
rect 184779 528886 184787 528920
rect 184735 528758 184787 528886
rect 184841 528920 184893 528932
rect 184841 528886 184849 528920
rect 184883 528886 184893 528920
rect 184841 528758 184893 528886
rect 185839 528920 185891 528932
rect 185839 528886 185849 528920
rect 185883 528886 185891 528920
rect 185839 528758 185891 528886
rect 185945 528920 185997 528932
rect 185945 528886 185953 528920
rect 185987 528886 185997 528920
rect 185945 528758 185997 528886
rect 186943 528920 186995 528932
rect 186943 528886 186953 528920
rect 186987 528886 186995 528920
rect 186943 528758 186995 528886
rect 187233 528920 187285 528932
rect 187233 528886 187241 528920
rect 187275 528886 187285 528920
rect 187233 528825 187285 528886
rect 187233 528791 187241 528825
rect 187275 528791 187285 528825
rect 187233 528758 187285 528791
rect 187403 528920 187455 528932
rect 187403 528886 187413 528920
rect 187447 528886 187455 528920
rect 187403 528825 187455 528886
rect 187403 528791 187413 528825
rect 187447 528791 187455 528825
rect 187403 528758 187455 528791
rect 172237 528079 172289 528112
rect 172237 528045 172245 528079
rect 172279 528045 172289 528079
rect 172237 527984 172289 528045
rect 172237 527950 172245 527984
rect 172279 527950 172289 527984
rect 172237 527938 172289 527950
rect 172407 528079 172459 528112
rect 172407 528045 172417 528079
rect 172451 528045 172459 528079
rect 172407 527984 172459 528045
rect 172407 527950 172417 527984
rect 172451 527950 172459 527984
rect 172407 527938 172459 527950
rect 172513 527984 172565 528112
rect 172513 527950 172521 527984
rect 172555 527950 172565 527984
rect 172513 527938 172565 527950
rect 173511 527984 173563 528112
rect 173511 527950 173521 527984
rect 173555 527950 173563 527984
rect 173511 527938 173563 527950
rect 173617 527984 173669 528112
rect 173617 527950 173625 527984
rect 173659 527950 173669 527984
rect 173617 527938 173669 527950
rect 174615 527984 174667 528112
rect 174615 527950 174625 527984
rect 174659 527950 174667 527984
rect 174905 527984 174957 528112
rect 174615 527938 174667 527950
rect 174905 527950 174913 527984
rect 174947 527950 174957 527984
rect 174905 527938 174957 527950
rect 175903 527984 175955 528112
rect 175903 527950 175913 527984
rect 175947 527950 175955 527984
rect 175903 527938 175955 527950
rect 176101 528060 176153 528072
rect 176101 528026 176109 528060
rect 176143 528026 176153 528060
rect 176101 527992 176153 528026
rect 176101 527958 176109 527992
rect 176143 527958 176153 527992
rect 176101 527944 176153 527958
rect 176183 528008 176237 528072
rect 176183 527974 176193 528008
rect 176227 527974 176237 528008
rect 176183 527944 176237 527974
rect 176267 528060 176319 528072
rect 176267 528026 176277 528060
rect 176311 528026 176319 528060
rect 176267 527992 176319 528026
rect 176267 527958 176277 527992
rect 176311 527958 176319 527992
rect 176267 527944 176319 527958
rect 176452 527984 176504 528022
rect 176452 527950 176460 527984
rect 176494 527950 176504 527984
rect 176452 527938 176504 527950
rect 176534 527992 176596 528022
rect 176534 527958 176544 527992
rect 176578 527958 176596 527992
rect 176534 527938 176596 527958
rect 176626 527986 176695 528022
rect 176626 527952 176637 527986
rect 176671 527952 176695 527986
rect 176626 527938 176695 527952
rect 176725 528010 176835 528022
rect 176725 527976 176791 528010
rect 176825 527976 176835 528010
rect 176725 527938 176835 527976
rect 176865 527994 176932 528022
rect 176865 527960 176888 527994
rect 176922 527960 176932 527994
rect 176865 527938 176932 527960
rect 176962 528010 177014 528022
rect 176962 527976 176972 528010
rect 177006 527976 177014 528010
rect 176962 527938 177014 527976
rect 177077 527984 177129 528106
rect 177077 527950 177085 527984
rect 177119 527950 177129 527984
rect 177077 527938 177129 527950
rect 177159 528022 177213 528106
rect 177755 528066 177805 528138
rect 177739 528052 177805 528066
rect 177159 527992 177228 528022
rect 177159 527958 177173 527992
rect 177207 527958 177228 527992
rect 177159 527938 177228 527958
rect 177258 527985 177314 528022
rect 177258 527951 177270 527985
rect 177304 527951 177314 527985
rect 177258 527938 177314 527951
rect 177344 527938 177398 528022
rect 177428 527984 177506 528022
rect 177428 527950 177462 527984
rect 177496 527950 177506 527984
rect 177428 527938 177506 527950
rect 177536 528010 177590 528022
rect 177536 527976 177546 528010
rect 177580 527976 177590 528010
rect 177536 527938 177590 527976
rect 177620 527984 177674 528022
rect 177620 527950 177632 527984
rect 177666 527950 177674 527984
rect 177620 527938 177674 527950
rect 177739 528018 177761 528052
rect 177795 528018 177805 528052
rect 177739 527984 177805 528018
rect 177739 527950 177761 527984
rect 177795 527950 177805 527984
rect 177739 527938 177805 527950
rect 177835 528088 177887 528138
rect 178953 528120 179005 528138
rect 177835 528054 177845 528088
rect 177879 528054 177887 528088
rect 177835 528020 177887 528054
rect 177835 527986 177845 528020
rect 177879 527986 177887 528020
rect 177835 527938 177887 527986
rect 177941 528073 177993 528096
rect 177941 528039 177949 528073
rect 177983 528039 177993 528073
rect 177941 527992 177993 528039
rect 177941 527958 177949 527992
rect 177983 527958 177993 527992
rect 177941 527938 177993 527958
rect 178023 528060 178081 528096
rect 178023 528026 178035 528060
rect 178069 528026 178081 528060
rect 178023 527992 178081 528026
rect 178023 527958 178035 527992
rect 178069 527958 178081 527992
rect 178023 527938 178081 527958
rect 178111 528060 178163 528096
rect 178111 528026 178121 528060
rect 178155 528026 178163 528060
rect 178111 527992 178163 528026
rect 178111 527958 178121 527992
rect 178155 527958 178163 527992
rect 178111 527938 178163 527958
rect 178217 528086 178269 528112
rect 178217 528052 178225 528086
rect 178259 528052 178269 528086
rect 178217 527984 178269 528052
rect 178217 527950 178225 527984
rect 178259 527950 178269 527984
rect 178217 527938 178269 527950
rect 178847 528086 178899 528112
rect 178847 528052 178857 528086
rect 178891 528052 178899 528086
rect 178847 527984 178899 528052
rect 178847 527950 178857 527984
rect 178891 527950 178899 527984
rect 178847 527938 178899 527950
rect 178953 528086 178961 528120
rect 178995 528086 179005 528120
rect 178953 528052 179005 528086
rect 178953 528018 178961 528052
rect 178995 528018 179005 528052
rect 178953 527984 179005 528018
rect 178953 527950 178961 527984
rect 178995 527950 179005 527984
rect 178953 527938 179005 527950
rect 179035 528120 179087 528138
rect 179035 528086 179045 528120
rect 179079 528086 179087 528120
rect 179035 528061 179087 528086
rect 180977 528120 181029 528138
rect 179035 528052 179114 528061
rect 179035 528018 179045 528052
rect 179079 528018 179114 528052
rect 179035 527984 179114 528018
rect 179035 527950 179045 527984
rect 179079 527977 179114 527984
rect 179144 527977 179217 528061
rect 179247 528044 179431 528061
rect 179247 528010 179281 528044
rect 179315 528010 179356 528044
rect 179390 528010 179431 528044
rect 179247 527977 179431 528010
rect 179461 527977 179503 528061
rect 179533 528044 179599 528061
rect 179533 528010 179553 528044
rect 179587 528010 179599 528044
rect 179533 527977 179599 528010
rect 179629 528044 179685 528061
rect 179629 528010 179639 528044
rect 179673 528010 179685 528044
rect 179629 527977 179685 528010
rect 179079 527950 179087 527977
rect 180057 528086 180109 528112
rect 180057 528052 180065 528086
rect 180099 528052 180109 528086
rect 180057 527984 180109 528052
rect 179035 527938 179087 527950
rect 180057 527950 180065 527984
rect 180099 527950 180109 527984
rect 180057 527938 180109 527950
rect 180687 528086 180739 528112
rect 180687 528052 180697 528086
rect 180731 528052 180739 528086
rect 180687 527984 180739 528052
rect 180687 527950 180697 527984
rect 180731 527950 180739 527984
rect 180687 527938 180739 527950
rect 180977 528086 180985 528120
rect 181019 528086 181029 528120
rect 180977 528052 181029 528086
rect 180977 528018 180985 528052
rect 181019 528018 181029 528052
rect 180977 527984 181029 528018
rect 180977 527950 180985 527984
rect 181019 527950 181029 527984
rect 180977 527938 181029 527950
rect 181059 528120 181111 528138
rect 181059 528086 181069 528120
rect 181103 528086 181111 528120
rect 181059 528061 181111 528086
rect 181059 528052 181138 528061
rect 181059 528018 181069 528052
rect 181103 528018 181138 528052
rect 181059 527984 181138 528018
rect 181059 527950 181069 527984
rect 181103 527977 181138 527984
rect 181168 527977 181241 528061
rect 181271 528044 181455 528061
rect 181271 528010 181305 528044
rect 181339 528010 181380 528044
rect 181414 528010 181455 528044
rect 181271 527977 181455 528010
rect 181485 527977 181527 528061
rect 181557 528044 181623 528061
rect 181557 528010 181577 528044
rect 181611 528010 181623 528044
rect 181557 527977 181623 528010
rect 181653 528044 181709 528061
rect 181653 528010 181663 528044
rect 181697 528010 181709 528044
rect 181653 527977 181709 528010
rect 181805 527984 181857 528112
rect 181103 527950 181111 527977
rect 181059 527938 181111 527950
rect 181805 527950 181813 527984
rect 181847 527950 181857 527984
rect 181805 527938 181857 527950
rect 182803 527984 182855 528112
rect 182803 527950 182813 527984
rect 182847 527950 182855 527984
rect 182803 527938 182855 527950
rect 182909 527984 182961 528112
rect 182909 527950 182917 527984
rect 182951 527950 182961 527984
rect 182909 527938 182961 527950
rect 183907 527984 183959 528112
rect 183907 527950 183917 527984
rect 183951 527950 183959 527984
rect 183907 527938 183959 527950
rect 184013 527984 184065 528112
rect 184013 527950 184021 527984
rect 184055 527950 184065 527984
rect 184013 527938 184065 527950
rect 185011 527984 185063 528112
rect 185011 527950 185021 527984
rect 185055 527950 185063 527984
rect 185209 527984 185261 528112
rect 185011 527938 185063 527950
rect 185209 527950 185217 527984
rect 185251 527950 185261 527984
rect 185209 527938 185261 527950
rect 186207 527984 186259 528112
rect 186207 527950 186217 527984
rect 186251 527950 186259 527984
rect 186207 527938 186259 527950
rect 186313 528086 186365 528112
rect 186313 528052 186321 528086
rect 186355 528052 186365 528086
rect 186313 527984 186365 528052
rect 186313 527950 186321 527984
rect 186355 527950 186365 527984
rect 186313 527938 186365 527950
rect 186943 528086 186995 528112
rect 186943 528052 186953 528086
rect 186987 528052 186995 528086
rect 186943 527984 186995 528052
rect 186943 527950 186953 527984
rect 186987 527950 186995 527984
rect 186943 527938 186995 527950
rect 187233 528079 187285 528112
rect 187233 528045 187241 528079
rect 187275 528045 187285 528079
rect 187233 527984 187285 528045
rect 187233 527950 187241 527984
rect 187275 527950 187285 527984
rect 187233 527938 187285 527950
rect 187403 528079 187455 528112
rect 187403 528045 187413 528079
rect 187447 528045 187455 528079
rect 187403 527984 187455 528045
rect 187403 527950 187413 527984
rect 187447 527950 187455 527984
rect 187403 527938 187455 527950
rect 172237 527832 172289 527844
rect 172237 527798 172245 527832
rect 172279 527798 172289 527832
rect 172237 527737 172289 527798
rect 172237 527703 172245 527737
rect 172279 527703 172289 527737
rect 172237 527670 172289 527703
rect 172407 527832 172459 527844
rect 172407 527798 172417 527832
rect 172451 527798 172459 527832
rect 172407 527737 172459 527798
rect 172407 527703 172417 527737
rect 172451 527703 172459 527737
rect 172407 527670 172459 527703
rect 172513 527832 172565 527844
rect 172513 527798 172521 527832
rect 172555 527798 172565 527832
rect 172513 527670 172565 527798
rect 173511 527832 173563 527844
rect 173511 527798 173521 527832
rect 173555 527798 173563 527832
rect 173511 527670 173563 527798
rect 173617 527832 173669 527844
rect 173617 527798 173625 527832
rect 173659 527798 173669 527832
rect 173617 527670 173669 527798
rect 174615 527832 174667 527844
rect 174615 527798 174625 527832
rect 174659 527798 174667 527832
rect 174615 527670 174667 527798
rect 174721 527832 174773 527844
rect 174721 527798 174729 527832
rect 174763 527798 174773 527832
rect 174721 527670 174773 527798
rect 175719 527832 175771 527844
rect 175719 527798 175729 527832
rect 175763 527798 175771 527832
rect 175719 527670 175771 527798
rect 175825 527832 175877 527844
rect 175825 527798 175833 527832
rect 175867 527798 175877 527832
rect 175825 527730 175877 527798
rect 175825 527696 175833 527730
rect 175867 527696 175877 527730
rect 175825 527670 175877 527696
rect 176271 527832 176323 527844
rect 176271 527798 176281 527832
rect 176315 527798 176323 527832
rect 176271 527730 176323 527798
rect 176271 527696 176281 527730
rect 176315 527696 176323 527730
rect 176271 527670 176323 527696
rect 176396 527806 176448 527844
rect 176396 527772 176404 527806
rect 176438 527772 176448 527806
rect 176396 527644 176448 527772
rect 176478 527832 176543 527844
rect 176478 527798 176494 527832
rect 176528 527798 176543 527832
rect 176478 527760 176543 527798
rect 176643 527806 176695 527844
rect 176643 527772 176653 527806
rect 176687 527772 176695 527806
rect 176643 527760 176695 527772
rect 176749 527806 176801 527844
rect 176749 527772 176757 527806
rect 176791 527772 176801 527806
rect 176749 527760 176801 527772
rect 176901 527832 176955 527844
rect 176901 527798 176911 527832
rect 176945 527798 176955 527832
rect 176901 527760 176955 527798
rect 176985 527806 177037 527844
rect 176985 527772 176995 527806
rect 177029 527772 177037 527806
rect 176985 527760 177037 527772
rect 177113 527832 177165 527844
rect 177113 527798 177121 527832
rect 177155 527798 177165 527832
rect 176478 527644 176528 527760
rect 177113 527737 177165 527798
rect 177113 527703 177121 527737
rect 177155 527703 177165 527737
rect 177113 527670 177165 527703
rect 177283 527832 177335 527844
rect 177283 527798 177293 527832
rect 177327 527798 177335 527832
rect 177481 527832 177533 527844
rect 177283 527737 177335 527798
rect 177283 527703 177293 527737
rect 177327 527703 177335 527737
rect 177283 527670 177335 527703
rect 177481 527798 177489 527832
rect 177523 527798 177533 527832
rect 177481 527670 177533 527798
rect 178479 527832 178531 527844
rect 178479 527798 178489 527832
rect 178523 527798 178531 527832
rect 178479 527670 178531 527798
rect 178585 527832 178637 527844
rect 178585 527798 178593 527832
rect 178627 527798 178637 527832
rect 178585 527730 178637 527798
rect 178585 527696 178593 527730
rect 178627 527696 178637 527730
rect 178585 527670 178637 527696
rect 178847 527832 178899 527844
rect 178847 527798 178857 527832
rect 178891 527798 178899 527832
rect 178847 527730 178899 527798
rect 178847 527696 178857 527730
rect 178891 527696 178899 527730
rect 178847 527670 178899 527696
rect 178972 527806 179024 527844
rect 178972 527772 178980 527806
rect 179014 527772 179024 527806
rect 178972 527644 179024 527772
rect 179054 527832 179119 527844
rect 179054 527798 179070 527832
rect 179104 527798 179119 527832
rect 179054 527760 179119 527798
rect 179219 527806 179271 527844
rect 179219 527772 179229 527806
rect 179263 527772 179271 527806
rect 179219 527760 179271 527772
rect 179325 527806 179377 527844
rect 179325 527772 179333 527806
rect 179367 527772 179377 527806
rect 179325 527760 179377 527772
rect 179477 527832 179531 527844
rect 179477 527798 179487 527832
rect 179521 527798 179531 527832
rect 179477 527760 179531 527798
rect 179561 527806 179613 527844
rect 179561 527772 179571 527806
rect 179605 527772 179613 527806
rect 179561 527760 179613 527772
rect 179689 527832 179741 527844
rect 179689 527798 179697 527832
rect 179731 527798 179741 527832
rect 179054 527644 179104 527760
rect 179689 527670 179741 527798
rect 180687 527832 180739 527844
rect 180687 527798 180697 527832
rect 180731 527798 180739 527832
rect 180687 527670 180739 527798
rect 180793 527832 180845 527844
rect 180793 527798 180801 527832
rect 180835 527798 180845 527832
rect 180793 527670 180845 527798
rect 181791 527832 181843 527844
rect 181791 527798 181801 527832
rect 181835 527798 181843 527832
rect 181791 527670 181843 527798
rect 181897 527832 181949 527844
rect 181897 527798 181905 527832
rect 181939 527798 181949 527832
rect 181897 527730 181949 527798
rect 181897 527696 181905 527730
rect 181939 527696 181949 527730
rect 181897 527670 181949 527696
rect 182343 527832 182395 527844
rect 182343 527798 182353 527832
rect 182387 527798 182395 527832
rect 182633 527832 182685 527844
rect 182343 527730 182395 527798
rect 182343 527696 182353 527730
rect 182387 527696 182395 527730
rect 182343 527670 182395 527696
rect 182633 527798 182641 527832
rect 182675 527798 182685 527832
rect 182633 527670 182685 527798
rect 183631 527832 183683 527844
rect 183631 527798 183641 527832
rect 183675 527798 183683 527832
rect 183631 527670 183683 527798
rect 183737 527832 183789 527844
rect 183737 527798 183745 527832
rect 183779 527798 183789 527832
rect 183737 527670 183789 527798
rect 184735 527832 184787 527844
rect 184735 527798 184745 527832
rect 184779 527798 184787 527832
rect 184735 527670 184787 527798
rect 184841 527832 184893 527844
rect 184841 527798 184849 527832
rect 184883 527798 184893 527832
rect 184841 527670 184893 527798
rect 185839 527832 185891 527844
rect 185839 527798 185849 527832
rect 185883 527798 185891 527832
rect 185839 527670 185891 527798
rect 185945 527832 185997 527844
rect 185945 527798 185953 527832
rect 185987 527798 185997 527832
rect 185945 527670 185997 527798
rect 186943 527832 186995 527844
rect 186943 527798 186953 527832
rect 186987 527798 186995 527832
rect 186943 527670 186995 527798
rect 187233 527832 187285 527844
rect 187233 527798 187241 527832
rect 187275 527798 187285 527832
rect 187233 527737 187285 527798
rect 187233 527703 187241 527737
rect 187275 527703 187285 527737
rect 187233 527670 187285 527703
rect 187403 527832 187455 527844
rect 187403 527798 187413 527832
rect 187447 527798 187455 527832
rect 187403 527737 187455 527798
rect 187403 527703 187413 527737
rect 187447 527703 187455 527737
rect 187403 527670 187455 527703
rect 172237 526991 172289 527024
rect 172237 526957 172245 526991
rect 172279 526957 172289 526991
rect 172237 526896 172289 526957
rect 172237 526862 172245 526896
rect 172279 526862 172289 526896
rect 172237 526850 172289 526862
rect 172407 526991 172459 527024
rect 172407 526957 172417 526991
rect 172451 526957 172459 526991
rect 172407 526896 172459 526957
rect 172407 526862 172417 526896
rect 172451 526862 172459 526896
rect 172407 526850 172459 526862
rect 172513 526896 172565 527024
rect 172513 526862 172521 526896
rect 172555 526862 172565 526896
rect 172513 526850 172565 526862
rect 173511 526896 173563 527024
rect 173511 526862 173521 526896
rect 173555 526862 173563 526896
rect 173511 526850 173563 526862
rect 173617 526896 173669 527024
rect 173617 526862 173625 526896
rect 173659 526862 173669 526896
rect 173617 526850 173669 526862
rect 174615 526896 174667 527024
rect 174615 526862 174625 526896
rect 174659 526862 174667 526896
rect 174905 526896 174957 527024
rect 174615 526850 174667 526862
rect 174905 526862 174913 526896
rect 174947 526862 174957 526896
rect 174905 526850 174957 526862
rect 175903 526896 175955 527024
rect 175903 526862 175913 526896
rect 175947 526862 175955 526896
rect 175903 526850 175955 526862
rect 176009 526896 176061 527024
rect 176009 526862 176017 526896
rect 176051 526862 176061 526896
rect 176009 526850 176061 526862
rect 177007 526896 177059 527024
rect 177007 526862 177017 526896
rect 177051 526862 177059 526896
rect 177007 526850 177059 526862
rect 177113 526896 177165 527024
rect 177113 526862 177121 526896
rect 177155 526862 177165 526896
rect 177113 526850 177165 526862
rect 178111 526896 178163 527024
rect 178111 526862 178121 526896
rect 178155 526862 178163 526896
rect 178111 526850 178163 526862
rect 178217 526896 178269 527024
rect 178217 526862 178225 526896
rect 178259 526862 178269 526896
rect 178217 526850 178269 526862
rect 179215 526896 179267 527024
rect 179215 526862 179225 526896
rect 179259 526862 179267 526896
rect 179215 526850 179267 526862
rect 179321 526998 179373 527024
rect 179321 526964 179329 526998
rect 179363 526964 179373 526998
rect 179321 526896 179373 526964
rect 179321 526862 179329 526896
rect 179363 526862 179373 526896
rect 179321 526850 179373 526862
rect 179767 526998 179819 527024
rect 179767 526964 179777 526998
rect 179811 526964 179819 526998
rect 179767 526896 179819 526964
rect 179767 526862 179777 526896
rect 179811 526862 179819 526896
rect 180057 526896 180109 527024
rect 179767 526850 179819 526862
rect 180057 526862 180065 526896
rect 180099 526862 180109 526896
rect 180057 526850 180109 526862
rect 181055 526896 181107 527024
rect 181055 526862 181065 526896
rect 181099 526862 181107 526896
rect 181055 526850 181107 526862
rect 181161 526896 181213 527024
rect 181161 526862 181169 526896
rect 181203 526862 181213 526896
rect 181161 526850 181213 526862
rect 182159 526896 182211 527024
rect 182159 526862 182169 526896
rect 182203 526862 182211 526896
rect 182159 526850 182211 526862
rect 182265 526896 182317 527024
rect 182265 526862 182273 526896
rect 182307 526862 182317 526896
rect 182265 526850 182317 526862
rect 183263 526896 183315 527024
rect 183263 526862 183273 526896
rect 183307 526862 183315 526896
rect 183263 526850 183315 526862
rect 183369 526896 183421 527024
rect 183369 526862 183377 526896
rect 183411 526862 183421 526896
rect 183369 526850 183421 526862
rect 184367 526896 184419 527024
rect 184367 526862 184377 526896
rect 184411 526862 184419 526896
rect 184367 526850 184419 526862
rect 184473 526998 184525 527024
rect 184473 526964 184481 526998
rect 184515 526964 184525 526998
rect 184473 526896 184525 526964
rect 184473 526862 184481 526896
rect 184515 526862 184525 526896
rect 184473 526850 184525 526862
rect 184919 526998 184971 527024
rect 184919 526964 184929 526998
rect 184963 526964 184971 526998
rect 184919 526896 184971 526964
rect 184919 526862 184929 526896
rect 184963 526862 184971 526896
rect 185209 526896 185261 527024
rect 184919 526850 184971 526862
rect 185209 526862 185217 526896
rect 185251 526862 185261 526896
rect 185209 526850 185261 526862
rect 186207 526896 186259 527024
rect 186207 526862 186217 526896
rect 186251 526862 186259 526896
rect 186207 526850 186259 526862
rect 186313 526998 186365 527024
rect 186313 526964 186321 526998
rect 186355 526964 186365 526998
rect 186313 526896 186365 526964
rect 186313 526862 186321 526896
rect 186355 526862 186365 526896
rect 186313 526850 186365 526862
rect 186943 526998 186995 527024
rect 186943 526964 186953 526998
rect 186987 526964 186995 526998
rect 186943 526896 186995 526964
rect 186943 526862 186953 526896
rect 186987 526862 186995 526896
rect 186943 526850 186995 526862
rect 187233 526991 187285 527024
rect 187233 526957 187241 526991
rect 187275 526957 187285 526991
rect 187233 526896 187285 526957
rect 187233 526862 187241 526896
rect 187275 526862 187285 526896
rect 187233 526850 187285 526862
rect 187403 526991 187455 527024
rect 187403 526957 187413 526991
rect 187447 526957 187455 526991
rect 187403 526896 187455 526957
rect 187403 526862 187413 526896
rect 187447 526862 187455 526896
rect 187403 526850 187455 526862
rect 172237 526744 172289 526756
rect 172237 526710 172245 526744
rect 172279 526710 172289 526744
rect 172237 526649 172289 526710
rect 172237 526615 172245 526649
rect 172279 526615 172289 526649
rect 172237 526582 172289 526615
rect 172407 526744 172459 526756
rect 172407 526710 172417 526744
rect 172451 526710 172459 526744
rect 172407 526649 172459 526710
rect 172407 526615 172417 526649
rect 172451 526615 172459 526649
rect 172407 526582 172459 526615
rect 172513 526744 172565 526756
rect 172513 526710 172521 526744
rect 172555 526710 172565 526744
rect 172513 526582 172565 526710
rect 173511 526744 173563 526756
rect 173511 526710 173521 526744
rect 173555 526710 173563 526744
rect 173511 526582 173563 526710
rect 173617 526744 173669 526756
rect 173617 526710 173625 526744
rect 173659 526710 173669 526744
rect 173617 526582 173669 526710
rect 174615 526744 174667 526756
rect 174615 526710 174625 526744
rect 174659 526710 174667 526744
rect 174615 526582 174667 526710
rect 174721 526744 174773 526756
rect 174721 526710 174729 526744
rect 174763 526710 174773 526744
rect 174721 526582 174773 526710
rect 175719 526744 175771 526756
rect 175719 526710 175729 526744
rect 175763 526710 175771 526744
rect 175719 526582 175771 526710
rect 175825 526744 175877 526756
rect 175825 526710 175833 526744
rect 175867 526710 175877 526744
rect 175825 526582 175877 526710
rect 176823 526744 176875 526756
rect 176823 526710 176833 526744
rect 176867 526710 176875 526744
rect 176823 526582 176875 526710
rect 176929 526744 176981 526756
rect 176929 526710 176937 526744
rect 176971 526710 176981 526744
rect 176929 526642 176981 526710
rect 176929 526608 176937 526642
rect 176971 526608 176981 526642
rect 176929 526582 176981 526608
rect 177191 526744 177243 526756
rect 177191 526710 177201 526744
rect 177235 526710 177243 526744
rect 177481 526744 177533 526756
rect 177191 526642 177243 526710
rect 177191 526608 177201 526642
rect 177235 526608 177243 526642
rect 177191 526582 177243 526608
rect 177481 526710 177489 526744
rect 177523 526710 177533 526744
rect 177481 526582 177533 526710
rect 178479 526744 178531 526756
rect 178479 526710 178489 526744
rect 178523 526710 178531 526744
rect 178479 526582 178531 526710
rect 178585 526744 178637 526756
rect 178585 526710 178593 526744
rect 178627 526710 178637 526744
rect 178585 526582 178637 526710
rect 179583 526744 179635 526756
rect 179583 526710 179593 526744
rect 179627 526710 179635 526744
rect 179583 526582 179635 526710
rect 179689 526744 179741 526756
rect 179689 526710 179697 526744
rect 179731 526710 179741 526744
rect 179689 526582 179741 526710
rect 180687 526744 180739 526756
rect 180687 526710 180697 526744
rect 180731 526710 180739 526744
rect 180687 526582 180739 526710
rect 180793 526744 180845 526756
rect 180793 526710 180801 526744
rect 180835 526710 180845 526744
rect 180793 526582 180845 526710
rect 181791 526744 181843 526756
rect 181791 526710 181801 526744
rect 181835 526710 181843 526744
rect 181791 526582 181843 526710
rect 181897 526744 181949 526756
rect 181897 526710 181905 526744
rect 181939 526710 181949 526744
rect 181897 526642 181949 526710
rect 181897 526608 181905 526642
rect 181939 526608 181949 526642
rect 181897 526582 181949 526608
rect 182343 526744 182395 526756
rect 182343 526710 182353 526744
rect 182387 526710 182395 526744
rect 182633 526744 182685 526756
rect 182343 526642 182395 526710
rect 182343 526608 182353 526642
rect 182387 526608 182395 526642
rect 182343 526582 182395 526608
rect 182633 526710 182641 526744
rect 182675 526710 182685 526744
rect 182633 526582 182685 526710
rect 183631 526744 183683 526756
rect 183631 526710 183641 526744
rect 183675 526710 183683 526744
rect 183631 526582 183683 526710
rect 183737 526744 183789 526756
rect 183737 526710 183745 526744
rect 183779 526710 183789 526744
rect 183737 526582 183789 526710
rect 184735 526744 184787 526756
rect 184735 526710 184745 526744
rect 184779 526710 184787 526744
rect 184735 526582 184787 526710
rect 184841 526744 184893 526756
rect 184841 526710 184849 526744
rect 184883 526710 184893 526744
rect 184841 526582 184893 526710
rect 185839 526744 185891 526756
rect 185839 526710 185849 526744
rect 185883 526710 185891 526744
rect 185839 526582 185891 526710
rect 185945 526744 185997 526756
rect 185945 526710 185953 526744
rect 185987 526710 185997 526744
rect 185945 526582 185997 526710
rect 186943 526744 186995 526756
rect 186943 526710 186953 526744
rect 186987 526710 186995 526744
rect 186943 526582 186995 526710
rect 187233 526744 187285 526756
rect 187233 526710 187241 526744
rect 187275 526710 187285 526744
rect 187233 526649 187285 526710
rect 187233 526615 187241 526649
rect 187275 526615 187285 526649
rect 187233 526582 187285 526615
rect 187403 526744 187455 526756
rect 187403 526710 187413 526744
rect 187447 526710 187455 526744
rect 187403 526649 187455 526710
rect 187403 526615 187413 526649
rect 187447 526615 187455 526649
rect 187403 526582 187455 526615
rect 172237 525903 172289 525936
rect 172237 525869 172245 525903
rect 172279 525869 172289 525903
rect 172237 525808 172289 525869
rect 172237 525774 172245 525808
rect 172279 525774 172289 525808
rect 172237 525762 172289 525774
rect 172407 525903 172459 525936
rect 172407 525869 172417 525903
rect 172451 525869 172459 525903
rect 172407 525808 172459 525869
rect 172407 525774 172417 525808
rect 172451 525774 172459 525808
rect 172407 525762 172459 525774
rect 172513 525808 172565 525936
rect 172513 525774 172521 525808
rect 172555 525774 172565 525808
rect 172513 525762 172565 525774
rect 173511 525808 173563 525936
rect 173511 525774 173521 525808
rect 173555 525774 173563 525808
rect 173511 525762 173563 525774
rect 173617 525808 173669 525936
rect 173617 525774 173625 525808
rect 173659 525774 173669 525808
rect 173617 525762 173669 525774
rect 174615 525808 174667 525936
rect 174615 525774 174625 525808
rect 174659 525774 174667 525808
rect 174905 525808 174957 525936
rect 174615 525762 174667 525774
rect 174905 525774 174913 525808
rect 174947 525774 174957 525808
rect 174905 525762 174957 525774
rect 175903 525808 175955 525936
rect 175903 525774 175913 525808
rect 175947 525774 175955 525808
rect 175903 525762 175955 525774
rect 176009 525808 176061 525936
rect 176009 525774 176017 525808
rect 176051 525774 176061 525808
rect 176009 525762 176061 525774
rect 177007 525808 177059 525936
rect 177007 525774 177017 525808
rect 177051 525774 177059 525808
rect 177007 525762 177059 525774
rect 177113 525808 177165 525936
rect 177113 525774 177121 525808
rect 177155 525774 177165 525808
rect 177113 525762 177165 525774
rect 178111 525808 178163 525936
rect 178111 525774 178121 525808
rect 178155 525774 178163 525808
rect 178111 525762 178163 525774
rect 178217 525808 178269 525936
rect 178217 525774 178225 525808
rect 178259 525774 178269 525808
rect 178217 525762 178269 525774
rect 179215 525808 179267 525936
rect 179215 525774 179225 525808
rect 179259 525774 179267 525808
rect 179215 525762 179267 525774
rect 179321 525910 179373 525936
rect 179321 525876 179329 525910
rect 179363 525876 179373 525910
rect 179321 525808 179373 525876
rect 179321 525774 179329 525808
rect 179363 525774 179373 525808
rect 179321 525762 179373 525774
rect 179767 525910 179819 525936
rect 179767 525876 179777 525910
rect 179811 525876 179819 525910
rect 179767 525808 179819 525876
rect 179767 525774 179777 525808
rect 179811 525774 179819 525808
rect 180057 525808 180109 525936
rect 179767 525762 179819 525774
rect 180057 525774 180065 525808
rect 180099 525774 180109 525808
rect 180057 525762 180109 525774
rect 181055 525808 181107 525936
rect 181055 525774 181065 525808
rect 181099 525774 181107 525808
rect 181055 525762 181107 525774
rect 181161 525808 181213 525936
rect 181161 525774 181169 525808
rect 181203 525774 181213 525808
rect 181161 525762 181213 525774
rect 182159 525808 182211 525936
rect 182159 525774 182169 525808
rect 182203 525774 182211 525808
rect 182159 525762 182211 525774
rect 182265 525808 182317 525936
rect 182265 525774 182273 525808
rect 182307 525774 182317 525808
rect 182265 525762 182317 525774
rect 183263 525808 183315 525936
rect 183263 525774 183273 525808
rect 183307 525774 183315 525808
rect 183263 525762 183315 525774
rect 183369 525808 183421 525936
rect 183369 525774 183377 525808
rect 183411 525774 183421 525808
rect 183369 525762 183421 525774
rect 184367 525808 184419 525936
rect 184367 525774 184377 525808
rect 184411 525774 184419 525808
rect 184367 525762 184419 525774
rect 184473 525910 184525 525936
rect 184473 525876 184481 525910
rect 184515 525876 184525 525910
rect 184473 525808 184525 525876
rect 184473 525774 184481 525808
rect 184515 525774 184525 525808
rect 184473 525762 184525 525774
rect 184919 525910 184971 525936
rect 184919 525876 184929 525910
rect 184963 525876 184971 525910
rect 184919 525808 184971 525876
rect 184919 525774 184929 525808
rect 184963 525774 184971 525808
rect 185209 525808 185261 525936
rect 184919 525762 184971 525774
rect 185209 525774 185217 525808
rect 185251 525774 185261 525808
rect 185209 525762 185261 525774
rect 186207 525808 186259 525936
rect 186207 525774 186217 525808
rect 186251 525774 186259 525808
rect 186207 525762 186259 525774
rect 186313 525910 186365 525936
rect 186313 525876 186321 525910
rect 186355 525876 186365 525910
rect 186313 525808 186365 525876
rect 186313 525774 186321 525808
rect 186355 525774 186365 525808
rect 186313 525762 186365 525774
rect 186943 525910 186995 525936
rect 186943 525876 186953 525910
rect 186987 525876 186995 525910
rect 186943 525808 186995 525876
rect 186943 525774 186953 525808
rect 186987 525774 186995 525808
rect 186943 525762 186995 525774
rect 187233 525903 187285 525936
rect 187233 525869 187241 525903
rect 187275 525869 187285 525903
rect 187233 525808 187285 525869
rect 187233 525774 187241 525808
rect 187275 525774 187285 525808
rect 187233 525762 187285 525774
rect 187403 525903 187455 525936
rect 187403 525869 187413 525903
rect 187447 525869 187455 525903
rect 187403 525808 187455 525869
rect 187403 525774 187413 525808
rect 187447 525774 187455 525808
rect 187403 525762 187455 525774
rect 172237 525656 172289 525668
rect 172237 525622 172245 525656
rect 172279 525622 172289 525656
rect 172237 525561 172289 525622
rect 172237 525527 172245 525561
rect 172279 525527 172289 525561
rect 172237 525494 172289 525527
rect 172407 525656 172459 525668
rect 172407 525622 172417 525656
rect 172451 525622 172459 525656
rect 172407 525561 172459 525622
rect 172407 525527 172417 525561
rect 172451 525527 172459 525561
rect 172407 525494 172459 525527
rect 172513 525656 172565 525668
rect 172513 525622 172521 525656
rect 172555 525622 172565 525656
rect 172513 525494 172565 525622
rect 173511 525656 173563 525668
rect 173511 525622 173521 525656
rect 173555 525622 173563 525656
rect 173511 525494 173563 525622
rect 173617 525656 173669 525668
rect 173617 525622 173625 525656
rect 173659 525622 173669 525656
rect 173617 525494 173669 525622
rect 174615 525656 174667 525668
rect 174615 525622 174625 525656
rect 174659 525622 174667 525656
rect 174615 525494 174667 525622
rect 174721 525656 174773 525668
rect 174721 525622 174729 525656
rect 174763 525622 174773 525656
rect 174721 525494 174773 525622
rect 175719 525656 175771 525668
rect 175719 525622 175729 525656
rect 175763 525622 175771 525656
rect 175719 525494 175771 525622
rect 175825 525656 175877 525668
rect 175825 525622 175833 525656
rect 175867 525622 175877 525656
rect 175825 525494 175877 525622
rect 176823 525656 176875 525668
rect 176823 525622 176833 525656
rect 176867 525622 176875 525656
rect 176823 525494 176875 525622
rect 176929 525656 176981 525668
rect 176929 525622 176937 525656
rect 176971 525622 176981 525656
rect 176929 525554 176981 525622
rect 176929 525520 176937 525554
rect 176971 525520 176981 525554
rect 176929 525494 176981 525520
rect 177191 525656 177243 525668
rect 177191 525622 177201 525656
rect 177235 525622 177243 525656
rect 177481 525656 177533 525668
rect 177191 525554 177243 525622
rect 177191 525520 177201 525554
rect 177235 525520 177243 525554
rect 177191 525494 177243 525520
rect 177481 525622 177489 525656
rect 177523 525622 177533 525656
rect 177481 525494 177533 525622
rect 178479 525656 178531 525668
rect 178479 525622 178489 525656
rect 178523 525622 178531 525656
rect 178479 525494 178531 525622
rect 178585 525656 178637 525668
rect 178585 525622 178593 525656
rect 178627 525622 178637 525656
rect 178585 525494 178637 525622
rect 179583 525656 179635 525668
rect 179583 525622 179593 525656
rect 179627 525622 179635 525656
rect 179583 525494 179635 525622
rect 179689 525656 179741 525668
rect 179689 525622 179697 525656
rect 179731 525622 179741 525656
rect 179689 525494 179741 525622
rect 180687 525656 180739 525668
rect 180687 525622 180697 525656
rect 180731 525622 180739 525656
rect 180687 525494 180739 525622
rect 180793 525656 180845 525668
rect 180793 525622 180801 525656
rect 180835 525622 180845 525656
rect 180793 525494 180845 525622
rect 181791 525656 181843 525668
rect 181791 525622 181801 525656
rect 181835 525622 181843 525656
rect 181791 525494 181843 525622
rect 181897 525656 181949 525668
rect 181897 525622 181905 525656
rect 181939 525622 181949 525656
rect 181897 525554 181949 525622
rect 181897 525520 181905 525554
rect 181939 525520 181949 525554
rect 181897 525494 181949 525520
rect 182343 525656 182395 525668
rect 182343 525622 182353 525656
rect 182387 525622 182395 525656
rect 182633 525656 182685 525668
rect 182343 525554 182395 525622
rect 182343 525520 182353 525554
rect 182387 525520 182395 525554
rect 182343 525494 182395 525520
rect 182633 525622 182641 525656
rect 182675 525622 182685 525656
rect 182633 525494 182685 525622
rect 183631 525656 183683 525668
rect 183631 525622 183641 525656
rect 183675 525622 183683 525656
rect 183631 525494 183683 525622
rect 183737 525656 183789 525668
rect 183737 525622 183745 525656
rect 183779 525622 183789 525656
rect 183737 525494 183789 525622
rect 184735 525656 184787 525668
rect 184735 525622 184745 525656
rect 184779 525622 184787 525656
rect 184735 525494 184787 525622
rect 184841 525656 184893 525668
rect 184841 525622 184849 525656
rect 184883 525622 184893 525656
rect 184841 525494 184893 525622
rect 185839 525656 185891 525668
rect 185839 525622 185849 525656
rect 185883 525622 185891 525656
rect 185839 525494 185891 525622
rect 185945 525656 185997 525668
rect 185945 525622 185953 525656
rect 185987 525622 185997 525656
rect 185945 525494 185997 525622
rect 186943 525656 186995 525668
rect 186943 525622 186953 525656
rect 186987 525622 186995 525656
rect 186943 525494 186995 525622
rect 187233 525656 187285 525668
rect 187233 525622 187241 525656
rect 187275 525622 187285 525656
rect 187233 525561 187285 525622
rect 187233 525527 187241 525561
rect 187275 525527 187285 525561
rect 187233 525494 187285 525527
rect 187403 525656 187455 525668
rect 187403 525622 187413 525656
rect 187447 525622 187455 525656
rect 187403 525561 187455 525622
rect 187403 525527 187413 525561
rect 187447 525527 187455 525561
rect 187403 525494 187455 525527
rect 172237 524815 172289 524848
rect 172237 524781 172245 524815
rect 172279 524781 172289 524815
rect 172237 524720 172289 524781
rect 172237 524686 172245 524720
rect 172279 524686 172289 524720
rect 172237 524674 172289 524686
rect 172407 524815 172459 524848
rect 172407 524781 172417 524815
rect 172451 524781 172459 524815
rect 172407 524720 172459 524781
rect 172407 524686 172417 524720
rect 172451 524686 172459 524720
rect 172407 524674 172459 524686
rect 172513 524720 172565 524848
rect 172513 524686 172521 524720
rect 172555 524686 172565 524720
rect 172513 524674 172565 524686
rect 173511 524720 173563 524848
rect 173511 524686 173521 524720
rect 173555 524686 173563 524720
rect 173511 524674 173563 524686
rect 173617 524720 173669 524848
rect 173617 524686 173625 524720
rect 173659 524686 173669 524720
rect 173617 524674 173669 524686
rect 174615 524720 174667 524848
rect 174615 524686 174625 524720
rect 174659 524686 174667 524720
rect 174905 524720 174957 524848
rect 174615 524674 174667 524686
rect 174905 524686 174913 524720
rect 174947 524686 174957 524720
rect 174905 524674 174957 524686
rect 175903 524720 175955 524848
rect 175903 524686 175913 524720
rect 175947 524686 175955 524720
rect 175903 524674 175955 524686
rect 176009 524720 176061 524848
rect 176009 524686 176017 524720
rect 176051 524686 176061 524720
rect 176009 524674 176061 524686
rect 177007 524720 177059 524848
rect 177007 524686 177017 524720
rect 177051 524686 177059 524720
rect 177007 524674 177059 524686
rect 177113 524720 177165 524848
rect 177113 524686 177121 524720
rect 177155 524686 177165 524720
rect 177113 524674 177165 524686
rect 178111 524720 178163 524848
rect 178111 524686 178121 524720
rect 178155 524686 178163 524720
rect 178111 524674 178163 524686
rect 178217 524720 178269 524848
rect 178217 524686 178225 524720
rect 178259 524686 178269 524720
rect 178217 524674 178269 524686
rect 179215 524720 179267 524848
rect 179215 524686 179225 524720
rect 179259 524686 179267 524720
rect 179215 524674 179267 524686
rect 179321 524822 179373 524848
rect 179321 524788 179329 524822
rect 179363 524788 179373 524822
rect 179321 524720 179373 524788
rect 179321 524686 179329 524720
rect 179363 524686 179373 524720
rect 179321 524674 179373 524686
rect 179767 524822 179819 524848
rect 179767 524788 179777 524822
rect 179811 524788 179819 524822
rect 179767 524720 179819 524788
rect 179767 524686 179777 524720
rect 179811 524686 179819 524720
rect 180057 524720 180109 524848
rect 179767 524674 179819 524686
rect 180057 524686 180065 524720
rect 180099 524686 180109 524720
rect 180057 524674 180109 524686
rect 181055 524720 181107 524848
rect 181055 524686 181065 524720
rect 181099 524686 181107 524720
rect 181055 524674 181107 524686
rect 181161 524720 181213 524848
rect 181161 524686 181169 524720
rect 181203 524686 181213 524720
rect 181161 524674 181213 524686
rect 182159 524720 182211 524848
rect 182159 524686 182169 524720
rect 182203 524686 182211 524720
rect 182159 524674 182211 524686
rect 182265 524720 182317 524848
rect 182265 524686 182273 524720
rect 182307 524686 182317 524720
rect 182265 524674 182317 524686
rect 183263 524720 183315 524848
rect 183263 524686 183273 524720
rect 183307 524686 183315 524720
rect 183263 524674 183315 524686
rect 183369 524720 183421 524848
rect 183369 524686 183377 524720
rect 183411 524686 183421 524720
rect 183369 524674 183421 524686
rect 184367 524720 184419 524848
rect 184367 524686 184377 524720
rect 184411 524686 184419 524720
rect 184367 524674 184419 524686
rect 184473 524822 184525 524848
rect 184473 524788 184481 524822
rect 184515 524788 184525 524822
rect 184473 524720 184525 524788
rect 184473 524686 184481 524720
rect 184515 524686 184525 524720
rect 184473 524674 184525 524686
rect 184919 524822 184971 524848
rect 184919 524788 184929 524822
rect 184963 524788 184971 524822
rect 184919 524720 184971 524788
rect 184919 524686 184929 524720
rect 184963 524686 184971 524720
rect 185209 524720 185261 524848
rect 184919 524674 184971 524686
rect 185209 524686 185217 524720
rect 185251 524686 185261 524720
rect 185209 524674 185261 524686
rect 186207 524720 186259 524848
rect 186207 524686 186217 524720
rect 186251 524686 186259 524720
rect 186207 524674 186259 524686
rect 186313 524822 186365 524848
rect 186313 524788 186321 524822
rect 186355 524788 186365 524822
rect 186313 524720 186365 524788
rect 186313 524686 186321 524720
rect 186355 524686 186365 524720
rect 186313 524674 186365 524686
rect 186943 524822 186995 524848
rect 186943 524788 186953 524822
rect 186987 524788 186995 524822
rect 186943 524720 186995 524788
rect 186943 524686 186953 524720
rect 186987 524686 186995 524720
rect 186943 524674 186995 524686
rect 187233 524815 187285 524848
rect 187233 524781 187241 524815
rect 187275 524781 187285 524815
rect 187233 524720 187285 524781
rect 187233 524686 187241 524720
rect 187275 524686 187285 524720
rect 187233 524674 187285 524686
rect 187403 524815 187455 524848
rect 187403 524781 187413 524815
rect 187447 524781 187455 524815
rect 187403 524720 187455 524781
rect 187403 524686 187413 524720
rect 187447 524686 187455 524720
rect 187403 524674 187455 524686
rect 172237 524568 172289 524580
rect 172237 524534 172245 524568
rect 172279 524534 172289 524568
rect 172237 524473 172289 524534
rect 172237 524439 172245 524473
rect 172279 524439 172289 524473
rect 172237 524406 172289 524439
rect 172407 524568 172459 524580
rect 172407 524534 172417 524568
rect 172451 524534 172459 524568
rect 172407 524473 172459 524534
rect 172407 524439 172417 524473
rect 172451 524439 172459 524473
rect 172407 524406 172459 524439
rect 172513 524568 172565 524580
rect 172513 524534 172521 524568
rect 172555 524534 172565 524568
rect 172513 524406 172565 524534
rect 173511 524568 173563 524580
rect 173511 524534 173521 524568
rect 173555 524534 173563 524568
rect 173511 524406 173563 524534
rect 173617 524568 173669 524580
rect 173617 524534 173625 524568
rect 173659 524534 173669 524568
rect 173617 524406 173669 524534
rect 174615 524568 174667 524580
rect 174615 524534 174625 524568
rect 174659 524534 174667 524568
rect 174615 524406 174667 524534
rect 174721 524568 174773 524580
rect 174721 524534 174729 524568
rect 174763 524534 174773 524568
rect 174721 524406 174773 524534
rect 175719 524568 175771 524580
rect 175719 524534 175729 524568
rect 175763 524534 175771 524568
rect 175719 524406 175771 524534
rect 175825 524568 175877 524580
rect 175825 524534 175833 524568
rect 175867 524534 175877 524568
rect 175825 524406 175877 524534
rect 176823 524568 176875 524580
rect 176823 524534 176833 524568
rect 176867 524534 176875 524568
rect 176823 524406 176875 524534
rect 176929 524568 176981 524580
rect 176929 524534 176937 524568
rect 176971 524534 176981 524568
rect 176929 524466 176981 524534
rect 176929 524432 176937 524466
rect 176971 524432 176981 524466
rect 176929 524406 176981 524432
rect 177191 524568 177243 524580
rect 177191 524534 177201 524568
rect 177235 524534 177243 524568
rect 177481 524568 177533 524580
rect 177191 524466 177243 524534
rect 177191 524432 177201 524466
rect 177235 524432 177243 524466
rect 177191 524406 177243 524432
rect 177481 524534 177489 524568
rect 177523 524534 177533 524568
rect 177481 524406 177533 524534
rect 178479 524568 178531 524580
rect 178479 524534 178489 524568
rect 178523 524534 178531 524568
rect 178479 524406 178531 524534
rect 178585 524568 178637 524580
rect 178585 524534 178593 524568
rect 178627 524534 178637 524568
rect 178585 524406 178637 524534
rect 179583 524568 179635 524580
rect 179583 524534 179593 524568
rect 179627 524534 179635 524568
rect 179583 524406 179635 524534
rect 179689 524568 179741 524580
rect 179689 524534 179697 524568
rect 179731 524534 179741 524568
rect 179689 524406 179741 524534
rect 180687 524568 180739 524580
rect 180687 524534 180697 524568
rect 180731 524534 180739 524568
rect 180687 524406 180739 524534
rect 180793 524568 180845 524580
rect 180793 524534 180801 524568
rect 180835 524534 180845 524568
rect 180793 524406 180845 524534
rect 181791 524568 181843 524580
rect 181791 524534 181801 524568
rect 181835 524534 181843 524568
rect 181791 524406 181843 524534
rect 181897 524568 181949 524580
rect 181897 524534 181905 524568
rect 181939 524534 181949 524568
rect 181897 524466 181949 524534
rect 181897 524432 181905 524466
rect 181939 524432 181949 524466
rect 181897 524406 181949 524432
rect 182343 524568 182395 524580
rect 182343 524534 182353 524568
rect 182387 524534 182395 524568
rect 182633 524568 182685 524580
rect 182343 524466 182395 524534
rect 182343 524432 182353 524466
rect 182387 524432 182395 524466
rect 182343 524406 182395 524432
rect 182633 524534 182641 524568
rect 182675 524534 182685 524568
rect 182633 524406 182685 524534
rect 183631 524568 183683 524580
rect 183631 524534 183641 524568
rect 183675 524534 183683 524568
rect 183631 524406 183683 524534
rect 183737 524568 183789 524580
rect 183737 524534 183745 524568
rect 183779 524534 183789 524568
rect 183737 524406 183789 524534
rect 184735 524568 184787 524580
rect 184735 524534 184745 524568
rect 184779 524534 184787 524568
rect 184735 524406 184787 524534
rect 184841 524568 184893 524580
rect 184841 524534 184849 524568
rect 184883 524534 184893 524568
rect 184841 524406 184893 524534
rect 185839 524568 185891 524580
rect 185839 524534 185849 524568
rect 185883 524534 185891 524568
rect 185839 524406 185891 524534
rect 185945 524568 185997 524580
rect 185945 524534 185953 524568
rect 185987 524534 185997 524568
rect 185945 524406 185997 524534
rect 186943 524568 186995 524580
rect 186943 524534 186953 524568
rect 186987 524534 186995 524568
rect 186943 524406 186995 524534
rect 187233 524568 187285 524580
rect 187233 524534 187241 524568
rect 187275 524534 187285 524568
rect 187233 524473 187285 524534
rect 187233 524439 187241 524473
rect 187275 524439 187285 524473
rect 187233 524406 187285 524439
rect 187403 524568 187455 524580
rect 187403 524534 187413 524568
rect 187447 524534 187455 524568
rect 187403 524473 187455 524534
rect 187403 524439 187413 524473
rect 187447 524439 187455 524473
rect 187403 524406 187455 524439
rect 172237 523727 172289 523760
rect 172237 523693 172245 523727
rect 172279 523693 172289 523727
rect 172237 523632 172289 523693
rect 172237 523598 172245 523632
rect 172279 523598 172289 523632
rect 172237 523586 172289 523598
rect 172407 523727 172459 523760
rect 172407 523693 172417 523727
rect 172451 523693 172459 523727
rect 172407 523632 172459 523693
rect 172407 523598 172417 523632
rect 172451 523598 172459 523632
rect 172407 523586 172459 523598
rect 172513 523632 172565 523760
rect 172513 523598 172521 523632
rect 172555 523598 172565 523632
rect 172513 523586 172565 523598
rect 173511 523632 173563 523760
rect 173511 523598 173521 523632
rect 173555 523598 173563 523632
rect 173511 523586 173563 523598
rect 173617 523632 173669 523760
rect 173617 523598 173625 523632
rect 173659 523598 173669 523632
rect 173617 523586 173669 523598
rect 174615 523632 174667 523760
rect 174615 523598 174625 523632
rect 174659 523598 174667 523632
rect 174905 523632 174957 523760
rect 174615 523586 174667 523598
rect 174905 523598 174913 523632
rect 174947 523598 174957 523632
rect 174905 523586 174957 523598
rect 175903 523632 175955 523760
rect 175903 523598 175913 523632
rect 175947 523598 175955 523632
rect 175903 523586 175955 523598
rect 176009 523632 176061 523760
rect 176009 523598 176017 523632
rect 176051 523598 176061 523632
rect 176009 523586 176061 523598
rect 177007 523632 177059 523760
rect 177007 523598 177017 523632
rect 177051 523598 177059 523632
rect 177007 523586 177059 523598
rect 177113 523632 177165 523760
rect 177113 523598 177121 523632
rect 177155 523598 177165 523632
rect 177113 523586 177165 523598
rect 178111 523632 178163 523760
rect 178111 523598 178121 523632
rect 178155 523598 178163 523632
rect 178111 523586 178163 523598
rect 178217 523632 178269 523760
rect 178217 523598 178225 523632
rect 178259 523598 178269 523632
rect 178217 523586 178269 523598
rect 179215 523632 179267 523760
rect 179215 523598 179225 523632
rect 179259 523598 179267 523632
rect 179215 523586 179267 523598
rect 179321 523734 179373 523760
rect 179321 523700 179329 523734
rect 179363 523700 179373 523734
rect 179321 523632 179373 523700
rect 179321 523598 179329 523632
rect 179363 523598 179373 523632
rect 179321 523586 179373 523598
rect 179767 523734 179819 523760
rect 179767 523700 179777 523734
rect 179811 523700 179819 523734
rect 179767 523632 179819 523700
rect 179767 523598 179777 523632
rect 179811 523598 179819 523632
rect 180057 523632 180109 523760
rect 179767 523586 179819 523598
rect 180057 523598 180065 523632
rect 180099 523598 180109 523632
rect 180057 523586 180109 523598
rect 181055 523632 181107 523760
rect 181055 523598 181065 523632
rect 181099 523598 181107 523632
rect 181055 523586 181107 523598
rect 181161 523632 181213 523760
rect 181161 523598 181169 523632
rect 181203 523598 181213 523632
rect 181161 523586 181213 523598
rect 182159 523632 182211 523760
rect 182159 523598 182169 523632
rect 182203 523598 182211 523632
rect 182159 523586 182211 523598
rect 182265 523632 182317 523760
rect 182265 523598 182273 523632
rect 182307 523598 182317 523632
rect 182265 523586 182317 523598
rect 183263 523632 183315 523760
rect 183263 523598 183273 523632
rect 183307 523598 183315 523632
rect 183263 523586 183315 523598
rect 183369 523632 183421 523760
rect 183369 523598 183377 523632
rect 183411 523598 183421 523632
rect 183369 523586 183421 523598
rect 184367 523632 184419 523760
rect 184367 523598 184377 523632
rect 184411 523598 184419 523632
rect 184367 523586 184419 523598
rect 184473 523734 184525 523760
rect 184473 523700 184481 523734
rect 184515 523700 184525 523734
rect 184473 523632 184525 523700
rect 184473 523598 184481 523632
rect 184515 523598 184525 523632
rect 184473 523586 184525 523598
rect 184919 523734 184971 523760
rect 184919 523700 184929 523734
rect 184963 523700 184971 523734
rect 184919 523632 184971 523700
rect 184919 523598 184929 523632
rect 184963 523598 184971 523632
rect 185209 523632 185261 523760
rect 184919 523586 184971 523598
rect 185209 523598 185217 523632
rect 185251 523598 185261 523632
rect 185209 523586 185261 523598
rect 186207 523632 186259 523760
rect 186207 523598 186217 523632
rect 186251 523598 186259 523632
rect 186207 523586 186259 523598
rect 186313 523734 186365 523760
rect 186313 523700 186321 523734
rect 186355 523700 186365 523734
rect 186313 523632 186365 523700
rect 186313 523598 186321 523632
rect 186355 523598 186365 523632
rect 186313 523586 186365 523598
rect 186943 523734 186995 523760
rect 186943 523700 186953 523734
rect 186987 523700 186995 523734
rect 186943 523632 186995 523700
rect 186943 523598 186953 523632
rect 186987 523598 186995 523632
rect 186943 523586 186995 523598
rect 187233 523727 187285 523760
rect 187233 523693 187241 523727
rect 187275 523693 187285 523727
rect 187233 523632 187285 523693
rect 187233 523598 187241 523632
rect 187275 523598 187285 523632
rect 187233 523586 187285 523598
rect 187403 523727 187455 523760
rect 187403 523693 187413 523727
rect 187447 523693 187455 523727
rect 187403 523632 187455 523693
rect 187403 523598 187413 523632
rect 187447 523598 187455 523632
rect 187403 523586 187455 523598
rect 172237 523480 172289 523492
rect 172237 523446 172245 523480
rect 172279 523446 172289 523480
rect 172237 523385 172289 523446
rect 172237 523351 172245 523385
rect 172279 523351 172289 523385
rect 172237 523318 172289 523351
rect 172407 523480 172459 523492
rect 172407 523446 172417 523480
rect 172451 523446 172459 523480
rect 172407 523385 172459 523446
rect 172407 523351 172417 523385
rect 172451 523351 172459 523385
rect 172407 523318 172459 523351
rect 172513 523480 172565 523492
rect 172513 523446 172521 523480
rect 172555 523446 172565 523480
rect 172513 523318 172565 523446
rect 173511 523480 173563 523492
rect 173511 523446 173521 523480
rect 173555 523446 173563 523480
rect 173511 523318 173563 523446
rect 173617 523480 173669 523492
rect 173617 523446 173625 523480
rect 173659 523446 173669 523480
rect 173617 523318 173669 523446
rect 174615 523480 174667 523492
rect 174615 523446 174625 523480
rect 174659 523446 174667 523480
rect 174615 523318 174667 523446
rect 174721 523480 174773 523492
rect 174721 523446 174729 523480
rect 174763 523446 174773 523480
rect 174721 523318 174773 523446
rect 175719 523480 175771 523492
rect 175719 523446 175729 523480
rect 175763 523446 175771 523480
rect 175719 523318 175771 523446
rect 175825 523480 175877 523492
rect 175825 523446 175833 523480
rect 175867 523446 175877 523480
rect 175825 523318 175877 523446
rect 176823 523480 176875 523492
rect 176823 523446 176833 523480
rect 176867 523446 176875 523480
rect 176823 523318 176875 523446
rect 176929 523480 176981 523492
rect 176929 523446 176937 523480
rect 176971 523446 176981 523480
rect 176929 523378 176981 523446
rect 176929 523344 176937 523378
rect 176971 523344 176981 523378
rect 176929 523318 176981 523344
rect 177191 523480 177243 523492
rect 177191 523446 177201 523480
rect 177235 523446 177243 523480
rect 177481 523480 177533 523492
rect 177191 523378 177243 523446
rect 177191 523344 177201 523378
rect 177235 523344 177243 523378
rect 177191 523318 177243 523344
rect 177481 523446 177489 523480
rect 177523 523446 177533 523480
rect 177481 523318 177533 523446
rect 178479 523480 178531 523492
rect 178479 523446 178489 523480
rect 178523 523446 178531 523480
rect 178479 523318 178531 523446
rect 178585 523480 178637 523492
rect 178585 523446 178593 523480
rect 178627 523446 178637 523480
rect 178585 523318 178637 523446
rect 179583 523480 179635 523492
rect 179583 523446 179593 523480
rect 179627 523446 179635 523480
rect 179583 523318 179635 523446
rect 179689 523480 179741 523492
rect 179689 523446 179697 523480
rect 179731 523446 179741 523480
rect 179689 523318 179741 523446
rect 180687 523480 180739 523492
rect 180687 523446 180697 523480
rect 180731 523446 180739 523480
rect 180687 523318 180739 523446
rect 180793 523480 180845 523492
rect 180793 523446 180801 523480
rect 180835 523446 180845 523480
rect 180793 523318 180845 523446
rect 181791 523480 181843 523492
rect 181791 523446 181801 523480
rect 181835 523446 181843 523480
rect 181791 523318 181843 523446
rect 181897 523480 181949 523492
rect 181897 523446 181905 523480
rect 181939 523446 181949 523480
rect 181897 523378 181949 523446
rect 181897 523344 181905 523378
rect 181939 523344 181949 523378
rect 181897 523318 181949 523344
rect 182343 523480 182395 523492
rect 182343 523446 182353 523480
rect 182387 523446 182395 523480
rect 182633 523480 182685 523492
rect 182343 523378 182395 523446
rect 182343 523344 182353 523378
rect 182387 523344 182395 523378
rect 182343 523318 182395 523344
rect 182633 523446 182641 523480
rect 182675 523446 182685 523480
rect 182633 523318 182685 523446
rect 183631 523480 183683 523492
rect 183631 523446 183641 523480
rect 183675 523446 183683 523480
rect 183631 523318 183683 523446
rect 183737 523480 183789 523492
rect 183737 523446 183745 523480
rect 183779 523446 183789 523480
rect 183737 523318 183789 523446
rect 184735 523480 184787 523492
rect 184735 523446 184745 523480
rect 184779 523446 184787 523480
rect 184735 523318 184787 523446
rect 184841 523480 184893 523492
rect 184841 523446 184849 523480
rect 184883 523446 184893 523480
rect 184841 523318 184893 523446
rect 185839 523480 185891 523492
rect 185839 523446 185849 523480
rect 185883 523446 185891 523480
rect 185839 523318 185891 523446
rect 185945 523480 185997 523492
rect 185945 523446 185953 523480
rect 185987 523446 185997 523480
rect 185945 523318 185997 523446
rect 186943 523480 186995 523492
rect 186943 523446 186953 523480
rect 186987 523446 186995 523480
rect 186943 523318 186995 523446
rect 187233 523480 187285 523492
rect 187233 523446 187241 523480
rect 187275 523446 187285 523480
rect 187233 523385 187285 523446
rect 187233 523351 187241 523385
rect 187275 523351 187285 523385
rect 187233 523318 187285 523351
rect 187403 523480 187455 523492
rect 187403 523446 187413 523480
rect 187447 523446 187455 523480
rect 187403 523385 187455 523446
rect 187403 523351 187413 523385
rect 187447 523351 187455 523385
rect 187403 523318 187455 523351
rect 172237 522639 172289 522672
rect 172237 522605 172245 522639
rect 172279 522605 172289 522639
rect 172237 522544 172289 522605
rect 172237 522510 172245 522544
rect 172279 522510 172289 522544
rect 172237 522498 172289 522510
rect 172407 522639 172459 522672
rect 172407 522605 172417 522639
rect 172451 522605 172459 522639
rect 172407 522544 172459 522605
rect 172407 522510 172417 522544
rect 172451 522510 172459 522544
rect 172407 522498 172459 522510
rect 172513 522544 172565 522672
rect 172513 522510 172521 522544
rect 172555 522510 172565 522544
rect 172513 522498 172565 522510
rect 173511 522544 173563 522672
rect 173511 522510 173521 522544
rect 173555 522510 173563 522544
rect 173511 522498 173563 522510
rect 173617 522544 173669 522672
rect 173617 522510 173625 522544
rect 173659 522510 173669 522544
rect 173617 522498 173669 522510
rect 174615 522544 174667 522672
rect 174615 522510 174625 522544
rect 174659 522510 174667 522544
rect 174905 522544 174957 522672
rect 174615 522498 174667 522510
rect 174905 522510 174913 522544
rect 174947 522510 174957 522544
rect 174905 522498 174957 522510
rect 175903 522544 175955 522672
rect 175903 522510 175913 522544
rect 175947 522510 175955 522544
rect 175903 522498 175955 522510
rect 176009 522544 176061 522672
rect 176009 522510 176017 522544
rect 176051 522510 176061 522544
rect 176009 522498 176061 522510
rect 177007 522544 177059 522672
rect 177007 522510 177017 522544
rect 177051 522510 177059 522544
rect 177007 522498 177059 522510
rect 177113 522544 177165 522672
rect 177113 522510 177121 522544
rect 177155 522510 177165 522544
rect 177113 522498 177165 522510
rect 178111 522544 178163 522672
rect 178111 522510 178121 522544
rect 178155 522510 178163 522544
rect 178111 522498 178163 522510
rect 178217 522544 178269 522672
rect 178217 522510 178225 522544
rect 178259 522510 178269 522544
rect 178217 522498 178269 522510
rect 179215 522544 179267 522672
rect 179215 522510 179225 522544
rect 179259 522510 179267 522544
rect 179215 522498 179267 522510
rect 179321 522646 179373 522672
rect 179321 522612 179329 522646
rect 179363 522612 179373 522646
rect 179321 522544 179373 522612
rect 179321 522510 179329 522544
rect 179363 522510 179373 522544
rect 179321 522498 179373 522510
rect 179767 522646 179819 522672
rect 179767 522612 179777 522646
rect 179811 522612 179819 522646
rect 179767 522544 179819 522612
rect 179767 522510 179777 522544
rect 179811 522510 179819 522544
rect 180057 522544 180109 522672
rect 179767 522498 179819 522510
rect 180057 522510 180065 522544
rect 180099 522510 180109 522544
rect 180057 522498 180109 522510
rect 181055 522544 181107 522672
rect 181055 522510 181065 522544
rect 181099 522510 181107 522544
rect 181055 522498 181107 522510
rect 181161 522544 181213 522672
rect 181161 522510 181169 522544
rect 181203 522510 181213 522544
rect 181161 522498 181213 522510
rect 182159 522544 182211 522672
rect 182159 522510 182169 522544
rect 182203 522510 182211 522544
rect 182159 522498 182211 522510
rect 182265 522544 182317 522672
rect 182265 522510 182273 522544
rect 182307 522510 182317 522544
rect 182265 522498 182317 522510
rect 183263 522544 183315 522672
rect 183263 522510 183273 522544
rect 183307 522510 183315 522544
rect 183263 522498 183315 522510
rect 183369 522544 183421 522672
rect 183369 522510 183377 522544
rect 183411 522510 183421 522544
rect 183369 522498 183421 522510
rect 184367 522544 184419 522672
rect 184367 522510 184377 522544
rect 184411 522510 184419 522544
rect 184367 522498 184419 522510
rect 184473 522646 184525 522672
rect 184473 522612 184481 522646
rect 184515 522612 184525 522646
rect 184473 522544 184525 522612
rect 184473 522510 184481 522544
rect 184515 522510 184525 522544
rect 184473 522498 184525 522510
rect 184919 522646 184971 522672
rect 184919 522612 184929 522646
rect 184963 522612 184971 522646
rect 184919 522544 184971 522612
rect 184919 522510 184929 522544
rect 184963 522510 184971 522544
rect 185209 522544 185261 522672
rect 184919 522498 184971 522510
rect 185209 522510 185217 522544
rect 185251 522510 185261 522544
rect 185209 522498 185261 522510
rect 186207 522544 186259 522672
rect 186207 522510 186217 522544
rect 186251 522510 186259 522544
rect 186207 522498 186259 522510
rect 186313 522646 186365 522672
rect 186313 522612 186321 522646
rect 186355 522612 186365 522646
rect 186313 522544 186365 522612
rect 186313 522510 186321 522544
rect 186355 522510 186365 522544
rect 186313 522498 186365 522510
rect 186943 522646 186995 522672
rect 186943 522612 186953 522646
rect 186987 522612 186995 522646
rect 186943 522544 186995 522612
rect 186943 522510 186953 522544
rect 186987 522510 186995 522544
rect 186943 522498 186995 522510
rect 187233 522639 187285 522672
rect 187233 522605 187241 522639
rect 187275 522605 187285 522639
rect 187233 522544 187285 522605
rect 187233 522510 187241 522544
rect 187275 522510 187285 522544
rect 187233 522498 187285 522510
rect 187403 522639 187455 522672
rect 187403 522605 187413 522639
rect 187447 522605 187455 522639
rect 187403 522544 187455 522605
rect 187403 522510 187413 522544
rect 187447 522510 187455 522544
rect 187403 522498 187455 522510
rect 172237 522392 172289 522404
rect 172237 522358 172245 522392
rect 172279 522358 172289 522392
rect 172237 522297 172289 522358
rect 172237 522263 172245 522297
rect 172279 522263 172289 522297
rect 172237 522230 172289 522263
rect 172407 522392 172459 522404
rect 172407 522358 172417 522392
rect 172451 522358 172459 522392
rect 172407 522297 172459 522358
rect 172407 522263 172417 522297
rect 172451 522263 172459 522297
rect 172407 522230 172459 522263
rect 172513 522392 172565 522404
rect 172513 522358 172521 522392
rect 172555 522358 172565 522392
rect 172513 522230 172565 522358
rect 173511 522392 173563 522404
rect 173511 522358 173521 522392
rect 173555 522358 173563 522392
rect 173511 522230 173563 522358
rect 173617 522392 173669 522404
rect 173617 522358 173625 522392
rect 173659 522358 173669 522392
rect 173617 522230 173669 522358
rect 174615 522392 174667 522404
rect 174615 522358 174625 522392
rect 174659 522358 174667 522392
rect 174615 522230 174667 522358
rect 174721 522392 174773 522404
rect 174721 522358 174729 522392
rect 174763 522358 174773 522392
rect 174721 522230 174773 522358
rect 175719 522392 175771 522404
rect 175719 522358 175729 522392
rect 175763 522358 175771 522392
rect 175719 522230 175771 522358
rect 175825 522392 175877 522404
rect 175825 522358 175833 522392
rect 175867 522358 175877 522392
rect 175825 522230 175877 522358
rect 176823 522392 176875 522404
rect 176823 522358 176833 522392
rect 176867 522358 176875 522392
rect 176823 522230 176875 522358
rect 176929 522392 176981 522404
rect 176929 522358 176937 522392
rect 176971 522358 176981 522392
rect 176929 522290 176981 522358
rect 176929 522256 176937 522290
rect 176971 522256 176981 522290
rect 176929 522230 176981 522256
rect 177191 522392 177243 522404
rect 177191 522358 177201 522392
rect 177235 522358 177243 522392
rect 177481 522392 177533 522404
rect 177191 522290 177243 522358
rect 177191 522256 177201 522290
rect 177235 522256 177243 522290
rect 177191 522230 177243 522256
rect 177481 522358 177489 522392
rect 177523 522358 177533 522392
rect 177481 522230 177533 522358
rect 178479 522392 178531 522404
rect 178479 522358 178489 522392
rect 178523 522358 178531 522392
rect 178479 522230 178531 522358
rect 178585 522392 178637 522404
rect 178585 522358 178593 522392
rect 178627 522358 178637 522392
rect 178585 522230 178637 522358
rect 179583 522392 179635 522404
rect 179583 522358 179593 522392
rect 179627 522358 179635 522392
rect 179583 522230 179635 522358
rect 179689 522392 179741 522404
rect 179689 522358 179697 522392
rect 179731 522358 179741 522392
rect 179689 522230 179741 522358
rect 180687 522392 180739 522404
rect 180687 522358 180697 522392
rect 180731 522358 180739 522392
rect 180687 522230 180739 522358
rect 180793 522392 180845 522404
rect 180793 522358 180801 522392
rect 180835 522358 180845 522392
rect 180793 522230 180845 522358
rect 181791 522392 181843 522404
rect 181791 522358 181801 522392
rect 181835 522358 181843 522392
rect 181791 522230 181843 522358
rect 181897 522392 181949 522404
rect 181897 522358 181905 522392
rect 181939 522358 181949 522392
rect 181897 522290 181949 522358
rect 181897 522256 181905 522290
rect 181939 522256 181949 522290
rect 181897 522230 181949 522256
rect 182343 522392 182395 522404
rect 182343 522358 182353 522392
rect 182387 522358 182395 522392
rect 182633 522392 182685 522404
rect 182343 522290 182395 522358
rect 182343 522256 182353 522290
rect 182387 522256 182395 522290
rect 182343 522230 182395 522256
rect 182633 522358 182641 522392
rect 182675 522358 182685 522392
rect 182633 522230 182685 522358
rect 183631 522392 183683 522404
rect 183631 522358 183641 522392
rect 183675 522358 183683 522392
rect 183631 522230 183683 522358
rect 183737 522392 183789 522404
rect 183737 522358 183745 522392
rect 183779 522358 183789 522392
rect 183737 522230 183789 522358
rect 184735 522392 184787 522404
rect 184735 522358 184745 522392
rect 184779 522358 184787 522392
rect 184735 522230 184787 522358
rect 184841 522392 184893 522404
rect 184841 522358 184849 522392
rect 184883 522358 184893 522392
rect 184841 522230 184893 522358
rect 185839 522392 185891 522404
rect 185839 522358 185849 522392
rect 185883 522358 185891 522392
rect 185839 522230 185891 522358
rect 185945 522392 185997 522404
rect 185945 522358 185953 522392
rect 185987 522358 185997 522392
rect 185945 522230 185997 522358
rect 186943 522392 186995 522404
rect 186943 522358 186953 522392
rect 186987 522358 186995 522392
rect 186943 522230 186995 522358
rect 187233 522392 187285 522404
rect 187233 522358 187241 522392
rect 187275 522358 187285 522392
rect 187233 522297 187285 522358
rect 187233 522263 187241 522297
rect 187275 522263 187285 522297
rect 187233 522230 187285 522263
rect 187403 522392 187455 522404
rect 187403 522358 187413 522392
rect 187447 522358 187455 522392
rect 187403 522297 187455 522358
rect 187403 522263 187413 522297
rect 187447 522263 187455 522297
rect 187403 522230 187455 522263
rect 172237 521551 172289 521584
rect 172237 521517 172245 521551
rect 172279 521517 172289 521551
rect 172237 521456 172289 521517
rect 172237 521422 172245 521456
rect 172279 521422 172289 521456
rect 172237 521410 172289 521422
rect 172407 521551 172459 521584
rect 172407 521517 172417 521551
rect 172451 521517 172459 521551
rect 172407 521456 172459 521517
rect 172407 521422 172417 521456
rect 172451 521422 172459 521456
rect 172407 521410 172459 521422
rect 172513 521456 172565 521584
rect 172513 521422 172521 521456
rect 172555 521422 172565 521456
rect 172513 521410 172565 521422
rect 173511 521456 173563 521584
rect 173511 521422 173521 521456
rect 173555 521422 173563 521456
rect 173511 521410 173563 521422
rect 173617 521456 173669 521584
rect 173617 521422 173625 521456
rect 173659 521422 173669 521456
rect 173617 521410 173669 521422
rect 174615 521456 174667 521584
rect 174615 521422 174625 521456
rect 174659 521422 174667 521456
rect 174905 521456 174957 521584
rect 174615 521410 174667 521422
rect 174905 521422 174913 521456
rect 174947 521422 174957 521456
rect 174905 521410 174957 521422
rect 175903 521456 175955 521584
rect 175903 521422 175913 521456
rect 175947 521422 175955 521456
rect 175903 521410 175955 521422
rect 176009 521456 176061 521584
rect 176009 521422 176017 521456
rect 176051 521422 176061 521456
rect 176009 521410 176061 521422
rect 177007 521456 177059 521584
rect 177007 521422 177017 521456
rect 177051 521422 177059 521456
rect 177007 521410 177059 521422
rect 177113 521456 177165 521584
rect 177113 521422 177121 521456
rect 177155 521422 177165 521456
rect 177113 521410 177165 521422
rect 178111 521456 178163 521584
rect 178111 521422 178121 521456
rect 178155 521422 178163 521456
rect 178111 521410 178163 521422
rect 178217 521456 178269 521584
rect 178217 521422 178225 521456
rect 178259 521422 178269 521456
rect 178217 521410 178269 521422
rect 179215 521456 179267 521584
rect 179215 521422 179225 521456
rect 179259 521422 179267 521456
rect 179215 521410 179267 521422
rect 179321 521558 179373 521584
rect 179321 521524 179329 521558
rect 179363 521524 179373 521558
rect 179321 521456 179373 521524
rect 179321 521422 179329 521456
rect 179363 521422 179373 521456
rect 179321 521410 179373 521422
rect 179767 521558 179819 521584
rect 179767 521524 179777 521558
rect 179811 521524 179819 521558
rect 179767 521456 179819 521524
rect 179767 521422 179777 521456
rect 179811 521422 179819 521456
rect 180057 521456 180109 521584
rect 179767 521410 179819 521422
rect 180057 521422 180065 521456
rect 180099 521422 180109 521456
rect 180057 521410 180109 521422
rect 181055 521456 181107 521584
rect 181055 521422 181065 521456
rect 181099 521422 181107 521456
rect 181055 521410 181107 521422
rect 181161 521456 181213 521584
rect 181161 521422 181169 521456
rect 181203 521422 181213 521456
rect 181161 521410 181213 521422
rect 182159 521456 182211 521584
rect 182159 521422 182169 521456
rect 182203 521422 182211 521456
rect 182159 521410 182211 521422
rect 182265 521456 182317 521584
rect 182265 521422 182273 521456
rect 182307 521422 182317 521456
rect 182265 521410 182317 521422
rect 183263 521456 183315 521584
rect 183263 521422 183273 521456
rect 183307 521422 183315 521456
rect 183263 521410 183315 521422
rect 183369 521456 183421 521584
rect 183369 521422 183377 521456
rect 183411 521422 183421 521456
rect 183369 521410 183421 521422
rect 184367 521456 184419 521584
rect 184367 521422 184377 521456
rect 184411 521422 184419 521456
rect 184367 521410 184419 521422
rect 184473 521558 184525 521584
rect 184473 521524 184481 521558
rect 184515 521524 184525 521558
rect 184473 521456 184525 521524
rect 184473 521422 184481 521456
rect 184515 521422 184525 521456
rect 184473 521410 184525 521422
rect 184919 521558 184971 521584
rect 184919 521524 184929 521558
rect 184963 521524 184971 521558
rect 184919 521456 184971 521524
rect 184919 521422 184929 521456
rect 184963 521422 184971 521456
rect 185209 521456 185261 521584
rect 184919 521410 184971 521422
rect 185209 521422 185217 521456
rect 185251 521422 185261 521456
rect 185209 521410 185261 521422
rect 186207 521456 186259 521584
rect 186207 521422 186217 521456
rect 186251 521422 186259 521456
rect 186207 521410 186259 521422
rect 186313 521558 186365 521584
rect 186313 521524 186321 521558
rect 186355 521524 186365 521558
rect 186313 521456 186365 521524
rect 186313 521422 186321 521456
rect 186355 521422 186365 521456
rect 186313 521410 186365 521422
rect 186943 521558 186995 521584
rect 186943 521524 186953 521558
rect 186987 521524 186995 521558
rect 186943 521456 186995 521524
rect 186943 521422 186953 521456
rect 186987 521422 186995 521456
rect 186943 521410 186995 521422
rect 187233 521551 187285 521584
rect 187233 521517 187241 521551
rect 187275 521517 187285 521551
rect 187233 521456 187285 521517
rect 187233 521422 187241 521456
rect 187275 521422 187285 521456
rect 187233 521410 187285 521422
rect 187403 521551 187455 521584
rect 187403 521517 187413 521551
rect 187447 521517 187455 521551
rect 187403 521456 187455 521517
rect 187403 521422 187413 521456
rect 187447 521422 187455 521456
rect 187403 521410 187455 521422
rect 172237 521304 172289 521316
rect 172237 521270 172245 521304
rect 172279 521270 172289 521304
rect 172237 521209 172289 521270
rect 172237 521175 172245 521209
rect 172279 521175 172289 521209
rect 172237 521142 172289 521175
rect 172407 521304 172459 521316
rect 172407 521270 172417 521304
rect 172451 521270 172459 521304
rect 172407 521209 172459 521270
rect 172407 521175 172417 521209
rect 172451 521175 172459 521209
rect 172407 521142 172459 521175
rect 172513 521304 172565 521316
rect 172513 521270 172521 521304
rect 172555 521270 172565 521304
rect 172513 521142 172565 521270
rect 173511 521304 173563 521316
rect 173511 521270 173521 521304
rect 173555 521270 173563 521304
rect 173511 521142 173563 521270
rect 173617 521304 173669 521316
rect 173617 521270 173625 521304
rect 173659 521270 173669 521304
rect 173617 521142 173669 521270
rect 174615 521304 174667 521316
rect 174615 521270 174625 521304
rect 174659 521270 174667 521304
rect 174615 521142 174667 521270
rect 174721 521304 174773 521316
rect 174721 521270 174729 521304
rect 174763 521270 174773 521304
rect 174721 521142 174773 521270
rect 175719 521304 175771 521316
rect 175719 521270 175729 521304
rect 175763 521270 175771 521304
rect 175719 521142 175771 521270
rect 175825 521304 175877 521316
rect 175825 521270 175833 521304
rect 175867 521270 175877 521304
rect 175825 521142 175877 521270
rect 176823 521304 176875 521316
rect 176823 521270 176833 521304
rect 176867 521270 176875 521304
rect 176823 521142 176875 521270
rect 176929 521304 176981 521316
rect 176929 521270 176937 521304
rect 176971 521270 176981 521304
rect 176929 521202 176981 521270
rect 176929 521168 176937 521202
rect 176971 521168 176981 521202
rect 176929 521142 176981 521168
rect 177191 521304 177243 521316
rect 177191 521270 177201 521304
rect 177235 521270 177243 521304
rect 177481 521304 177533 521316
rect 177191 521202 177243 521270
rect 177191 521168 177201 521202
rect 177235 521168 177243 521202
rect 177191 521142 177243 521168
rect 177481 521270 177489 521304
rect 177523 521270 177533 521304
rect 177481 521142 177533 521270
rect 178479 521304 178531 521316
rect 178479 521270 178489 521304
rect 178523 521270 178531 521304
rect 178479 521142 178531 521270
rect 178585 521304 178637 521316
rect 178585 521270 178593 521304
rect 178627 521270 178637 521304
rect 178585 521142 178637 521270
rect 179583 521304 179635 521316
rect 179583 521270 179593 521304
rect 179627 521270 179635 521304
rect 179583 521142 179635 521270
rect 179689 521304 179741 521316
rect 179689 521270 179697 521304
rect 179731 521270 179741 521304
rect 179689 521142 179741 521270
rect 180687 521304 180739 521316
rect 180687 521270 180697 521304
rect 180731 521270 180739 521304
rect 180687 521142 180739 521270
rect 180793 521304 180845 521316
rect 180793 521270 180801 521304
rect 180835 521270 180845 521304
rect 180793 521142 180845 521270
rect 181791 521304 181843 521316
rect 181791 521270 181801 521304
rect 181835 521270 181843 521304
rect 181791 521142 181843 521270
rect 181897 521304 181949 521316
rect 181897 521270 181905 521304
rect 181939 521270 181949 521304
rect 181897 521202 181949 521270
rect 181897 521168 181905 521202
rect 181939 521168 181949 521202
rect 181897 521142 181949 521168
rect 182343 521304 182395 521316
rect 182343 521270 182353 521304
rect 182387 521270 182395 521304
rect 182633 521304 182685 521316
rect 182343 521202 182395 521270
rect 182343 521168 182353 521202
rect 182387 521168 182395 521202
rect 182343 521142 182395 521168
rect 182633 521270 182641 521304
rect 182675 521270 182685 521304
rect 182633 521142 182685 521270
rect 183631 521304 183683 521316
rect 183631 521270 183641 521304
rect 183675 521270 183683 521304
rect 183631 521142 183683 521270
rect 183737 521304 183789 521316
rect 183737 521270 183745 521304
rect 183779 521270 183789 521304
rect 183737 521142 183789 521270
rect 184735 521304 184787 521316
rect 184735 521270 184745 521304
rect 184779 521270 184787 521304
rect 184735 521142 184787 521270
rect 184841 521304 184893 521316
rect 184841 521270 184849 521304
rect 184883 521270 184893 521304
rect 184841 521142 184893 521270
rect 185839 521304 185891 521316
rect 185839 521270 185849 521304
rect 185883 521270 185891 521304
rect 185839 521142 185891 521270
rect 185945 521304 185997 521316
rect 185945 521270 185953 521304
rect 185987 521270 185997 521304
rect 185945 521142 185997 521270
rect 186943 521304 186995 521316
rect 186943 521270 186953 521304
rect 186987 521270 186995 521304
rect 186943 521142 186995 521270
rect 187233 521304 187285 521316
rect 187233 521270 187241 521304
rect 187275 521270 187285 521304
rect 187233 521209 187285 521270
rect 187233 521175 187241 521209
rect 187275 521175 187285 521209
rect 187233 521142 187285 521175
rect 187403 521304 187455 521316
rect 187403 521270 187413 521304
rect 187447 521270 187455 521304
rect 187403 521209 187455 521270
rect 187403 521175 187413 521209
rect 187447 521175 187455 521209
rect 187403 521142 187455 521175
rect 172237 520463 172289 520496
rect 172237 520429 172245 520463
rect 172279 520429 172289 520463
rect 172237 520368 172289 520429
rect 172237 520334 172245 520368
rect 172279 520334 172289 520368
rect 172237 520322 172289 520334
rect 172407 520463 172459 520496
rect 172407 520429 172417 520463
rect 172451 520429 172459 520463
rect 172407 520368 172459 520429
rect 172407 520334 172417 520368
rect 172451 520334 172459 520368
rect 172407 520322 172459 520334
rect 172513 520368 172565 520496
rect 172513 520334 172521 520368
rect 172555 520334 172565 520368
rect 172513 520322 172565 520334
rect 173511 520368 173563 520496
rect 173511 520334 173521 520368
rect 173555 520334 173563 520368
rect 173511 520322 173563 520334
rect 173617 520368 173669 520496
rect 173617 520334 173625 520368
rect 173659 520334 173669 520368
rect 173617 520322 173669 520334
rect 174615 520368 174667 520496
rect 174615 520334 174625 520368
rect 174659 520334 174667 520368
rect 174905 520368 174957 520496
rect 174615 520322 174667 520334
rect 174905 520334 174913 520368
rect 174947 520334 174957 520368
rect 174905 520322 174957 520334
rect 175903 520368 175955 520496
rect 175903 520334 175913 520368
rect 175947 520334 175955 520368
rect 175903 520322 175955 520334
rect 176009 520368 176061 520496
rect 176009 520334 176017 520368
rect 176051 520334 176061 520368
rect 176009 520322 176061 520334
rect 177007 520368 177059 520496
rect 177007 520334 177017 520368
rect 177051 520334 177059 520368
rect 177007 520322 177059 520334
rect 177113 520368 177165 520496
rect 177113 520334 177121 520368
rect 177155 520334 177165 520368
rect 177113 520322 177165 520334
rect 178111 520368 178163 520496
rect 178111 520334 178121 520368
rect 178155 520334 178163 520368
rect 178111 520322 178163 520334
rect 178217 520368 178269 520496
rect 178217 520334 178225 520368
rect 178259 520334 178269 520368
rect 178217 520322 178269 520334
rect 179215 520368 179267 520496
rect 179215 520334 179225 520368
rect 179259 520334 179267 520368
rect 179215 520322 179267 520334
rect 179321 520470 179373 520496
rect 179321 520436 179329 520470
rect 179363 520436 179373 520470
rect 179321 520368 179373 520436
rect 179321 520334 179329 520368
rect 179363 520334 179373 520368
rect 179321 520322 179373 520334
rect 179767 520470 179819 520496
rect 179767 520436 179777 520470
rect 179811 520436 179819 520470
rect 179767 520368 179819 520436
rect 179767 520334 179777 520368
rect 179811 520334 179819 520368
rect 180057 520368 180109 520496
rect 179767 520322 179819 520334
rect 180057 520334 180065 520368
rect 180099 520334 180109 520368
rect 180057 520322 180109 520334
rect 181055 520368 181107 520496
rect 181055 520334 181065 520368
rect 181099 520334 181107 520368
rect 181055 520322 181107 520334
rect 181161 520368 181213 520496
rect 181161 520334 181169 520368
rect 181203 520334 181213 520368
rect 181161 520322 181213 520334
rect 182159 520368 182211 520496
rect 182159 520334 182169 520368
rect 182203 520334 182211 520368
rect 182159 520322 182211 520334
rect 182265 520368 182317 520496
rect 182265 520334 182273 520368
rect 182307 520334 182317 520368
rect 182265 520322 182317 520334
rect 183263 520368 183315 520496
rect 183263 520334 183273 520368
rect 183307 520334 183315 520368
rect 183263 520322 183315 520334
rect 183369 520368 183421 520496
rect 183369 520334 183377 520368
rect 183411 520334 183421 520368
rect 183369 520322 183421 520334
rect 184367 520368 184419 520496
rect 184367 520334 184377 520368
rect 184411 520334 184419 520368
rect 184367 520322 184419 520334
rect 184473 520470 184525 520496
rect 184473 520436 184481 520470
rect 184515 520436 184525 520470
rect 184473 520368 184525 520436
rect 184473 520334 184481 520368
rect 184515 520334 184525 520368
rect 184473 520322 184525 520334
rect 184919 520470 184971 520496
rect 184919 520436 184929 520470
rect 184963 520436 184971 520470
rect 184919 520368 184971 520436
rect 184919 520334 184929 520368
rect 184963 520334 184971 520368
rect 185209 520368 185261 520496
rect 184919 520322 184971 520334
rect 185209 520334 185217 520368
rect 185251 520334 185261 520368
rect 185209 520322 185261 520334
rect 186207 520368 186259 520496
rect 186207 520334 186217 520368
rect 186251 520334 186259 520368
rect 186207 520322 186259 520334
rect 186313 520470 186365 520496
rect 186313 520436 186321 520470
rect 186355 520436 186365 520470
rect 186313 520368 186365 520436
rect 186313 520334 186321 520368
rect 186355 520334 186365 520368
rect 186313 520322 186365 520334
rect 186943 520470 186995 520496
rect 186943 520436 186953 520470
rect 186987 520436 186995 520470
rect 186943 520368 186995 520436
rect 186943 520334 186953 520368
rect 186987 520334 186995 520368
rect 186943 520322 186995 520334
rect 187233 520463 187285 520496
rect 187233 520429 187241 520463
rect 187275 520429 187285 520463
rect 187233 520368 187285 520429
rect 187233 520334 187241 520368
rect 187275 520334 187285 520368
rect 187233 520322 187285 520334
rect 187403 520463 187455 520496
rect 187403 520429 187413 520463
rect 187447 520429 187455 520463
rect 187403 520368 187455 520429
rect 187403 520334 187413 520368
rect 187447 520334 187455 520368
rect 187403 520322 187455 520334
rect 172237 520216 172289 520228
rect 172237 520182 172245 520216
rect 172279 520182 172289 520216
rect 172237 520121 172289 520182
rect 172237 520087 172245 520121
rect 172279 520087 172289 520121
rect 172237 520054 172289 520087
rect 172407 520216 172459 520228
rect 172407 520182 172417 520216
rect 172451 520182 172459 520216
rect 172407 520121 172459 520182
rect 172407 520087 172417 520121
rect 172451 520087 172459 520121
rect 172407 520054 172459 520087
rect 172513 520216 172565 520228
rect 172513 520182 172521 520216
rect 172555 520182 172565 520216
rect 172513 520054 172565 520182
rect 173511 520216 173563 520228
rect 173511 520182 173521 520216
rect 173555 520182 173563 520216
rect 173511 520054 173563 520182
rect 173617 520216 173669 520228
rect 173617 520182 173625 520216
rect 173659 520182 173669 520216
rect 173617 520054 173669 520182
rect 174615 520216 174667 520228
rect 174615 520182 174625 520216
rect 174659 520182 174667 520216
rect 174615 520054 174667 520182
rect 174721 520216 174773 520228
rect 174721 520182 174729 520216
rect 174763 520182 174773 520216
rect 174721 520054 174773 520182
rect 175719 520216 175771 520228
rect 175719 520182 175729 520216
rect 175763 520182 175771 520216
rect 175719 520054 175771 520182
rect 175825 520216 175877 520228
rect 175825 520182 175833 520216
rect 175867 520182 175877 520216
rect 175825 520054 175877 520182
rect 176823 520216 176875 520228
rect 176823 520182 176833 520216
rect 176867 520182 176875 520216
rect 176823 520054 176875 520182
rect 176929 520216 176981 520228
rect 176929 520182 176937 520216
rect 176971 520182 176981 520216
rect 176929 520114 176981 520182
rect 176929 520080 176937 520114
rect 176971 520080 176981 520114
rect 176929 520054 176981 520080
rect 177191 520216 177243 520228
rect 177191 520182 177201 520216
rect 177235 520182 177243 520216
rect 177481 520216 177533 520228
rect 177191 520114 177243 520182
rect 177191 520080 177201 520114
rect 177235 520080 177243 520114
rect 177191 520054 177243 520080
rect 177481 520182 177489 520216
rect 177523 520182 177533 520216
rect 177481 520054 177533 520182
rect 178479 520216 178531 520228
rect 178479 520182 178489 520216
rect 178523 520182 178531 520216
rect 178479 520054 178531 520182
rect 178585 520216 178637 520228
rect 178585 520182 178593 520216
rect 178627 520182 178637 520216
rect 178585 520054 178637 520182
rect 179583 520216 179635 520228
rect 179583 520182 179593 520216
rect 179627 520182 179635 520216
rect 179583 520054 179635 520182
rect 179689 520216 179741 520228
rect 179689 520182 179697 520216
rect 179731 520182 179741 520216
rect 179689 520054 179741 520182
rect 180687 520216 180739 520228
rect 180687 520182 180697 520216
rect 180731 520182 180739 520216
rect 180687 520054 180739 520182
rect 180793 520216 180845 520228
rect 180793 520182 180801 520216
rect 180835 520182 180845 520216
rect 180793 520054 180845 520182
rect 181791 520216 181843 520228
rect 181791 520182 181801 520216
rect 181835 520182 181843 520216
rect 181791 520054 181843 520182
rect 181897 520216 181949 520228
rect 181897 520182 181905 520216
rect 181939 520182 181949 520216
rect 181897 520114 181949 520182
rect 181897 520080 181905 520114
rect 181939 520080 181949 520114
rect 181897 520054 181949 520080
rect 182343 520216 182395 520228
rect 182343 520182 182353 520216
rect 182387 520182 182395 520216
rect 182633 520216 182685 520228
rect 182343 520114 182395 520182
rect 182343 520080 182353 520114
rect 182387 520080 182395 520114
rect 182343 520054 182395 520080
rect 182633 520182 182641 520216
rect 182675 520182 182685 520216
rect 182633 520054 182685 520182
rect 183631 520216 183683 520228
rect 183631 520182 183641 520216
rect 183675 520182 183683 520216
rect 183631 520054 183683 520182
rect 183737 520216 183789 520228
rect 183737 520182 183745 520216
rect 183779 520182 183789 520216
rect 183737 520054 183789 520182
rect 184735 520216 184787 520228
rect 184735 520182 184745 520216
rect 184779 520182 184787 520216
rect 184735 520054 184787 520182
rect 184841 520216 184893 520228
rect 184841 520182 184849 520216
rect 184883 520182 184893 520216
rect 184841 520054 184893 520182
rect 185839 520216 185891 520228
rect 185839 520182 185849 520216
rect 185883 520182 185891 520216
rect 185839 520054 185891 520182
rect 185945 520216 185997 520228
rect 185945 520182 185953 520216
rect 185987 520182 185997 520216
rect 185945 520054 185997 520182
rect 186943 520216 186995 520228
rect 186943 520182 186953 520216
rect 186987 520182 186995 520216
rect 186943 520054 186995 520182
rect 187233 520216 187285 520228
rect 187233 520182 187241 520216
rect 187275 520182 187285 520216
rect 187233 520121 187285 520182
rect 187233 520087 187241 520121
rect 187275 520087 187285 520121
rect 187233 520054 187285 520087
rect 187403 520216 187455 520228
rect 187403 520182 187413 520216
rect 187447 520182 187455 520216
rect 187403 520121 187455 520182
rect 187403 520087 187413 520121
rect 187447 520087 187455 520121
rect 187403 520054 187455 520087
rect 172237 519375 172289 519408
rect 172237 519341 172245 519375
rect 172279 519341 172289 519375
rect 172237 519280 172289 519341
rect 172237 519246 172245 519280
rect 172279 519246 172289 519280
rect 172237 519234 172289 519246
rect 172407 519375 172459 519408
rect 172407 519341 172417 519375
rect 172451 519341 172459 519375
rect 172407 519280 172459 519341
rect 172407 519246 172417 519280
rect 172451 519246 172459 519280
rect 172407 519234 172459 519246
rect 172513 519280 172565 519408
rect 172513 519246 172521 519280
rect 172555 519246 172565 519280
rect 172513 519234 172565 519246
rect 173511 519280 173563 519408
rect 173511 519246 173521 519280
rect 173555 519246 173563 519280
rect 173511 519234 173563 519246
rect 173617 519280 173669 519408
rect 173617 519246 173625 519280
rect 173659 519246 173669 519280
rect 173617 519234 173669 519246
rect 174615 519280 174667 519408
rect 174615 519246 174625 519280
rect 174659 519246 174667 519280
rect 174905 519280 174957 519408
rect 174615 519234 174667 519246
rect 174905 519246 174913 519280
rect 174947 519246 174957 519280
rect 174905 519234 174957 519246
rect 175903 519280 175955 519408
rect 175903 519246 175913 519280
rect 175947 519246 175955 519280
rect 175903 519234 175955 519246
rect 176009 519280 176061 519408
rect 176009 519246 176017 519280
rect 176051 519246 176061 519280
rect 176009 519234 176061 519246
rect 177007 519280 177059 519408
rect 177007 519246 177017 519280
rect 177051 519246 177059 519280
rect 177007 519234 177059 519246
rect 177113 519280 177165 519408
rect 177113 519246 177121 519280
rect 177155 519246 177165 519280
rect 177113 519234 177165 519246
rect 178111 519280 178163 519408
rect 178111 519246 178121 519280
rect 178155 519246 178163 519280
rect 178111 519234 178163 519246
rect 178217 519280 178269 519408
rect 178217 519246 178225 519280
rect 178259 519246 178269 519280
rect 178217 519234 178269 519246
rect 179215 519280 179267 519408
rect 179215 519246 179225 519280
rect 179259 519246 179267 519280
rect 179215 519234 179267 519246
rect 179321 519382 179373 519408
rect 179321 519348 179329 519382
rect 179363 519348 179373 519382
rect 179321 519280 179373 519348
rect 179321 519246 179329 519280
rect 179363 519246 179373 519280
rect 179321 519234 179373 519246
rect 179767 519382 179819 519408
rect 179767 519348 179777 519382
rect 179811 519348 179819 519382
rect 179767 519280 179819 519348
rect 179767 519246 179777 519280
rect 179811 519246 179819 519280
rect 180057 519280 180109 519408
rect 179767 519234 179819 519246
rect 180057 519246 180065 519280
rect 180099 519246 180109 519280
rect 180057 519234 180109 519246
rect 181055 519280 181107 519408
rect 181055 519246 181065 519280
rect 181099 519246 181107 519280
rect 181055 519234 181107 519246
rect 181161 519280 181213 519408
rect 181161 519246 181169 519280
rect 181203 519246 181213 519280
rect 181161 519234 181213 519246
rect 182159 519280 182211 519408
rect 182159 519246 182169 519280
rect 182203 519246 182211 519280
rect 182159 519234 182211 519246
rect 182265 519280 182317 519408
rect 182265 519246 182273 519280
rect 182307 519246 182317 519280
rect 182265 519234 182317 519246
rect 183263 519280 183315 519408
rect 183263 519246 183273 519280
rect 183307 519246 183315 519280
rect 183263 519234 183315 519246
rect 183369 519280 183421 519408
rect 183369 519246 183377 519280
rect 183411 519246 183421 519280
rect 183369 519234 183421 519246
rect 184367 519280 184419 519408
rect 184367 519246 184377 519280
rect 184411 519246 184419 519280
rect 184367 519234 184419 519246
rect 184473 519382 184525 519408
rect 184473 519348 184481 519382
rect 184515 519348 184525 519382
rect 184473 519280 184525 519348
rect 184473 519246 184481 519280
rect 184515 519246 184525 519280
rect 184473 519234 184525 519246
rect 184919 519382 184971 519408
rect 184919 519348 184929 519382
rect 184963 519348 184971 519382
rect 184919 519280 184971 519348
rect 184919 519246 184929 519280
rect 184963 519246 184971 519280
rect 185209 519280 185261 519408
rect 184919 519234 184971 519246
rect 185209 519246 185217 519280
rect 185251 519246 185261 519280
rect 185209 519234 185261 519246
rect 186207 519280 186259 519408
rect 186207 519246 186217 519280
rect 186251 519246 186259 519280
rect 186207 519234 186259 519246
rect 186313 519382 186365 519408
rect 186313 519348 186321 519382
rect 186355 519348 186365 519382
rect 186313 519280 186365 519348
rect 186313 519246 186321 519280
rect 186355 519246 186365 519280
rect 186313 519234 186365 519246
rect 186943 519382 186995 519408
rect 186943 519348 186953 519382
rect 186987 519348 186995 519382
rect 186943 519280 186995 519348
rect 186943 519246 186953 519280
rect 186987 519246 186995 519280
rect 186943 519234 186995 519246
rect 187233 519375 187285 519408
rect 187233 519341 187241 519375
rect 187275 519341 187285 519375
rect 187233 519280 187285 519341
rect 187233 519246 187241 519280
rect 187275 519246 187285 519280
rect 187233 519234 187285 519246
rect 187403 519375 187455 519408
rect 187403 519341 187413 519375
rect 187447 519341 187455 519375
rect 187403 519280 187455 519341
rect 187403 519246 187413 519280
rect 187447 519246 187455 519280
rect 187403 519234 187455 519246
rect 172237 519128 172289 519140
rect 172237 519094 172245 519128
rect 172279 519094 172289 519128
rect 172237 519033 172289 519094
rect 172237 518999 172245 519033
rect 172279 518999 172289 519033
rect 172237 518966 172289 518999
rect 172407 519128 172459 519140
rect 172407 519094 172417 519128
rect 172451 519094 172459 519128
rect 172407 519033 172459 519094
rect 172407 518999 172417 519033
rect 172451 518999 172459 519033
rect 172407 518966 172459 518999
rect 172513 519128 172565 519140
rect 172513 519094 172521 519128
rect 172555 519094 172565 519128
rect 172513 518966 172565 519094
rect 173511 519128 173563 519140
rect 173511 519094 173521 519128
rect 173555 519094 173563 519128
rect 173511 518966 173563 519094
rect 173617 519128 173669 519140
rect 173617 519094 173625 519128
rect 173659 519094 173669 519128
rect 173617 518966 173669 519094
rect 174615 519128 174667 519140
rect 174615 519094 174625 519128
rect 174659 519094 174667 519128
rect 174615 518966 174667 519094
rect 174721 519128 174773 519140
rect 174721 519094 174729 519128
rect 174763 519094 174773 519128
rect 174721 518966 174773 519094
rect 175719 519128 175771 519140
rect 175719 519094 175729 519128
rect 175763 519094 175771 519128
rect 175719 518966 175771 519094
rect 175825 519128 175877 519140
rect 175825 519094 175833 519128
rect 175867 519094 175877 519128
rect 175825 518966 175877 519094
rect 176823 519128 176875 519140
rect 176823 519094 176833 519128
rect 176867 519094 176875 519128
rect 176823 518966 176875 519094
rect 176929 519128 176981 519140
rect 176929 519094 176937 519128
rect 176971 519094 176981 519128
rect 176929 519026 176981 519094
rect 176929 518992 176937 519026
rect 176971 518992 176981 519026
rect 176929 518966 176981 518992
rect 177191 519128 177243 519140
rect 177191 519094 177201 519128
rect 177235 519094 177243 519128
rect 177481 519128 177533 519140
rect 177191 519026 177243 519094
rect 177191 518992 177201 519026
rect 177235 518992 177243 519026
rect 177191 518966 177243 518992
rect 177481 519094 177489 519128
rect 177523 519094 177533 519128
rect 177481 518966 177533 519094
rect 178479 519128 178531 519140
rect 178479 519094 178489 519128
rect 178523 519094 178531 519128
rect 178479 518966 178531 519094
rect 178585 519128 178637 519140
rect 178585 519094 178593 519128
rect 178627 519094 178637 519128
rect 178585 518966 178637 519094
rect 179583 519128 179635 519140
rect 179583 519094 179593 519128
rect 179627 519094 179635 519128
rect 179583 518966 179635 519094
rect 179689 519128 179741 519140
rect 179689 519094 179697 519128
rect 179731 519094 179741 519128
rect 179689 518966 179741 519094
rect 180687 519128 180739 519140
rect 180687 519094 180697 519128
rect 180731 519094 180739 519128
rect 180687 518966 180739 519094
rect 180793 519128 180845 519140
rect 180793 519094 180801 519128
rect 180835 519094 180845 519128
rect 180793 518966 180845 519094
rect 181791 519128 181843 519140
rect 181791 519094 181801 519128
rect 181835 519094 181843 519128
rect 181791 518966 181843 519094
rect 181897 519128 181949 519140
rect 181897 519094 181905 519128
rect 181939 519094 181949 519128
rect 181897 519026 181949 519094
rect 181897 518992 181905 519026
rect 181939 518992 181949 519026
rect 181897 518966 181949 518992
rect 182343 519128 182395 519140
rect 182343 519094 182353 519128
rect 182387 519094 182395 519128
rect 182633 519128 182685 519140
rect 182343 519026 182395 519094
rect 182343 518992 182353 519026
rect 182387 518992 182395 519026
rect 182343 518966 182395 518992
rect 182633 519094 182641 519128
rect 182675 519094 182685 519128
rect 182633 518966 182685 519094
rect 183631 519128 183683 519140
rect 183631 519094 183641 519128
rect 183675 519094 183683 519128
rect 183631 518966 183683 519094
rect 183737 519128 183789 519140
rect 183737 519094 183745 519128
rect 183779 519094 183789 519128
rect 183737 518966 183789 519094
rect 184735 519128 184787 519140
rect 184735 519094 184745 519128
rect 184779 519094 184787 519128
rect 184735 518966 184787 519094
rect 184841 519128 184893 519140
rect 184841 519094 184849 519128
rect 184883 519094 184893 519128
rect 184841 518966 184893 519094
rect 185839 519128 185891 519140
rect 185839 519094 185849 519128
rect 185883 519094 185891 519128
rect 185839 518966 185891 519094
rect 185945 519128 185997 519140
rect 185945 519094 185953 519128
rect 185987 519094 185997 519128
rect 185945 518966 185997 519094
rect 186943 519128 186995 519140
rect 186943 519094 186953 519128
rect 186987 519094 186995 519128
rect 186943 518966 186995 519094
rect 187233 519128 187285 519140
rect 187233 519094 187241 519128
rect 187275 519094 187285 519128
rect 187233 519033 187285 519094
rect 187233 518999 187241 519033
rect 187275 518999 187285 519033
rect 187233 518966 187285 518999
rect 187403 519128 187455 519140
rect 187403 519094 187413 519128
rect 187447 519094 187455 519128
rect 187403 519033 187455 519094
rect 187403 518999 187413 519033
rect 187447 518999 187455 519033
rect 187403 518966 187455 518999
rect 172237 518287 172289 518320
rect 172237 518253 172245 518287
rect 172279 518253 172289 518287
rect 172237 518192 172289 518253
rect 172237 518158 172245 518192
rect 172279 518158 172289 518192
rect 172237 518146 172289 518158
rect 172407 518287 172459 518320
rect 172407 518253 172417 518287
rect 172451 518253 172459 518287
rect 172407 518192 172459 518253
rect 172407 518158 172417 518192
rect 172451 518158 172459 518192
rect 172407 518146 172459 518158
rect 172513 518192 172565 518320
rect 172513 518158 172521 518192
rect 172555 518158 172565 518192
rect 172513 518146 172565 518158
rect 173511 518192 173563 518320
rect 173511 518158 173521 518192
rect 173555 518158 173563 518192
rect 173511 518146 173563 518158
rect 173617 518192 173669 518320
rect 173617 518158 173625 518192
rect 173659 518158 173669 518192
rect 173617 518146 173669 518158
rect 174615 518192 174667 518320
rect 174615 518158 174625 518192
rect 174659 518158 174667 518192
rect 174905 518192 174957 518320
rect 174615 518146 174667 518158
rect 174905 518158 174913 518192
rect 174947 518158 174957 518192
rect 174905 518146 174957 518158
rect 175903 518192 175955 518320
rect 175903 518158 175913 518192
rect 175947 518158 175955 518192
rect 175903 518146 175955 518158
rect 176009 518192 176061 518320
rect 176009 518158 176017 518192
rect 176051 518158 176061 518192
rect 176009 518146 176061 518158
rect 177007 518192 177059 518320
rect 177007 518158 177017 518192
rect 177051 518158 177059 518192
rect 177007 518146 177059 518158
rect 177113 518192 177165 518320
rect 177113 518158 177121 518192
rect 177155 518158 177165 518192
rect 177113 518146 177165 518158
rect 178111 518192 178163 518320
rect 178111 518158 178121 518192
rect 178155 518158 178163 518192
rect 178111 518146 178163 518158
rect 178217 518192 178269 518320
rect 178217 518158 178225 518192
rect 178259 518158 178269 518192
rect 178217 518146 178269 518158
rect 179215 518192 179267 518320
rect 179215 518158 179225 518192
rect 179259 518158 179267 518192
rect 179215 518146 179267 518158
rect 179321 518294 179373 518320
rect 179321 518260 179329 518294
rect 179363 518260 179373 518294
rect 179321 518192 179373 518260
rect 179321 518158 179329 518192
rect 179363 518158 179373 518192
rect 179321 518146 179373 518158
rect 179767 518294 179819 518320
rect 179767 518260 179777 518294
rect 179811 518260 179819 518294
rect 179767 518192 179819 518260
rect 179767 518158 179777 518192
rect 179811 518158 179819 518192
rect 180057 518192 180109 518320
rect 179767 518146 179819 518158
rect 180057 518158 180065 518192
rect 180099 518158 180109 518192
rect 180057 518146 180109 518158
rect 181055 518192 181107 518320
rect 181055 518158 181065 518192
rect 181099 518158 181107 518192
rect 181055 518146 181107 518158
rect 181161 518192 181213 518320
rect 181161 518158 181169 518192
rect 181203 518158 181213 518192
rect 181161 518146 181213 518158
rect 182159 518192 182211 518320
rect 182159 518158 182169 518192
rect 182203 518158 182211 518192
rect 182159 518146 182211 518158
rect 182265 518192 182317 518320
rect 182265 518158 182273 518192
rect 182307 518158 182317 518192
rect 182265 518146 182317 518158
rect 183263 518192 183315 518320
rect 183263 518158 183273 518192
rect 183307 518158 183315 518192
rect 183263 518146 183315 518158
rect 183369 518192 183421 518320
rect 183369 518158 183377 518192
rect 183411 518158 183421 518192
rect 183369 518146 183421 518158
rect 184367 518192 184419 518320
rect 184367 518158 184377 518192
rect 184411 518158 184419 518192
rect 184367 518146 184419 518158
rect 184473 518294 184525 518320
rect 184473 518260 184481 518294
rect 184515 518260 184525 518294
rect 184473 518192 184525 518260
rect 184473 518158 184481 518192
rect 184515 518158 184525 518192
rect 184473 518146 184525 518158
rect 184919 518294 184971 518320
rect 184919 518260 184929 518294
rect 184963 518260 184971 518294
rect 184919 518192 184971 518260
rect 184919 518158 184929 518192
rect 184963 518158 184971 518192
rect 185209 518192 185261 518320
rect 184919 518146 184971 518158
rect 185209 518158 185217 518192
rect 185251 518158 185261 518192
rect 185209 518146 185261 518158
rect 186207 518192 186259 518320
rect 186207 518158 186217 518192
rect 186251 518158 186259 518192
rect 186207 518146 186259 518158
rect 186313 518294 186365 518320
rect 186313 518260 186321 518294
rect 186355 518260 186365 518294
rect 186313 518192 186365 518260
rect 186313 518158 186321 518192
rect 186355 518158 186365 518192
rect 186313 518146 186365 518158
rect 186943 518294 186995 518320
rect 186943 518260 186953 518294
rect 186987 518260 186995 518294
rect 186943 518192 186995 518260
rect 186943 518158 186953 518192
rect 186987 518158 186995 518192
rect 186943 518146 186995 518158
rect 187233 518287 187285 518320
rect 187233 518253 187241 518287
rect 187275 518253 187285 518287
rect 187233 518192 187285 518253
rect 187233 518158 187241 518192
rect 187275 518158 187285 518192
rect 187233 518146 187285 518158
rect 187403 518287 187455 518320
rect 187403 518253 187413 518287
rect 187447 518253 187455 518287
rect 187403 518192 187455 518253
rect 187403 518158 187413 518192
rect 187447 518158 187455 518192
rect 187403 518146 187455 518158
rect 172237 518040 172289 518052
rect 172237 518006 172245 518040
rect 172279 518006 172289 518040
rect 172237 517945 172289 518006
rect 172237 517911 172245 517945
rect 172279 517911 172289 517945
rect 172237 517878 172289 517911
rect 172407 518040 172459 518052
rect 172407 518006 172417 518040
rect 172451 518006 172459 518040
rect 172407 517945 172459 518006
rect 172407 517911 172417 517945
rect 172451 517911 172459 517945
rect 172407 517878 172459 517911
rect 172513 518040 172565 518052
rect 172513 518006 172521 518040
rect 172555 518006 172565 518040
rect 172513 517878 172565 518006
rect 173511 518040 173563 518052
rect 173511 518006 173521 518040
rect 173555 518006 173563 518040
rect 173511 517878 173563 518006
rect 173617 518040 173669 518052
rect 173617 518006 173625 518040
rect 173659 518006 173669 518040
rect 173617 517878 173669 518006
rect 174615 518040 174667 518052
rect 174615 518006 174625 518040
rect 174659 518006 174667 518040
rect 174615 517878 174667 518006
rect 174721 518040 174773 518052
rect 174721 518006 174729 518040
rect 174763 518006 174773 518040
rect 174721 517878 174773 518006
rect 175719 518040 175771 518052
rect 175719 518006 175729 518040
rect 175763 518006 175771 518040
rect 175719 517878 175771 518006
rect 175825 518040 175877 518052
rect 175825 518006 175833 518040
rect 175867 518006 175877 518040
rect 175825 517878 175877 518006
rect 176823 518040 176875 518052
rect 176823 518006 176833 518040
rect 176867 518006 176875 518040
rect 176823 517878 176875 518006
rect 176929 518040 176981 518052
rect 176929 518006 176937 518040
rect 176971 518006 176981 518040
rect 176929 517938 176981 518006
rect 176929 517904 176937 517938
rect 176971 517904 176981 517938
rect 176929 517878 176981 517904
rect 177191 518040 177243 518052
rect 177191 518006 177201 518040
rect 177235 518006 177243 518040
rect 177481 518040 177533 518052
rect 177191 517938 177243 518006
rect 177191 517904 177201 517938
rect 177235 517904 177243 517938
rect 177191 517878 177243 517904
rect 177481 518006 177489 518040
rect 177523 518006 177533 518040
rect 177481 517878 177533 518006
rect 178479 518040 178531 518052
rect 178479 518006 178489 518040
rect 178523 518006 178531 518040
rect 178479 517878 178531 518006
rect 178585 518040 178637 518052
rect 178585 518006 178593 518040
rect 178627 518006 178637 518040
rect 178585 517878 178637 518006
rect 179583 518040 179635 518052
rect 179583 518006 179593 518040
rect 179627 518006 179635 518040
rect 179583 517878 179635 518006
rect 179689 518040 179741 518052
rect 179689 518006 179697 518040
rect 179731 518006 179741 518040
rect 179689 517878 179741 518006
rect 180687 518040 180739 518052
rect 180687 518006 180697 518040
rect 180731 518006 180739 518040
rect 180687 517878 180739 518006
rect 180793 518040 180845 518052
rect 180793 518006 180801 518040
rect 180835 518006 180845 518040
rect 180793 517878 180845 518006
rect 181791 518040 181843 518052
rect 181791 518006 181801 518040
rect 181835 518006 181843 518040
rect 181791 517878 181843 518006
rect 181897 518040 181949 518052
rect 181897 518006 181905 518040
rect 181939 518006 181949 518040
rect 181897 517938 181949 518006
rect 181897 517904 181905 517938
rect 181939 517904 181949 517938
rect 181897 517878 181949 517904
rect 182343 518040 182395 518052
rect 182343 518006 182353 518040
rect 182387 518006 182395 518040
rect 182633 518040 182685 518052
rect 182343 517938 182395 518006
rect 182343 517904 182353 517938
rect 182387 517904 182395 517938
rect 182343 517878 182395 517904
rect 182633 518006 182641 518040
rect 182675 518006 182685 518040
rect 182633 517878 182685 518006
rect 183631 518040 183683 518052
rect 183631 518006 183641 518040
rect 183675 518006 183683 518040
rect 183631 517878 183683 518006
rect 183737 518040 183789 518052
rect 183737 518006 183745 518040
rect 183779 518006 183789 518040
rect 183737 517878 183789 518006
rect 184735 518040 184787 518052
rect 184735 518006 184745 518040
rect 184779 518006 184787 518040
rect 184735 517878 184787 518006
rect 184841 518040 184893 518052
rect 184841 518006 184849 518040
rect 184883 518006 184893 518040
rect 184841 517878 184893 518006
rect 185839 518040 185891 518052
rect 185839 518006 185849 518040
rect 185883 518006 185891 518040
rect 185839 517878 185891 518006
rect 185945 518040 185997 518052
rect 185945 518006 185953 518040
rect 185987 518006 185997 518040
rect 185945 517878 185997 518006
rect 186943 518040 186995 518052
rect 186943 518006 186953 518040
rect 186987 518006 186995 518040
rect 186943 517878 186995 518006
rect 187233 518040 187285 518052
rect 187233 518006 187241 518040
rect 187275 518006 187285 518040
rect 187233 517945 187285 518006
rect 187233 517911 187241 517945
rect 187275 517911 187285 517945
rect 187233 517878 187285 517911
rect 187403 518040 187455 518052
rect 187403 518006 187413 518040
rect 187447 518006 187455 518040
rect 187403 517945 187455 518006
rect 187403 517911 187413 517945
rect 187447 517911 187455 517945
rect 187403 517878 187455 517911
rect 172237 517199 172289 517232
rect 172237 517165 172245 517199
rect 172279 517165 172289 517199
rect 172237 517104 172289 517165
rect 172237 517070 172245 517104
rect 172279 517070 172289 517104
rect 172237 517058 172289 517070
rect 172407 517199 172459 517232
rect 172407 517165 172417 517199
rect 172451 517165 172459 517199
rect 172407 517104 172459 517165
rect 172407 517070 172417 517104
rect 172451 517070 172459 517104
rect 172407 517058 172459 517070
rect 172513 517104 172565 517232
rect 172513 517070 172521 517104
rect 172555 517070 172565 517104
rect 172513 517058 172565 517070
rect 173511 517104 173563 517232
rect 173511 517070 173521 517104
rect 173555 517070 173563 517104
rect 173511 517058 173563 517070
rect 173617 517104 173669 517232
rect 173617 517070 173625 517104
rect 173659 517070 173669 517104
rect 173617 517058 173669 517070
rect 174615 517104 174667 517232
rect 174615 517070 174625 517104
rect 174659 517070 174667 517104
rect 174905 517104 174957 517232
rect 174615 517058 174667 517070
rect 174905 517070 174913 517104
rect 174947 517070 174957 517104
rect 174905 517058 174957 517070
rect 175903 517104 175955 517232
rect 175903 517070 175913 517104
rect 175947 517070 175955 517104
rect 175903 517058 175955 517070
rect 176009 517104 176061 517232
rect 176009 517070 176017 517104
rect 176051 517070 176061 517104
rect 176009 517058 176061 517070
rect 177007 517104 177059 517232
rect 177007 517070 177017 517104
rect 177051 517070 177059 517104
rect 177007 517058 177059 517070
rect 177113 517104 177165 517232
rect 177113 517070 177121 517104
rect 177155 517070 177165 517104
rect 177113 517058 177165 517070
rect 178111 517104 178163 517232
rect 178111 517070 178121 517104
rect 178155 517070 178163 517104
rect 178111 517058 178163 517070
rect 178217 517104 178269 517232
rect 178217 517070 178225 517104
rect 178259 517070 178269 517104
rect 178217 517058 178269 517070
rect 179215 517104 179267 517232
rect 179215 517070 179225 517104
rect 179259 517070 179267 517104
rect 179215 517058 179267 517070
rect 179321 517206 179373 517232
rect 179321 517172 179329 517206
rect 179363 517172 179373 517206
rect 179321 517104 179373 517172
rect 179321 517070 179329 517104
rect 179363 517070 179373 517104
rect 179321 517058 179373 517070
rect 179767 517206 179819 517232
rect 179767 517172 179777 517206
rect 179811 517172 179819 517206
rect 179767 517104 179819 517172
rect 179767 517070 179777 517104
rect 179811 517070 179819 517104
rect 180057 517104 180109 517232
rect 179767 517058 179819 517070
rect 180057 517070 180065 517104
rect 180099 517070 180109 517104
rect 180057 517058 180109 517070
rect 181055 517104 181107 517232
rect 181055 517070 181065 517104
rect 181099 517070 181107 517104
rect 181055 517058 181107 517070
rect 181161 517104 181213 517232
rect 181161 517070 181169 517104
rect 181203 517070 181213 517104
rect 181161 517058 181213 517070
rect 182159 517104 182211 517232
rect 182159 517070 182169 517104
rect 182203 517070 182211 517104
rect 182159 517058 182211 517070
rect 182265 517104 182317 517232
rect 182265 517070 182273 517104
rect 182307 517070 182317 517104
rect 182265 517058 182317 517070
rect 183263 517104 183315 517232
rect 183263 517070 183273 517104
rect 183307 517070 183315 517104
rect 183263 517058 183315 517070
rect 183369 517104 183421 517232
rect 183369 517070 183377 517104
rect 183411 517070 183421 517104
rect 183369 517058 183421 517070
rect 184367 517104 184419 517232
rect 184367 517070 184377 517104
rect 184411 517070 184419 517104
rect 184367 517058 184419 517070
rect 184473 517206 184525 517232
rect 184473 517172 184481 517206
rect 184515 517172 184525 517206
rect 184473 517104 184525 517172
rect 184473 517070 184481 517104
rect 184515 517070 184525 517104
rect 184473 517058 184525 517070
rect 184919 517206 184971 517232
rect 184919 517172 184929 517206
rect 184963 517172 184971 517206
rect 184919 517104 184971 517172
rect 184919 517070 184929 517104
rect 184963 517070 184971 517104
rect 185209 517104 185261 517232
rect 184919 517058 184971 517070
rect 185209 517070 185217 517104
rect 185251 517070 185261 517104
rect 185209 517058 185261 517070
rect 186207 517104 186259 517232
rect 186207 517070 186217 517104
rect 186251 517070 186259 517104
rect 186207 517058 186259 517070
rect 186313 517206 186365 517232
rect 186313 517172 186321 517206
rect 186355 517172 186365 517206
rect 186313 517104 186365 517172
rect 186313 517070 186321 517104
rect 186355 517070 186365 517104
rect 186313 517058 186365 517070
rect 186943 517206 186995 517232
rect 186943 517172 186953 517206
rect 186987 517172 186995 517206
rect 186943 517104 186995 517172
rect 186943 517070 186953 517104
rect 186987 517070 186995 517104
rect 186943 517058 186995 517070
rect 187233 517199 187285 517232
rect 187233 517165 187241 517199
rect 187275 517165 187285 517199
rect 187233 517104 187285 517165
rect 187233 517070 187241 517104
rect 187275 517070 187285 517104
rect 187233 517058 187285 517070
rect 187403 517199 187455 517232
rect 187403 517165 187413 517199
rect 187447 517165 187455 517199
rect 187403 517104 187455 517165
rect 187403 517070 187413 517104
rect 187447 517070 187455 517104
rect 187403 517058 187455 517070
rect 172237 516952 172289 516964
rect 172237 516918 172245 516952
rect 172279 516918 172289 516952
rect 172237 516857 172289 516918
rect 172237 516823 172245 516857
rect 172279 516823 172289 516857
rect 172237 516790 172289 516823
rect 172407 516952 172459 516964
rect 172407 516918 172417 516952
rect 172451 516918 172459 516952
rect 172407 516857 172459 516918
rect 172407 516823 172417 516857
rect 172451 516823 172459 516857
rect 172407 516790 172459 516823
rect 172513 516952 172565 516964
rect 172513 516918 172521 516952
rect 172555 516918 172565 516952
rect 172513 516790 172565 516918
rect 173511 516952 173563 516964
rect 173511 516918 173521 516952
rect 173555 516918 173563 516952
rect 173511 516790 173563 516918
rect 173617 516952 173669 516964
rect 173617 516918 173625 516952
rect 173659 516918 173669 516952
rect 173617 516790 173669 516918
rect 174615 516952 174667 516964
rect 174615 516918 174625 516952
rect 174659 516918 174667 516952
rect 174615 516790 174667 516918
rect 174721 516952 174773 516964
rect 174721 516918 174729 516952
rect 174763 516918 174773 516952
rect 174721 516790 174773 516918
rect 175719 516952 175771 516964
rect 175719 516918 175729 516952
rect 175763 516918 175771 516952
rect 175719 516790 175771 516918
rect 175825 516952 175877 516964
rect 175825 516918 175833 516952
rect 175867 516918 175877 516952
rect 175825 516790 175877 516918
rect 176823 516952 176875 516964
rect 176823 516918 176833 516952
rect 176867 516918 176875 516952
rect 176823 516790 176875 516918
rect 176929 516952 176981 516964
rect 176929 516918 176937 516952
rect 176971 516918 176981 516952
rect 176929 516850 176981 516918
rect 176929 516816 176937 516850
rect 176971 516816 176981 516850
rect 176929 516790 176981 516816
rect 177191 516952 177243 516964
rect 177191 516918 177201 516952
rect 177235 516918 177243 516952
rect 177481 516952 177533 516964
rect 177191 516850 177243 516918
rect 177191 516816 177201 516850
rect 177235 516816 177243 516850
rect 177191 516790 177243 516816
rect 177481 516918 177489 516952
rect 177523 516918 177533 516952
rect 177481 516790 177533 516918
rect 178479 516952 178531 516964
rect 178479 516918 178489 516952
rect 178523 516918 178531 516952
rect 178479 516790 178531 516918
rect 178585 516952 178637 516964
rect 178585 516918 178593 516952
rect 178627 516918 178637 516952
rect 178585 516790 178637 516918
rect 179583 516952 179635 516964
rect 179583 516918 179593 516952
rect 179627 516918 179635 516952
rect 179583 516790 179635 516918
rect 179689 516952 179741 516964
rect 179689 516918 179697 516952
rect 179731 516918 179741 516952
rect 179689 516790 179741 516918
rect 180687 516952 180739 516964
rect 180687 516918 180697 516952
rect 180731 516918 180739 516952
rect 180687 516790 180739 516918
rect 180793 516952 180845 516964
rect 180793 516918 180801 516952
rect 180835 516918 180845 516952
rect 180793 516790 180845 516918
rect 181791 516952 181843 516964
rect 181791 516918 181801 516952
rect 181835 516918 181843 516952
rect 181791 516790 181843 516918
rect 181897 516952 181949 516964
rect 181897 516918 181905 516952
rect 181939 516918 181949 516952
rect 181897 516850 181949 516918
rect 181897 516816 181905 516850
rect 181939 516816 181949 516850
rect 181897 516790 181949 516816
rect 182343 516952 182395 516964
rect 182343 516918 182353 516952
rect 182387 516918 182395 516952
rect 182633 516952 182685 516964
rect 182343 516850 182395 516918
rect 182343 516816 182353 516850
rect 182387 516816 182395 516850
rect 182343 516790 182395 516816
rect 182633 516918 182641 516952
rect 182675 516918 182685 516952
rect 182633 516790 182685 516918
rect 183631 516952 183683 516964
rect 183631 516918 183641 516952
rect 183675 516918 183683 516952
rect 183631 516790 183683 516918
rect 183737 516952 183789 516964
rect 183737 516918 183745 516952
rect 183779 516918 183789 516952
rect 183737 516790 183789 516918
rect 184735 516952 184787 516964
rect 184735 516918 184745 516952
rect 184779 516918 184787 516952
rect 184735 516790 184787 516918
rect 184841 516952 184893 516964
rect 184841 516918 184849 516952
rect 184883 516918 184893 516952
rect 184841 516790 184893 516918
rect 185839 516952 185891 516964
rect 185839 516918 185849 516952
rect 185883 516918 185891 516952
rect 185839 516790 185891 516918
rect 185945 516952 185997 516964
rect 185945 516918 185953 516952
rect 185987 516918 185997 516952
rect 185945 516790 185997 516918
rect 186943 516952 186995 516964
rect 186943 516918 186953 516952
rect 186987 516918 186995 516952
rect 186943 516790 186995 516918
rect 187233 516952 187285 516964
rect 187233 516918 187241 516952
rect 187275 516918 187285 516952
rect 187233 516857 187285 516918
rect 187233 516823 187241 516857
rect 187275 516823 187285 516857
rect 187233 516790 187285 516823
rect 187403 516952 187455 516964
rect 187403 516918 187413 516952
rect 187447 516918 187455 516952
rect 187403 516857 187455 516918
rect 187403 516823 187413 516857
rect 187447 516823 187455 516857
rect 187403 516790 187455 516823
rect 172237 516111 172289 516144
rect 172237 516077 172245 516111
rect 172279 516077 172289 516111
rect 172237 516016 172289 516077
rect 172237 515982 172245 516016
rect 172279 515982 172289 516016
rect 172237 515970 172289 515982
rect 172407 516111 172459 516144
rect 172407 516077 172417 516111
rect 172451 516077 172459 516111
rect 172407 516016 172459 516077
rect 172407 515982 172417 516016
rect 172451 515982 172459 516016
rect 172407 515970 172459 515982
rect 172513 516016 172565 516144
rect 172513 515982 172521 516016
rect 172555 515982 172565 516016
rect 172513 515970 172565 515982
rect 173511 516016 173563 516144
rect 173511 515982 173521 516016
rect 173555 515982 173563 516016
rect 173511 515970 173563 515982
rect 173617 516016 173669 516144
rect 173617 515982 173625 516016
rect 173659 515982 173669 516016
rect 173617 515970 173669 515982
rect 174615 516016 174667 516144
rect 174615 515982 174625 516016
rect 174659 515982 174667 516016
rect 174905 516016 174957 516144
rect 174615 515970 174667 515982
rect 174905 515982 174913 516016
rect 174947 515982 174957 516016
rect 174905 515970 174957 515982
rect 175903 516016 175955 516144
rect 175903 515982 175913 516016
rect 175947 515982 175955 516016
rect 175903 515970 175955 515982
rect 176009 516016 176061 516144
rect 176009 515982 176017 516016
rect 176051 515982 176061 516016
rect 176009 515970 176061 515982
rect 177007 516016 177059 516144
rect 177007 515982 177017 516016
rect 177051 515982 177059 516016
rect 177007 515970 177059 515982
rect 177113 516016 177165 516144
rect 177113 515982 177121 516016
rect 177155 515982 177165 516016
rect 177113 515970 177165 515982
rect 178111 516016 178163 516144
rect 178111 515982 178121 516016
rect 178155 515982 178163 516016
rect 178111 515970 178163 515982
rect 178217 516016 178269 516144
rect 178217 515982 178225 516016
rect 178259 515982 178269 516016
rect 178217 515970 178269 515982
rect 179215 516016 179267 516144
rect 179215 515982 179225 516016
rect 179259 515982 179267 516016
rect 179215 515970 179267 515982
rect 179321 516118 179373 516144
rect 179321 516084 179329 516118
rect 179363 516084 179373 516118
rect 179321 516016 179373 516084
rect 179321 515982 179329 516016
rect 179363 515982 179373 516016
rect 179321 515970 179373 515982
rect 179767 516118 179819 516144
rect 179767 516084 179777 516118
rect 179811 516084 179819 516118
rect 179767 516016 179819 516084
rect 179767 515982 179777 516016
rect 179811 515982 179819 516016
rect 180057 516016 180109 516144
rect 179767 515970 179819 515982
rect 180057 515982 180065 516016
rect 180099 515982 180109 516016
rect 180057 515970 180109 515982
rect 181055 516016 181107 516144
rect 181055 515982 181065 516016
rect 181099 515982 181107 516016
rect 181055 515970 181107 515982
rect 181161 516016 181213 516144
rect 181161 515982 181169 516016
rect 181203 515982 181213 516016
rect 181161 515970 181213 515982
rect 182159 516016 182211 516144
rect 182159 515982 182169 516016
rect 182203 515982 182211 516016
rect 182159 515970 182211 515982
rect 182265 516016 182317 516144
rect 182265 515982 182273 516016
rect 182307 515982 182317 516016
rect 182265 515970 182317 515982
rect 183263 516016 183315 516144
rect 183263 515982 183273 516016
rect 183307 515982 183315 516016
rect 183263 515970 183315 515982
rect 183369 516016 183421 516144
rect 183369 515982 183377 516016
rect 183411 515982 183421 516016
rect 183369 515970 183421 515982
rect 184367 516016 184419 516144
rect 184367 515982 184377 516016
rect 184411 515982 184419 516016
rect 184367 515970 184419 515982
rect 184473 516118 184525 516144
rect 184473 516084 184481 516118
rect 184515 516084 184525 516118
rect 184473 516016 184525 516084
rect 184473 515982 184481 516016
rect 184515 515982 184525 516016
rect 184473 515970 184525 515982
rect 184919 516118 184971 516144
rect 184919 516084 184929 516118
rect 184963 516084 184971 516118
rect 184919 516016 184971 516084
rect 184919 515982 184929 516016
rect 184963 515982 184971 516016
rect 185209 516016 185261 516144
rect 184919 515970 184971 515982
rect 185209 515982 185217 516016
rect 185251 515982 185261 516016
rect 185209 515970 185261 515982
rect 186207 516016 186259 516144
rect 186207 515982 186217 516016
rect 186251 515982 186259 516016
rect 186207 515970 186259 515982
rect 186313 516118 186365 516144
rect 186313 516084 186321 516118
rect 186355 516084 186365 516118
rect 186313 516016 186365 516084
rect 186313 515982 186321 516016
rect 186355 515982 186365 516016
rect 186313 515970 186365 515982
rect 186943 516118 186995 516144
rect 186943 516084 186953 516118
rect 186987 516084 186995 516118
rect 186943 516016 186995 516084
rect 186943 515982 186953 516016
rect 186987 515982 186995 516016
rect 186943 515970 186995 515982
rect 187233 516111 187285 516144
rect 187233 516077 187241 516111
rect 187275 516077 187285 516111
rect 187233 516016 187285 516077
rect 187233 515982 187241 516016
rect 187275 515982 187285 516016
rect 187233 515970 187285 515982
rect 187403 516111 187455 516144
rect 187403 516077 187413 516111
rect 187447 516077 187455 516111
rect 187403 516016 187455 516077
rect 187403 515982 187413 516016
rect 187447 515982 187455 516016
rect 187403 515970 187455 515982
rect 172237 515864 172289 515876
rect 172237 515830 172245 515864
rect 172279 515830 172289 515864
rect 172237 515769 172289 515830
rect 172237 515735 172245 515769
rect 172279 515735 172289 515769
rect 172237 515702 172289 515735
rect 172407 515864 172459 515876
rect 172407 515830 172417 515864
rect 172451 515830 172459 515864
rect 172407 515769 172459 515830
rect 172407 515735 172417 515769
rect 172451 515735 172459 515769
rect 172407 515702 172459 515735
rect 172513 515864 172565 515876
rect 172513 515830 172521 515864
rect 172555 515830 172565 515864
rect 172513 515762 172565 515830
rect 172513 515728 172521 515762
rect 172555 515728 172565 515762
rect 172513 515702 172565 515728
rect 173143 515864 173195 515876
rect 173143 515830 173153 515864
rect 173187 515830 173195 515864
rect 173143 515762 173195 515830
rect 173143 515728 173153 515762
rect 173187 515728 173195 515762
rect 173143 515702 173195 515728
rect 173433 515856 173486 515876
rect 173433 515822 173441 515856
rect 173475 515822 173486 515856
rect 173433 515734 173486 515822
rect 173433 515700 173441 515734
rect 173475 515700 173486 515734
rect 173433 515676 173486 515700
rect 173516 515864 173582 515876
rect 173516 515830 173527 515864
rect 173561 515830 173582 515864
rect 173516 515796 173582 515830
rect 173516 515762 173527 515796
rect 173561 515762 173582 515796
rect 173516 515676 173582 515762
rect 173612 515829 173668 515876
rect 173612 515795 173623 515829
rect 173657 515795 173668 515829
rect 173612 515676 173668 515795
rect 173698 515864 173754 515876
rect 173698 515830 173709 515864
rect 173743 515830 173754 515864
rect 173698 515676 173754 515830
rect 173784 515856 173840 515876
rect 173784 515822 173795 515856
rect 173829 515822 173840 515856
rect 173784 515788 173840 515822
rect 173784 515754 173795 515788
rect 173829 515754 173840 515788
rect 173784 515720 173840 515754
rect 173784 515686 173795 515720
rect 173829 515686 173840 515720
rect 173784 515676 173840 515686
rect 173870 515850 173930 515876
rect 173870 515816 173881 515850
rect 173915 515816 173930 515850
rect 173870 515782 173930 515816
rect 173870 515748 173881 515782
rect 173915 515748 173930 515782
rect 173870 515676 173930 515748
rect 173985 515864 174037 515876
rect 173985 515830 173993 515864
rect 174027 515830 174037 515864
rect 173985 515762 174037 515830
rect 173985 515728 173993 515762
rect 174027 515728 174037 515762
rect 173985 515702 174037 515728
rect 174615 515864 174667 515876
rect 174615 515830 174625 515864
rect 174659 515830 174667 515864
rect 174905 515864 174957 515876
rect 174615 515762 174667 515830
rect 174615 515728 174625 515762
rect 174659 515728 174667 515762
rect 174615 515702 174667 515728
rect 174905 515830 174913 515864
rect 174947 515830 174957 515864
rect 174905 515702 174957 515830
rect 175903 515864 175955 515876
rect 175903 515830 175913 515864
rect 175947 515830 175955 515864
rect 175903 515702 175955 515830
rect 176009 515864 176061 515876
rect 176009 515830 176017 515864
rect 176051 515830 176061 515864
rect 176009 515702 176061 515830
rect 177007 515864 177059 515876
rect 177007 515830 177017 515864
rect 177051 515830 177059 515864
rect 177007 515702 177059 515830
rect 177113 515864 177165 515876
rect 177113 515830 177121 515864
rect 177155 515830 177165 515864
rect 177113 515769 177165 515830
rect 177113 515735 177121 515769
rect 177155 515735 177165 515769
rect 177113 515702 177165 515735
rect 177283 515864 177335 515876
rect 177283 515830 177293 515864
rect 177327 515830 177335 515864
rect 177481 515864 177533 515876
rect 177283 515769 177335 515830
rect 177283 515735 177293 515769
rect 177327 515735 177335 515769
rect 177283 515702 177335 515735
rect 177481 515830 177489 515864
rect 177523 515830 177533 515864
rect 177481 515702 177533 515830
rect 178479 515864 178531 515876
rect 178479 515830 178489 515864
rect 178523 515830 178531 515864
rect 178479 515702 178531 515830
rect 178585 515864 178637 515876
rect 178585 515830 178593 515864
rect 178627 515830 178637 515864
rect 178585 515702 178637 515830
rect 179583 515864 179635 515876
rect 179583 515830 179593 515864
rect 179627 515830 179635 515864
rect 179583 515702 179635 515830
rect 179689 515864 179741 515876
rect 179689 515830 179697 515864
rect 179731 515830 179741 515864
rect 179689 515769 179741 515830
rect 179689 515735 179697 515769
rect 179731 515735 179741 515769
rect 179689 515702 179741 515735
rect 179859 515864 179911 515876
rect 179859 515830 179869 515864
rect 179903 515830 179911 515864
rect 180057 515864 180109 515876
rect 179859 515769 179911 515830
rect 179859 515735 179869 515769
rect 179903 515735 179911 515769
rect 179859 515702 179911 515735
rect 180057 515830 180065 515864
rect 180099 515830 180109 515864
rect 180057 515702 180109 515830
rect 181055 515864 181107 515876
rect 181055 515830 181065 515864
rect 181099 515830 181107 515864
rect 181055 515702 181107 515830
rect 181161 515864 181213 515876
rect 181161 515830 181169 515864
rect 181203 515830 181213 515864
rect 181161 515762 181213 515830
rect 181161 515728 181169 515762
rect 181203 515728 181213 515762
rect 181161 515702 181213 515728
rect 181791 515864 181843 515876
rect 181791 515830 181801 515864
rect 181835 515830 181843 515864
rect 181791 515762 181843 515830
rect 181791 515728 181801 515762
rect 181835 515728 181843 515762
rect 181791 515702 181843 515728
rect 182081 515856 182133 515876
rect 182081 515822 182089 515856
rect 182123 515822 182133 515856
rect 182081 515775 182133 515822
rect 182081 515741 182089 515775
rect 182123 515741 182133 515775
rect 182081 515718 182133 515741
rect 182163 515856 182221 515876
rect 182163 515822 182175 515856
rect 182209 515822 182221 515856
rect 182163 515788 182221 515822
rect 182163 515754 182175 515788
rect 182209 515754 182221 515788
rect 182163 515718 182221 515754
rect 182251 515856 182303 515876
rect 182633 515864 182685 515876
rect 182251 515822 182261 515856
rect 182295 515822 182303 515856
rect 182251 515788 182303 515822
rect 182251 515754 182261 515788
rect 182295 515754 182303 515788
rect 182251 515718 182303 515754
rect 182633 515830 182641 515864
rect 182675 515830 182685 515864
rect 182633 515702 182685 515830
rect 183631 515864 183683 515876
rect 183631 515830 183641 515864
rect 183675 515830 183683 515864
rect 183631 515702 183683 515830
rect 183737 515864 183789 515876
rect 183737 515830 183745 515864
rect 183779 515830 183789 515864
rect 183737 515702 183789 515830
rect 184735 515864 184787 515876
rect 184735 515830 184745 515864
rect 184779 515830 184787 515864
rect 184735 515702 184787 515830
rect 184841 515864 184893 515876
rect 184841 515830 184849 515864
rect 184883 515830 184893 515864
rect 184841 515769 184893 515830
rect 184841 515735 184849 515769
rect 184883 515735 184893 515769
rect 184841 515702 184893 515735
rect 185011 515864 185063 515876
rect 185011 515830 185021 515864
rect 185055 515830 185063 515864
rect 185209 515864 185261 515876
rect 185011 515769 185063 515830
rect 185011 515735 185021 515769
rect 185055 515735 185063 515769
rect 185011 515702 185063 515735
rect 185209 515830 185217 515864
rect 185251 515830 185261 515864
rect 185209 515702 185261 515830
rect 186207 515864 186259 515876
rect 186207 515830 186217 515864
rect 186251 515830 186259 515864
rect 186207 515702 186259 515830
rect 186405 515856 186458 515876
rect 186405 515822 186413 515856
rect 186447 515822 186458 515856
rect 186405 515734 186458 515822
rect 186405 515700 186413 515734
rect 186447 515700 186458 515734
rect 186405 515676 186458 515700
rect 186488 515864 186554 515876
rect 186488 515830 186499 515864
rect 186533 515830 186554 515864
rect 186488 515796 186554 515830
rect 186488 515762 186499 515796
rect 186533 515762 186554 515796
rect 186488 515676 186554 515762
rect 186584 515829 186640 515876
rect 186584 515795 186595 515829
rect 186629 515795 186640 515829
rect 186584 515676 186640 515795
rect 186670 515864 186726 515876
rect 186670 515830 186681 515864
rect 186715 515830 186726 515864
rect 186670 515676 186726 515830
rect 186756 515856 186812 515876
rect 186756 515822 186767 515856
rect 186801 515822 186812 515856
rect 186756 515788 186812 515822
rect 186756 515754 186767 515788
rect 186801 515754 186812 515788
rect 186756 515720 186812 515754
rect 186756 515686 186767 515720
rect 186801 515686 186812 515720
rect 186756 515676 186812 515686
rect 186842 515850 186902 515876
rect 186842 515816 186853 515850
rect 186887 515816 186902 515850
rect 186842 515782 186902 515816
rect 186842 515748 186853 515782
rect 186887 515748 186902 515782
rect 186842 515676 186902 515748
rect 186957 515864 187009 515876
rect 186957 515830 186965 515864
rect 186999 515830 187009 515864
rect 186957 515769 187009 515830
rect 186957 515735 186965 515769
rect 186999 515735 187009 515769
rect 186957 515702 187009 515735
rect 187127 515864 187179 515876
rect 187127 515830 187137 515864
rect 187171 515830 187179 515864
rect 187127 515769 187179 515830
rect 187127 515735 187137 515769
rect 187171 515735 187179 515769
rect 187127 515702 187179 515735
rect 187233 515864 187285 515876
rect 187233 515830 187241 515864
rect 187275 515830 187285 515864
rect 187233 515769 187285 515830
rect 187233 515735 187241 515769
rect 187275 515735 187285 515769
rect 187233 515702 187285 515735
rect 187403 515864 187455 515876
rect 187403 515830 187413 515864
rect 187447 515830 187455 515864
rect 187403 515769 187455 515830
rect 187403 515735 187413 515769
rect 187447 515735 187455 515769
rect 187403 515702 187455 515735
<< ndiffc >>
rect 164686 540091 164720 541067
rect 164774 540091 164808 541067
rect 164889 540098 164923 541074
rect 164985 540098 165019 541074
rect 165081 540098 165115 541074
rect 165177 540098 165211 541074
rect 165273 540098 165307 541074
rect 165369 540098 165403 541074
rect 165465 540098 165499 541074
rect 165561 540098 165595 541074
rect 165657 540098 165691 541074
rect 165753 540098 165787 541074
rect 165849 540098 165883 541074
rect 165945 540098 165979 541074
rect 166041 540098 166075 541074
rect 166166 540091 166200 540267
rect 166254 540091 166288 540267
rect 166366 540091 166400 541067
rect 166454 540091 166488 541067
rect 168486 540091 168520 541067
rect 168574 540091 168608 541067
rect 168689 540098 168723 541074
rect 168785 540098 168819 541074
rect 168881 540098 168915 541074
rect 168977 540098 169011 541074
rect 169073 540098 169107 541074
rect 169169 540098 169203 541074
rect 169265 540098 169299 541074
rect 169361 540098 169395 541074
rect 169457 540098 169491 541074
rect 169553 540098 169587 541074
rect 169649 540098 169683 541074
rect 169745 540098 169779 541074
rect 169841 540098 169875 541074
rect 169966 540091 170000 540267
rect 170054 540091 170088 540267
rect 170166 540091 170200 541067
rect 170254 540091 170288 541067
rect 172186 540091 172220 541067
rect 172274 540091 172308 541067
rect 172389 540098 172423 541074
rect 172485 540098 172519 541074
rect 172581 540098 172615 541074
rect 172677 540098 172711 541074
rect 172773 540098 172807 541074
rect 172869 540098 172903 541074
rect 172965 540098 172999 541074
rect 173061 540098 173095 541074
rect 173157 540098 173191 541074
rect 173253 540098 173287 541074
rect 173349 540098 173383 541074
rect 173445 540098 173479 541074
rect 173541 540098 173575 541074
rect 173666 540091 173700 540267
rect 173754 540091 173788 540267
rect 173866 540091 173900 541067
rect 173954 540091 173988 541067
rect 175686 540091 175720 541067
rect 175774 540091 175808 541067
rect 175889 540098 175923 541074
rect 175985 540098 176019 541074
rect 176081 540098 176115 541074
rect 176177 540098 176211 541074
rect 176273 540098 176307 541074
rect 176369 540098 176403 541074
rect 176465 540098 176499 541074
rect 176561 540098 176595 541074
rect 176657 540098 176691 541074
rect 176753 540098 176787 541074
rect 176849 540098 176883 541074
rect 176945 540098 176979 541074
rect 177041 540098 177075 541074
rect 177166 540091 177200 540267
rect 177254 540091 177288 540267
rect 177366 540091 177400 541067
rect 177454 540091 177488 541067
rect 179286 540091 179320 541067
rect 179374 540091 179408 541067
rect 179489 540098 179523 541074
rect 179585 540098 179619 541074
rect 179681 540098 179715 541074
rect 179777 540098 179811 541074
rect 179873 540098 179907 541074
rect 179969 540098 180003 541074
rect 180065 540098 180099 541074
rect 180161 540098 180195 541074
rect 180257 540098 180291 541074
rect 180353 540098 180387 541074
rect 180449 540098 180483 541074
rect 180545 540098 180579 541074
rect 180641 540098 180675 541074
rect 180766 540091 180800 540267
rect 180854 540091 180888 540267
rect 180966 540091 181000 541067
rect 181054 540091 181088 541067
rect 182586 540091 182620 541067
rect 182674 540091 182708 541067
rect 182789 540098 182823 541074
rect 182885 540098 182919 541074
rect 182981 540098 183015 541074
rect 183077 540098 183111 541074
rect 183173 540098 183207 541074
rect 183269 540098 183303 541074
rect 183365 540098 183399 541074
rect 183461 540098 183495 541074
rect 183557 540098 183591 541074
rect 183653 540098 183687 541074
rect 183749 540098 183783 541074
rect 183845 540098 183879 541074
rect 183941 540098 183975 541074
rect 184066 540091 184100 540267
rect 184154 540091 184188 540267
rect 184266 540091 184300 541067
rect 184354 540091 184388 541067
rect 185886 540091 185920 541067
rect 185974 540091 186008 541067
rect 186089 540098 186123 541074
rect 186185 540098 186219 541074
rect 186281 540098 186315 541074
rect 186377 540098 186411 541074
rect 186473 540098 186507 541074
rect 186569 540098 186603 541074
rect 186665 540098 186699 541074
rect 186761 540098 186795 541074
rect 186857 540098 186891 541074
rect 186953 540098 186987 541074
rect 187049 540098 187083 541074
rect 187145 540098 187179 541074
rect 187241 540098 187275 541074
rect 187366 540091 187400 540267
rect 187454 540091 187488 540267
rect 187566 540091 187600 541067
rect 187654 540091 187688 541067
rect 189186 540091 189220 541067
rect 189274 540091 189308 541067
rect 189389 540098 189423 541074
rect 189485 540098 189519 541074
rect 189581 540098 189615 541074
rect 189677 540098 189711 541074
rect 189773 540098 189807 541074
rect 189869 540098 189903 541074
rect 189965 540098 189999 541074
rect 190061 540098 190095 541074
rect 190157 540098 190191 541074
rect 190253 540098 190287 541074
rect 190349 540098 190383 541074
rect 190445 540098 190479 541074
rect 190541 540098 190575 541074
rect 190666 540091 190700 540267
rect 190754 540091 190788 540267
rect 190866 540091 190900 541067
rect 190954 540091 190988 541067
rect 158666 538241 158700 538417
rect 158924 538241 158958 538417
rect 159042 538241 159076 538417
rect 159300 538241 159334 538417
rect 159558 538241 159592 538417
rect 159816 538241 159850 538417
rect 160074 538241 160108 538417
rect 160332 538241 160366 538417
rect 160590 538241 160624 538417
rect 160848 538241 160882 538417
rect 161106 538241 161140 538417
rect 161364 538241 161398 538417
rect 161486 538241 161520 538417
rect 161744 538241 161778 538417
rect 161886 538241 161920 538417
rect 162144 538241 162178 538417
rect 162266 538241 162300 538417
rect 162524 538241 162558 538417
rect 172245 530497 172279 530531
rect 172417 530497 172451 530531
rect 172528 530514 172562 530548
rect 172614 530492 172648 530526
rect 172700 530514 172734 530548
rect 172786 530492 172820 530526
rect 172883 530514 172917 530548
rect 172969 530510 173003 530544
rect 173073 530499 173107 530533
rect 174073 530499 174107 530533
rect 174177 530499 174211 530533
rect 174625 530499 174659 530533
rect 174920 530514 174954 530548
rect 175006 530492 175040 530526
rect 175092 530514 175126 530548
rect 175178 530492 175212 530526
rect 175275 530514 175309 530548
rect 175361 530510 175395 530544
rect 175557 530468 175591 530502
rect 175641 530518 175675 530552
rect 175765 530502 175799 530536
rect 175983 530522 176017 530556
rect 176195 530518 176229 530552
rect 176305 530522 176339 530556
rect 176417 530518 176451 530552
rect 176763 530516 176797 530550
rect 176870 530516 176904 530550
rect 177003 530522 177037 530556
rect 177125 530492 177159 530526
rect 177209 530518 177243 530552
rect 177293 530492 177327 530526
rect 177692 530492 177726 530526
rect 177782 530518 177816 530552
rect 177941 530492 177975 530526
rect 178045 530492 178079 530526
rect 178199 530518 178233 530552
rect 178283 530492 178317 530526
rect 178409 530488 178443 530522
rect 178495 530518 178529 530552
rect 178581 530505 178615 530539
rect 178692 530514 178726 530548
rect 178778 530492 178812 530526
rect 178864 530514 178898 530548
rect 178950 530492 178984 530526
rect 179047 530514 179081 530548
rect 179133 530510 179167 530544
rect 179237 530510 179271 530544
rect 179323 530514 179357 530548
rect 179420 530492 179454 530526
rect 179506 530514 179540 530548
rect 179592 530492 179626 530526
rect 179678 530514 179712 530548
rect 180249 530499 180283 530533
rect 180333 530518 180367 530552
rect 180540 530503 180574 530537
rect 180775 530503 180809 530537
rect 180843 530503 180877 530537
rect 180927 530503 180961 530537
rect 181215 530503 181249 530537
rect 181299 530503 181333 530537
rect 181367 530503 181401 530537
rect 181602 530503 181636 530537
rect 181809 530518 181843 530552
rect 181893 530499 181927 530533
rect 181997 530510 182031 530544
rect 182083 530514 182117 530548
rect 182180 530492 182214 530526
rect 182266 530514 182300 530548
rect 182352 530492 182386 530526
rect 182438 530514 182472 530548
rect 182641 530492 182675 530526
rect 182905 530492 182939 530526
rect 183101 530510 183135 530544
rect 183187 530514 183221 530548
rect 183284 530492 183318 530526
rect 183370 530514 183404 530548
rect 183456 530492 183490 530526
rect 183542 530514 183576 530548
rect 183653 530499 183687 530533
rect 184653 530499 184687 530533
rect 184757 530492 184791 530526
rect 185021 530492 185055 530526
rect 185217 530510 185251 530544
rect 185303 530514 185337 530548
rect 185400 530492 185434 530526
rect 185486 530514 185520 530548
rect 185572 530492 185606 530526
rect 185658 530514 185692 530548
rect 185769 530499 185803 530533
rect 186769 530499 186803 530533
rect 187241 530497 187275 530531
rect 187413 530497 187447 530531
rect 172245 529603 172279 529637
rect 172417 529603 172451 529637
rect 172521 529601 172555 529635
rect 173521 529601 173555 529635
rect 173625 529601 173659 529635
rect 174625 529601 174659 529635
rect 174843 529608 174877 529642
rect 174927 529582 174961 529616
rect 175081 529608 175115 529642
rect 175185 529608 175219 529642
rect 175344 529582 175378 529616
rect 175434 529608 175468 529642
rect 175557 529608 175591 529642
rect 175641 529582 175675 529616
rect 175725 529608 175759 529642
rect 175847 529578 175881 529612
rect 175980 529584 176014 529618
rect 176087 529584 176121 529618
rect 176433 529582 176467 529616
rect 176545 529578 176579 529612
rect 176655 529582 176689 529616
rect 176867 529578 176901 529612
rect 177085 529598 177119 529632
rect 177209 529582 177243 529616
rect 177293 529632 177327 529666
rect 177627 529597 177661 529631
rect 177711 529597 177745 529631
rect 177779 529597 177813 529631
rect 178014 529597 178048 529631
rect 178221 529582 178255 529616
rect 178305 529601 178339 529635
rect 178409 529632 178443 529666
rect 178493 529582 178527 529616
rect 178617 529598 178651 529632
rect 178835 529578 178869 529612
rect 179047 529582 179081 529616
rect 179157 529578 179191 529612
rect 179269 529582 179303 529616
rect 179615 529584 179649 529618
rect 179722 529584 179756 529618
rect 179855 529578 179889 529612
rect 179977 529608 180011 529642
rect 180061 529582 180095 529616
rect 180145 529608 180179 529642
rect 180249 529608 180283 529642
rect 180333 529582 180367 529616
rect 180417 529608 180451 529642
rect 180539 529578 180573 529612
rect 180672 529584 180706 529618
rect 180779 529584 180813 529618
rect 181125 529582 181159 529616
rect 181237 529578 181271 529612
rect 181347 529582 181381 529616
rect 181559 529578 181593 529612
rect 181777 529598 181811 529632
rect 181901 529582 181935 529616
rect 181985 529632 182019 529666
rect 182089 529608 182123 529642
rect 182353 529608 182387 529642
rect 182660 529608 182694 529642
rect 182750 529582 182784 529616
rect 182909 529608 182943 529642
rect 183013 529608 183047 529642
rect 183167 529582 183201 529616
rect 183251 529608 183285 529642
rect 183377 529601 183411 529635
rect 184377 529601 184411 529635
rect 184481 529601 184515 529635
rect 185481 529601 185515 529635
rect 185585 529601 185619 529635
rect 186585 529601 186619 529635
rect 186689 529601 186723 529635
rect 187137 529601 187171 529635
rect 187241 529603 187275 529637
rect 187413 529603 187447 529637
rect 172245 529409 172279 529443
rect 172417 529409 172451 529443
rect 172521 529411 172555 529445
rect 173521 529411 173555 529445
rect 173625 529411 173659 529445
rect 174625 529411 174659 529445
rect 175143 529415 175177 529449
rect 175227 529415 175261 529449
rect 175295 529415 175329 529449
rect 175530 529415 175564 529449
rect 175737 529430 175771 529464
rect 175821 529411 175855 529445
rect 175942 529426 175976 529460
rect 176028 529417 176062 529451
rect 176114 529426 176148 529460
rect 176200 529417 176234 529451
rect 176286 529426 176320 529460
rect 176372 529417 176406 529451
rect 176458 529426 176492 529460
rect 176544 529417 176578 529451
rect 176629 529426 176663 529460
rect 176715 529417 176749 529451
rect 176801 529426 176835 529460
rect 176887 529417 176921 529451
rect 176973 529426 177007 529460
rect 177059 529417 177093 529451
rect 177145 529426 177179 529460
rect 177231 529417 177265 529451
rect 177317 529417 177351 529451
rect 177403 529417 177437 529451
rect 177489 529417 177523 529451
rect 177575 529417 177609 529451
rect 177661 529430 177695 529464
rect 177765 529404 177799 529438
rect 177849 529430 177883 529464
rect 177933 529404 177967 529438
rect 178055 529434 178089 529468
rect 178188 529428 178222 529462
rect 178295 529428 178329 529462
rect 178641 529430 178675 529464
rect 178753 529434 178787 529468
rect 178863 529430 178897 529464
rect 179075 529434 179109 529468
rect 179293 529414 179327 529448
rect 179417 529430 179451 529464
rect 179501 529380 179535 529414
rect 179697 529417 179731 529451
rect 179783 529430 179817 529464
rect 179869 529400 179903 529434
rect 180065 529411 180099 529445
rect 180513 529411 180547 529445
rect 180709 529430 180743 529464
rect 180795 529417 180829 529451
rect 180881 529417 180915 529451
rect 180967 529417 181001 529451
rect 181053 529417 181087 529451
rect 181139 529417 181173 529451
rect 181225 529426 181259 529460
rect 181311 529417 181345 529451
rect 181397 529426 181431 529460
rect 181483 529417 181517 529451
rect 181569 529426 181603 529460
rect 181655 529417 181689 529451
rect 181741 529426 181775 529460
rect 181826 529417 181860 529451
rect 181912 529426 181946 529460
rect 181998 529417 182032 529451
rect 182084 529426 182118 529460
rect 182170 529417 182204 529451
rect 182256 529426 182290 529460
rect 182342 529417 182376 529451
rect 182428 529426 182462 529460
rect 182549 529400 182583 529434
rect 182635 529430 182669 529464
rect 182721 529417 182755 529451
rect 182825 529411 182859 529445
rect 183825 529411 183859 529445
rect 183929 529411 183963 529445
rect 184929 529411 184963 529445
rect 185217 529411 185251 529445
rect 186217 529411 186251 529445
rect 186321 529411 186355 529445
rect 186953 529411 186987 529445
rect 187241 529409 187275 529443
rect 187413 529409 187447 529443
rect 172245 528515 172279 528549
rect 172417 528515 172451 528549
rect 172521 528513 172555 528547
rect 173521 528513 173555 528547
rect 173625 528513 173659 528547
rect 174625 528513 174659 528547
rect 174729 528513 174763 528547
rect 175729 528513 175763 528547
rect 175925 528507 175959 528541
rect 176011 528494 176045 528528
rect 176097 528524 176131 528558
rect 176201 528507 176235 528541
rect 176287 528494 176321 528528
rect 176373 528524 176407 528558
rect 176523 528509 176557 528543
rect 176607 528509 176641 528543
rect 176675 528509 176709 528543
rect 176910 528509 176944 528543
rect 177117 528494 177151 528528
rect 177201 528513 177235 528547
rect 177508 528520 177542 528554
rect 177598 528494 177632 528528
rect 177757 528520 177791 528554
rect 177861 528520 177895 528554
rect 178015 528494 178049 528528
rect 178099 528520 178133 528554
rect 178409 528494 178443 528528
rect 178495 528507 178529 528541
rect 178581 528507 178615 528541
rect 178667 528507 178701 528541
rect 178753 528507 178787 528541
rect 178839 528507 178873 528541
rect 178925 528498 178959 528532
rect 179011 528507 179045 528541
rect 179097 528498 179131 528532
rect 179183 528507 179217 528541
rect 179269 528498 179303 528532
rect 179355 528507 179389 528541
rect 179441 528498 179475 528532
rect 179526 528507 179560 528541
rect 179612 528498 179646 528532
rect 179698 528507 179732 528541
rect 179784 528498 179818 528532
rect 179870 528507 179904 528541
rect 179956 528498 179990 528532
rect 180042 528507 180076 528541
rect 180128 528498 180162 528532
rect 180249 528507 180283 528541
rect 180335 528494 180369 528528
rect 180421 528524 180455 528558
rect 180525 528520 180559 528554
rect 180609 528494 180643 528528
rect 180693 528520 180727 528554
rect 180815 528490 180849 528524
rect 180948 528496 180982 528530
rect 181055 528496 181089 528530
rect 181401 528494 181435 528528
rect 181513 528490 181547 528524
rect 181623 528494 181657 528528
rect 181835 528490 181869 528524
rect 182053 528510 182087 528544
rect 182177 528494 182211 528528
rect 182261 528544 182295 528578
rect 182641 528513 182675 528547
rect 183641 528513 183675 528547
rect 183745 528513 183779 528547
rect 184745 528513 184779 528547
rect 184849 528513 184883 528547
rect 185849 528513 185883 528547
rect 185953 528513 185987 528547
rect 186953 528513 186987 528547
rect 187241 528515 187275 528549
rect 187413 528515 187447 528549
rect 172245 528321 172279 528355
rect 172417 528321 172451 528355
rect 172521 528323 172555 528357
rect 173521 528323 173555 528357
rect 173625 528323 173659 528357
rect 174625 528323 174659 528357
rect 174913 528323 174947 528357
rect 175913 528323 175947 528357
rect 176109 528316 176143 528350
rect 176193 528342 176227 528376
rect 176277 528316 176311 528350
rect 176399 528346 176433 528380
rect 176532 528340 176566 528374
rect 176639 528340 176673 528374
rect 176985 528342 177019 528376
rect 177097 528346 177131 528380
rect 177207 528342 177241 528376
rect 177419 528346 177453 528380
rect 177637 528326 177671 528360
rect 177761 528342 177795 528376
rect 177845 528292 177879 528326
rect 177949 528312 177983 528346
rect 178035 528342 178069 528376
rect 178121 528329 178155 528363
rect 178225 528323 178259 528357
rect 178857 528323 178891 528357
rect 178961 528323 178995 528357
rect 179045 528342 179079 528376
rect 179252 528327 179286 528361
rect 179487 528327 179521 528361
rect 179555 528327 179589 528361
rect 179639 528327 179673 528361
rect 180065 528323 180099 528357
rect 180697 528323 180731 528357
rect 180985 528323 181019 528357
rect 181069 528342 181103 528376
rect 181276 528327 181310 528361
rect 181511 528327 181545 528361
rect 181579 528327 181613 528361
rect 181663 528327 181697 528361
rect 181813 528323 181847 528357
rect 182813 528323 182847 528357
rect 182917 528323 182951 528357
rect 183917 528323 183951 528357
rect 184021 528323 184055 528357
rect 185021 528323 185055 528357
rect 185217 528323 185251 528357
rect 186217 528323 186251 528357
rect 186321 528323 186355 528357
rect 186953 528323 186987 528357
rect 187241 528321 187275 528355
rect 187413 528321 187447 528355
rect 172245 527427 172279 527461
rect 172417 527427 172451 527461
rect 172521 527425 172555 527459
rect 173521 527425 173555 527459
rect 173625 527425 173659 527459
rect 174625 527425 174659 527459
rect 174729 527425 174763 527459
rect 175729 527425 175763 527459
rect 175833 527425 175867 527459
rect 176281 527425 176315 527459
rect 176404 527432 176438 527466
rect 176494 527406 176528 527440
rect 176653 527432 176687 527466
rect 176757 527432 176791 527466
rect 176911 527406 176945 527440
rect 176995 527432 177029 527466
rect 177121 527427 177155 527461
rect 177293 527427 177327 527461
rect 177489 527425 177523 527459
rect 178489 527425 178523 527459
rect 178593 527432 178627 527466
rect 178857 527432 178891 527466
rect 178980 527432 179014 527466
rect 179070 527406 179104 527440
rect 179229 527432 179263 527466
rect 179333 527432 179367 527466
rect 179487 527406 179521 527440
rect 179571 527432 179605 527466
rect 179697 527425 179731 527459
rect 180697 527425 180731 527459
rect 180801 527425 180835 527459
rect 181801 527425 181835 527459
rect 181905 527425 181939 527459
rect 182353 527425 182387 527459
rect 182641 527425 182675 527459
rect 183641 527425 183675 527459
rect 183745 527425 183779 527459
rect 184745 527425 184779 527459
rect 184849 527425 184883 527459
rect 185849 527425 185883 527459
rect 185953 527425 185987 527459
rect 186953 527425 186987 527459
rect 187241 527427 187275 527461
rect 187413 527427 187447 527461
rect 172245 527233 172279 527267
rect 172417 527233 172451 527267
rect 172521 527235 172555 527269
rect 173521 527235 173555 527269
rect 173625 527235 173659 527269
rect 174625 527235 174659 527269
rect 174913 527235 174947 527269
rect 175913 527235 175947 527269
rect 176017 527235 176051 527269
rect 177017 527235 177051 527269
rect 177121 527235 177155 527269
rect 178121 527235 178155 527269
rect 178225 527235 178259 527269
rect 179225 527235 179259 527269
rect 179329 527235 179363 527269
rect 179777 527235 179811 527269
rect 180065 527235 180099 527269
rect 181065 527235 181099 527269
rect 181169 527235 181203 527269
rect 182169 527235 182203 527269
rect 182273 527235 182307 527269
rect 183273 527235 183307 527269
rect 183377 527235 183411 527269
rect 184377 527235 184411 527269
rect 184481 527235 184515 527269
rect 184929 527235 184963 527269
rect 185217 527235 185251 527269
rect 186217 527235 186251 527269
rect 186321 527235 186355 527269
rect 186953 527235 186987 527269
rect 187241 527233 187275 527267
rect 187413 527233 187447 527267
rect 172245 526339 172279 526373
rect 172417 526339 172451 526373
rect 172521 526337 172555 526371
rect 173521 526337 173555 526371
rect 173625 526337 173659 526371
rect 174625 526337 174659 526371
rect 174729 526337 174763 526371
rect 175729 526337 175763 526371
rect 175833 526337 175867 526371
rect 176833 526337 176867 526371
rect 176937 526344 176971 526378
rect 177201 526344 177235 526378
rect 177489 526337 177523 526371
rect 178489 526337 178523 526371
rect 178593 526337 178627 526371
rect 179593 526337 179627 526371
rect 179697 526337 179731 526371
rect 180697 526337 180731 526371
rect 180801 526337 180835 526371
rect 181801 526337 181835 526371
rect 181905 526337 181939 526371
rect 182353 526337 182387 526371
rect 182641 526337 182675 526371
rect 183641 526337 183675 526371
rect 183745 526337 183779 526371
rect 184745 526337 184779 526371
rect 184849 526337 184883 526371
rect 185849 526337 185883 526371
rect 185953 526337 185987 526371
rect 186953 526337 186987 526371
rect 187241 526339 187275 526373
rect 187413 526339 187447 526373
rect 172245 526145 172279 526179
rect 172417 526145 172451 526179
rect 172521 526147 172555 526181
rect 173521 526147 173555 526181
rect 173625 526147 173659 526181
rect 174625 526147 174659 526181
rect 174913 526147 174947 526181
rect 175913 526147 175947 526181
rect 176017 526147 176051 526181
rect 177017 526147 177051 526181
rect 177121 526147 177155 526181
rect 178121 526147 178155 526181
rect 178225 526147 178259 526181
rect 179225 526147 179259 526181
rect 179329 526147 179363 526181
rect 179777 526147 179811 526181
rect 180065 526147 180099 526181
rect 181065 526147 181099 526181
rect 181169 526147 181203 526181
rect 182169 526147 182203 526181
rect 182273 526147 182307 526181
rect 183273 526147 183307 526181
rect 183377 526147 183411 526181
rect 184377 526147 184411 526181
rect 184481 526147 184515 526181
rect 184929 526147 184963 526181
rect 185217 526147 185251 526181
rect 186217 526147 186251 526181
rect 186321 526147 186355 526181
rect 186953 526147 186987 526181
rect 187241 526145 187275 526179
rect 187413 526145 187447 526179
rect 172245 525251 172279 525285
rect 172417 525251 172451 525285
rect 172521 525249 172555 525283
rect 173521 525249 173555 525283
rect 173625 525249 173659 525283
rect 174625 525249 174659 525283
rect 174729 525249 174763 525283
rect 175729 525249 175763 525283
rect 175833 525249 175867 525283
rect 176833 525249 176867 525283
rect 176937 525256 176971 525290
rect 177201 525256 177235 525290
rect 177489 525249 177523 525283
rect 178489 525249 178523 525283
rect 178593 525249 178627 525283
rect 179593 525249 179627 525283
rect 179697 525249 179731 525283
rect 180697 525249 180731 525283
rect 180801 525249 180835 525283
rect 181801 525249 181835 525283
rect 181905 525249 181939 525283
rect 182353 525249 182387 525283
rect 182641 525249 182675 525283
rect 183641 525249 183675 525283
rect 183745 525249 183779 525283
rect 184745 525249 184779 525283
rect 184849 525249 184883 525283
rect 185849 525249 185883 525283
rect 185953 525249 185987 525283
rect 186953 525249 186987 525283
rect 187241 525251 187275 525285
rect 187413 525251 187447 525285
rect 172245 525057 172279 525091
rect 172417 525057 172451 525091
rect 172521 525059 172555 525093
rect 173521 525059 173555 525093
rect 173625 525059 173659 525093
rect 174625 525059 174659 525093
rect 174913 525059 174947 525093
rect 175913 525059 175947 525093
rect 176017 525059 176051 525093
rect 177017 525059 177051 525093
rect 177121 525059 177155 525093
rect 178121 525059 178155 525093
rect 178225 525059 178259 525093
rect 179225 525059 179259 525093
rect 179329 525059 179363 525093
rect 179777 525059 179811 525093
rect 180065 525059 180099 525093
rect 181065 525059 181099 525093
rect 181169 525059 181203 525093
rect 182169 525059 182203 525093
rect 182273 525059 182307 525093
rect 183273 525059 183307 525093
rect 183377 525059 183411 525093
rect 184377 525059 184411 525093
rect 184481 525059 184515 525093
rect 184929 525059 184963 525093
rect 185217 525059 185251 525093
rect 186217 525059 186251 525093
rect 186321 525059 186355 525093
rect 186953 525059 186987 525093
rect 187241 525057 187275 525091
rect 187413 525057 187447 525091
rect 172245 524163 172279 524197
rect 172417 524163 172451 524197
rect 172521 524161 172555 524195
rect 173521 524161 173555 524195
rect 173625 524161 173659 524195
rect 174625 524161 174659 524195
rect 174729 524161 174763 524195
rect 175729 524161 175763 524195
rect 175833 524161 175867 524195
rect 176833 524161 176867 524195
rect 176937 524168 176971 524202
rect 177201 524168 177235 524202
rect 177489 524161 177523 524195
rect 178489 524161 178523 524195
rect 178593 524161 178627 524195
rect 179593 524161 179627 524195
rect 179697 524161 179731 524195
rect 180697 524161 180731 524195
rect 180801 524161 180835 524195
rect 181801 524161 181835 524195
rect 181905 524161 181939 524195
rect 182353 524161 182387 524195
rect 182641 524161 182675 524195
rect 183641 524161 183675 524195
rect 183745 524161 183779 524195
rect 184745 524161 184779 524195
rect 184849 524161 184883 524195
rect 185849 524161 185883 524195
rect 185953 524161 185987 524195
rect 186953 524161 186987 524195
rect 187241 524163 187275 524197
rect 187413 524163 187447 524197
rect 172245 523969 172279 524003
rect 172417 523969 172451 524003
rect 172521 523971 172555 524005
rect 173521 523971 173555 524005
rect 173625 523971 173659 524005
rect 174625 523971 174659 524005
rect 174913 523971 174947 524005
rect 175913 523971 175947 524005
rect 176017 523971 176051 524005
rect 177017 523971 177051 524005
rect 177121 523971 177155 524005
rect 178121 523971 178155 524005
rect 178225 523971 178259 524005
rect 179225 523971 179259 524005
rect 179329 523971 179363 524005
rect 179777 523971 179811 524005
rect 180065 523971 180099 524005
rect 181065 523971 181099 524005
rect 181169 523971 181203 524005
rect 182169 523971 182203 524005
rect 182273 523971 182307 524005
rect 183273 523971 183307 524005
rect 183377 523971 183411 524005
rect 184377 523971 184411 524005
rect 184481 523971 184515 524005
rect 184929 523971 184963 524005
rect 185217 523971 185251 524005
rect 186217 523971 186251 524005
rect 186321 523971 186355 524005
rect 186953 523971 186987 524005
rect 187241 523969 187275 524003
rect 187413 523969 187447 524003
rect 172245 523075 172279 523109
rect 172417 523075 172451 523109
rect 172521 523073 172555 523107
rect 173521 523073 173555 523107
rect 173625 523073 173659 523107
rect 174625 523073 174659 523107
rect 174729 523073 174763 523107
rect 175729 523073 175763 523107
rect 175833 523073 175867 523107
rect 176833 523073 176867 523107
rect 176937 523080 176971 523114
rect 177201 523080 177235 523114
rect 177489 523073 177523 523107
rect 178489 523073 178523 523107
rect 178593 523073 178627 523107
rect 179593 523073 179627 523107
rect 179697 523073 179731 523107
rect 180697 523073 180731 523107
rect 180801 523073 180835 523107
rect 181801 523073 181835 523107
rect 181905 523073 181939 523107
rect 182353 523073 182387 523107
rect 182641 523073 182675 523107
rect 183641 523073 183675 523107
rect 183745 523073 183779 523107
rect 184745 523073 184779 523107
rect 184849 523073 184883 523107
rect 185849 523073 185883 523107
rect 185953 523073 185987 523107
rect 186953 523073 186987 523107
rect 187241 523075 187275 523109
rect 187413 523075 187447 523109
rect 172245 522881 172279 522915
rect 172417 522881 172451 522915
rect 172521 522883 172555 522917
rect 173521 522883 173555 522917
rect 173625 522883 173659 522917
rect 174625 522883 174659 522917
rect 174913 522883 174947 522917
rect 175913 522883 175947 522917
rect 176017 522883 176051 522917
rect 177017 522883 177051 522917
rect 177121 522883 177155 522917
rect 178121 522883 178155 522917
rect 178225 522883 178259 522917
rect 179225 522883 179259 522917
rect 179329 522883 179363 522917
rect 179777 522883 179811 522917
rect 180065 522883 180099 522917
rect 181065 522883 181099 522917
rect 181169 522883 181203 522917
rect 182169 522883 182203 522917
rect 182273 522883 182307 522917
rect 183273 522883 183307 522917
rect 183377 522883 183411 522917
rect 184377 522883 184411 522917
rect 184481 522883 184515 522917
rect 184929 522883 184963 522917
rect 185217 522883 185251 522917
rect 186217 522883 186251 522917
rect 186321 522883 186355 522917
rect 186953 522883 186987 522917
rect 187241 522881 187275 522915
rect 187413 522881 187447 522915
rect 172245 521987 172279 522021
rect 172417 521987 172451 522021
rect 172521 521985 172555 522019
rect 173521 521985 173555 522019
rect 173625 521985 173659 522019
rect 174625 521985 174659 522019
rect 174729 521985 174763 522019
rect 175729 521985 175763 522019
rect 175833 521985 175867 522019
rect 176833 521985 176867 522019
rect 176937 521992 176971 522026
rect 177201 521992 177235 522026
rect 177489 521985 177523 522019
rect 178489 521985 178523 522019
rect 178593 521985 178627 522019
rect 179593 521985 179627 522019
rect 179697 521985 179731 522019
rect 180697 521985 180731 522019
rect 180801 521985 180835 522019
rect 181801 521985 181835 522019
rect 181905 521985 181939 522019
rect 182353 521985 182387 522019
rect 182641 521985 182675 522019
rect 183641 521985 183675 522019
rect 183745 521985 183779 522019
rect 184745 521985 184779 522019
rect 184849 521985 184883 522019
rect 185849 521985 185883 522019
rect 185953 521985 185987 522019
rect 186953 521985 186987 522019
rect 187241 521987 187275 522021
rect 187413 521987 187447 522021
rect 172245 521793 172279 521827
rect 172417 521793 172451 521827
rect 172521 521795 172555 521829
rect 173521 521795 173555 521829
rect 173625 521795 173659 521829
rect 174625 521795 174659 521829
rect 174913 521795 174947 521829
rect 175913 521795 175947 521829
rect 176017 521795 176051 521829
rect 177017 521795 177051 521829
rect 177121 521795 177155 521829
rect 178121 521795 178155 521829
rect 178225 521795 178259 521829
rect 179225 521795 179259 521829
rect 179329 521795 179363 521829
rect 179777 521795 179811 521829
rect 180065 521795 180099 521829
rect 181065 521795 181099 521829
rect 181169 521795 181203 521829
rect 182169 521795 182203 521829
rect 182273 521795 182307 521829
rect 183273 521795 183307 521829
rect 183377 521795 183411 521829
rect 184377 521795 184411 521829
rect 184481 521795 184515 521829
rect 184929 521795 184963 521829
rect 185217 521795 185251 521829
rect 186217 521795 186251 521829
rect 186321 521795 186355 521829
rect 186953 521795 186987 521829
rect 187241 521793 187275 521827
rect 187413 521793 187447 521827
rect 172245 520899 172279 520933
rect 172417 520899 172451 520933
rect 172521 520897 172555 520931
rect 173521 520897 173555 520931
rect 173625 520897 173659 520931
rect 174625 520897 174659 520931
rect 174729 520897 174763 520931
rect 175729 520897 175763 520931
rect 175833 520897 175867 520931
rect 176833 520897 176867 520931
rect 176937 520904 176971 520938
rect 177201 520904 177235 520938
rect 177489 520897 177523 520931
rect 178489 520897 178523 520931
rect 178593 520897 178627 520931
rect 179593 520897 179627 520931
rect 179697 520897 179731 520931
rect 180697 520897 180731 520931
rect 180801 520897 180835 520931
rect 181801 520897 181835 520931
rect 181905 520897 181939 520931
rect 182353 520897 182387 520931
rect 182641 520897 182675 520931
rect 183641 520897 183675 520931
rect 183745 520897 183779 520931
rect 184745 520897 184779 520931
rect 184849 520897 184883 520931
rect 185849 520897 185883 520931
rect 185953 520897 185987 520931
rect 186953 520897 186987 520931
rect 187241 520899 187275 520933
rect 187413 520899 187447 520933
rect 172245 520705 172279 520739
rect 172417 520705 172451 520739
rect 172521 520707 172555 520741
rect 173521 520707 173555 520741
rect 173625 520707 173659 520741
rect 174625 520707 174659 520741
rect 174913 520707 174947 520741
rect 175913 520707 175947 520741
rect 176017 520707 176051 520741
rect 177017 520707 177051 520741
rect 177121 520707 177155 520741
rect 178121 520707 178155 520741
rect 178225 520707 178259 520741
rect 179225 520707 179259 520741
rect 179329 520707 179363 520741
rect 179777 520707 179811 520741
rect 180065 520707 180099 520741
rect 181065 520707 181099 520741
rect 181169 520707 181203 520741
rect 182169 520707 182203 520741
rect 182273 520707 182307 520741
rect 183273 520707 183307 520741
rect 183377 520707 183411 520741
rect 184377 520707 184411 520741
rect 184481 520707 184515 520741
rect 184929 520707 184963 520741
rect 185217 520707 185251 520741
rect 186217 520707 186251 520741
rect 186321 520707 186355 520741
rect 186953 520707 186987 520741
rect 187241 520705 187275 520739
rect 187413 520705 187447 520739
rect 172245 519811 172279 519845
rect 172417 519811 172451 519845
rect 172521 519809 172555 519843
rect 173521 519809 173555 519843
rect 173625 519809 173659 519843
rect 174625 519809 174659 519843
rect 174729 519809 174763 519843
rect 175729 519809 175763 519843
rect 175833 519809 175867 519843
rect 176833 519809 176867 519843
rect 176937 519816 176971 519850
rect 177201 519816 177235 519850
rect 177489 519809 177523 519843
rect 178489 519809 178523 519843
rect 178593 519809 178627 519843
rect 179593 519809 179627 519843
rect 179697 519809 179731 519843
rect 180697 519809 180731 519843
rect 180801 519809 180835 519843
rect 181801 519809 181835 519843
rect 181905 519809 181939 519843
rect 182353 519809 182387 519843
rect 182641 519809 182675 519843
rect 183641 519809 183675 519843
rect 183745 519809 183779 519843
rect 184745 519809 184779 519843
rect 184849 519809 184883 519843
rect 185849 519809 185883 519843
rect 185953 519809 185987 519843
rect 186953 519809 186987 519843
rect 187241 519811 187275 519845
rect 187413 519811 187447 519845
rect 172245 519617 172279 519651
rect 172417 519617 172451 519651
rect 172521 519619 172555 519653
rect 173521 519619 173555 519653
rect 173625 519619 173659 519653
rect 174625 519619 174659 519653
rect 174913 519619 174947 519653
rect 175913 519619 175947 519653
rect 176017 519619 176051 519653
rect 177017 519619 177051 519653
rect 177121 519619 177155 519653
rect 178121 519619 178155 519653
rect 178225 519619 178259 519653
rect 179225 519619 179259 519653
rect 179329 519619 179363 519653
rect 179777 519619 179811 519653
rect 180065 519619 180099 519653
rect 181065 519619 181099 519653
rect 181169 519619 181203 519653
rect 182169 519619 182203 519653
rect 182273 519619 182307 519653
rect 183273 519619 183307 519653
rect 183377 519619 183411 519653
rect 184377 519619 184411 519653
rect 184481 519619 184515 519653
rect 184929 519619 184963 519653
rect 185217 519619 185251 519653
rect 186217 519619 186251 519653
rect 186321 519619 186355 519653
rect 186953 519619 186987 519653
rect 187241 519617 187275 519651
rect 187413 519617 187447 519651
rect 172245 518723 172279 518757
rect 172417 518723 172451 518757
rect 172521 518721 172555 518755
rect 173521 518721 173555 518755
rect 173625 518721 173659 518755
rect 174625 518721 174659 518755
rect 174729 518721 174763 518755
rect 175729 518721 175763 518755
rect 175833 518721 175867 518755
rect 176833 518721 176867 518755
rect 176937 518728 176971 518762
rect 177201 518728 177235 518762
rect 177489 518721 177523 518755
rect 178489 518721 178523 518755
rect 178593 518721 178627 518755
rect 179593 518721 179627 518755
rect 179697 518721 179731 518755
rect 180697 518721 180731 518755
rect 180801 518721 180835 518755
rect 181801 518721 181835 518755
rect 181905 518721 181939 518755
rect 182353 518721 182387 518755
rect 182641 518721 182675 518755
rect 183641 518721 183675 518755
rect 183745 518721 183779 518755
rect 184745 518721 184779 518755
rect 184849 518721 184883 518755
rect 185849 518721 185883 518755
rect 185953 518721 185987 518755
rect 186953 518721 186987 518755
rect 187241 518723 187275 518757
rect 187413 518723 187447 518757
rect 172245 518529 172279 518563
rect 172417 518529 172451 518563
rect 172521 518531 172555 518565
rect 173521 518531 173555 518565
rect 173625 518531 173659 518565
rect 174625 518531 174659 518565
rect 174913 518531 174947 518565
rect 175913 518531 175947 518565
rect 176017 518531 176051 518565
rect 177017 518531 177051 518565
rect 177121 518531 177155 518565
rect 178121 518531 178155 518565
rect 178225 518531 178259 518565
rect 179225 518531 179259 518565
rect 179329 518531 179363 518565
rect 179777 518531 179811 518565
rect 180065 518531 180099 518565
rect 181065 518531 181099 518565
rect 181169 518531 181203 518565
rect 182169 518531 182203 518565
rect 182273 518531 182307 518565
rect 183273 518531 183307 518565
rect 183377 518531 183411 518565
rect 184377 518531 184411 518565
rect 184481 518531 184515 518565
rect 184929 518531 184963 518565
rect 185217 518531 185251 518565
rect 186217 518531 186251 518565
rect 186321 518531 186355 518565
rect 186953 518531 186987 518565
rect 187241 518529 187275 518563
rect 187413 518529 187447 518563
rect 172245 517635 172279 517669
rect 172417 517635 172451 517669
rect 172521 517633 172555 517667
rect 173521 517633 173555 517667
rect 173625 517633 173659 517667
rect 174625 517633 174659 517667
rect 174729 517633 174763 517667
rect 175729 517633 175763 517667
rect 175833 517633 175867 517667
rect 176833 517633 176867 517667
rect 176937 517640 176971 517674
rect 177201 517640 177235 517674
rect 177489 517633 177523 517667
rect 178489 517633 178523 517667
rect 178593 517633 178627 517667
rect 179593 517633 179627 517667
rect 179697 517633 179731 517667
rect 180697 517633 180731 517667
rect 180801 517633 180835 517667
rect 181801 517633 181835 517667
rect 181905 517633 181939 517667
rect 182353 517633 182387 517667
rect 182641 517633 182675 517667
rect 183641 517633 183675 517667
rect 183745 517633 183779 517667
rect 184745 517633 184779 517667
rect 184849 517633 184883 517667
rect 185849 517633 185883 517667
rect 185953 517633 185987 517667
rect 186953 517633 186987 517667
rect 187241 517635 187275 517669
rect 187413 517635 187447 517669
rect 172245 517441 172279 517475
rect 172417 517441 172451 517475
rect 172521 517443 172555 517477
rect 173521 517443 173555 517477
rect 173625 517443 173659 517477
rect 174625 517443 174659 517477
rect 174913 517443 174947 517477
rect 175913 517443 175947 517477
rect 176017 517443 176051 517477
rect 177017 517443 177051 517477
rect 177121 517443 177155 517477
rect 178121 517443 178155 517477
rect 178225 517443 178259 517477
rect 179225 517443 179259 517477
rect 179329 517443 179363 517477
rect 179777 517443 179811 517477
rect 180065 517443 180099 517477
rect 181065 517443 181099 517477
rect 181169 517443 181203 517477
rect 182169 517443 182203 517477
rect 182273 517443 182307 517477
rect 183273 517443 183307 517477
rect 183377 517443 183411 517477
rect 184377 517443 184411 517477
rect 184481 517443 184515 517477
rect 184929 517443 184963 517477
rect 185217 517443 185251 517477
rect 186217 517443 186251 517477
rect 186321 517443 186355 517477
rect 186953 517443 186987 517477
rect 187241 517441 187275 517475
rect 187413 517441 187447 517475
rect 172245 516547 172279 516581
rect 172417 516547 172451 516581
rect 172521 516545 172555 516579
rect 173521 516545 173555 516579
rect 173625 516545 173659 516579
rect 174625 516545 174659 516579
rect 174729 516545 174763 516579
rect 175729 516545 175763 516579
rect 175833 516545 175867 516579
rect 176833 516545 176867 516579
rect 176937 516552 176971 516586
rect 177201 516552 177235 516586
rect 177489 516545 177523 516579
rect 178489 516545 178523 516579
rect 178593 516545 178627 516579
rect 179593 516545 179627 516579
rect 179697 516545 179731 516579
rect 180697 516545 180731 516579
rect 180801 516545 180835 516579
rect 181801 516545 181835 516579
rect 181905 516545 181939 516579
rect 182353 516545 182387 516579
rect 182641 516545 182675 516579
rect 183641 516545 183675 516579
rect 183745 516545 183779 516579
rect 184745 516545 184779 516579
rect 184849 516545 184883 516579
rect 185849 516545 185883 516579
rect 185953 516545 185987 516579
rect 186953 516545 186987 516579
rect 187241 516547 187275 516581
rect 187413 516547 187447 516581
rect 172245 516353 172279 516387
rect 172417 516353 172451 516387
rect 172521 516355 172555 516389
rect 173521 516355 173555 516389
rect 173625 516355 173659 516389
rect 174625 516355 174659 516389
rect 174913 516355 174947 516389
rect 175913 516355 175947 516389
rect 176017 516355 176051 516389
rect 177017 516355 177051 516389
rect 177121 516355 177155 516389
rect 178121 516355 178155 516389
rect 178225 516355 178259 516389
rect 179225 516355 179259 516389
rect 179329 516355 179363 516389
rect 179777 516355 179811 516389
rect 180065 516355 180099 516389
rect 181065 516355 181099 516389
rect 181169 516355 181203 516389
rect 182169 516355 182203 516389
rect 182273 516355 182307 516389
rect 183273 516355 183307 516389
rect 183377 516355 183411 516389
rect 184377 516355 184411 516389
rect 184481 516355 184515 516389
rect 184929 516355 184963 516389
rect 185217 516355 185251 516389
rect 186217 516355 186251 516389
rect 186321 516355 186355 516389
rect 186953 516355 186987 516389
rect 187241 516353 187275 516387
rect 187413 516353 187447 516387
rect 172245 515459 172279 515493
rect 172417 515459 172451 515493
rect 172521 515457 172555 515491
rect 173153 515457 173187 515491
rect 173441 515446 173475 515480
rect 173527 515442 173561 515476
rect 173624 515464 173658 515498
rect 173710 515442 173744 515476
rect 173796 515464 173830 515498
rect 173882 515442 173916 515476
rect 173993 515457 174027 515491
rect 174625 515457 174659 515491
rect 174913 515457 174947 515491
rect 175913 515457 175947 515491
rect 176017 515457 176051 515491
rect 177017 515457 177051 515491
rect 177121 515459 177155 515493
rect 177293 515459 177327 515493
rect 177489 515457 177523 515491
rect 178489 515457 178523 515491
rect 178593 515457 178627 515491
rect 179593 515457 179627 515491
rect 179697 515459 179731 515493
rect 179869 515459 179903 515493
rect 180065 515457 180099 515491
rect 181065 515457 181099 515491
rect 181169 515457 181203 515491
rect 181801 515457 181835 515491
rect 182089 515468 182123 515502
rect 182175 515438 182209 515472
rect 182261 515451 182295 515485
rect 182641 515457 182675 515491
rect 183641 515457 183675 515491
rect 183745 515457 183779 515491
rect 184745 515457 184779 515491
rect 184849 515459 184883 515493
rect 185021 515459 185055 515493
rect 185217 515457 185251 515491
rect 186217 515457 186251 515491
rect 186413 515446 186447 515480
rect 186499 515442 186533 515476
rect 186596 515464 186630 515498
rect 186682 515442 186716 515476
rect 186768 515464 186802 515498
rect 186854 515442 186888 515476
rect 186965 515459 186999 515493
rect 187137 515459 187171 515493
rect 187241 515459 187275 515493
rect 187413 515459 187447 515493
<< pdiffc >>
rect 164670 538569 164704 539545
rect 164758 538569 164792 539545
rect 164893 538576 164927 539552
rect 164989 538576 165023 539552
rect 165085 538576 165119 539552
rect 165181 538576 165215 539552
rect 165277 538576 165311 539552
rect 165373 538576 165407 539552
rect 165469 538576 165503 539552
rect 165565 538576 165599 539552
rect 165661 538576 165695 539552
rect 165757 538576 165791 539552
rect 165853 538576 165887 539552
rect 165949 538576 165983 539552
rect 166045 538576 166079 539552
rect 166170 538969 166204 539545
rect 166258 538969 166292 539545
rect 166370 538569 166404 539545
rect 166458 538569 166492 539545
rect 168470 538569 168504 539545
rect 168558 538569 168592 539545
rect 168693 538576 168727 539552
rect 168789 538576 168823 539552
rect 168885 538576 168919 539552
rect 168981 538576 169015 539552
rect 169077 538576 169111 539552
rect 169173 538576 169207 539552
rect 169269 538576 169303 539552
rect 169365 538576 169399 539552
rect 169461 538576 169495 539552
rect 169557 538576 169591 539552
rect 169653 538576 169687 539552
rect 169749 538576 169783 539552
rect 169845 538576 169879 539552
rect 169970 538969 170004 539545
rect 170058 538969 170092 539545
rect 170170 538569 170204 539545
rect 170258 538569 170292 539545
rect 172170 538569 172204 539545
rect 172258 538569 172292 539545
rect 172393 538576 172427 539552
rect 172489 538576 172523 539552
rect 172585 538576 172619 539552
rect 172681 538576 172715 539552
rect 172777 538576 172811 539552
rect 172873 538576 172907 539552
rect 172969 538576 173003 539552
rect 173065 538576 173099 539552
rect 173161 538576 173195 539552
rect 173257 538576 173291 539552
rect 173353 538576 173387 539552
rect 173449 538576 173483 539552
rect 173545 538576 173579 539552
rect 173670 538969 173704 539545
rect 173758 538969 173792 539545
rect 173870 538569 173904 539545
rect 173958 538569 173992 539545
rect 175670 538569 175704 539545
rect 175758 538569 175792 539545
rect 175893 538576 175927 539552
rect 175989 538576 176023 539552
rect 176085 538576 176119 539552
rect 176181 538576 176215 539552
rect 176277 538576 176311 539552
rect 176373 538576 176407 539552
rect 176469 538576 176503 539552
rect 176565 538576 176599 539552
rect 176661 538576 176695 539552
rect 176757 538576 176791 539552
rect 176853 538576 176887 539552
rect 176949 538576 176983 539552
rect 177045 538576 177079 539552
rect 177170 538969 177204 539545
rect 177258 538969 177292 539545
rect 177370 538569 177404 539545
rect 177458 538569 177492 539545
rect 179270 538569 179304 539545
rect 179358 538569 179392 539545
rect 179493 538576 179527 539552
rect 179589 538576 179623 539552
rect 179685 538576 179719 539552
rect 179781 538576 179815 539552
rect 179877 538576 179911 539552
rect 179973 538576 180007 539552
rect 180069 538576 180103 539552
rect 180165 538576 180199 539552
rect 180261 538576 180295 539552
rect 180357 538576 180391 539552
rect 180453 538576 180487 539552
rect 180549 538576 180583 539552
rect 180645 538576 180679 539552
rect 180770 538969 180804 539545
rect 180858 538969 180892 539545
rect 180970 538569 181004 539545
rect 181058 538569 181092 539545
rect 182570 538569 182604 539545
rect 182658 538569 182692 539545
rect 182793 538576 182827 539552
rect 182889 538576 182923 539552
rect 182985 538576 183019 539552
rect 183081 538576 183115 539552
rect 183177 538576 183211 539552
rect 183273 538576 183307 539552
rect 183369 538576 183403 539552
rect 183465 538576 183499 539552
rect 183561 538576 183595 539552
rect 183657 538576 183691 539552
rect 183753 538576 183787 539552
rect 183849 538576 183883 539552
rect 183945 538576 183979 539552
rect 184070 538969 184104 539545
rect 184158 538969 184192 539545
rect 184270 538569 184304 539545
rect 184358 538569 184392 539545
rect 185870 538569 185904 539545
rect 185958 538569 185992 539545
rect 186093 538576 186127 539552
rect 186189 538576 186223 539552
rect 186285 538576 186319 539552
rect 186381 538576 186415 539552
rect 186477 538576 186511 539552
rect 186573 538576 186607 539552
rect 186669 538576 186703 539552
rect 186765 538576 186799 539552
rect 186861 538576 186895 539552
rect 186957 538576 186991 539552
rect 187053 538576 187087 539552
rect 187149 538576 187183 539552
rect 187245 538576 187279 539552
rect 187370 538969 187404 539545
rect 187458 538969 187492 539545
rect 187570 538569 187604 539545
rect 187658 538569 187692 539545
rect 189170 538569 189204 539545
rect 189258 538569 189292 539545
rect 189393 538576 189427 539552
rect 189489 538576 189523 539552
rect 189585 538576 189619 539552
rect 189681 538576 189715 539552
rect 189777 538576 189811 539552
rect 189873 538576 189907 539552
rect 189969 538576 190003 539552
rect 190065 538576 190099 539552
rect 190161 538576 190195 539552
rect 190257 538576 190291 539552
rect 190353 538576 190387 539552
rect 190449 538576 190483 539552
rect 190545 538576 190579 539552
rect 190670 538969 190704 539545
rect 190758 538969 190792 539545
rect 190870 538569 190904 539545
rect 190958 538569 190992 539545
rect 161260 537069 161294 537645
rect 161348 537069 161382 537645
rect 161460 537069 161494 537645
rect 161556 537069 161590 537645
rect 161652 537069 161686 537645
rect 161748 537069 161782 537645
rect 161860 537069 161894 537645
rect 161956 537069 161990 537645
rect 162052 537069 162086 537645
rect 162148 537069 162182 537645
rect 162280 537069 162314 537645
rect 162368 537069 162402 537645
rect 157750 536049 157784 536625
rect 158008 536049 158042 536625
rect 158128 536049 158162 536625
rect 158386 536049 158420 536625
rect 158644 536049 158678 536625
rect 158902 536049 158936 536625
rect 159160 536049 159194 536625
rect 159418 536049 159452 536625
rect 159676 536049 159710 536625
rect 159934 536049 159968 536625
rect 160192 536049 160226 536625
rect 160450 536049 160484 536625
rect 160708 536049 160742 536625
rect 160834 536049 160868 536625
rect 161092 536049 161126 536625
rect 161350 536049 161384 536625
rect 161608 536049 161642 536625
rect 161732 536049 161766 536625
rect 161990 536049 162024 536625
rect 162248 536049 162282 536625
rect 162370 536049 162404 536625
rect 162628 536049 162662 536625
rect 172245 530221 172279 530255
rect 172245 530126 172279 530160
rect 172417 530221 172451 530255
rect 172417 530126 172451 530160
rect 172529 530208 172563 530242
rect 172529 530140 172563 530174
rect 172615 530270 172649 530304
rect 172615 530202 172649 530236
rect 172615 530134 172649 530168
rect 172701 530126 172735 530160
rect 172787 530161 172821 530195
rect 172883 530194 172917 530228
rect 172883 530126 172917 530160
rect 172969 530256 173003 530290
rect 172969 530134 173003 530168
rect 173073 530126 173107 530160
rect 174073 530126 174107 530160
rect 174177 530228 174211 530262
rect 174177 530126 174211 530160
rect 174625 530228 174659 530262
rect 174625 530126 174659 530160
rect 174921 530208 174955 530242
rect 174921 530140 174955 530174
rect 175007 530270 175041 530304
rect 175007 530202 175041 530236
rect 175007 530134 175041 530168
rect 175093 530126 175127 530160
rect 175179 530161 175213 530195
rect 175275 530194 175309 530228
rect 175275 530126 175309 530160
rect 175361 530256 175395 530290
rect 175361 530134 175395 530168
rect 175557 530230 175591 530264
rect 175557 530162 175591 530196
rect 175641 530194 175675 530228
rect 175641 530126 175675 530160
rect 175770 530126 175804 530160
rect 175856 530152 175890 530186
rect 175940 530126 175974 530160
rect 176132 530127 176166 530161
rect 176229 530134 176263 530168
rect 177125 530202 177159 530236
rect 176317 530126 176351 530160
rect 176430 530152 176464 530186
rect 176514 530136 176548 530170
rect 176611 530152 176645 530186
rect 176765 530128 176799 530162
rect 176858 530134 176892 530168
rect 176942 530126 176976 530160
rect 177125 530134 177159 530168
rect 177209 530150 177243 530184
rect 177293 530202 177327 530236
rect 177293 530134 177327 530168
rect 177692 530152 177726 530186
rect 178409 530215 178443 530249
rect 177782 530126 177816 530160
rect 177941 530152 177975 530186
rect 178045 530152 178079 530186
rect 178199 530126 178233 530160
rect 178283 530152 178317 530186
rect 178409 530134 178443 530168
rect 178495 530202 178529 530236
rect 178495 530134 178529 530168
rect 178581 530202 178615 530236
rect 178581 530134 178615 530168
rect 178693 530208 178727 530242
rect 178693 530140 178727 530174
rect 178779 530270 178813 530304
rect 178779 530202 178813 530236
rect 178779 530134 178813 530168
rect 178865 530126 178899 530160
rect 178951 530161 178985 530195
rect 179047 530194 179081 530228
rect 179047 530126 179081 530160
rect 179133 530256 179167 530290
rect 179133 530134 179167 530168
rect 179237 530256 179271 530290
rect 179237 530134 179271 530168
rect 179323 530194 179357 530228
rect 179323 530126 179357 530160
rect 179419 530161 179453 530195
rect 179505 530126 179539 530160
rect 179591 530270 179625 530304
rect 179591 530202 179625 530236
rect 179591 530134 179625 530168
rect 179677 530208 179711 530242
rect 179677 530140 179711 530174
rect 180249 530262 180283 530296
rect 180249 530194 180283 530228
rect 180249 530126 180283 530160
rect 180333 530262 180367 530296
rect 181809 530262 181843 530296
rect 180333 530194 180367 530228
rect 180333 530126 180367 530160
rect 180569 530186 180603 530220
rect 180644 530186 180678 530220
rect 180841 530186 180875 530220
rect 180927 530186 180961 530220
rect 181215 530186 181249 530220
rect 181301 530186 181335 530220
rect 181498 530186 181532 530220
rect 181573 530186 181607 530220
rect 181809 530194 181843 530228
rect 181809 530126 181843 530160
rect 181893 530262 181927 530296
rect 181893 530194 181927 530228
rect 181893 530126 181927 530160
rect 181997 530256 182031 530290
rect 181997 530134 182031 530168
rect 182083 530194 182117 530228
rect 182083 530126 182117 530160
rect 182179 530161 182213 530195
rect 182265 530126 182299 530160
rect 182351 530270 182385 530304
rect 182351 530202 182385 530236
rect 182351 530134 182385 530168
rect 182437 530208 182471 530242
rect 182437 530140 182471 530174
rect 182641 530228 182675 530262
rect 182641 530126 182675 530160
rect 182905 530228 182939 530262
rect 182905 530126 182939 530160
rect 183101 530256 183135 530290
rect 183101 530134 183135 530168
rect 183187 530194 183221 530228
rect 183187 530126 183221 530160
rect 183283 530161 183317 530195
rect 183369 530126 183403 530160
rect 183455 530270 183489 530304
rect 183455 530202 183489 530236
rect 183455 530134 183489 530168
rect 183541 530208 183575 530242
rect 183541 530140 183575 530174
rect 183653 530126 183687 530160
rect 184653 530126 184687 530160
rect 184757 530228 184791 530262
rect 184757 530126 184791 530160
rect 185021 530228 185055 530262
rect 185021 530126 185055 530160
rect 185217 530256 185251 530290
rect 185217 530134 185251 530168
rect 185303 530194 185337 530228
rect 185303 530126 185337 530160
rect 185399 530161 185433 530195
rect 185485 530126 185519 530160
rect 185571 530270 185605 530304
rect 185571 530202 185605 530236
rect 185571 530134 185605 530168
rect 185657 530208 185691 530242
rect 185657 530140 185691 530174
rect 185769 530126 185803 530160
rect 186769 530126 186803 530160
rect 187241 530221 187275 530255
rect 187241 530126 187275 530160
rect 187413 530221 187447 530255
rect 187413 530126 187447 530160
rect 172245 529974 172279 530008
rect 172245 529879 172279 529913
rect 172417 529974 172451 530008
rect 172417 529879 172451 529913
rect 172521 529974 172555 530008
rect 173521 529974 173555 530008
rect 173625 529974 173659 530008
rect 174625 529974 174659 530008
rect 174843 529948 174877 529982
rect 174927 529974 174961 530008
rect 175081 529948 175115 529982
rect 175185 529948 175219 529982
rect 175344 529974 175378 530008
rect 175434 529948 175468 529982
rect 175557 529966 175591 530000
rect 175557 529898 175591 529932
rect 175641 529950 175675 529984
rect 175725 529966 175759 530000
rect 175908 529974 175942 530008
rect 175992 529966 176026 530000
rect 176085 529972 176119 530006
rect 176239 529948 176273 529982
rect 176336 529964 176370 529998
rect 176420 529948 176454 529982
rect 176533 529974 176567 530008
rect 175725 529898 175759 529932
rect 176621 529966 176655 530000
rect 176718 529973 176752 530007
rect 176910 529974 176944 530008
rect 176994 529948 177028 529982
rect 177080 529974 177114 530008
rect 177209 529974 177243 530008
rect 177209 529906 177243 529940
rect 177293 529938 177327 529972
rect 177293 529870 177327 529904
rect 177627 529914 177661 529948
rect 177713 529914 177747 529948
rect 177910 529914 177944 529948
rect 177985 529914 178019 529948
rect 178221 529974 178255 530008
rect 178221 529906 178255 529940
rect 178221 529838 178255 529872
rect 178305 529974 178339 530008
rect 178305 529906 178339 529940
rect 178305 529838 178339 529872
rect 178409 529938 178443 529972
rect 178409 529870 178443 529904
rect 178493 529974 178527 530008
rect 178493 529906 178527 529940
rect 178622 529974 178656 530008
rect 178708 529948 178742 529982
rect 178792 529974 178826 530008
rect 178984 529973 179018 530007
rect 179081 529966 179115 530000
rect 179169 529974 179203 530008
rect 179282 529948 179316 529982
rect 179366 529964 179400 529998
rect 179463 529948 179497 529982
rect 179617 529972 179651 530006
rect 179710 529966 179744 530000
rect 179794 529974 179828 530008
rect 179977 529966 180011 530000
rect 179977 529898 180011 529932
rect 180061 529950 180095 529984
rect 180145 529966 180179 530000
rect 180145 529898 180179 529932
rect 180249 529966 180283 530000
rect 180249 529898 180283 529932
rect 180333 529950 180367 529984
rect 180417 529966 180451 530000
rect 180600 529974 180634 530008
rect 180684 529966 180718 530000
rect 180777 529972 180811 530006
rect 180931 529948 180965 529982
rect 181028 529964 181062 529998
rect 181112 529948 181146 529982
rect 181225 529974 181259 530008
rect 180417 529898 180451 529932
rect 181313 529966 181347 530000
rect 181410 529973 181444 530007
rect 181602 529974 181636 530008
rect 181686 529948 181720 529982
rect 181772 529974 181806 530008
rect 181901 529974 181935 530008
rect 181901 529906 181935 529940
rect 181985 529938 182019 529972
rect 181985 529870 182019 529904
rect 182089 529974 182123 530008
rect 182089 529872 182123 529906
rect 182353 529974 182387 530008
rect 182353 529872 182387 529906
rect 182660 529948 182694 529982
rect 182750 529974 182784 530008
rect 182909 529948 182943 529982
rect 183013 529948 183047 529982
rect 183167 529974 183201 530008
rect 183251 529948 183285 529982
rect 183377 529974 183411 530008
rect 184377 529974 184411 530008
rect 184481 529974 184515 530008
rect 185481 529974 185515 530008
rect 185585 529974 185619 530008
rect 186585 529974 186619 530008
rect 186689 529974 186723 530008
rect 186689 529872 186723 529906
rect 187137 529974 187171 530008
rect 187137 529872 187171 529906
rect 187241 529974 187275 530008
rect 187241 529879 187275 529913
rect 187413 529974 187447 530008
rect 187413 529879 187447 529913
rect 172245 529133 172279 529167
rect 172245 529038 172279 529072
rect 172417 529133 172451 529167
rect 172417 529038 172451 529072
rect 172521 529038 172555 529072
rect 173521 529038 173555 529072
rect 173625 529038 173659 529072
rect 174625 529038 174659 529072
rect 175737 529174 175771 529208
rect 175143 529098 175177 529132
rect 175229 529098 175263 529132
rect 175426 529098 175460 529132
rect 175501 529098 175535 529132
rect 175737 529106 175771 529140
rect 175737 529038 175771 529072
rect 175821 529174 175855 529208
rect 175821 529106 175855 529140
rect 175821 529038 175855 529072
rect 175942 529062 175976 529096
rect 176028 529168 176062 529202
rect 176028 529082 176062 529116
rect 176114 529062 176148 529096
rect 176200 529168 176234 529202
rect 176200 529082 176234 529116
rect 176286 529062 176320 529096
rect 176372 529168 176406 529202
rect 176372 529082 176406 529116
rect 176458 529062 176492 529096
rect 176544 529168 176578 529202
rect 176544 529082 176578 529116
rect 176629 529062 176663 529096
rect 176715 529168 176749 529202
rect 176715 529082 176749 529116
rect 176801 529062 176835 529096
rect 176887 529168 176921 529202
rect 176887 529082 176921 529116
rect 176973 529062 177007 529096
rect 177059 529168 177093 529202
rect 177059 529082 177093 529116
rect 177145 529062 177179 529096
rect 177231 529168 177265 529202
rect 177231 529082 177265 529116
rect 177317 529106 177351 529140
rect 177317 529038 177351 529072
rect 177403 529122 177437 529156
rect 177403 529054 177437 529088
rect 177489 529106 177523 529140
rect 177489 529038 177523 529072
rect 177575 529114 177609 529148
rect 177575 529046 177609 529080
rect 177661 529106 177695 529140
rect 177661 529038 177695 529072
rect 177765 529114 177799 529148
rect 177765 529046 177799 529080
rect 177849 529062 177883 529096
rect 177933 529114 177967 529148
rect 177933 529046 177967 529080
rect 178116 529038 178150 529072
rect 178200 529046 178234 529080
rect 178293 529040 178327 529074
rect 178447 529064 178481 529098
rect 178544 529048 178578 529082
rect 178628 529064 178662 529098
rect 178741 529038 178775 529072
rect 178829 529046 178863 529080
rect 178926 529039 178960 529073
rect 179118 529038 179152 529072
rect 179202 529064 179236 529098
rect 179288 529038 179322 529072
rect 179417 529106 179451 529140
rect 179417 529038 179451 529072
rect 179501 529142 179535 529176
rect 179501 529074 179535 529108
rect 179697 529114 179731 529148
rect 179697 529046 179731 529080
rect 179783 529114 179817 529148
rect 179783 529046 179817 529080
rect 179869 529127 179903 529161
rect 179869 529046 179903 529080
rect 180065 529140 180099 529174
rect 180065 529038 180099 529072
rect 180513 529140 180547 529174
rect 180513 529038 180547 529072
rect 180709 529106 180743 529140
rect 180709 529038 180743 529072
rect 180795 529114 180829 529148
rect 180795 529046 180829 529080
rect 180881 529106 180915 529140
rect 180881 529038 180915 529072
rect 180967 529122 181001 529156
rect 180967 529054 181001 529088
rect 181053 529106 181087 529140
rect 181053 529038 181087 529072
rect 181139 529168 181173 529202
rect 181139 529082 181173 529116
rect 181225 529062 181259 529096
rect 181311 529168 181345 529202
rect 181311 529082 181345 529116
rect 181397 529062 181431 529096
rect 181483 529168 181517 529202
rect 181483 529082 181517 529116
rect 181569 529062 181603 529096
rect 181655 529168 181689 529202
rect 181655 529082 181689 529116
rect 181741 529062 181775 529096
rect 181826 529168 181860 529202
rect 181826 529082 181860 529116
rect 181912 529062 181946 529096
rect 181998 529168 182032 529202
rect 181998 529082 182032 529116
rect 182084 529062 182118 529096
rect 182170 529168 182204 529202
rect 182170 529082 182204 529116
rect 182256 529062 182290 529096
rect 182342 529168 182376 529202
rect 182342 529082 182376 529116
rect 182428 529062 182462 529096
rect 182549 529127 182583 529161
rect 182549 529046 182583 529080
rect 182635 529114 182669 529148
rect 182635 529046 182669 529080
rect 182721 529114 182755 529148
rect 182721 529046 182755 529080
rect 182825 529038 182859 529072
rect 183825 529038 183859 529072
rect 183929 529038 183963 529072
rect 184929 529038 184963 529072
rect 185217 529038 185251 529072
rect 186217 529038 186251 529072
rect 186321 529140 186355 529174
rect 186321 529038 186355 529072
rect 186953 529140 186987 529174
rect 186953 529038 186987 529072
rect 187241 529133 187275 529167
rect 187241 529038 187275 529072
rect 187413 529133 187447 529167
rect 187413 529038 187447 529072
rect 172245 528886 172279 528920
rect 172245 528791 172279 528825
rect 172417 528886 172451 528920
rect 172417 528791 172451 528825
rect 172521 528886 172555 528920
rect 173521 528886 173555 528920
rect 173625 528886 173659 528920
rect 174625 528886 174659 528920
rect 174729 528886 174763 528920
rect 175729 528886 175763 528920
rect 175925 528878 175959 528912
rect 175925 528810 175959 528844
rect 176011 528878 176045 528912
rect 176011 528810 176045 528844
rect 176097 528878 176131 528912
rect 176097 528797 176131 528831
rect 176201 528878 176235 528912
rect 176201 528810 176235 528844
rect 176287 528878 176321 528912
rect 176287 528810 176321 528844
rect 176373 528878 176407 528912
rect 176373 528797 176407 528831
rect 176523 528826 176557 528860
rect 176609 528826 176643 528860
rect 176806 528826 176840 528860
rect 176881 528826 176915 528860
rect 177117 528886 177151 528920
rect 177117 528818 177151 528852
rect 177117 528750 177151 528784
rect 177201 528886 177235 528920
rect 177201 528818 177235 528852
rect 177201 528750 177235 528784
rect 177508 528860 177542 528894
rect 177598 528886 177632 528920
rect 177757 528860 177791 528894
rect 177861 528860 177895 528894
rect 178015 528886 178049 528920
rect 178099 528860 178133 528894
rect 178409 528886 178443 528920
rect 178409 528818 178443 528852
rect 178495 528878 178529 528912
rect 178495 528810 178529 528844
rect 178581 528886 178615 528920
rect 178581 528818 178615 528852
rect 178667 528870 178701 528904
rect 178667 528802 178701 528836
rect 178753 528886 178787 528920
rect 178753 528818 178787 528852
rect 178839 528842 178873 528876
rect 178839 528756 178873 528790
rect 178925 528862 178959 528896
rect 179011 528842 179045 528876
rect 179011 528756 179045 528790
rect 179097 528862 179131 528896
rect 179183 528842 179217 528876
rect 179183 528756 179217 528790
rect 179269 528862 179303 528896
rect 179355 528842 179389 528876
rect 179355 528756 179389 528790
rect 179441 528862 179475 528896
rect 179526 528842 179560 528876
rect 179526 528756 179560 528790
rect 179612 528862 179646 528896
rect 179698 528842 179732 528876
rect 179698 528756 179732 528790
rect 179784 528862 179818 528896
rect 179870 528842 179904 528876
rect 179870 528756 179904 528790
rect 179956 528862 179990 528896
rect 180042 528842 180076 528876
rect 180042 528756 180076 528790
rect 180128 528862 180162 528896
rect 180249 528878 180283 528912
rect 180249 528810 180283 528844
rect 180335 528878 180369 528912
rect 180335 528810 180369 528844
rect 180421 528878 180455 528912
rect 180421 528797 180455 528831
rect 180525 528878 180559 528912
rect 180525 528810 180559 528844
rect 180609 528862 180643 528896
rect 180693 528878 180727 528912
rect 180876 528886 180910 528920
rect 180960 528878 180994 528912
rect 181053 528884 181087 528918
rect 181207 528860 181241 528894
rect 181304 528876 181338 528910
rect 181388 528860 181422 528894
rect 181501 528886 181535 528920
rect 180693 528810 180727 528844
rect 181589 528878 181623 528912
rect 181686 528885 181720 528919
rect 181878 528886 181912 528920
rect 181962 528860 181996 528894
rect 182048 528886 182082 528920
rect 182177 528886 182211 528920
rect 182177 528818 182211 528852
rect 182261 528850 182295 528884
rect 182261 528782 182295 528816
rect 182641 528886 182675 528920
rect 183641 528886 183675 528920
rect 183745 528886 183779 528920
rect 184745 528886 184779 528920
rect 184849 528886 184883 528920
rect 185849 528886 185883 528920
rect 185953 528886 185987 528920
rect 186953 528886 186987 528920
rect 187241 528886 187275 528920
rect 187241 528791 187275 528825
rect 187413 528886 187447 528920
rect 187413 528791 187447 528825
rect 172245 528045 172279 528079
rect 172245 527950 172279 527984
rect 172417 528045 172451 528079
rect 172417 527950 172451 527984
rect 172521 527950 172555 527984
rect 173521 527950 173555 527984
rect 173625 527950 173659 527984
rect 174625 527950 174659 527984
rect 174913 527950 174947 527984
rect 175913 527950 175947 527984
rect 176109 528026 176143 528060
rect 176109 527958 176143 527992
rect 176193 527974 176227 528008
rect 176277 528026 176311 528060
rect 176277 527958 176311 527992
rect 176460 527950 176494 527984
rect 176544 527958 176578 527992
rect 176637 527952 176671 527986
rect 176791 527976 176825 528010
rect 176888 527960 176922 527994
rect 176972 527976 177006 528010
rect 177085 527950 177119 527984
rect 177173 527958 177207 527992
rect 177270 527951 177304 527985
rect 177462 527950 177496 527984
rect 177546 527976 177580 528010
rect 177632 527950 177666 527984
rect 177761 528018 177795 528052
rect 177761 527950 177795 527984
rect 177845 528054 177879 528088
rect 177845 527986 177879 528020
rect 177949 528039 177983 528073
rect 177949 527958 177983 527992
rect 178035 528026 178069 528060
rect 178035 527958 178069 527992
rect 178121 528026 178155 528060
rect 178121 527958 178155 527992
rect 178225 528052 178259 528086
rect 178225 527950 178259 527984
rect 178857 528052 178891 528086
rect 178857 527950 178891 527984
rect 178961 528086 178995 528120
rect 178961 528018 178995 528052
rect 178961 527950 178995 527984
rect 179045 528086 179079 528120
rect 179045 528018 179079 528052
rect 179045 527950 179079 527984
rect 179281 528010 179315 528044
rect 179356 528010 179390 528044
rect 179553 528010 179587 528044
rect 179639 528010 179673 528044
rect 180065 528052 180099 528086
rect 180065 527950 180099 527984
rect 180697 528052 180731 528086
rect 180697 527950 180731 527984
rect 180985 528086 181019 528120
rect 180985 528018 181019 528052
rect 180985 527950 181019 527984
rect 181069 528086 181103 528120
rect 181069 528018 181103 528052
rect 181069 527950 181103 527984
rect 181305 528010 181339 528044
rect 181380 528010 181414 528044
rect 181577 528010 181611 528044
rect 181663 528010 181697 528044
rect 181813 527950 181847 527984
rect 182813 527950 182847 527984
rect 182917 527950 182951 527984
rect 183917 527950 183951 527984
rect 184021 527950 184055 527984
rect 185021 527950 185055 527984
rect 185217 527950 185251 527984
rect 186217 527950 186251 527984
rect 186321 528052 186355 528086
rect 186321 527950 186355 527984
rect 186953 528052 186987 528086
rect 186953 527950 186987 527984
rect 187241 528045 187275 528079
rect 187241 527950 187275 527984
rect 187413 528045 187447 528079
rect 187413 527950 187447 527984
rect 172245 527798 172279 527832
rect 172245 527703 172279 527737
rect 172417 527798 172451 527832
rect 172417 527703 172451 527737
rect 172521 527798 172555 527832
rect 173521 527798 173555 527832
rect 173625 527798 173659 527832
rect 174625 527798 174659 527832
rect 174729 527798 174763 527832
rect 175729 527798 175763 527832
rect 175833 527798 175867 527832
rect 175833 527696 175867 527730
rect 176281 527798 176315 527832
rect 176281 527696 176315 527730
rect 176404 527772 176438 527806
rect 176494 527798 176528 527832
rect 176653 527772 176687 527806
rect 176757 527772 176791 527806
rect 176911 527798 176945 527832
rect 176995 527772 177029 527806
rect 177121 527798 177155 527832
rect 177121 527703 177155 527737
rect 177293 527798 177327 527832
rect 177293 527703 177327 527737
rect 177489 527798 177523 527832
rect 178489 527798 178523 527832
rect 178593 527798 178627 527832
rect 178593 527696 178627 527730
rect 178857 527798 178891 527832
rect 178857 527696 178891 527730
rect 178980 527772 179014 527806
rect 179070 527798 179104 527832
rect 179229 527772 179263 527806
rect 179333 527772 179367 527806
rect 179487 527798 179521 527832
rect 179571 527772 179605 527806
rect 179697 527798 179731 527832
rect 180697 527798 180731 527832
rect 180801 527798 180835 527832
rect 181801 527798 181835 527832
rect 181905 527798 181939 527832
rect 181905 527696 181939 527730
rect 182353 527798 182387 527832
rect 182353 527696 182387 527730
rect 182641 527798 182675 527832
rect 183641 527798 183675 527832
rect 183745 527798 183779 527832
rect 184745 527798 184779 527832
rect 184849 527798 184883 527832
rect 185849 527798 185883 527832
rect 185953 527798 185987 527832
rect 186953 527798 186987 527832
rect 187241 527798 187275 527832
rect 187241 527703 187275 527737
rect 187413 527798 187447 527832
rect 187413 527703 187447 527737
rect 172245 526957 172279 526991
rect 172245 526862 172279 526896
rect 172417 526957 172451 526991
rect 172417 526862 172451 526896
rect 172521 526862 172555 526896
rect 173521 526862 173555 526896
rect 173625 526862 173659 526896
rect 174625 526862 174659 526896
rect 174913 526862 174947 526896
rect 175913 526862 175947 526896
rect 176017 526862 176051 526896
rect 177017 526862 177051 526896
rect 177121 526862 177155 526896
rect 178121 526862 178155 526896
rect 178225 526862 178259 526896
rect 179225 526862 179259 526896
rect 179329 526964 179363 526998
rect 179329 526862 179363 526896
rect 179777 526964 179811 526998
rect 179777 526862 179811 526896
rect 180065 526862 180099 526896
rect 181065 526862 181099 526896
rect 181169 526862 181203 526896
rect 182169 526862 182203 526896
rect 182273 526862 182307 526896
rect 183273 526862 183307 526896
rect 183377 526862 183411 526896
rect 184377 526862 184411 526896
rect 184481 526964 184515 526998
rect 184481 526862 184515 526896
rect 184929 526964 184963 526998
rect 184929 526862 184963 526896
rect 185217 526862 185251 526896
rect 186217 526862 186251 526896
rect 186321 526964 186355 526998
rect 186321 526862 186355 526896
rect 186953 526964 186987 526998
rect 186953 526862 186987 526896
rect 187241 526957 187275 526991
rect 187241 526862 187275 526896
rect 187413 526957 187447 526991
rect 187413 526862 187447 526896
rect 172245 526710 172279 526744
rect 172245 526615 172279 526649
rect 172417 526710 172451 526744
rect 172417 526615 172451 526649
rect 172521 526710 172555 526744
rect 173521 526710 173555 526744
rect 173625 526710 173659 526744
rect 174625 526710 174659 526744
rect 174729 526710 174763 526744
rect 175729 526710 175763 526744
rect 175833 526710 175867 526744
rect 176833 526710 176867 526744
rect 176937 526710 176971 526744
rect 176937 526608 176971 526642
rect 177201 526710 177235 526744
rect 177201 526608 177235 526642
rect 177489 526710 177523 526744
rect 178489 526710 178523 526744
rect 178593 526710 178627 526744
rect 179593 526710 179627 526744
rect 179697 526710 179731 526744
rect 180697 526710 180731 526744
rect 180801 526710 180835 526744
rect 181801 526710 181835 526744
rect 181905 526710 181939 526744
rect 181905 526608 181939 526642
rect 182353 526710 182387 526744
rect 182353 526608 182387 526642
rect 182641 526710 182675 526744
rect 183641 526710 183675 526744
rect 183745 526710 183779 526744
rect 184745 526710 184779 526744
rect 184849 526710 184883 526744
rect 185849 526710 185883 526744
rect 185953 526710 185987 526744
rect 186953 526710 186987 526744
rect 187241 526710 187275 526744
rect 187241 526615 187275 526649
rect 187413 526710 187447 526744
rect 187413 526615 187447 526649
rect 172245 525869 172279 525903
rect 172245 525774 172279 525808
rect 172417 525869 172451 525903
rect 172417 525774 172451 525808
rect 172521 525774 172555 525808
rect 173521 525774 173555 525808
rect 173625 525774 173659 525808
rect 174625 525774 174659 525808
rect 174913 525774 174947 525808
rect 175913 525774 175947 525808
rect 176017 525774 176051 525808
rect 177017 525774 177051 525808
rect 177121 525774 177155 525808
rect 178121 525774 178155 525808
rect 178225 525774 178259 525808
rect 179225 525774 179259 525808
rect 179329 525876 179363 525910
rect 179329 525774 179363 525808
rect 179777 525876 179811 525910
rect 179777 525774 179811 525808
rect 180065 525774 180099 525808
rect 181065 525774 181099 525808
rect 181169 525774 181203 525808
rect 182169 525774 182203 525808
rect 182273 525774 182307 525808
rect 183273 525774 183307 525808
rect 183377 525774 183411 525808
rect 184377 525774 184411 525808
rect 184481 525876 184515 525910
rect 184481 525774 184515 525808
rect 184929 525876 184963 525910
rect 184929 525774 184963 525808
rect 185217 525774 185251 525808
rect 186217 525774 186251 525808
rect 186321 525876 186355 525910
rect 186321 525774 186355 525808
rect 186953 525876 186987 525910
rect 186953 525774 186987 525808
rect 187241 525869 187275 525903
rect 187241 525774 187275 525808
rect 187413 525869 187447 525903
rect 187413 525774 187447 525808
rect 172245 525622 172279 525656
rect 172245 525527 172279 525561
rect 172417 525622 172451 525656
rect 172417 525527 172451 525561
rect 172521 525622 172555 525656
rect 173521 525622 173555 525656
rect 173625 525622 173659 525656
rect 174625 525622 174659 525656
rect 174729 525622 174763 525656
rect 175729 525622 175763 525656
rect 175833 525622 175867 525656
rect 176833 525622 176867 525656
rect 176937 525622 176971 525656
rect 176937 525520 176971 525554
rect 177201 525622 177235 525656
rect 177201 525520 177235 525554
rect 177489 525622 177523 525656
rect 178489 525622 178523 525656
rect 178593 525622 178627 525656
rect 179593 525622 179627 525656
rect 179697 525622 179731 525656
rect 180697 525622 180731 525656
rect 180801 525622 180835 525656
rect 181801 525622 181835 525656
rect 181905 525622 181939 525656
rect 181905 525520 181939 525554
rect 182353 525622 182387 525656
rect 182353 525520 182387 525554
rect 182641 525622 182675 525656
rect 183641 525622 183675 525656
rect 183745 525622 183779 525656
rect 184745 525622 184779 525656
rect 184849 525622 184883 525656
rect 185849 525622 185883 525656
rect 185953 525622 185987 525656
rect 186953 525622 186987 525656
rect 187241 525622 187275 525656
rect 187241 525527 187275 525561
rect 187413 525622 187447 525656
rect 187413 525527 187447 525561
rect 172245 524781 172279 524815
rect 172245 524686 172279 524720
rect 172417 524781 172451 524815
rect 172417 524686 172451 524720
rect 172521 524686 172555 524720
rect 173521 524686 173555 524720
rect 173625 524686 173659 524720
rect 174625 524686 174659 524720
rect 174913 524686 174947 524720
rect 175913 524686 175947 524720
rect 176017 524686 176051 524720
rect 177017 524686 177051 524720
rect 177121 524686 177155 524720
rect 178121 524686 178155 524720
rect 178225 524686 178259 524720
rect 179225 524686 179259 524720
rect 179329 524788 179363 524822
rect 179329 524686 179363 524720
rect 179777 524788 179811 524822
rect 179777 524686 179811 524720
rect 180065 524686 180099 524720
rect 181065 524686 181099 524720
rect 181169 524686 181203 524720
rect 182169 524686 182203 524720
rect 182273 524686 182307 524720
rect 183273 524686 183307 524720
rect 183377 524686 183411 524720
rect 184377 524686 184411 524720
rect 184481 524788 184515 524822
rect 184481 524686 184515 524720
rect 184929 524788 184963 524822
rect 184929 524686 184963 524720
rect 185217 524686 185251 524720
rect 186217 524686 186251 524720
rect 186321 524788 186355 524822
rect 186321 524686 186355 524720
rect 186953 524788 186987 524822
rect 186953 524686 186987 524720
rect 187241 524781 187275 524815
rect 187241 524686 187275 524720
rect 187413 524781 187447 524815
rect 187413 524686 187447 524720
rect 172245 524534 172279 524568
rect 172245 524439 172279 524473
rect 172417 524534 172451 524568
rect 172417 524439 172451 524473
rect 172521 524534 172555 524568
rect 173521 524534 173555 524568
rect 173625 524534 173659 524568
rect 174625 524534 174659 524568
rect 174729 524534 174763 524568
rect 175729 524534 175763 524568
rect 175833 524534 175867 524568
rect 176833 524534 176867 524568
rect 176937 524534 176971 524568
rect 176937 524432 176971 524466
rect 177201 524534 177235 524568
rect 177201 524432 177235 524466
rect 177489 524534 177523 524568
rect 178489 524534 178523 524568
rect 178593 524534 178627 524568
rect 179593 524534 179627 524568
rect 179697 524534 179731 524568
rect 180697 524534 180731 524568
rect 180801 524534 180835 524568
rect 181801 524534 181835 524568
rect 181905 524534 181939 524568
rect 181905 524432 181939 524466
rect 182353 524534 182387 524568
rect 182353 524432 182387 524466
rect 182641 524534 182675 524568
rect 183641 524534 183675 524568
rect 183745 524534 183779 524568
rect 184745 524534 184779 524568
rect 184849 524534 184883 524568
rect 185849 524534 185883 524568
rect 185953 524534 185987 524568
rect 186953 524534 186987 524568
rect 187241 524534 187275 524568
rect 187241 524439 187275 524473
rect 187413 524534 187447 524568
rect 187413 524439 187447 524473
rect 172245 523693 172279 523727
rect 172245 523598 172279 523632
rect 172417 523693 172451 523727
rect 172417 523598 172451 523632
rect 172521 523598 172555 523632
rect 173521 523598 173555 523632
rect 173625 523598 173659 523632
rect 174625 523598 174659 523632
rect 174913 523598 174947 523632
rect 175913 523598 175947 523632
rect 176017 523598 176051 523632
rect 177017 523598 177051 523632
rect 177121 523598 177155 523632
rect 178121 523598 178155 523632
rect 178225 523598 178259 523632
rect 179225 523598 179259 523632
rect 179329 523700 179363 523734
rect 179329 523598 179363 523632
rect 179777 523700 179811 523734
rect 179777 523598 179811 523632
rect 180065 523598 180099 523632
rect 181065 523598 181099 523632
rect 181169 523598 181203 523632
rect 182169 523598 182203 523632
rect 182273 523598 182307 523632
rect 183273 523598 183307 523632
rect 183377 523598 183411 523632
rect 184377 523598 184411 523632
rect 184481 523700 184515 523734
rect 184481 523598 184515 523632
rect 184929 523700 184963 523734
rect 184929 523598 184963 523632
rect 185217 523598 185251 523632
rect 186217 523598 186251 523632
rect 186321 523700 186355 523734
rect 186321 523598 186355 523632
rect 186953 523700 186987 523734
rect 186953 523598 186987 523632
rect 187241 523693 187275 523727
rect 187241 523598 187275 523632
rect 187413 523693 187447 523727
rect 187413 523598 187447 523632
rect 172245 523446 172279 523480
rect 172245 523351 172279 523385
rect 172417 523446 172451 523480
rect 172417 523351 172451 523385
rect 172521 523446 172555 523480
rect 173521 523446 173555 523480
rect 173625 523446 173659 523480
rect 174625 523446 174659 523480
rect 174729 523446 174763 523480
rect 175729 523446 175763 523480
rect 175833 523446 175867 523480
rect 176833 523446 176867 523480
rect 176937 523446 176971 523480
rect 176937 523344 176971 523378
rect 177201 523446 177235 523480
rect 177201 523344 177235 523378
rect 177489 523446 177523 523480
rect 178489 523446 178523 523480
rect 178593 523446 178627 523480
rect 179593 523446 179627 523480
rect 179697 523446 179731 523480
rect 180697 523446 180731 523480
rect 180801 523446 180835 523480
rect 181801 523446 181835 523480
rect 181905 523446 181939 523480
rect 181905 523344 181939 523378
rect 182353 523446 182387 523480
rect 182353 523344 182387 523378
rect 182641 523446 182675 523480
rect 183641 523446 183675 523480
rect 183745 523446 183779 523480
rect 184745 523446 184779 523480
rect 184849 523446 184883 523480
rect 185849 523446 185883 523480
rect 185953 523446 185987 523480
rect 186953 523446 186987 523480
rect 187241 523446 187275 523480
rect 187241 523351 187275 523385
rect 187413 523446 187447 523480
rect 187413 523351 187447 523385
rect 172245 522605 172279 522639
rect 172245 522510 172279 522544
rect 172417 522605 172451 522639
rect 172417 522510 172451 522544
rect 172521 522510 172555 522544
rect 173521 522510 173555 522544
rect 173625 522510 173659 522544
rect 174625 522510 174659 522544
rect 174913 522510 174947 522544
rect 175913 522510 175947 522544
rect 176017 522510 176051 522544
rect 177017 522510 177051 522544
rect 177121 522510 177155 522544
rect 178121 522510 178155 522544
rect 178225 522510 178259 522544
rect 179225 522510 179259 522544
rect 179329 522612 179363 522646
rect 179329 522510 179363 522544
rect 179777 522612 179811 522646
rect 179777 522510 179811 522544
rect 180065 522510 180099 522544
rect 181065 522510 181099 522544
rect 181169 522510 181203 522544
rect 182169 522510 182203 522544
rect 182273 522510 182307 522544
rect 183273 522510 183307 522544
rect 183377 522510 183411 522544
rect 184377 522510 184411 522544
rect 184481 522612 184515 522646
rect 184481 522510 184515 522544
rect 184929 522612 184963 522646
rect 184929 522510 184963 522544
rect 185217 522510 185251 522544
rect 186217 522510 186251 522544
rect 186321 522612 186355 522646
rect 186321 522510 186355 522544
rect 186953 522612 186987 522646
rect 186953 522510 186987 522544
rect 187241 522605 187275 522639
rect 187241 522510 187275 522544
rect 187413 522605 187447 522639
rect 187413 522510 187447 522544
rect 172245 522358 172279 522392
rect 172245 522263 172279 522297
rect 172417 522358 172451 522392
rect 172417 522263 172451 522297
rect 172521 522358 172555 522392
rect 173521 522358 173555 522392
rect 173625 522358 173659 522392
rect 174625 522358 174659 522392
rect 174729 522358 174763 522392
rect 175729 522358 175763 522392
rect 175833 522358 175867 522392
rect 176833 522358 176867 522392
rect 176937 522358 176971 522392
rect 176937 522256 176971 522290
rect 177201 522358 177235 522392
rect 177201 522256 177235 522290
rect 177489 522358 177523 522392
rect 178489 522358 178523 522392
rect 178593 522358 178627 522392
rect 179593 522358 179627 522392
rect 179697 522358 179731 522392
rect 180697 522358 180731 522392
rect 180801 522358 180835 522392
rect 181801 522358 181835 522392
rect 181905 522358 181939 522392
rect 181905 522256 181939 522290
rect 182353 522358 182387 522392
rect 182353 522256 182387 522290
rect 182641 522358 182675 522392
rect 183641 522358 183675 522392
rect 183745 522358 183779 522392
rect 184745 522358 184779 522392
rect 184849 522358 184883 522392
rect 185849 522358 185883 522392
rect 185953 522358 185987 522392
rect 186953 522358 186987 522392
rect 187241 522358 187275 522392
rect 187241 522263 187275 522297
rect 187413 522358 187447 522392
rect 187413 522263 187447 522297
rect 172245 521517 172279 521551
rect 172245 521422 172279 521456
rect 172417 521517 172451 521551
rect 172417 521422 172451 521456
rect 172521 521422 172555 521456
rect 173521 521422 173555 521456
rect 173625 521422 173659 521456
rect 174625 521422 174659 521456
rect 174913 521422 174947 521456
rect 175913 521422 175947 521456
rect 176017 521422 176051 521456
rect 177017 521422 177051 521456
rect 177121 521422 177155 521456
rect 178121 521422 178155 521456
rect 178225 521422 178259 521456
rect 179225 521422 179259 521456
rect 179329 521524 179363 521558
rect 179329 521422 179363 521456
rect 179777 521524 179811 521558
rect 179777 521422 179811 521456
rect 180065 521422 180099 521456
rect 181065 521422 181099 521456
rect 181169 521422 181203 521456
rect 182169 521422 182203 521456
rect 182273 521422 182307 521456
rect 183273 521422 183307 521456
rect 183377 521422 183411 521456
rect 184377 521422 184411 521456
rect 184481 521524 184515 521558
rect 184481 521422 184515 521456
rect 184929 521524 184963 521558
rect 184929 521422 184963 521456
rect 185217 521422 185251 521456
rect 186217 521422 186251 521456
rect 186321 521524 186355 521558
rect 186321 521422 186355 521456
rect 186953 521524 186987 521558
rect 186953 521422 186987 521456
rect 187241 521517 187275 521551
rect 187241 521422 187275 521456
rect 187413 521517 187447 521551
rect 187413 521422 187447 521456
rect 172245 521270 172279 521304
rect 172245 521175 172279 521209
rect 172417 521270 172451 521304
rect 172417 521175 172451 521209
rect 172521 521270 172555 521304
rect 173521 521270 173555 521304
rect 173625 521270 173659 521304
rect 174625 521270 174659 521304
rect 174729 521270 174763 521304
rect 175729 521270 175763 521304
rect 175833 521270 175867 521304
rect 176833 521270 176867 521304
rect 176937 521270 176971 521304
rect 176937 521168 176971 521202
rect 177201 521270 177235 521304
rect 177201 521168 177235 521202
rect 177489 521270 177523 521304
rect 178489 521270 178523 521304
rect 178593 521270 178627 521304
rect 179593 521270 179627 521304
rect 179697 521270 179731 521304
rect 180697 521270 180731 521304
rect 180801 521270 180835 521304
rect 181801 521270 181835 521304
rect 181905 521270 181939 521304
rect 181905 521168 181939 521202
rect 182353 521270 182387 521304
rect 182353 521168 182387 521202
rect 182641 521270 182675 521304
rect 183641 521270 183675 521304
rect 183745 521270 183779 521304
rect 184745 521270 184779 521304
rect 184849 521270 184883 521304
rect 185849 521270 185883 521304
rect 185953 521270 185987 521304
rect 186953 521270 186987 521304
rect 187241 521270 187275 521304
rect 187241 521175 187275 521209
rect 187413 521270 187447 521304
rect 187413 521175 187447 521209
rect 172245 520429 172279 520463
rect 172245 520334 172279 520368
rect 172417 520429 172451 520463
rect 172417 520334 172451 520368
rect 172521 520334 172555 520368
rect 173521 520334 173555 520368
rect 173625 520334 173659 520368
rect 174625 520334 174659 520368
rect 174913 520334 174947 520368
rect 175913 520334 175947 520368
rect 176017 520334 176051 520368
rect 177017 520334 177051 520368
rect 177121 520334 177155 520368
rect 178121 520334 178155 520368
rect 178225 520334 178259 520368
rect 179225 520334 179259 520368
rect 179329 520436 179363 520470
rect 179329 520334 179363 520368
rect 179777 520436 179811 520470
rect 179777 520334 179811 520368
rect 180065 520334 180099 520368
rect 181065 520334 181099 520368
rect 181169 520334 181203 520368
rect 182169 520334 182203 520368
rect 182273 520334 182307 520368
rect 183273 520334 183307 520368
rect 183377 520334 183411 520368
rect 184377 520334 184411 520368
rect 184481 520436 184515 520470
rect 184481 520334 184515 520368
rect 184929 520436 184963 520470
rect 184929 520334 184963 520368
rect 185217 520334 185251 520368
rect 186217 520334 186251 520368
rect 186321 520436 186355 520470
rect 186321 520334 186355 520368
rect 186953 520436 186987 520470
rect 186953 520334 186987 520368
rect 187241 520429 187275 520463
rect 187241 520334 187275 520368
rect 187413 520429 187447 520463
rect 187413 520334 187447 520368
rect 172245 520182 172279 520216
rect 172245 520087 172279 520121
rect 172417 520182 172451 520216
rect 172417 520087 172451 520121
rect 172521 520182 172555 520216
rect 173521 520182 173555 520216
rect 173625 520182 173659 520216
rect 174625 520182 174659 520216
rect 174729 520182 174763 520216
rect 175729 520182 175763 520216
rect 175833 520182 175867 520216
rect 176833 520182 176867 520216
rect 176937 520182 176971 520216
rect 176937 520080 176971 520114
rect 177201 520182 177235 520216
rect 177201 520080 177235 520114
rect 177489 520182 177523 520216
rect 178489 520182 178523 520216
rect 178593 520182 178627 520216
rect 179593 520182 179627 520216
rect 179697 520182 179731 520216
rect 180697 520182 180731 520216
rect 180801 520182 180835 520216
rect 181801 520182 181835 520216
rect 181905 520182 181939 520216
rect 181905 520080 181939 520114
rect 182353 520182 182387 520216
rect 182353 520080 182387 520114
rect 182641 520182 182675 520216
rect 183641 520182 183675 520216
rect 183745 520182 183779 520216
rect 184745 520182 184779 520216
rect 184849 520182 184883 520216
rect 185849 520182 185883 520216
rect 185953 520182 185987 520216
rect 186953 520182 186987 520216
rect 187241 520182 187275 520216
rect 187241 520087 187275 520121
rect 187413 520182 187447 520216
rect 187413 520087 187447 520121
rect 172245 519341 172279 519375
rect 172245 519246 172279 519280
rect 172417 519341 172451 519375
rect 172417 519246 172451 519280
rect 172521 519246 172555 519280
rect 173521 519246 173555 519280
rect 173625 519246 173659 519280
rect 174625 519246 174659 519280
rect 174913 519246 174947 519280
rect 175913 519246 175947 519280
rect 176017 519246 176051 519280
rect 177017 519246 177051 519280
rect 177121 519246 177155 519280
rect 178121 519246 178155 519280
rect 178225 519246 178259 519280
rect 179225 519246 179259 519280
rect 179329 519348 179363 519382
rect 179329 519246 179363 519280
rect 179777 519348 179811 519382
rect 179777 519246 179811 519280
rect 180065 519246 180099 519280
rect 181065 519246 181099 519280
rect 181169 519246 181203 519280
rect 182169 519246 182203 519280
rect 182273 519246 182307 519280
rect 183273 519246 183307 519280
rect 183377 519246 183411 519280
rect 184377 519246 184411 519280
rect 184481 519348 184515 519382
rect 184481 519246 184515 519280
rect 184929 519348 184963 519382
rect 184929 519246 184963 519280
rect 185217 519246 185251 519280
rect 186217 519246 186251 519280
rect 186321 519348 186355 519382
rect 186321 519246 186355 519280
rect 186953 519348 186987 519382
rect 186953 519246 186987 519280
rect 187241 519341 187275 519375
rect 187241 519246 187275 519280
rect 187413 519341 187447 519375
rect 187413 519246 187447 519280
rect 172245 519094 172279 519128
rect 172245 518999 172279 519033
rect 172417 519094 172451 519128
rect 172417 518999 172451 519033
rect 172521 519094 172555 519128
rect 173521 519094 173555 519128
rect 173625 519094 173659 519128
rect 174625 519094 174659 519128
rect 174729 519094 174763 519128
rect 175729 519094 175763 519128
rect 175833 519094 175867 519128
rect 176833 519094 176867 519128
rect 176937 519094 176971 519128
rect 176937 518992 176971 519026
rect 177201 519094 177235 519128
rect 177201 518992 177235 519026
rect 177489 519094 177523 519128
rect 178489 519094 178523 519128
rect 178593 519094 178627 519128
rect 179593 519094 179627 519128
rect 179697 519094 179731 519128
rect 180697 519094 180731 519128
rect 180801 519094 180835 519128
rect 181801 519094 181835 519128
rect 181905 519094 181939 519128
rect 181905 518992 181939 519026
rect 182353 519094 182387 519128
rect 182353 518992 182387 519026
rect 182641 519094 182675 519128
rect 183641 519094 183675 519128
rect 183745 519094 183779 519128
rect 184745 519094 184779 519128
rect 184849 519094 184883 519128
rect 185849 519094 185883 519128
rect 185953 519094 185987 519128
rect 186953 519094 186987 519128
rect 187241 519094 187275 519128
rect 187241 518999 187275 519033
rect 187413 519094 187447 519128
rect 187413 518999 187447 519033
rect 172245 518253 172279 518287
rect 172245 518158 172279 518192
rect 172417 518253 172451 518287
rect 172417 518158 172451 518192
rect 172521 518158 172555 518192
rect 173521 518158 173555 518192
rect 173625 518158 173659 518192
rect 174625 518158 174659 518192
rect 174913 518158 174947 518192
rect 175913 518158 175947 518192
rect 176017 518158 176051 518192
rect 177017 518158 177051 518192
rect 177121 518158 177155 518192
rect 178121 518158 178155 518192
rect 178225 518158 178259 518192
rect 179225 518158 179259 518192
rect 179329 518260 179363 518294
rect 179329 518158 179363 518192
rect 179777 518260 179811 518294
rect 179777 518158 179811 518192
rect 180065 518158 180099 518192
rect 181065 518158 181099 518192
rect 181169 518158 181203 518192
rect 182169 518158 182203 518192
rect 182273 518158 182307 518192
rect 183273 518158 183307 518192
rect 183377 518158 183411 518192
rect 184377 518158 184411 518192
rect 184481 518260 184515 518294
rect 184481 518158 184515 518192
rect 184929 518260 184963 518294
rect 184929 518158 184963 518192
rect 185217 518158 185251 518192
rect 186217 518158 186251 518192
rect 186321 518260 186355 518294
rect 186321 518158 186355 518192
rect 186953 518260 186987 518294
rect 186953 518158 186987 518192
rect 187241 518253 187275 518287
rect 187241 518158 187275 518192
rect 187413 518253 187447 518287
rect 187413 518158 187447 518192
rect 172245 518006 172279 518040
rect 172245 517911 172279 517945
rect 172417 518006 172451 518040
rect 172417 517911 172451 517945
rect 172521 518006 172555 518040
rect 173521 518006 173555 518040
rect 173625 518006 173659 518040
rect 174625 518006 174659 518040
rect 174729 518006 174763 518040
rect 175729 518006 175763 518040
rect 175833 518006 175867 518040
rect 176833 518006 176867 518040
rect 176937 518006 176971 518040
rect 176937 517904 176971 517938
rect 177201 518006 177235 518040
rect 177201 517904 177235 517938
rect 177489 518006 177523 518040
rect 178489 518006 178523 518040
rect 178593 518006 178627 518040
rect 179593 518006 179627 518040
rect 179697 518006 179731 518040
rect 180697 518006 180731 518040
rect 180801 518006 180835 518040
rect 181801 518006 181835 518040
rect 181905 518006 181939 518040
rect 181905 517904 181939 517938
rect 182353 518006 182387 518040
rect 182353 517904 182387 517938
rect 182641 518006 182675 518040
rect 183641 518006 183675 518040
rect 183745 518006 183779 518040
rect 184745 518006 184779 518040
rect 184849 518006 184883 518040
rect 185849 518006 185883 518040
rect 185953 518006 185987 518040
rect 186953 518006 186987 518040
rect 187241 518006 187275 518040
rect 187241 517911 187275 517945
rect 187413 518006 187447 518040
rect 187413 517911 187447 517945
rect 172245 517165 172279 517199
rect 172245 517070 172279 517104
rect 172417 517165 172451 517199
rect 172417 517070 172451 517104
rect 172521 517070 172555 517104
rect 173521 517070 173555 517104
rect 173625 517070 173659 517104
rect 174625 517070 174659 517104
rect 174913 517070 174947 517104
rect 175913 517070 175947 517104
rect 176017 517070 176051 517104
rect 177017 517070 177051 517104
rect 177121 517070 177155 517104
rect 178121 517070 178155 517104
rect 178225 517070 178259 517104
rect 179225 517070 179259 517104
rect 179329 517172 179363 517206
rect 179329 517070 179363 517104
rect 179777 517172 179811 517206
rect 179777 517070 179811 517104
rect 180065 517070 180099 517104
rect 181065 517070 181099 517104
rect 181169 517070 181203 517104
rect 182169 517070 182203 517104
rect 182273 517070 182307 517104
rect 183273 517070 183307 517104
rect 183377 517070 183411 517104
rect 184377 517070 184411 517104
rect 184481 517172 184515 517206
rect 184481 517070 184515 517104
rect 184929 517172 184963 517206
rect 184929 517070 184963 517104
rect 185217 517070 185251 517104
rect 186217 517070 186251 517104
rect 186321 517172 186355 517206
rect 186321 517070 186355 517104
rect 186953 517172 186987 517206
rect 186953 517070 186987 517104
rect 187241 517165 187275 517199
rect 187241 517070 187275 517104
rect 187413 517165 187447 517199
rect 187413 517070 187447 517104
rect 172245 516918 172279 516952
rect 172245 516823 172279 516857
rect 172417 516918 172451 516952
rect 172417 516823 172451 516857
rect 172521 516918 172555 516952
rect 173521 516918 173555 516952
rect 173625 516918 173659 516952
rect 174625 516918 174659 516952
rect 174729 516918 174763 516952
rect 175729 516918 175763 516952
rect 175833 516918 175867 516952
rect 176833 516918 176867 516952
rect 176937 516918 176971 516952
rect 176937 516816 176971 516850
rect 177201 516918 177235 516952
rect 177201 516816 177235 516850
rect 177489 516918 177523 516952
rect 178489 516918 178523 516952
rect 178593 516918 178627 516952
rect 179593 516918 179627 516952
rect 179697 516918 179731 516952
rect 180697 516918 180731 516952
rect 180801 516918 180835 516952
rect 181801 516918 181835 516952
rect 181905 516918 181939 516952
rect 181905 516816 181939 516850
rect 182353 516918 182387 516952
rect 182353 516816 182387 516850
rect 182641 516918 182675 516952
rect 183641 516918 183675 516952
rect 183745 516918 183779 516952
rect 184745 516918 184779 516952
rect 184849 516918 184883 516952
rect 185849 516918 185883 516952
rect 185953 516918 185987 516952
rect 186953 516918 186987 516952
rect 187241 516918 187275 516952
rect 187241 516823 187275 516857
rect 187413 516918 187447 516952
rect 187413 516823 187447 516857
rect 172245 516077 172279 516111
rect 172245 515982 172279 516016
rect 172417 516077 172451 516111
rect 172417 515982 172451 516016
rect 172521 515982 172555 516016
rect 173521 515982 173555 516016
rect 173625 515982 173659 516016
rect 174625 515982 174659 516016
rect 174913 515982 174947 516016
rect 175913 515982 175947 516016
rect 176017 515982 176051 516016
rect 177017 515982 177051 516016
rect 177121 515982 177155 516016
rect 178121 515982 178155 516016
rect 178225 515982 178259 516016
rect 179225 515982 179259 516016
rect 179329 516084 179363 516118
rect 179329 515982 179363 516016
rect 179777 516084 179811 516118
rect 179777 515982 179811 516016
rect 180065 515982 180099 516016
rect 181065 515982 181099 516016
rect 181169 515982 181203 516016
rect 182169 515982 182203 516016
rect 182273 515982 182307 516016
rect 183273 515982 183307 516016
rect 183377 515982 183411 516016
rect 184377 515982 184411 516016
rect 184481 516084 184515 516118
rect 184481 515982 184515 516016
rect 184929 516084 184963 516118
rect 184929 515982 184963 516016
rect 185217 515982 185251 516016
rect 186217 515982 186251 516016
rect 186321 516084 186355 516118
rect 186321 515982 186355 516016
rect 186953 516084 186987 516118
rect 186953 515982 186987 516016
rect 187241 516077 187275 516111
rect 187241 515982 187275 516016
rect 187413 516077 187447 516111
rect 187413 515982 187447 516016
rect 172245 515830 172279 515864
rect 172245 515735 172279 515769
rect 172417 515830 172451 515864
rect 172417 515735 172451 515769
rect 172521 515830 172555 515864
rect 172521 515728 172555 515762
rect 173153 515830 173187 515864
rect 173153 515728 173187 515762
rect 173441 515822 173475 515856
rect 173441 515700 173475 515734
rect 173527 515830 173561 515864
rect 173527 515762 173561 515796
rect 173623 515795 173657 515829
rect 173709 515830 173743 515864
rect 173795 515822 173829 515856
rect 173795 515754 173829 515788
rect 173795 515686 173829 515720
rect 173881 515816 173915 515850
rect 173881 515748 173915 515782
rect 173993 515830 174027 515864
rect 173993 515728 174027 515762
rect 174625 515830 174659 515864
rect 174625 515728 174659 515762
rect 174913 515830 174947 515864
rect 175913 515830 175947 515864
rect 176017 515830 176051 515864
rect 177017 515830 177051 515864
rect 177121 515830 177155 515864
rect 177121 515735 177155 515769
rect 177293 515830 177327 515864
rect 177293 515735 177327 515769
rect 177489 515830 177523 515864
rect 178489 515830 178523 515864
rect 178593 515830 178627 515864
rect 179593 515830 179627 515864
rect 179697 515830 179731 515864
rect 179697 515735 179731 515769
rect 179869 515830 179903 515864
rect 179869 515735 179903 515769
rect 180065 515830 180099 515864
rect 181065 515830 181099 515864
rect 181169 515830 181203 515864
rect 181169 515728 181203 515762
rect 181801 515830 181835 515864
rect 181801 515728 181835 515762
rect 182089 515822 182123 515856
rect 182089 515741 182123 515775
rect 182175 515822 182209 515856
rect 182175 515754 182209 515788
rect 182261 515822 182295 515856
rect 182261 515754 182295 515788
rect 182641 515830 182675 515864
rect 183641 515830 183675 515864
rect 183745 515830 183779 515864
rect 184745 515830 184779 515864
rect 184849 515830 184883 515864
rect 184849 515735 184883 515769
rect 185021 515830 185055 515864
rect 185021 515735 185055 515769
rect 185217 515830 185251 515864
rect 186217 515830 186251 515864
rect 186413 515822 186447 515856
rect 186413 515700 186447 515734
rect 186499 515830 186533 515864
rect 186499 515762 186533 515796
rect 186595 515795 186629 515829
rect 186681 515830 186715 515864
rect 186767 515822 186801 515856
rect 186767 515754 186801 515788
rect 186767 515686 186801 515720
rect 186853 515816 186887 515850
rect 186853 515748 186887 515782
rect 186965 515830 186999 515864
rect 186965 515735 186999 515769
rect 187137 515830 187171 515864
rect 187137 515735 187171 515769
rect 187241 515830 187275 515864
rect 187241 515735 187275 515769
rect 187413 515830 187447 515864
rect 187413 515735 187447 515769
<< psubdiff >>
rect 164520 541287 166650 541307
rect 164520 541277 164620 541287
rect 164520 539897 164540 541277
rect 164580 541247 164620 541277
rect 166540 541267 166650 541287
rect 166540 541247 166580 541267
rect 164580 541217 166580 541247
rect 164580 539947 164600 541217
rect 166560 539947 166580 541217
rect 164580 539927 166580 539947
rect 164580 539897 164620 539927
rect 164520 539887 164620 539897
rect 166540 539887 166580 539927
rect 166620 539887 166650 541267
rect 164520 539857 166650 539887
rect 168320 541287 170450 541307
rect 168320 541277 168420 541287
rect 168320 539897 168340 541277
rect 168380 541247 168420 541277
rect 170340 541267 170450 541287
rect 170340 541247 170380 541267
rect 168380 541217 170380 541247
rect 168380 539947 168400 541217
rect 170360 539947 170380 541217
rect 168380 539927 170380 539947
rect 168380 539897 168420 539927
rect 168320 539887 168420 539897
rect 170340 539887 170380 539927
rect 170420 539887 170450 541267
rect 168320 539857 170450 539887
rect 172020 541287 174150 541307
rect 172020 541277 172120 541287
rect 172020 539897 172040 541277
rect 172080 541247 172120 541277
rect 174040 541267 174150 541287
rect 174040 541247 174080 541267
rect 172080 541217 174080 541247
rect 172080 539947 172100 541217
rect 174060 539947 174080 541217
rect 172080 539927 174080 539947
rect 172080 539897 172120 539927
rect 172020 539887 172120 539897
rect 174040 539887 174080 539927
rect 174120 539887 174150 541267
rect 172020 539857 174150 539887
rect 175520 541287 177650 541307
rect 175520 541277 175620 541287
rect 175520 539897 175540 541277
rect 175580 541247 175620 541277
rect 177540 541267 177650 541287
rect 177540 541247 177580 541267
rect 175580 541217 177580 541247
rect 175580 539947 175600 541217
rect 177560 539947 177580 541217
rect 175580 539927 177580 539947
rect 175580 539897 175620 539927
rect 175520 539887 175620 539897
rect 177540 539887 177580 539927
rect 177620 539887 177650 541267
rect 175520 539857 177650 539887
rect 179120 541287 181250 541307
rect 179120 541277 179220 541287
rect 179120 539897 179140 541277
rect 179180 541247 179220 541277
rect 181140 541267 181250 541287
rect 181140 541247 181180 541267
rect 179180 541217 181180 541247
rect 179180 539947 179200 541217
rect 181160 539947 181180 541217
rect 179180 539927 181180 539947
rect 179180 539897 179220 539927
rect 179120 539887 179220 539897
rect 181140 539887 181180 539927
rect 181220 539887 181250 541267
rect 179120 539857 181250 539887
rect 182420 541287 184550 541307
rect 182420 541277 182520 541287
rect 182420 539897 182440 541277
rect 182480 541247 182520 541277
rect 184440 541267 184550 541287
rect 184440 541247 184480 541267
rect 182480 541217 184480 541247
rect 182480 539947 182500 541217
rect 184460 539947 184480 541217
rect 182480 539927 184480 539947
rect 182480 539897 182520 539927
rect 182420 539887 182520 539897
rect 184440 539887 184480 539927
rect 184520 539887 184550 541267
rect 182420 539857 184550 539887
rect 185720 541287 187850 541307
rect 185720 541277 185820 541287
rect 185720 539897 185740 541277
rect 185780 541247 185820 541277
rect 187740 541267 187850 541287
rect 187740 541247 187780 541267
rect 185780 541217 187780 541247
rect 185780 539947 185800 541217
rect 187760 539947 187780 541217
rect 185780 539927 187780 539947
rect 185780 539897 185820 539927
rect 185720 539887 185820 539897
rect 187740 539887 187780 539927
rect 187820 539887 187850 541267
rect 185720 539857 187850 539887
rect 189020 541287 191150 541307
rect 189020 541277 189120 541287
rect 189020 539897 189040 541277
rect 189080 541247 189120 541277
rect 191040 541267 191150 541287
rect 191040 541247 191080 541267
rect 189080 541217 191080 541247
rect 189080 539947 189100 541217
rect 191060 539947 191080 541217
rect 189080 539927 191080 539947
rect 189080 539897 189120 539927
rect 189020 539887 189120 539897
rect 191040 539887 191080 539927
rect 191120 539887 191150 541267
rect 191810 540277 191990 540301
rect 191810 540073 191990 540097
rect 189020 539857 191150 539887
rect 157630 538737 162870 538757
rect 157630 538697 157710 538737
rect 162770 538697 162870 538737
rect 157630 538677 162870 538697
rect 157630 538657 157710 538677
rect 157630 537997 157650 538657
rect 157690 538037 157710 538657
rect 162790 538037 162810 538677
rect 162850 538037 162870 538677
rect 157690 538017 162870 538037
rect 157690 537997 157730 538017
rect 157630 537977 157730 537997
rect 162770 537977 162870 538017
rect 157630 537957 162870 537977
rect 164188 538077 164284 538111
rect 166648 538077 166744 538111
rect 164188 538015 164222 538077
rect 166710 538015 166744 538077
rect 164188 535937 164222 535999
rect 166710 535937 166744 535999
rect 164188 535903 164284 535937
rect 166648 535903 166744 535937
rect 167960 538077 168056 538111
rect 169148 538077 169244 538111
rect 167960 538015 167994 538077
rect 169210 538015 169244 538077
rect 167960 535937 167994 535999
rect 169210 535937 169244 535999
rect 167960 535903 168056 535937
rect 169148 535903 169244 535937
rect 171696 538077 171792 538111
rect 172248 538077 172344 538111
rect 171696 538015 171730 538077
rect 172310 538015 172344 538077
rect 171696 535937 171730 535999
rect 172310 535937 172344 535999
rect 171696 535903 171792 535937
rect 172248 535903 172344 535937
rect 175214 538077 175310 538111
rect 175448 538077 175544 538111
rect 175214 538015 175248 538077
rect 175510 538015 175544 538077
rect 175214 535937 175248 535999
rect 178814 538077 178910 538111
rect 179048 538077 179144 538111
rect 178814 538015 178848 538077
rect 179110 538015 179144 538077
rect 178814 536497 178848 536559
rect 182114 538077 182210 538111
rect 182348 538077 182444 538111
rect 182114 538015 182148 538077
rect 182410 538015 182444 538077
rect 182114 536777 182148 536839
rect 185414 538077 185510 538111
rect 185648 538077 185744 538111
rect 185414 538015 185448 538077
rect 185710 538015 185744 538077
rect 185414 536917 185448 536979
rect 185710 536917 185744 536979
rect 185414 536883 185510 536917
rect 185648 536883 185744 536917
rect 188714 538077 188810 538111
rect 188948 538077 189044 538111
rect 188714 538015 188748 538077
rect 189010 538015 189044 538077
rect 182410 536777 182444 536839
rect 188714 536821 188748 536883
rect 189010 536821 189044 536883
rect 188714 536787 188810 536821
rect 188948 536787 189044 536821
rect 182114 536743 182210 536777
rect 182348 536743 182444 536777
rect 179110 536497 179144 536559
rect 178814 536463 178910 536497
rect 179048 536463 179144 536497
rect 175510 535937 175544 535999
rect 175214 535903 175310 535937
rect 175448 535903 175544 535937
rect 164158 535737 164254 535771
rect 166618 535737 166714 535771
rect 164158 535675 164192 535737
rect 166680 535675 166714 535737
rect 164158 533597 164192 533659
rect 166680 533597 166714 533659
rect 164158 533563 164254 533597
rect 166618 533563 166714 533597
rect 174815 530500 174849 530547
rect 174815 530442 174849 530466
rect 177391 530500 177425 530547
rect 177391 530442 177425 530466
rect 179967 530500 180001 530547
rect 179967 530442 180001 530466
rect 182543 530500 182577 530547
rect 182543 530442 182577 530466
rect 185119 530500 185153 530547
rect 185119 530442 185153 530466
rect 177391 529668 177425 529692
rect 177391 529587 177425 529634
rect 182543 529668 182577 529692
rect 182543 529587 182577 529634
rect 174815 529412 174849 529459
rect 174815 529354 174849 529378
rect 179967 529412 180001 529459
rect 179967 529354 180001 529378
rect 185119 529412 185153 529459
rect 185119 529354 185153 529378
rect 177391 528580 177425 528604
rect 177391 528499 177425 528546
rect 182543 528580 182577 528604
rect 182543 528499 182577 528546
rect 174815 528324 174849 528371
rect 174815 528266 174849 528290
rect 179967 528324 180001 528371
rect 179967 528266 180001 528290
rect 185119 528324 185153 528371
rect 185119 528266 185153 528290
rect 177391 527492 177425 527516
rect 177391 527411 177425 527458
rect 182543 527492 182577 527516
rect 182543 527411 182577 527458
rect 174815 527236 174849 527283
rect 174815 527178 174849 527202
rect 179967 527236 180001 527283
rect 179967 527178 180001 527202
rect 185119 527236 185153 527283
rect 185119 527178 185153 527202
rect 177391 526404 177425 526428
rect 177391 526323 177425 526370
rect 182543 526404 182577 526428
rect 182543 526323 182577 526370
rect 174815 526148 174849 526195
rect 174815 526090 174849 526114
rect 179967 526148 180001 526195
rect 179967 526090 180001 526114
rect 185119 526148 185153 526195
rect 185119 526090 185153 526114
rect 177391 525316 177425 525340
rect 177391 525235 177425 525282
rect 182543 525316 182577 525340
rect 182543 525235 182577 525282
rect 174815 525060 174849 525107
rect 174815 525002 174849 525026
rect 179967 525060 180001 525107
rect 179967 525002 180001 525026
rect 185119 525060 185153 525107
rect 185119 525002 185153 525026
rect 177391 524228 177425 524252
rect 177391 524147 177425 524194
rect 182543 524228 182577 524252
rect 182543 524147 182577 524194
rect 174815 523972 174849 524019
rect 174815 523914 174849 523938
rect 179967 523972 180001 524019
rect 179967 523914 180001 523938
rect 185119 523972 185153 524019
rect 185119 523914 185153 523938
rect 177391 523140 177425 523164
rect 177391 523059 177425 523106
rect 182543 523140 182577 523164
rect 182543 523059 182577 523106
rect 174815 522884 174849 522931
rect 174815 522826 174849 522850
rect 179967 522884 180001 522931
rect 179967 522826 180001 522850
rect 185119 522884 185153 522931
rect 185119 522826 185153 522850
rect 177391 522052 177425 522076
rect 177391 521971 177425 522018
rect 182543 522052 182577 522076
rect 182543 521971 182577 522018
rect 174815 521796 174849 521843
rect 174815 521738 174849 521762
rect 179967 521796 180001 521843
rect 179967 521738 180001 521762
rect 185119 521796 185153 521843
rect 185119 521738 185153 521762
rect 177391 520964 177425 520988
rect 177391 520883 177425 520930
rect 182543 520964 182577 520988
rect 182543 520883 182577 520930
rect 174815 520708 174849 520755
rect 174815 520650 174849 520674
rect 179967 520708 180001 520755
rect 179967 520650 180001 520674
rect 185119 520708 185153 520755
rect 185119 520650 185153 520674
rect 177391 519876 177425 519900
rect 177391 519795 177425 519842
rect 182543 519876 182577 519900
rect 182543 519795 182577 519842
rect 174815 519620 174849 519667
rect 174815 519562 174849 519586
rect 179967 519620 180001 519667
rect 179967 519562 180001 519586
rect 185119 519620 185153 519667
rect 185119 519562 185153 519586
rect 177391 518788 177425 518812
rect 177391 518707 177425 518754
rect 182543 518788 182577 518812
rect 182543 518707 182577 518754
rect 174815 518532 174849 518579
rect 174815 518474 174849 518498
rect 179967 518532 180001 518579
rect 179967 518474 180001 518498
rect 185119 518532 185153 518579
rect 185119 518474 185153 518498
rect 177391 517700 177425 517724
rect 177391 517619 177425 517666
rect 182543 517700 182577 517724
rect 182543 517619 182577 517666
rect 174815 517444 174849 517491
rect 174815 517386 174849 517410
rect 179967 517444 180001 517491
rect 179967 517386 180001 517410
rect 185119 517444 185153 517491
rect 185119 517386 185153 517410
rect 177391 516612 177425 516636
rect 177391 516531 177425 516578
rect 182543 516612 182577 516636
rect 182543 516531 182577 516578
rect 174815 516356 174849 516403
rect 174815 516298 174849 516322
rect 179967 516356 180001 516403
rect 179967 516298 180001 516322
rect 185119 516356 185153 516403
rect 185119 516298 185153 516322
rect 174815 515524 174849 515548
rect 174815 515443 174849 515490
rect 177391 515524 177425 515548
rect 177391 515443 177425 515490
rect 179967 515524 180001 515548
rect 179967 515443 180001 515490
rect 182543 515524 182577 515548
rect 182543 515443 182577 515490
rect 185119 515524 185153 515548
rect 185119 515443 185153 515490
<< nsubdiff >>
rect 164520 539767 166640 539787
rect 164520 539747 164620 539767
rect 164520 538347 164540 539747
rect 164580 539727 164620 539747
rect 166540 539747 166640 539767
rect 166540 539727 166580 539747
rect 164580 539707 166580 539727
rect 164580 538387 164600 539707
rect 166540 539687 166580 539707
rect 166560 538387 166580 539687
rect 164580 538367 166580 538387
rect 164580 538347 164620 538367
rect 164520 538327 164620 538347
rect 166540 538347 166580 538367
rect 166620 538347 166640 539747
rect 166540 538327 166640 538347
rect 164520 538307 166640 538327
rect 168320 539767 170440 539787
rect 168320 539747 168420 539767
rect 168320 538347 168340 539747
rect 168380 539727 168420 539747
rect 170340 539747 170440 539767
rect 170340 539727 170380 539747
rect 168380 539707 170380 539727
rect 168380 538387 168400 539707
rect 170340 539687 170380 539707
rect 170360 538387 170380 539687
rect 168380 538367 170380 538387
rect 168380 538347 168420 538367
rect 168320 538327 168420 538347
rect 170340 538347 170380 538367
rect 170420 538347 170440 539747
rect 170340 538327 170440 538347
rect 168320 538307 170440 538327
rect 172020 539767 174140 539787
rect 172020 539747 172120 539767
rect 172020 538347 172040 539747
rect 172080 539727 172120 539747
rect 174040 539747 174140 539767
rect 174040 539727 174080 539747
rect 172080 539707 174080 539727
rect 172080 538387 172100 539707
rect 174040 539687 174080 539707
rect 174060 538387 174080 539687
rect 172080 538367 174080 538387
rect 172080 538347 172120 538367
rect 172020 538327 172120 538347
rect 174040 538347 174080 538367
rect 174120 538347 174140 539747
rect 174040 538327 174140 538347
rect 172020 538307 174140 538327
rect 175520 539767 177640 539787
rect 175520 539747 175620 539767
rect 175520 538347 175540 539747
rect 175580 539727 175620 539747
rect 177540 539747 177640 539767
rect 177540 539727 177580 539747
rect 175580 539707 177580 539727
rect 175580 538387 175600 539707
rect 177540 539687 177580 539707
rect 177560 538387 177580 539687
rect 175580 538367 177580 538387
rect 175580 538347 175620 538367
rect 175520 538327 175620 538347
rect 177540 538347 177580 538367
rect 177620 538347 177640 539747
rect 177540 538327 177640 538347
rect 175520 538307 177640 538327
rect 179120 539767 181240 539787
rect 179120 539747 179220 539767
rect 179120 538347 179140 539747
rect 179180 539727 179220 539747
rect 181140 539747 181240 539767
rect 181140 539727 181180 539747
rect 179180 539707 181180 539727
rect 179180 538387 179200 539707
rect 181140 539687 181180 539707
rect 181160 538387 181180 539687
rect 179180 538367 181180 538387
rect 179180 538347 179220 538367
rect 179120 538327 179220 538347
rect 181140 538347 181180 538367
rect 181220 538347 181240 539747
rect 181140 538327 181240 538347
rect 179120 538307 181240 538327
rect 182420 539767 184540 539787
rect 182420 539747 182520 539767
rect 182420 538347 182440 539747
rect 182480 539727 182520 539747
rect 184440 539747 184540 539767
rect 184440 539727 184480 539747
rect 182480 539707 184480 539727
rect 182480 538387 182500 539707
rect 184440 539687 184480 539707
rect 184460 538387 184480 539687
rect 182480 538367 184480 538387
rect 182480 538347 182520 538367
rect 182420 538327 182520 538347
rect 184440 538347 184480 538367
rect 184520 538347 184540 539747
rect 184440 538327 184540 538347
rect 182420 538307 184540 538327
rect 185720 539767 187840 539787
rect 185720 539747 185820 539767
rect 185720 538347 185740 539747
rect 185780 539727 185820 539747
rect 187740 539747 187840 539767
rect 187740 539727 187780 539747
rect 185780 539707 187780 539727
rect 185780 538387 185800 539707
rect 187740 539687 187780 539707
rect 187760 538387 187780 539687
rect 185780 538367 187780 538387
rect 185780 538347 185820 538367
rect 185720 538327 185820 538347
rect 187740 538347 187780 538367
rect 187820 538347 187840 539747
rect 187740 538327 187840 538347
rect 185720 538307 187840 538327
rect 189020 539767 191140 539787
rect 189020 539747 189120 539767
rect 189020 538347 189040 539747
rect 189080 539727 189120 539747
rect 191040 539747 191140 539767
rect 191040 539727 191080 539747
rect 189080 539707 191080 539727
rect 189080 538387 189100 539707
rect 191040 539687 191080 539707
rect 191060 538387 191080 539687
rect 189080 538367 191080 538387
rect 189080 538347 189120 538367
rect 189020 538327 189120 538347
rect 191040 538347 191080 538367
rect 191120 538347 191140 539747
rect 191040 538327 191140 538347
rect 189020 538307 191140 538327
rect 157590 537857 162850 537877
rect 157590 537817 157650 537857
rect 162750 537817 162850 537857
rect 157590 537797 162790 537817
rect 157590 537757 157670 537797
rect 157590 535817 157610 537757
rect 157650 535817 157670 537757
rect 157590 535797 157670 535817
rect 162770 535797 162790 537797
rect 162830 535797 162850 537817
rect 157590 535777 162850 535797
rect 157590 535737 157670 535777
rect 162750 535737 162850 535777
rect 157590 535717 162850 535737
rect 174815 530282 174849 530306
rect 174815 530189 174849 530248
rect 174815 530131 174849 530155
rect 177391 530282 177425 530306
rect 177391 530189 177425 530248
rect 177391 530131 177425 530155
rect 179967 530282 180001 530306
rect 179967 530189 180001 530248
rect 179967 530131 180001 530155
rect 182543 530282 182577 530306
rect 182543 530189 182577 530248
rect 182543 530131 182577 530155
rect 185119 530282 185153 530306
rect 185119 530189 185153 530248
rect 185119 530131 185153 530155
rect 177391 529979 177425 530003
rect 177391 529886 177425 529945
rect 177391 529828 177425 529852
rect 182543 529979 182577 530003
rect 182543 529886 182577 529945
rect 182543 529828 182577 529852
rect 174815 529194 174849 529218
rect 174815 529101 174849 529160
rect 174815 529043 174849 529067
rect 179967 529194 180001 529218
rect 179967 529101 180001 529160
rect 179967 529043 180001 529067
rect 185119 529194 185153 529218
rect 185119 529101 185153 529160
rect 185119 529043 185153 529067
rect 177391 528891 177425 528915
rect 177391 528798 177425 528857
rect 177391 528740 177425 528764
rect 182543 528891 182577 528915
rect 182543 528798 182577 528857
rect 182543 528740 182577 528764
rect 174815 528106 174849 528130
rect 174815 528013 174849 528072
rect 174815 527955 174849 527979
rect 179967 528106 180001 528130
rect 179967 528013 180001 528072
rect 179967 527955 180001 527979
rect 185119 528106 185153 528130
rect 185119 528013 185153 528072
rect 185119 527955 185153 527979
rect 177391 527803 177425 527827
rect 177391 527710 177425 527769
rect 177391 527652 177425 527676
rect 182543 527803 182577 527827
rect 182543 527710 182577 527769
rect 182543 527652 182577 527676
rect 174815 527018 174849 527042
rect 174815 526925 174849 526984
rect 174815 526867 174849 526891
rect 179967 527018 180001 527042
rect 179967 526925 180001 526984
rect 179967 526867 180001 526891
rect 185119 527018 185153 527042
rect 185119 526925 185153 526984
rect 185119 526867 185153 526891
rect 177391 526715 177425 526739
rect 177391 526622 177425 526681
rect 177391 526564 177425 526588
rect 182543 526715 182577 526739
rect 182543 526622 182577 526681
rect 182543 526564 182577 526588
rect 174815 525930 174849 525954
rect 174815 525837 174849 525896
rect 174815 525779 174849 525803
rect 179967 525930 180001 525954
rect 179967 525837 180001 525896
rect 179967 525779 180001 525803
rect 185119 525930 185153 525954
rect 185119 525837 185153 525896
rect 185119 525779 185153 525803
rect 177391 525627 177425 525651
rect 177391 525534 177425 525593
rect 177391 525476 177425 525500
rect 182543 525627 182577 525651
rect 182543 525534 182577 525593
rect 182543 525476 182577 525500
rect 174815 524842 174849 524866
rect 174815 524749 174849 524808
rect 174815 524691 174849 524715
rect 179967 524842 180001 524866
rect 179967 524749 180001 524808
rect 179967 524691 180001 524715
rect 185119 524842 185153 524866
rect 185119 524749 185153 524808
rect 185119 524691 185153 524715
rect 177391 524539 177425 524563
rect 177391 524446 177425 524505
rect 177391 524388 177425 524412
rect 182543 524539 182577 524563
rect 182543 524446 182577 524505
rect 182543 524388 182577 524412
rect 174815 523754 174849 523778
rect 174815 523661 174849 523720
rect 174815 523603 174849 523627
rect 179967 523754 180001 523778
rect 179967 523661 180001 523720
rect 179967 523603 180001 523627
rect 185119 523754 185153 523778
rect 185119 523661 185153 523720
rect 185119 523603 185153 523627
rect 177391 523451 177425 523475
rect 177391 523358 177425 523417
rect 177391 523300 177425 523324
rect 182543 523451 182577 523475
rect 182543 523358 182577 523417
rect 182543 523300 182577 523324
rect 174815 522666 174849 522690
rect 174815 522573 174849 522632
rect 174815 522515 174849 522539
rect 179967 522666 180001 522690
rect 179967 522573 180001 522632
rect 179967 522515 180001 522539
rect 185119 522666 185153 522690
rect 185119 522573 185153 522632
rect 185119 522515 185153 522539
rect 177391 522363 177425 522387
rect 177391 522270 177425 522329
rect 177391 522212 177425 522236
rect 182543 522363 182577 522387
rect 182543 522270 182577 522329
rect 182543 522212 182577 522236
rect 174815 521578 174849 521602
rect 174815 521485 174849 521544
rect 174815 521427 174849 521451
rect 179967 521578 180001 521602
rect 179967 521485 180001 521544
rect 179967 521427 180001 521451
rect 185119 521578 185153 521602
rect 185119 521485 185153 521544
rect 185119 521427 185153 521451
rect 177391 521275 177425 521299
rect 177391 521182 177425 521241
rect 177391 521124 177425 521148
rect 182543 521275 182577 521299
rect 182543 521182 182577 521241
rect 182543 521124 182577 521148
rect 174815 520490 174849 520514
rect 174815 520397 174849 520456
rect 174815 520339 174849 520363
rect 179967 520490 180001 520514
rect 179967 520397 180001 520456
rect 179967 520339 180001 520363
rect 185119 520490 185153 520514
rect 185119 520397 185153 520456
rect 185119 520339 185153 520363
rect 177391 520187 177425 520211
rect 177391 520094 177425 520153
rect 177391 520036 177425 520060
rect 182543 520187 182577 520211
rect 182543 520094 182577 520153
rect 182543 520036 182577 520060
rect 174815 519402 174849 519426
rect 174815 519309 174849 519368
rect 174815 519251 174849 519275
rect 179967 519402 180001 519426
rect 179967 519309 180001 519368
rect 179967 519251 180001 519275
rect 185119 519402 185153 519426
rect 185119 519309 185153 519368
rect 185119 519251 185153 519275
rect 177391 519099 177425 519123
rect 177391 519006 177425 519065
rect 177391 518948 177425 518972
rect 182543 519099 182577 519123
rect 182543 519006 182577 519065
rect 182543 518948 182577 518972
rect 174815 518314 174849 518338
rect 174815 518221 174849 518280
rect 174815 518163 174849 518187
rect 179967 518314 180001 518338
rect 179967 518221 180001 518280
rect 179967 518163 180001 518187
rect 185119 518314 185153 518338
rect 185119 518221 185153 518280
rect 185119 518163 185153 518187
rect 177391 518011 177425 518035
rect 177391 517918 177425 517977
rect 177391 517860 177425 517884
rect 182543 518011 182577 518035
rect 182543 517918 182577 517977
rect 182543 517860 182577 517884
rect 174815 517226 174849 517250
rect 174815 517133 174849 517192
rect 174815 517075 174849 517099
rect 179967 517226 180001 517250
rect 179967 517133 180001 517192
rect 179967 517075 180001 517099
rect 185119 517226 185153 517250
rect 185119 517133 185153 517192
rect 185119 517075 185153 517099
rect 177391 516923 177425 516947
rect 177391 516830 177425 516889
rect 177391 516772 177425 516796
rect 182543 516923 182577 516947
rect 182543 516830 182577 516889
rect 182543 516772 182577 516796
rect 174815 516138 174849 516162
rect 174815 516045 174849 516104
rect 174815 515987 174849 516011
rect 179967 516138 180001 516162
rect 179967 516045 180001 516104
rect 179967 515987 180001 516011
rect 185119 516138 185153 516162
rect 185119 516045 185153 516104
rect 185119 515987 185153 516011
rect 174815 515835 174849 515859
rect 174815 515742 174849 515801
rect 174815 515684 174849 515708
rect 177391 515835 177425 515859
rect 177391 515742 177425 515801
rect 177391 515684 177425 515708
rect 179967 515835 180001 515859
rect 179967 515742 180001 515801
rect 179967 515684 180001 515708
rect 182543 515835 182577 515859
rect 182543 515742 182577 515801
rect 182543 515684 182577 515708
rect 185119 515835 185153 515859
rect 185119 515742 185153 515801
rect 185119 515684 185153 515708
<< psubdiffcont >>
rect 164540 539897 164580 541277
rect 164620 541247 166540 541287
rect 164620 539887 166540 539927
rect 166580 539887 166620 541267
rect 168340 539897 168380 541277
rect 168420 541247 170340 541287
rect 168420 539887 170340 539927
rect 170380 539887 170420 541267
rect 172040 539897 172080 541277
rect 172120 541247 174040 541287
rect 172120 539887 174040 539927
rect 174080 539887 174120 541267
rect 175540 539897 175580 541277
rect 175620 541247 177540 541287
rect 175620 539887 177540 539927
rect 177580 539887 177620 541267
rect 179140 539897 179180 541277
rect 179220 541247 181140 541287
rect 179220 539887 181140 539927
rect 181180 539887 181220 541267
rect 182440 539897 182480 541277
rect 182520 541247 184440 541287
rect 182520 539887 184440 539927
rect 184480 539887 184520 541267
rect 185740 539897 185780 541277
rect 185820 541247 187740 541287
rect 185820 539887 187740 539927
rect 187780 539887 187820 541267
rect 189040 539897 189080 541277
rect 189120 541247 191040 541287
rect 189120 539887 191040 539927
rect 191080 539887 191120 541267
rect 191810 540097 191990 540277
rect 157710 538697 162770 538737
rect 157650 537997 157690 538657
rect 162810 538037 162850 538677
rect 157730 537977 162770 538017
rect 164284 538077 166648 538111
rect 164188 535999 164222 538015
rect 166710 535999 166744 538015
rect 164284 535903 166648 535937
rect 168056 538077 169148 538111
rect 167960 535999 167994 538015
rect 169210 535999 169244 538015
rect 168056 535903 169148 535937
rect 171792 538077 172248 538111
rect 171696 535999 171730 538015
rect 172310 535999 172344 538015
rect 171792 535903 172248 535937
rect 175310 538077 175448 538111
rect 175214 535999 175248 538015
rect 175510 535999 175544 538015
rect 178910 538077 179048 538111
rect 178814 536559 178848 538015
rect 179110 536559 179144 538015
rect 182210 538077 182348 538111
rect 182114 536839 182148 538015
rect 182410 536839 182444 538015
rect 185510 538077 185648 538111
rect 185414 536979 185448 538015
rect 185710 536979 185744 538015
rect 185510 536883 185648 536917
rect 188810 538077 188948 538111
rect 188714 536883 188748 538015
rect 189010 536883 189044 538015
rect 188810 536787 188948 536821
rect 182210 536743 182348 536777
rect 178910 536463 179048 536497
rect 175310 535903 175448 535937
rect 164254 535737 166618 535771
rect 164158 533659 164192 535675
rect 166680 533659 166714 535675
rect 164254 533563 166618 533597
rect 174815 530466 174849 530500
rect 177391 530466 177425 530500
rect 179967 530466 180001 530500
rect 182543 530466 182577 530500
rect 185119 530466 185153 530500
rect 177391 529634 177425 529668
rect 182543 529634 182577 529668
rect 174815 529378 174849 529412
rect 179967 529378 180001 529412
rect 185119 529378 185153 529412
rect 177391 528546 177425 528580
rect 182543 528546 182577 528580
rect 174815 528290 174849 528324
rect 179967 528290 180001 528324
rect 185119 528290 185153 528324
rect 177391 527458 177425 527492
rect 182543 527458 182577 527492
rect 174815 527202 174849 527236
rect 179967 527202 180001 527236
rect 185119 527202 185153 527236
rect 177391 526370 177425 526404
rect 182543 526370 182577 526404
rect 174815 526114 174849 526148
rect 179967 526114 180001 526148
rect 185119 526114 185153 526148
rect 177391 525282 177425 525316
rect 182543 525282 182577 525316
rect 174815 525026 174849 525060
rect 179967 525026 180001 525060
rect 185119 525026 185153 525060
rect 177391 524194 177425 524228
rect 182543 524194 182577 524228
rect 174815 523938 174849 523972
rect 179967 523938 180001 523972
rect 185119 523938 185153 523972
rect 177391 523106 177425 523140
rect 182543 523106 182577 523140
rect 174815 522850 174849 522884
rect 179967 522850 180001 522884
rect 185119 522850 185153 522884
rect 177391 522018 177425 522052
rect 182543 522018 182577 522052
rect 174815 521762 174849 521796
rect 179967 521762 180001 521796
rect 185119 521762 185153 521796
rect 177391 520930 177425 520964
rect 182543 520930 182577 520964
rect 174815 520674 174849 520708
rect 179967 520674 180001 520708
rect 185119 520674 185153 520708
rect 177391 519842 177425 519876
rect 182543 519842 182577 519876
rect 174815 519586 174849 519620
rect 179967 519586 180001 519620
rect 185119 519586 185153 519620
rect 177391 518754 177425 518788
rect 182543 518754 182577 518788
rect 174815 518498 174849 518532
rect 179967 518498 180001 518532
rect 185119 518498 185153 518532
rect 177391 517666 177425 517700
rect 182543 517666 182577 517700
rect 174815 517410 174849 517444
rect 179967 517410 180001 517444
rect 185119 517410 185153 517444
rect 177391 516578 177425 516612
rect 182543 516578 182577 516612
rect 174815 516322 174849 516356
rect 179967 516322 180001 516356
rect 185119 516322 185153 516356
rect 174815 515490 174849 515524
rect 177391 515490 177425 515524
rect 179967 515490 180001 515524
rect 182543 515490 182577 515524
rect 185119 515490 185153 515524
<< nsubdiffcont >>
rect 164540 538347 164580 539747
rect 164620 539727 166540 539767
rect 164620 538327 166540 538367
rect 166580 538347 166620 539747
rect 168340 538347 168380 539747
rect 168420 539727 170340 539767
rect 168420 538327 170340 538367
rect 170380 538347 170420 539747
rect 172040 538347 172080 539747
rect 172120 539727 174040 539767
rect 172120 538327 174040 538367
rect 174080 538347 174120 539747
rect 175540 538347 175580 539747
rect 175620 539727 177540 539767
rect 175620 538327 177540 538367
rect 177580 538347 177620 539747
rect 179140 538347 179180 539747
rect 179220 539727 181140 539767
rect 179220 538327 181140 538367
rect 181180 538347 181220 539747
rect 182440 538347 182480 539747
rect 182520 539727 184440 539767
rect 182520 538327 184440 538367
rect 184480 538347 184520 539747
rect 185740 538347 185780 539747
rect 185820 539727 187740 539767
rect 185820 538327 187740 538367
rect 187780 538347 187820 539747
rect 189040 538347 189080 539747
rect 189120 539727 191040 539767
rect 189120 538327 191040 538367
rect 191080 538347 191120 539747
rect 157650 537817 162750 537857
rect 157610 535817 157650 537757
rect 162790 535797 162830 537817
rect 157670 535737 162750 535777
rect 174815 530248 174849 530282
rect 174815 530155 174849 530189
rect 177391 530248 177425 530282
rect 177391 530155 177425 530189
rect 179967 530248 180001 530282
rect 179967 530155 180001 530189
rect 182543 530248 182577 530282
rect 182543 530155 182577 530189
rect 185119 530248 185153 530282
rect 185119 530155 185153 530189
rect 177391 529945 177425 529979
rect 177391 529852 177425 529886
rect 182543 529945 182577 529979
rect 182543 529852 182577 529886
rect 174815 529160 174849 529194
rect 174815 529067 174849 529101
rect 179967 529160 180001 529194
rect 179967 529067 180001 529101
rect 185119 529160 185153 529194
rect 185119 529067 185153 529101
rect 177391 528857 177425 528891
rect 177391 528764 177425 528798
rect 182543 528857 182577 528891
rect 182543 528764 182577 528798
rect 174815 528072 174849 528106
rect 174815 527979 174849 528013
rect 179967 528072 180001 528106
rect 179967 527979 180001 528013
rect 185119 528072 185153 528106
rect 185119 527979 185153 528013
rect 177391 527769 177425 527803
rect 177391 527676 177425 527710
rect 182543 527769 182577 527803
rect 182543 527676 182577 527710
rect 174815 526984 174849 527018
rect 174815 526891 174849 526925
rect 179967 526984 180001 527018
rect 179967 526891 180001 526925
rect 185119 526984 185153 527018
rect 185119 526891 185153 526925
rect 177391 526681 177425 526715
rect 177391 526588 177425 526622
rect 182543 526681 182577 526715
rect 182543 526588 182577 526622
rect 174815 525896 174849 525930
rect 174815 525803 174849 525837
rect 179967 525896 180001 525930
rect 179967 525803 180001 525837
rect 185119 525896 185153 525930
rect 185119 525803 185153 525837
rect 177391 525593 177425 525627
rect 177391 525500 177425 525534
rect 182543 525593 182577 525627
rect 182543 525500 182577 525534
rect 174815 524808 174849 524842
rect 174815 524715 174849 524749
rect 179967 524808 180001 524842
rect 179967 524715 180001 524749
rect 185119 524808 185153 524842
rect 185119 524715 185153 524749
rect 177391 524505 177425 524539
rect 177391 524412 177425 524446
rect 182543 524505 182577 524539
rect 182543 524412 182577 524446
rect 174815 523720 174849 523754
rect 174815 523627 174849 523661
rect 179967 523720 180001 523754
rect 179967 523627 180001 523661
rect 185119 523720 185153 523754
rect 185119 523627 185153 523661
rect 177391 523417 177425 523451
rect 177391 523324 177425 523358
rect 182543 523417 182577 523451
rect 182543 523324 182577 523358
rect 174815 522632 174849 522666
rect 174815 522539 174849 522573
rect 179967 522632 180001 522666
rect 179967 522539 180001 522573
rect 185119 522632 185153 522666
rect 185119 522539 185153 522573
rect 177391 522329 177425 522363
rect 177391 522236 177425 522270
rect 182543 522329 182577 522363
rect 182543 522236 182577 522270
rect 174815 521544 174849 521578
rect 174815 521451 174849 521485
rect 179967 521544 180001 521578
rect 179967 521451 180001 521485
rect 185119 521544 185153 521578
rect 185119 521451 185153 521485
rect 177391 521241 177425 521275
rect 177391 521148 177425 521182
rect 182543 521241 182577 521275
rect 182543 521148 182577 521182
rect 174815 520456 174849 520490
rect 174815 520363 174849 520397
rect 179967 520456 180001 520490
rect 179967 520363 180001 520397
rect 185119 520456 185153 520490
rect 185119 520363 185153 520397
rect 177391 520153 177425 520187
rect 177391 520060 177425 520094
rect 182543 520153 182577 520187
rect 182543 520060 182577 520094
rect 174815 519368 174849 519402
rect 174815 519275 174849 519309
rect 179967 519368 180001 519402
rect 179967 519275 180001 519309
rect 185119 519368 185153 519402
rect 185119 519275 185153 519309
rect 177391 519065 177425 519099
rect 177391 518972 177425 519006
rect 182543 519065 182577 519099
rect 182543 518972 182577 519006
rect 174815 518280 174849 518314
rect 174815 518187 174849 518221
rect 179967 518280 180001 518314
rect 179967 518187 180001 518221
rect 185119 518280 185153 518314
rect 185119 518187 185153 518221
rect 177391 517977 177425 518011
rect 177391 517884 177425 517918
rect 182543 517977 182577 518011
rect 182543 517884 182577 517918
rect 174815 517192 174849 517226
rect 174815 517099 174849 517133
rect 179967 517192 180001 517226
rect 179967 517099 180001 517133
rect 185119 517192 185153 517226
rect 185119 517099 185153 517133
rect 177391 516889 177425 516923
rect 177391 516796 177425 516830
rect 182543 516889 182577 516923
rect 182543 516796 182577 516830
rect 174815 516104 174849 516138
rect 174815 516011 174849 516045
rect 179967 516104 180001 516138
rect 179967 516011 180001 516045
rect 185119 516104 185153 516138
rect 185119 516011 185153 516045
rect 174815 515801 174849 515835
rect 174815 515708 174849 515742
rect 177391 515801 177425 515835
rect 177391 515708 177425 515742
rect 179967 515801 180001 515835
rect 179967 515708 180001 515742
rect 182543 515801 182577 515835
rect 182543 515708 182577 515742
rect 185119 515801 185153 515835
rect 185119 515708 185153 515742
<< poly >>
rect 164940 541174 166030 541177
rect 164940 541167 166043 541174
rect 164714 541151 164780 541167
rect 164714 541117 164730 541151
rect 164764 541117 164780 541151
rect 164714 541101 164780 541117
rect 164939 541158 166043 541167
rect 164939 541124 165033 541158
rect 165067 541124 165225 541158
rect 165259 541124 165417 541158
rect 165451 541124 165609 541158
rect 165643 541124 165801 541158
rect 165835 541124 165993 541158
rect 166027 541124 166043 541158
rect 164939 541117 166043 541124
rect 164732 541079 164762 541101
rect 164939 541086 164969 541117
rect 165017 541108 166043 541117
rect 166394 541151 166460 541167
rect 166394 541117 166410 541151
rect 166444 541117 166460 541151
rect 165034 541107 166030 541108
rect 165035 541086 165065 541107
rect 165131 541086 165161 541107
rect 165227 541086 165257 541107
rect 165323 541086 165353 541107
rect 165419 541086 165449 541107
rect 165515 541086 165545 541107
rect 165611 541086 165641 541107
rect 165707 541086 165737 541107
rect 165803 541086 165833 541107
rect 165899 541086 165929 541107
rect 165995 541086 166025 541107
rect 166394 541101 166460 541117
rect 166412 541079 166442 541101
rect 166194 540351 166260 540367
rect 166194 540317 166210 540351
rect 166244 540317 166260 540351
rect 166194 540301 166260 540317
rect 166212 540279 166242 540301
rect 164732 540057 164762 540079
rect 164939 540064 164969 540086
rect 164714 540041 164780 540057
rect 164714 540007 164730 540041
rect 164764 540007 164780 540041
rect 164714 539991 164780 540007
rect 164921 540048 164987 540064
rect 165035 540060 165065 540086
rect 165131 540064 165161 540086
rect 164921 540014 164937 540048
rect 164971 540014 164987 540048
rect 164921 539998 164987 540014
rect 165113 540048 165179 540064
rect 165227 540060 165257 540086
rect 165323 540064 165353 540086
rect 165113 540014 165129 540048
rect 165163 540014 165179 540048
rect 165113 539998 165179 540014
rect 165305 540048 165371 540064
rect 165419 540060 165449 540086
rect 165515 540064 165545 540086
rect 165305 540014 165321 540048
rect 165355 540014 165371 540048
rect 165305 539998 165371 540014
rect 165497 540048 165563 540064
rect 165611 540060 165641 540086
rect 165707 540064 165737 540086
rect 165497 540014 165513 540048
rect 165547 540014 165563 540048
rect 165497 539998 165563 540014
rect 165689 540048 165755 540064
rect 165803 540060 165833 540086
rect 165899 540064 165929 540086
rect 165689 540014 165705 540048
rect 165739 540014 165755 540048
rect 165689 539998 165755 540014
rect 165881 540048 165947 540064
rect 165995 540060 166025 540086
rect 166212 540057 166242 540079
rect 166412 540057 166442 540079
rect 165881 540014 165897 540048
rect 165931 540014 165947 540048
rect 165881 539998 165947 540014
rect 166194 540041 166260 540057
rect 166194 540007 166210 540041
rect 166244 540007 166260 540041
rect 166194 539991 166260 540007
rect 166394 540041 166460 540057
rect 166394 540007 166410 540041
rect 166444 540007 166460 540041
rect 166394 539991 166460 540007
rect 168740 541174 169830 541177
rect 168740 541167 169843 541174
rect 168514 541151 168580 541167
rect 168514 541117 168530 541151
rect 168564 541117 168580 541151
rect 168514 541101 168580 541117
rect 168739 541158 169843 541167
rect 168739 541124 168833 541158
rect 168867 541124 169025 541158
rect 169059 541124 169217 541158
rect 169251 541124 169409 541158
rect 169443 541124 169601 541158
rect 169635 541124 169793 541158
rect 169827 541124 169843 541158
rect 168739 541117 169843 541124
rect 168532 541079 168562 541101
rect 168739 541086 168769 541117
rect 168817 541108 169843 541117
rect 170194 541151 170260 541167
rect 170194 541117 170210 541151
rect 170244 541117 170260 541151
rect 168834 541107 169830 541108
rect 168835 541086 168865 541107
rect 168931 541086 168961 541107
rect 169027 541086 169057 541107
rect 169123 541086 169153 541107
rect 169219 541086 169249 541107
rect 169315 541086 169345 541107
rect 169411 541086 169441 541107
rect 169507 541086 169537 541107
rect 169603 541086 169633 541107
rect 169699 541086 169729 541107
rect 169795 541086 169825 541107
rect 170194 541101 170260 541117
rect 170212 541079 170242 541101
rect 169994 540351 170060 540367
rect 169994 540317 170010 540351
rect 170044 540317 170060 540351
rect 169994 540301 170060 540317
rect 170012 540279 170042 540301
rect 168532 540057 168562 540079
rect 168739 540064 168769 540086
rect 168514 540041 168580 540057
rect 168514 540007 168530 540041
rect 168564 540007 168580 540041
rect 168514 539991 168580 540007
rect 168721 540048 168787 540064
rect 168835 540060 168865 540086
rect 168931 540064 168961 540086
rect 168721 540014 168737 540048
rect 168771 540014 168787 540048
rect 168721 539998 168787 540014
rect 168913 540048 168979 540064
rect 169027 540060 169057 540086
rect 169123 540064 169153 540086
rect 168913 540014 168929 540048
rect 168963 540014 168979 540048
rect 168913 539998 168979 540014
rect 169105 540048 169171 540064
rect 169219 540060 169249 540086
rect 169315 540064 169345 540086
rect 169105 540014 169121 540048
rect 169155 540014 169171 540048
rect 169105 539998 169171 540014
rect 169297 540048 169363 540064
rect 169411 540060 169441 540086
rect 169507 540064 169537 540086
rect 169297 540014 169313 540048
rect 169347 540014 169363 540048
rect 169297 539998 169363 540014
rect 169489 540048 169555 540064
rect 169603 540060 169633 540086
rect 169699 540064 169729 540086
rect 169489 540014 169505 540048
rect 169539 540014 169555 540048
rect 169489 539998 169555 540014
rect 169681 540048 169747 540064
rect 169795 540060 169825 540086
rect 170012 540057 170042 540079
rect 170212 540057 170242 540079
rect 169681 540014 169697 540048
rect 169731 540014 169747 540048
rect 169681 539998 169747 540014
rect 169994 540041 170060 540057
rect 169994 540007 170010 540041
rect 170044 540007 170060 540041
rect 169994 539991 170060 540007
rect 170194 540041 170260 540057
rect 170194 540007 170210 540041
rect 170244 540007 170260 540041
rect 170194 539991 170260 540007
rect 172440 541174 173530 541177
rect 172440 541167 173543 541174
rect 172214 541151 172280 541167
rect 172214 541117 172230 541151
rect 172264 541117 172280 541151
rect 172214 541101 172280 541117
rect 172439 541158 173543 541167
rect 172439 541124 172533 541158
rect 172567 541124 172725 541158
rect 172759 541124 172917 541158
rect 172951 541124 173109 541158
rect 173143 541124 173301 541158
rect 173335 541124 173493 541158
rect 173527 541124 173543 541158
rect 172439 541117 173543 541124
rect 172232 541079 172262 541101
rect 172439 541086 172469 541117
rect 172517 541108 173543 541117
rect 173894 541151 173960 541167
rect 173894 541117 173910 541151
rect 173944 541117 173960 541151
rect 172534 541107 173530 541108
rect 172535 541086 172565 541107
rect 172631 541086 172661 541107
rect 172727 541086 172757 541107
rect 172823 541086 172853 541107
rect 172919 541086 172949 541107
rect 173015 541086 173045 541107
rect 173111 541086 173141 541107
rect 173207 541086 173237 541107
rect 173303 541086 173333 541107
rect 173399 541086 173429 541107
rect 173495 541086 173525 541107
rect 173894 541101 173960 541117
rect 173912 541079 173942 541101
rect 173694 540351 173760 540367
rect 173694 540317 173710 540351
rect 173744 540317 173760 540351
rect 173694 540301 173760 540317
rect 173712 540279 173742 540301
rect 172232 540057 172262 540079
rect 172439 540064 172469 540086
rect 172214 540041 172280 540057
rect 172214 540007 172230 540041
rect 172264 540007 172280 540041
rect 172214 539991 172280 540007
rect 172421 540048 172487 540064
rect 172535 540060 172565 540086
rect 172631 540064 172661 540086
rect 172421 540014 172437 540048
rect 172471 540014 172487 540048
rect 172421 539998 172487 540014
rect 172613 540048 172679 540064
rect 172727 540060 172757 540086
rect 172823 540064 172853 540086
rect 172613 540014 172629 540048
rect 172663 540014 172679 540048
rect 172613 539998 172679 540014
rect 172805 540048 172871 540064
rect 172919 540060 172949 540086
rect 173015 540064 173045 540086
rect 172805 540014 172821 540048
rect 172855 540014 172871 540048
rect 172805 539998 172871 540014
rect 172997 540048 173063 540064
rect 173111 540060 173141 540086
rect 173207 540064 173237 540086
rect 172997 540014 173013 540048
rect 173047 540014 173063 540048
rect 172997 539998 173063 540014
rect 173189 540048 173255 540064
rect 173303 540060 173333 540086
rect 173399 540064 173429 540086
rect 173189 540014 173205 540048
rect 173239 540014 173255 540048
rect 173189 539998 173255 540014
rect 173381 540048 173447 540064
rect 173495 540060 173525 540086
rect 173712 540057 173742 540079
rect 173912 540057 173942 540079
rect 173381 540014 173397 540048
rect 173431 540014 173447 540048
rect 173381 539998 173447 540014
rect 173694 540041 173760 540057
rect 173694 540007 173710 540041
rect 173744 540007 173760 540041
rect 173694 539991 173760 540007
rect 173894 540041 173960 540057
rect 173894 540007 173910 540041
rect 173944 540007 173960 540041
rect 173894 539991 173960 540007
rect 175940 541174 177030 541177
rect 175940 541167 177043 541174
rect 175714 541151 175780 541167
rect 175714 541117 175730 541151
rect 175764 541117 175780 541151
rect 175714 541101 175780 541117
rect 175939 541158 177043 541167
rect 175939 541124 176033 541158
rect 176067 541124 176225 541158
rect 176259 541124 176417 541158
rect 176451 541124 176609 541158
rect 176643 541124 176801 541158
rect 176835 541124 176993 541158
rect 177027 541124 177043 541158
rect 175939 541117 177043 541124
rect 175732 541079 175762 541101
rect 175939 541086 175969 541117
rect 176017 541108 177043 541117
rect 177394 541151 177460 541167
rect 177394 541117 177410 541151
rect 177444 541117 177460 541151
rect 176034 541107 177030 541108
rect 176035 541086 176065 541107
rect 176131 541086 176161 541107
rect 176227 541086 176257 541107
rect 176323 541086 176353 541107
rect 176419 541086 176449 541107
rect 176515 541086 176545 541107
rect 176611 541086 176641 541107
rect 176707 541086 176737 541107
rect 176803 541086 176833 541107
rect 176899 541086 176929 541107
rect 176995 541086 177025 541107
rect 177394 541101 177460 541117
rect 177412 541079 177442 541101
rect 177194 540351 177260 540367
rect 177194 540317 177210 540351
rect 177244 540317 177260 540351
rect 177194 540301 177260 540317
rect 177212 540279 177242 540301
rect 175732 540057 175762 540079
rect 175939 540064 175969 540086
rect 175714 540041 175780 540057
rect 175714 540007 175730 540041
rect 175764 540007 175780 540041
rect 175714 539991 175780 540007
rect 175921 540048 175987 540064
rect 176035 540060 176065 540086
rect 176131 540064 176161 540086
rect 175921 540014 175937 540048
rect 175971 540014 175987 540048
rect 175921 539998 175987 540014
rect 176113 540048 176179 540064
rect 176227 540060 176257 540086
rect 176323 540064 176353 540086
rect 176113 540014 176129 540048
rect 176163 540014 176179 540048
rect 176113 539998 176179 540014
rect 176305 540048 176371 540064
rect 176419 540060 176449 540086
rect 176515 540064 176545 540086
rect 176305 540014 176321 540048
rect 176355 540014 176371 540048
rect 176305 539998 176371 540014
rect 176497 540048 176563 540064
rect 176611 540060 176641 540086
rect 176707 540064 176737 540086
rect 176497 540014 176513 540048
rect 176547 540014 176563 540048
rect 176497 539998 176563 540014
rect 176689 540048 176755 540064
rect 176803 540060 176833 540086
rect 176899 540064 176929 540086
rect 176689 540014 176705 540048
rect 176739 540014 176755 540048
rect 176689 539998 176755 540014
rect 176881 540048 176947 540064
rect 176995 540060 177025 540086
rect 177212 540057 177242 540079
rect 177412 540057 177442 540079
rect 176881 540014 176897 540048
rect 176931 540014 176947 540048
rect 176881 539998 176947 540014
rect 177194 540041 177260 540057
rect 177194 540007 177210 540041
rect 177244 540007 177260 540041
rect 177194 539991 177260 540007
rect 177394 540041 177460 540057
rect 177394 540007 177410 540041
rect 177444 540007 177460 540041
rect 177394 539991 177460 540007
rect 179540 541174 180630 541177
rect 179540 541167 180643 541174
rect 179314 541151 179380 541167
rect 179314 541117 179330 541151
rect 179364 541117 179380 541151
rect 179314 541101 179380 541117
rect 179539 541158 180643 541167
rect 179539 541124 179633 541158
rect 179667 541124 179825 541158
rect 179859 541124 180017 541158
rect 180051 541124 180209 541158
rect 180243 541124 180401 541158
rect 180435 541124 180593 541158
rect 180627 541124 180643 541158
rect 179539 541117 180643 541124
rect 179332 541079 179362 541101
rect 179539 541086 179569 541117
rect 179617 541108 180643 541117
rect 180994 541151 181060 541167
rect 180994 541117 181010 541151
rect 181044 541117 181060 541151
rect 179634 541107 180630 541108
rect 179635 541086 179665 541107
rect 179731 541086 179761 541107
rect 179827 541086 179857 541107
rect 179923 541086 179953 541107
rect 180019 541086 180049 541107
rect 180115 541086 180145 541107
rect 180211 541086 180241 541107
rect 180307 541086 180337 541107
rect 180403 541086 180433 541107
rect 180499 541086 180529 541107
rect 180595 541086 180625 541107
rect 180994 541101 181060 541117
rect 181012 541079 181042 541101
rect 180794 540351 180860 540367
rect 180794 540317 180810 540351
rect 180844 540317 180860 540351
rect 180794 540301 180860 540317
rect 180812 540279 180842 540301
rect 179332 540057 179362 540079
rect 179539 540064 179569 540086
rect 179314 540041 179380 540057
rect 179314 540007 179330 540041
rect 179364 540007 179380 540041
rect 179314 539991 179380 540007
rect 179521 540048 179587 540064
rect 179635 540060 179665 540086
rect 179731 540064 179761 540086
rect 179521 540014 179537 540048
rect 179571 540014 179587 540048
rect 179521 539998 179587 540014
rect 179713 540048 179779 540064
rect 179827 540060 179857 540086
rect 179923 540064 179953 540086
rect 179713 540014 179729 540048
rect 179763 540014 179779 540048
rect 179713 539998 179779 540014
rect 179905 540048 179971 540064
rect 180019 540060 180049 540086
rect 180115 540064 180145 540086
rect 179905 540014 179921 540048
rect 179955 540014 179971 540048
rect 179905 539998 179971 540014
rect 180097 540048 180163 540064
rect 180211 540060 180241 540086
rect 180307 540064 180337 540086
rect 180097 540014 180113 540048
rect 180147 540014 180163 540048
rect 180097 539998 180163 540014
rect 180289 540048 180355 540064
rect 180403 540060 180433 540086
rect 180499 540064 180529 540086
rect 180289 540014 180305 540048
rect 180339 540014 180355 540048
rect 180289 539998 180355 540014
rect 180481 540048 180547 540064
rect 180595 540060 180625 540086
rect 180812 540057 180842 540079
rect 181012 540057 181042 540079
rect 180481 540014 180497 540048
rect 180531 540014 180547 540048
rect 180481 539998 180547 540014
rect 180794 540041 180860 540057
rect 180794 540007 180810 540041
rect 180844 540007 180860 540041
rect 180794 539991 180860 540007
rect 180994 540041 181060 540057
rect 180994 540007 181010 540041
rect 181044 540007 181060 540041
rect 180994 539991 181060 540007
rect 182840 541174 183930 541177
rect 182840 541167 183943 541174
rect 182614 541151 182680 541167
rect 182614 541117 182630 541151
rect 182664 541117 182680 541151
rect 182614 541101 182680 541117
rect 182839 541158 183943 541167
rect 182839 541124 182933 541158
rect 182967 541124 183125 541158
rect 183159 541124 183317 541158
rect 183351 541124 183509 541158
rect 183543 541124 183701 541158
rect 183735 541124 183893 541158
rect 183927 541124 183943 541158
rect 182839 541117 183943 541124
rect 182632 541079 182662 541101
rect 182839 541086 182869 541117
rect 182917 541108 183943 541117
rect 184294 541151 184360 541167
rect 184294 541117 184310 541151
rect 184344 541117 184360 541151
rect 182934 541107 183930 541108
rect 182935 541086 182965 541107
rect 183031 541086 183061 541107
rect 183127 541086 183157 541107
rect 183223 541086 183253 541107
rect 183319 541086 183349 541107
rect 183415 541086 183445 541107
rect 183511 541086 183541 541107
rect 183607 541086 183637 541107
rect 183703 541086 183733 541107
rect 183799 541086 183829 541107
rect 183895 541086 183925 541107
rect 184294 541101 184360 541117
rect 184312 541079 184342 541101
rect 184094 540351 184160 540367
rect 184094 540317 184110 540351
rect 184144 540317 184160 540351
rect 184094 540301 184160 540317
rect 184112 540279 184142 540301
rect 182632 540057 182662 540079
rect 182839 540064 182869 540086
rect 182614 540041 182680 540057
rect 182614 540007 182630 540041
rect 182664 540007 182680 540041
rect 182614 539991 182680 540007
rect 182821 540048 182887 540064
rect 182935 540060 182965 540086
rect 183031 540064 183061 540086
rect 182821 540014 182837 540048
rect 182871 540014 182887 540048
rect 182821 539998 182887 540014
rect 183013 540048 183079 540064
rect 183127 540060 183157 540086
rect 183223 540064 183253 540086
rect 183013 540014 183029 540048
rect 183063 540014 183079 540048
rect 183013 539998 183079 540014
rect 183205 540048 183271 540064
rect 183319 540060 183349 540086
rect 183415 540064 183445 540086
rect 183205 540014 183221 540048
rect 183255 540014 183271 540048
rect 183205 539998 183271 540014
rect 183397 540048 183463 540064
rect 183511 540060 183541 540086
rect 183607 540064 183637 540086
rect 183397 540014 183413 540048
rect 183447 540014 183463 540048
rect 183397 539998 183463 540014
rect 183589 540048 183655 540064
rect 183703 540060 183733 540086
rect 183799 540064 183829 540086
rect 183589 540014 183605 540048
rect 183639 540014 183655 540048
rect 183589 539998 183655 540014
rect 183781 540048 183847 540064
rect 183895 540060 183925 540086
rect 184112 540057 184142 540079
rect 184312 540057 184342 540079
rect 183781 540014 183797 540048
rect 183831 540014 183847 540048
rect 183781 539998 183847 540014
rect 184094 540041 184160 540057
rect 184094 540007 184110 540041
rect 184144 540007 184160 540041
rect 184094 539991 184160 540007
rect 184294 540041 184360 540057
rect 184294 540007 184310 540041
rect 184344 540007 184360 540041
rect 184294 539991 184360 540007
rect 186140 541174 187230 541177
rect 186140 541167 187243 541174
rect 185914 541151 185980 541167
rect 185914 541117 185930 541151
rect 185964 541117 185980 541151
rect 185914 541101 185980 541117
rect 186139 541158 187243 541167
rect 186139 541124 186233 541158
rect 186267 541124 186425 541158
rect 186459 541124 186617 541158
rect 186651 541124 186809 541158
rect 186843 541124 187001 541158
rect 187035 541124 187193 541158
rect 187227 541124 187243 541158
rect 186139 541117 187243 541124
rect 185932 541079 185962 541101
rect 186139 541086 186169 541117
rect 186217 541108 187243 541117
rect 187594 541151 187660 541167
rect 187594 541117 187610 541151
rect 187644 541117 187660 541151
rect 186234 541107 187230 541108
rect 186235 541086 186265 541107
rect 186331 541086 186361 541107
rect 186427 541086 186457 541107
rect 186523 541086 186553 541107
rect 186619 541086 186649 541107
rect 186715 541086 186745 541107
rect 186811 541086 186841 541107
rect 186907 541086 186937 541107
rect 187003 541086 187033 541107
rect 187099 541086 187129 541107
rect 187195 541086 187225 541107
rect 187594 541101 187660 541117
rect 187612 541079 187642 541101
rect 187394 540351 187460 540367
rect 187394 540317 187410 540351
rect 187444 540317 187460 540351
rect 187394 540301 187460 540317
rect 187412 540279 187442 540301
rect 185932 540057 185962 540079
rect 186139 540064 186169 540086
rect 185914 540041 185980 540057
rect 185914 540007 185930 540041
rect 185964 540007 185980 540041
rect 185914 539991 185980 540007
rect 186121 540048 186187 540064
rect 186235 540060 186265 540086
rect 186331 540064 186361 540086
rect 186121 540014 186137 540048
rect 186171 540014 186187 540048
rect 186121 539998 186187 540014
rect 186313 540048 186379 540064
rect 186427 540060 186457 540086
rect 186523 540064 186553 540086
rect 186313 540014 186329 540048
rect 186363 540014 186379 540048
rect 186313 539998 186379 540014
rect 186505 540048 186571 540064
rect 186619 540060 186649 540086
rect 186715 540064 186745 540086
rect 186505 540014 186521 540048
rect 186555 540014 186571 540048
rect 186505 539998 186571 540014
rect 186697 540048 186763 540064
rect 186811 540060 186841 540086
rect 186907 540064 186937 540086
rect 186697 540014 186713 540048
rect 186747 540014 186763 540048
rect 186697 539998 186763 540014
rect 186889 540048 186955 540064
rect 187003 540060 187033 540086
rect 187099 540064 187129 540086
rect 186889 540014 186905 540048
rect 186939 540014 186955 540048
rect 186889 539998 186955 540014
rect 187081 540048 187147 540064
rect 187195 540060 187225 540086
rect 187412 540057 187442 540079
rect 187612 540057 187642 540079
rect 187081 540014 187097 540048
rect 187131 540014 187147 540048
rect 187081 539998 187147 540014
rect 187394 540041 187460 540057
rect 187394 540007 187410 540041
rect 187444 540007 187460 540041
rect 187394 539991 187460 540007
rect 187594 540041 187660 540057
rect 187594 540007 187610 540041
rect 187644 540007 187660 540041
rect 187594 539991 187660 540007
rect 189440 541174 190530 541177
rect 189440 541167 190543 541174
rect 189214 541151 189280 541167
rect 189214 541117 189230 541151
rect 189264 541117 189280 541151
rect 189214 541101 189280 541117
rect 189439 541158 190543 541167
rect 189439 541124 189533 541158
rect 189567 541124 189725 541158
rect 189759 541124 189917 541158
rect 189951 541124 190109 541158
rect 190143 541124 190301 541158
rect 190335 541124 190493 541158
rect 190527 541124 190543 541158
rect 189439 541117 190543 541124
rect 189232 541079 189262 541101
rect 189439 541086 189469 541117
rect 189517 541108 190543 541117
rect 190894 541151 190960 541167
rect 190894 541117 190910 541151
rect 190944 541117 190960 541151
rect 189534 541107 190530 541108
rect 189535 541086 189565 541107
rect 189631 541086 189661 541107
rect 189727 541086 189757 541107
rect 189823 541086 189853 541107
rect 189919 541086 189949 541107
rect 190015 541086 190045 541107
rect 190111 541086 190141 541107
rect 190207 541086 190237 541107
rect 190303 541086 190333 541107
rect 190399 541086 190429 541107
rect 190495 541086 190525 541107
rect 190894 541101 190960 541117
rect 190912 541079 190942 541101
rect 190694 540351 190760 540367
rect 190694 540317 190710 540351
rect 190744 540317 190760 540351
rect 190694 540301 190760 540317
rect 190712 540279 190742 540301
rect 189232 540057 189262 540079
rect 189439 540064 189469 540086
rect 189214 540041 189280 540057
rect 189214 540007 189230 540041
rect 189264 540007 189280 540041
rect 189214 539991 189280 540007
rect 189421 540048 189487 540064
rect 189535 540060 189565 540086
rect 189631 540064 189661 540086
rect 189421 540014 189437 540048
rect 189471 540014 189487 540048
rect 189421 539998 189487 540014
rect 189613 540048 189679 540064
rect 189727 540060 189757 540086
rect 189823 540064 189853 540086
rect 189613 540014 189629 540048
rect 189663 540014 189679 540048
rect 189613 539998 189679 540014
rect 189805 540048 189871 540064
rect 189919 540060 189949 540086
rect 190015 540064 190045 540086
rect 189805 540014 189821 540048
rect 189855 540014 189871 540048
rect 189805 539998 189871 540014
rect 189997 540048 190063 540064
rect 190111 540060 190141 540086
rect 190207 540064 190237 540086
rect 189997 540014 190013 540048
rect 190047 540014 190063 540048
rect 189997 539998 190063 540014
rect 190189 540048 190255 540064
rect 190303 540060 190333 540086
rect 190399 540064 190429 540086
rect 190189 540014 190205 540048
rect 190239 540014 190255 540048
rect 190189 539998 190255 540014
rect 190381 540048 190447 540064
rect 190495 540060 190525 540086
rect 190712 540057 190742 540079
rect 190912 540057 190942 540079
rect 190381 540014 190397 540048
rect 190431 540014 190447 540048
rect 190381 539998 190447 540014
rect 190694 540041 190760 540057
rect 190694 540007 190710 540041
rect 190744 540007 190760 540041
rect 190694 539991 190760 540007
rect 190894 540041 190960 540057
rect 190894 540007 190910 540041
rect 190944 540007 190960 540041
rect 190894 539991 190960 540007
rect 158712 538501 158912 538517
rect 158712 538467 158728 538501
rect 158896 538467 158912 538501
rect 158712 538429 158912 538467
rect 159088 538501 159288 538517
rect 159088 538467 159104 538501
rect 159272 538467 159288 538501
rect 159088 538429 159288 538467
rect 159346 538501 159546 538517
rect 159346 538467 159362 538501
rect 159530 538467 159546 538501
rect 159346 538429 159546 538467
rect 159604 538501 159804 538517
rect 159604 538467 159620 538501
rect 159788 538467 159804 538501
rect 159604 538429 159804 538467
rect 159862 538501 160062 538517
rect 159862 538467 159878 538501
rect 160046 538467 160062 538501
rect 159862 538429 160062 538467
rect 160120 538501 160320 538517
rect 160120 538467 160136 538501
rect 160304 538467 160320 538501
rect 160120 538429 160320 538467
rect 160378 538501 160578 538517
rect 160378 538467 160394 538501
rect 160562 538467 160578 538501
rect 160378 538429 160578 538467
rect 160636 538501 160836 538517
rect 160636 538467 160652 538501
rect 160820 538467 160836 538501
rect 160636 538429 160836 538467
rect 160894 538501 161094 538517
rect 160894 538467 160910 538501
rect 161078 538467 161094 538501
rect 160894 538429 161094 538467
rect 161152 538501 161352 538517
rect 161152 538467 161168 538501
rect 161336 538467 161352 538501
rect 161152 538429 161352 538467
rect 161532 538501 161732 538517
rect 161532 538467 161548 538501
rect 161716 538467 161732 538501
rect 161532 538429 161732 538467
rect 161932 538501 162132 538517
rect 161932 538467 161948 538501
rect 162116 538467 162132 538501
rect 161932 538429 162132 538467
rect 162312 538501 162512 538517
rect 162312 538467 162328 538501
rect 162496 538467 162512 538501
rect 162312 538429 162512 538467
rect 158712 538191 158912 538229
rect 158712 538157 158728 538191
rect 158896 538157 158912 538191
rect 158712 538141 158912 538157
rect 159088 538191 159288 538229
rect 159088 538157 159104 538191
rect 159272 538157 159288 538191
rect 159088 538141 159288 538157
rect 159346 538191 159546 538229
rect 159346 538157 159362 538191
rect 159530 538157 159546 538191
rect 159346 538141 159546 538157
rect 159604 538191 159804 538229
rect 159604 538157 159620 538191
rect 159788 538157 159804 538191
rect 159604 538141 159804 538157
rect 159862 538191 160062 538229
rect 159862 538157 159878 538191
rect 160046 538157 160062 538191
rect 159862 538141 160062 538157
rect 160120 538191 160320 538229
rect 160120 538157 160136 538191
rect 160304 538157 160320 538191
rect 160120 538141 160320 538157
rect 160378 538191 160578 538229
rect 160378 538157 160394 538191
rect 160562 538157 160578 538191
rect 160378 538141 160578 538157
rect 160636 538191 160836 538229
rect 160636 538157 160652 538191
rect 160820 538157 160836 538191
rect 160636 538141 160836 538157
rect 160894 538191 161094 538229
rect 160894 538157 160910 538191
rect 161078 538157 161094 538191
rect 160894 538141 161094 538157
rect 161152 538191 161352 538229
rect 161152 538157 161168 538191
rect 161336 538157 161352 538191
rect 161152 538141 161352 538157
rect 161532 538191 161732 538229
rect 161532 538157 161548 538191
rect 161716 538157 161732 538191
rect 161532 538141 161732 538157
rect 161932 538191 162132 538229
rect 161932 538157 161948 538191
rect 162116 538157 162132 538191
rect 161932 538141 162132 538157
rect 162312 538191 162512 538229
rect 162312 538157 162328 538191
rect 162496 538157 162512 538191
rect 162312 538141 162512 538157
rect 164698 539638 164764 539654
rect 164698 539604 164714 539638
rect 164748 539604 164764 539638
rect 164698 539588 164764 539604
rect 165021 539645 165087 539661
rect 165021 539611 165037 539645
rect 165071 539611 165087 539645
rect 165021 539595 165087 539611
rect 165213 539645 165279 539661
rect 165213 539611 165229 539645
rect 165263 539611 165279 539645
rect 165213 539595 165279 539611
rect 165405 539645 165471 539661
rect 165405 539611 165421 539645
rect 165455 539611 165471 539645
rect 165405 539595 165471 539611
rect 165597 539645 165663 539661
rect 165597 539611 165613 539645
rect 165647 539611 165663 539645
rect 165597 539595 165663 539611
rect 165789 539645 165855 539661
rect 165789 539611 165805 539645
rect 165839 539611 165855 539645
rect 165789 539595 165855 539611
rect 165981 539645 166047 539661
rect 165981 539611 165997 539645
rect 166031 539611 166047 539645
rect 165981 539595 166047 539611
rect 166198 539638 166264 539654
rect 166198 539604 166214 539638
rect 166248 539604 166264 539638
rect 164716 539557 164746 539588
rect 164943 539564 164973 539590
rect 165039 539564 165069 539595
rect 165135 539564 165165 539590
rect 165231 539564 165261 539595
rect 165327 539564 165357 539590
rect 165423 539564 165453 539595
rect 165519 539564 165549 539590
rect 165615 539564 165645 539595
rect 165711 539564 165741 539590
rect 165807 539564 165837 539595
rect 165903 539564 165933 539590
rect 165999 539564 166029 539595
rect 166198 539588 166264 539604
rect 166398 539638 166464 539654
rect 166398 539604 166414 539638
rect 166448 539604 166464 539638
rect 166398 539588 166464 539604
rect 166216 539557 166246 539588
rect 166416 539557 166446 539588
rect 166216 538926 166246 538957
rect 166198 538910 166264 538926
rect 166198 538876 166214 538910
rect 166248 538876 166264 538910
rect 166198 538860 166264 538876
rect 164716 538526 164746 538557
rect 164943 538533 164973 538564
rect 164925 538527 164991 538533
rect 165039 538527 165069 538564
rect 165135 538533 165165 538564
rect 165117 538527 165183 538533
rect 165231 538527 165261 538564
rect 165327 538533 165357 538564
rect 165309 538527 165375 538533
rect 165423 538527 165453 538564
rect 165519 538533 165549 538564
rect 165501 538527 165567 538533
rect 165615 538527 165645 538564
rect 165711 538533 165741 538564
rect 165693 538527 165759 538533
rect 165807 538527 165837 538564
rect 165903 538533 165933 538564
rect 165999 538547 166029 538564
rect 165885 538527 165951 538533
rect 165996 538527 166030 538547
rect 164698 538510 164764 538526
rect 164698 538476 164714 538510
rect 164748 538476 164764 538510
rect 164698 538460 164764 538476
rect 164925 538517 166030 538527
rect 166416 538526 166446 538557
rect 164925 538483 164941 538517
rect 164975 538483 165133 538517
rect 165167 538483 165325 538517
rect 165359 538483 165517 538517
rect 165551 538483 165709 538517
rect 165743 538483 165901 538517
rect 165935 538483 166030 538517
rect 164925 538477 166030 538483
rect 166398 538510 166464 538526
rect 164925 538467 164991 538477
rect 165117 538467 165183 538477
rect 165309 538467 165375 538477
rect 165501 538467 165567 538477
rect 165693 538467 165759 538477
rect 165885 538467 165951 538477
rect 166398 538476 166414 538510
rect 166448 538476 166464 538510
rect 166398 538460 166464 538476
rect 168498 539638 168564 539654
rect 168498 539604 168514 539638
rect 168548 539604 168564 539638
rect 168498 539588 168564 539604
rect 168821 539645 168887 539661
rect 168821 539611 168837 539645
rect 168871 539611 168887 539645
rect 168821 539595 168887 539611
rect 169013 539645 169079 539661
rect 169013 539611 169029 539645
rect 169063 539611 169079 539645
rect 169013 539595 169079 539611
rect 169205 539645 169271 539661
rect 169205 539611 169221 539645
rect 169255 539611 169271 539645
rect 169205 539595 169271 539611
rect 169397 539645 169463 539661
rect 169397 539611 169413 539645
rect 169447 539611 169463 539645
rect 169397 539595 169463 539611
rect 169589 539645 169655 539661
rect 169589 539611 169605 539645
rect 169639 539611 169655 539645
rect 169589 539595 169655 539611
rect 169781 539645 169847 539661
rect 169781 539611 169797 539645
rect 169831 539611 169847 539645
rect 169781 539595 169847 539611
rect 169998 539638 170064 539654
rect 169998 539604 170014 539638
rect 170048 539604 170064 539638
rect 168516 539557 168546 539588
rect 168743 539564 168773 539590
rect 168839 539564 168869 539595
rect 168935 539564 168965 539590
rect 169031 539564 169061 539595
rect 169127 539564 169157 539590
rect 169223 539564 169253 539595
rect 169319 539564 169349 539590
rect 169415 539564 169445 539595
rect 169511 539564 169541 539590
rect 169607 539564 169637 539595
rect 169703 539564 169733 539590
rect 169799 539564 169829 539595
rect 169998 539588 170064 539604
rect 170198 539638 170264 539654
rect 170198 539604 170214 539638
rect 170248 539604 170264 539638
rect 170198 539588 170264 539604
rect 170016 539557 170046 539588
rect 170216 539557 170246 539588
rect 170016 538926 170046 538957
rect 169998 538910 170064 538926
rect 169998 538876 170014 538910
rect 170048 538876 170064 538910
rect 169998 538860 170064 538876
rect 168516 538526 168546 538557
rect 168743 538533 168773 538564
rect 168725 538527 168791 538533
rect 168839 538527 168869 538564
rect 168935 538533 168965 538564
rect 168917 538527 168983 538533
rect 169031 538527 169061 538564
rect 169127 538533 169157 538564
rect 169109 538527 169175 538533
rect 169223 538527 169253 538564
rect 169319 538533 169349 538564
rect 169301 538527 169367 538533
rect 169415 538527 169445 538564
rect 169511 538533 169541 538564
rect 169493 538527 169559 538533
rect 169607 538527 169637 538564
rect 169703 538533 169733 538564
rect 169799 538547 169829 538564
rect 169685 538527 169751 538533
rect 169796 538527 169830 538547
rect 168498 538510 168564 538526
rect 168498 538476 168514 538510
rect 168548 538476 168564 538510
rect 168498 538460 168564 538476
rect 168725 538517 169830 538527
rect 170216 538526 170246 538557
rect 168725 538483 168741 538517
rect 168775 538483 168933 538517
rect 168967 538483 169125 538517
rect 169159 538483 169317 538517
rect 169351 538483 169509 538517
rect 169543 538483 169701 538517
rect 169735 538483 169830 538517
rect 168725 538477 169830 538483
rect 170198 538510 170264 538526
rect 168725 538467 168791 538477
rect 168917 538467 168983 538477
rect 169109 538467 169175 538477
rect 169301 538467 169367 538477
rect 169493 538467 169559 538477
rect 169685 538467 169751 538477
rect 170198 538476 170214 538510
rect 170248 538476 170264 538510
rect 170198 538460 170264 538476
rect 172198 539638 172264 539654
rect 172198 539604 172214 539638
rect 172248 539604 172264 539638
rect 172198 539588 172264 539604
rect 172521 539645 172587 539661
rect 172521 539611 172537 539645
rect 172571 539611 172587 539645
rect 172521 539595 172587 539611
rect 172713 539645 172779 539661
rect 172713 539611 172729 539645
rect 172763 539611 172779 539645
rect 172713 539595 172779 539611
rect 172905 539645 172971 539661
rect 172905 539611 172921 539645
rect 172955 539611 172971 539645
rect 172905 539595 172971 539611
rect 173097 539645 173163 539661
rect 173097 539611 173113 539645
rect 173147 539611 173163 539645
rect 173097 539595 173163 539611
rect 173289 539645 173355 539661
rect 173289 539611 173305 539645
rect 173339 539611 173355 539645
rect 173289 539595 173355 539611
rect 173481 539645 173547 539661
rect 173481 539611 173497 539645
rect 173531 539611 173547 539645
rect 173481 539595 173547 539611
rect 173698 539638 173764 539654
rect 173698 539604 173714 539638
rect 173748 539604 173764 539638
rect 172216 539557 172246 539588
rect 172443 539564 172473 539590
rect 172539 539564 172569 539595
rect 172635 539564 172665 539590
rect 172731 539564 172761 539595
rect 172827 539564 172857 539590
rect 172923 539564 172953 539595
rect 173019 539564 173049 539590
rect 173115 539564 173145 539595
rect 173211 539564 173241 539590
rect 173307 539564 173337 539595
rect 173403 539564 173433 539590
rect 173499 539564 173529 539595
rect 173698 539588 173764 539604
rect 173898 539638 173964 539654
rect 173898 539604 173914 539638
rect 173948 539604 173964 539638
rect 173898 539588 173964 539604
rect 173716 539557 173746 539588
rect 173916 539557 173946 539588
rect 173716 538926 173746 538957
rect 173698 538910 173764 538926
rect 173698 538876 173714 538910
rect 173748 538876 173764 538910
rect 173698 538860 173764 538876
rect 172216 538526 172246 538557
rect 172443 538533 172473 538564
rect 172425 538527 172491 538533
rect 172539 538527 172569 538564
rect 172635 538533 172665 538564
rect 172617 538527 172683 538533
rect 172731 538527 172761 538564
rect 172827 538533 172857 538564
rect 172809 538527 172875 538533
rect 172923 538527 172953 538564
rect 173019 538533 173049 538564
rect 173001 538527 173067 538533
rect 173115 538527 173145 538564
rect 173211 538533 173241 538564
rect 173193 538527 173259 538533
rect 173307 538527 173337 538564
rect 173403 538533 173433 538564
rect 173499 538547 173529 538564
rect 173385 538527 173451 538533
rect 173496 538527 173530 538547
rect 172198 538510 172264 538526
rect 172198 538476 172214 538510
rect 172248 538476 172264 538510
rect 172198 538460 172264 538476
rect 172425 538517 173530 538527
rect 173916 538526 173946 538557
rect 172425 538483 172441 538517
rect 172475 538483 172633 538517
rect 172667 538483 172825 538517
rect 172859 538483 173017 538517
rect 173051 538483 173209 538517
rect 173243 538483 173401 538517
rect 173435 538483 173530 538517
rect 172425 538477 173530 538483
rect 173898 538510 173964 538526
rect 172425 538467 172491 538477
rect 172617 538467 172683 538477
rect 172809 538467 172875 538477
rect 173001 538467 173067 538477
rect 173193 538467 173259 538477
rect 173385 538467 173451 538477
rect 173898 538476 173914 538510
rect 173948 538476 173964 538510
rect 173898 538460 173964 538476
rect 175698 539638 175764 539654
rect 175698 539604 175714 539638
rect 175748 539604 175764 539638
rect 175698 539588 175764 539604
rect 176021 539645 176087 539661
rect 176021 539611 176037 539645
rect 176071 539611 176087 539645
rect 176021 539595 176087 539611
rect 176213 539645 176279 539661
rect 176213 539611 176229 539645
rect 176263 539611 176279 539645
rect 176213 539595 176279 539611
rect 176405 539645 176471 539661
rect 176405 539611 176421 539645
rect 176455 539611 176471 539645
rect 176405 539595 176471 539611
rect 176597 539645 176663 539661
rect 176597 539611 176613 539645
rect 176647 539611 176663 539645
rect 176597 539595 176663 539611
rect 176789 539645 176855 539661
rect 176789 539611 176805 539645
rect 176839 539611 176855 539645
rect 176789 539595 176855 539611
rect 176981 539645 177047 539661
rect 176981 539611 176997 539645
rect 177031 539611 177047 539645
rect 176981 539595 177047 539611
rect 177198 539638 177264 539654
rect 177198 539604 177214 539638
rect 177248 539604 177264 539638
rect 175716 539557 175746 539588
rect 175943 539564 175973 539590
rect 176039 539564 176069 539595
rect 176135 539564 176165 539590
rect 176231 539564 176261 539595
rect 176327 539564 176357 539590
rect 176423 539564 176453 539595
rect 176519 539564 176549 539590
rect 176615 539564 176645 539595
rect 176711 539564 176741 539590
rect 176807 539564 176837 539595
rect 176903 539564 176933 539590
rect 176999 539564 177029 539595
rect 177198 539588 177264 539604
rect 177398 539638 177464 539654
rect 177398 539604 177414 539638
rect 177448 539604 177464 539638
rect 177398 539588 177464 539604
rect 177216 539557 177246 539588
rect 177416 539557 177446 539588
rect 177216 538926 177246 538957
rect 177198 538910 177264 538926
rect 177198 538876 177214 538910
rect 177248 538876 177264 538910
rect 177198 538860 177264 538876
rect 175716 538526 175746 538557
rect 175943 538533 175973 538564
rect 175925 538527 175991 538533
rect 176039 538527 176069 538564
rect 176135 538533 176165 538564
rect 176117 538527 176183 538533
rect 176231 538527 176261 538564
rect 176327 538533 176357 538564
rect 176309 538527 176375 538533
rect 176423 538527 176453 538564
rect 176519 538533 176549 538564
rect 176501 538527 176567 538533
rect 176615 538527 176645 538564
rect 176711 538533 176741 538564
rect 176693 538527 176759 538533
rect 176807 538527 176837 538564
rect 176903 538533 176933 538564
rect 176999 538547 177029 538564
rect 176885 538527 176951 538533
rect 176996 538527 177030 538547
rect 175698 538510 175764 538526
rect 175698 538476 175714 538510
rect 175748 538476 175764 538510
rect 175698 538460 175764 538476
rect 175925 538517 177030 538527
rect 177416 538526 177446 538557
rect 175925 538483 175941 538517
rect 175975 538483 176133 538517
rect 176167 538483 176325 538517
rect 176359 538483 176517 538517
rect 176551 538483 176709 538517
rect 176743 538483 176901 538517
rect 176935 538483 177030 538517
rect 175925 538477 177030 538483
rect 177398 538510 177464 538526
rect 175925 538467 175991 538477
rect 176117 538467 176183 538477
rect 176309 538467 176375 538477
rect 176501 538467 176567 538477
rect 176693 538467 176759 538477
rect 176885 538467 176951 538477
rect 177398 538476 177414 538510
rect 177448 538476 177464 538510
rect 177398 538460 177464 538476
rect 179298 539638 179364 539654
rect 179298 539604 179314 539638
rect 179348 539604 179364 539638
rect 179298 539588 179364 539604
rect 179621 539645 179687 539661
rect 179621 539611 179637 539645
rect 179671 539611 179687 539645
rect 179621 539595 179687 539611
rect 179813 539645 179879 539661
rect 179813 539611 179829 539645
rect 179863 539611 179879 539645
rect 179813 539595 179879 539611
rect 180005 539645 180071 539661
rect 180005 539611 180021 539645
rect 180055 539611 180071 539645
rect 180005 539595 180071 539611
rect 180197 539645 180263 539661
rect 180197 539611 180213 539645
rect 180247 539611 180263 539645
rect 180197 539595 180263 539611
rect 180389 539645 180455 539661
rect 180389 539611 180405 539645
rect 180439 539611 180455 539645
rect 180389 539595 180455 539611
rect 180581 539645 180647 539661
rect 180581 539611 180597 539645
rect 180631 539611 180647 539645
rect 180581 539595 180647 539611
rect 180798 539638 180864 539654
rect 180798 539604 180814 539638
rect 180848 539604 180864 539638
rect 179316 539557 179346 539588
rect 179543 539564 179573 539590
rect 179639 539564 179669 539595
rect 179735 539564 179765 539590
rect 179831 539564 179861 539595
rect 179927 539564 179957 539590
rect 180023 539564 180053 539595
rect 180119 539564 180149 539590
rect 180215 539564 180245 539595
rect 180311 539564 180341 539590
rect 180407 539564 180437 539595
rect 180503 539564 180533 539590
rect 180599 539564 180629 539595
rect 180798 539588 180864 539604
rect 180998 539638 181064 539654
rect 180998 539604 181014 539638
rect 181048 539604 181064 539638
rect 180998 539588 181064 539604
rect 180816 539557 180846 539588
rect 181016 539557 181046 539588
rect 180816 538926 180846 538957
rect 180798 538910 180864 538926
rect 180798 538876 180814 538910
rect 180848 538876 180864 538910
rect 180798 538860 180864 538876
rect 179316 538526 179346 538557
rect 179543 538533 179573 538564
rect 179525 538527 179591 538533
rect 179639 538527 179669 538564
rect 179735 538533 179765 538564
rect 179717 538527 179783 538533
rect 179831 538527 179861 538564
rect 179927 538533 179957 538564
rect 179909 538527 179975 538533
rect 180023 538527 180053 538564
rect 180119 538533 180149 538564
rect 180101 538527 180167 538533
rect 180215 538527 180245 538564
rect 180311 538533 180341 538564
rect 180293 538527 180359 538533
rect 180407 538527 180437 538564
rect 180503 538533 180533 538564
rect 180599 538547 180629 538564
rect 180485 538527 180551 538533
rect 180596 538527 180630 538547
rect 179298 538510 179364 538526
rect 179298 538476 179314 538510
rect 179348 538476 179364 538510
rect 179298 538460 179364 538476
rect 179525 538517 180630 538527
rect 181016 538526 181046 538557
rect 179525 538483 179541 538517
rect 179575 538483 179733 538517
rect 179767 538483 179925 538517
rect 179959 538483 180117 538517
rect 180151 538483 180309 538517
rect 180343 538483 180501 538517
rect 180535 538483 180630 538517
rect 179525 538477 180630 538483
rect 180998 538510 181064 538526
rect 179525 538467 179591 538477
rect 179717 538467 179783 538477
rect 179909 538467 179975 538477
rect 180101 538467 180167 538477
rect 180293 538467 180359 538477
rect 180485 538467 180551 538477
rect 180998 538476 181014 538510
rect 181048 538476 181064 538510
rect 180998 538460 181064 538476
rect 182598 539638 182664 539654
rect 182598 539604 182614 539638
rect 182648 539604 182664 539638
rect 182598 539588 182664 539604
rect 182921 539645 182987 539661
rect 182921 539611 182937 539645
rect 182971 539611 182987 539645
rect 182921 539595 182987 539611
rect 183113 539645 183179 539661
rect 183113 539611 183129 539645
rect 183163 539611 183179 539645
rect 183113 539595 183179 539611
rect 183305 539645 183371 539661
rect 183305 539611 183321 539645
rect 183355 539611 183371 539645
rect 183305 539595 183371 539611
rect 183497 539645 183563 539661
rect 183497 539611 183513 539645
rect 183547 539611 183563 539645
rect 183497 539595 183563 539611
rect 183689 539645 183755 539661
rect 183689 539611 183705 539645
rect 183739 539611 183755 539645
rect 183689 539595 183755 539611
rect 183881 539645 183947 539661
rect 183881 539611 183897 539645
rect 183931 539611 183947 539645
rect 183881 539595 183947 539611
rect 184098 539638 184164 539654
rect 184098 539604 184114 539638
rect 184148 539604 184164 539638
rect 182616 539557 182646 539588
rect 182843 539564 182873 539590
rect 182939 539564 182969 539595
rect 183035 539564 183065 539590
rect 183131 539564 183161 539595
rect 183227 539564 183257 539590
rect 183323 539564 183353 539595
rect 183419 539564 183449 539590
rect 183515 539564 183545 539595
rect 183611 539564 183641 539590
rect 183707 539564 183737 539595
rect 183803 539564 183833 539590
rect 183899 539564 183929 539595
rect 184098 539588 184164 539604
rect 184298 539638 184364 539654
rect 184298 539604 184314 539638
rect 184348 539604 184364 539638
rect 184298 539588 184364 539604
rect 184116 539557 184146 539588
rect 184316 539557 184346 539588
rect 184116 538926 184146 538957
rect 184098 538910 184164 538926
rect 184098 538876 184114 538910
rect 184148 538876 184164 538910
rect 184098 538860 184164 538876
rect 182616 538526 182646 538557
rect 182843 538533 182873 538564
rect 182825 538527 182891 538533
rect 182939 538527 182969 538564
rect 183035 538533 183065 538564
rect 183017 538527 183083 538533
rect 183131 538527 183161 538564
rect 183227 538533 183257 538564
rect 183209 538527 183275 538533
rect 183323 538527 183353 538564
rect 183419 538533 183449 538564
rect 183401 538527 183467 538533
rect 183515 538527 183545 538564
rect 183611 538533 183641 538564
rect 183593 538527 183659 538533
rect 183707 538527 183737 538564
rect 183803 538533 183833 538564
rect 183899 538547 183929 538564
rect 183785 538527 183851 538533
rect 183896 538527 183930 538547
rect 182598 538510 182664 538526
rect 182598 538476 182614 538510
rect 182648 538476 182664 538510
rect 182598 538460 182664 538476
rect 182825 538517 183930 538527
rect 184316 538526 184346 538557
rect 182825 538483 182841 538517
rect 182875 538483 183033 538517
rect 183067 538483 183225 538517
rect 183259 538483 183417 538517
rect 183451 538483 183609 538517
rect 183643 538483 183801 538517
rect 183835 538483 183930 538517
rect 182825 538477 183930 538483
rect 184298 538510 184364 538526
rect 182825 538467 182891 538477
rect 183017 538467 183083 538477
rect 183209 538467 183275 538477
rect 183401 538467 183467 538477
rect 183593 538467 183659 538477
rect 183785 538467 183851 538477
rect 184298 538476 184314 538510
rect 184348 538476 184364 538510
rect 184298 538460 184364 538476
rect 185898 539638 185964 539654
rect 185898 539604 185914 539638
rect 185948 539604 185964 539638
rect 185898 539588 185964 539604
rect 186221 539645 186287 539661
rect 186221 539611 186237 539645
rect 186271 539611 186287 539645
rect 186221 539595 186287 539611
rect 186413 539645 186479 539661
rect 186413 539611 186429 539645
rect 186463 539611 186479 539645
rect 186413 539595 186479 539611
rect 186605 539645 186671 539661
rect 186605 539611 186621 539645
rect 186655 539611 186671 539645
rect 186605 539595 186671 539611
rect 186797 539645 186863 539661
rect 186797 539611 186813 539645
rect 186847 539611 186863 539645
rect 186797 539595 186863 539611
rect 186989 539645 187055 539661
rect 186989 539611 187005 539645
rect 187039 539611 187055 539645
rect 186989 539595 187055 539611
rect 187181 539645 187247 539661
rect 187181 539611 187197 539645
rect 187231 539611 187247 539645
rect 187181 539595 187247 539611
rect 187398 539638 187464 539654
rect 187398 539604 187414 539638
rect 187448 539604 187464 539638
rect 185916 539557 185946 539588
rect 186143 539564 186173 539590
rect 186239 539564 186269 539595
rect 186335 539564 186365 539590
rect 186431 539564 186461 539595
rect 186527 539564 186557 539590
rect 186623 539564 186653 539595
rect 186719 539564 186749 539590
rect 186815 539564 186845 539595
rect 186911 539564 186941 539590
rect 187007 539564 187037 539595
rect 187103 539564 187133 539590
rect 187199 539564 187229 539595
rect 187398 539588 187464 539604
rect 187598 539638 187664 539654
rect 187598 539604 187614 539638
rect 187648 539604 187664 539638
rect 187598 539588 187664 539604
rect 187416 539557 187446 539588
rect 187616 539557 187646 539588
rect 187416 538926 187446 538957
rect 187398 538910 187464 538926
rect 187398 538876 187414 538910
rect 187448 538876 187464 538910
rect 187398 538860 187464 538876
rect 185916 538526 185946 538557
rect 186143 538533 186173 538564
rect 186125 538527 186191 538533
rect 186239 538527 186269 538564
rect 186335 538533 186365 538564
rect 186317 538527 186383 538533
rect 186431 538527 186461 538564
rect 186527 538533 186557 538564
rect 186509 538527 186575 538533
rect 186623 538527 186653 538564
rect 186719 538533 186749 538564
rect 186701 538527 186767 538533
rect 186815 538527 186845 538564
rect 186911 538533 186941 538564
rect 186893 538527 186959 538533
rect 187007 538527 187037 538564
rect 187103 538533 187133 538564
rect 187199 538547 187229 538564
rect 187085 538527 187151 538533
rect 187196 538527 187230 538547
rect 185898 538510 185964 538526
rect 185898 538476 185914 538510
rect 185948 538476 185964 538510
rect 185898 538460 185964 538476
rect 186125 538517 187230 538527
rect 187616 538526 187646 538557
rect 186125 538483 186141 538517
rect 186175 538483 186333 538517
rect 186367 538483 186525 538517
rect 186559 538483 186717 538517
rect 186751 538483 186909 538517
rect 186943 538483 187101 538517
rect 187135 538483 187230 538517
rect 186125 538477 187230 538483
rect 187598 538510 187664 538526
rect 186125 538467 186191 538477
rect 186317 538467 186383 538477
rect 186509 538467 186575 538477
rect 186701 538467 186767 538477
rect 186893 538467 186959 538477
rect 187085 538467 187151 538477
rect 187598 538476 187614 538510
rect 187648 538476 187664 538510
rect 187598 538460 187664 538476
rect 189198 539638 189264 539654
rect 189198 539604 189214 539638
rect 189248 539604 189264 539638
rect 189198 539588 189264 539604
rect 189521 539645 189587 539661
rect 189521 539611 189537 539645
rect 189571 539611 189587 539645
rect 189521 539595 189587 539611
rect 189713 539645 189779 539661
rect 189713 539611 189729 539645
rect 189763 539611 189779 539645
rect 189713 539595 189779 539611
rect 189905 539645 189971 539661
rect 189905 539611 189921 539645
rect 189955 539611 189971 539645
rect 189905 539595 189971 539611
rect 190097 539645 190163 539661
rect 190097 539611 190113 539645
rect 190147 539611 190163 539645
rect 190097 539595 190163 539611
rect 190289 539645 190355 539661
rect 190289 539611 190305 539645
rect 190339 539611 190355 539645
rect 190289 539595 190355 539611
rect 190481 539645 190547 539661
rect 190481 539611 190497 539645
rect 190531 539611 190547 539645
rect 190481 539595 190547 539611
rect 190698 539638 190764 539654
rect 190698 539604 190714 539638
rect 190748 539604 190764 539638
rect 189216 539557 189246 539588
rect 189443 539564 189473 539590
rect 189539 539564 189569 539595
rect 189635 539564 189665 539590
rect 189731 539564 189761 539595
rect 189827 539564 189857 539590
rect 189923 539564 189953 539595
rect 190019 539564 190049 539590
rect 190115 539564 190145 539595
rect 190211 539564 190241 539590
rect 190307 539564 190337 539595
rect 190403 539564 190433 539590
rect 190499 539564 190529 539595
rect 190698 539588 190764 539604
rect 190898 539638 190964 539654
rect 190898 539604 190914 539638
rect 190948 539604 190964 539638
rect 190898 539588 190964 539604
rect 190716 539557 190746 539588
rect 190916 539557 190946 539588
rect 190716 538926 190746 538957
rect 190698 538910 190764 538926
rect 190698 538876 190714 538910
rect 190748 538876 190764 538910
rect 190698 538860 190764 538876
rect 189216 538526 189246 538557
rect 189443 538533 189473 538564
rect 189425 538527 189491 538533
rect 189539 538527 189569 538564
rect 189635 538533 189665 538564
rect 189617 538527 189683 538533
rect 189731 538527 189761 538564
rect 189827 538533 189857 538564
rect 189809 538527 189875 538533
rect 189923 538527 189953 538564
rect 190019 538533 190049 538564
rect 190001 538527 190067 538533
rect 190115 538527 190145 538564
rect 190211 538533 190241 538564
rect 190193 538527 190259 538533
rect 190307 538527 190337 538564
rect 190403 538533 190433 538564
rect 190499 538547 190529 538564
rect 190385 538527 190451 538533
rect 190496 538527 190530 538547
rect 189198 538510 189264 538526
rect 189198 538476 189214 538510
rect 189248 538476 189264 538510
rect 189198 538460 189264 538476
rect 189425 538517 190530 538527
rect 190916 538526 190946 538557
rect 189425 538483 189441 538517
rect 189475 538483 189633 538517
rect 189667 538483 189825 538517
rect 189859 538483 190017 538517
rect 190051 538483 190209 538517
rect 190243 538483 190401 538517
rect 190435 538483 190530 538517
rect 189425 538477 190530 538483
rect 190898 538510 190964 538526
rect 189425 538467 189491 538477
rect 189617 538467 189683 538477
rect 189809 538467 189875 538477
rect 190001 538467 190067 538477
rect 190193 538467 190259 538477
rect 190385 538467 190451 538477
rect 190898 538476 190914 538510
rect 190948 538476 190964 538510
rect 190898 538460 190964 538476
rect 161288 537738 161354 537754
rect 161288 537704 161304 537738
rect 161338 537704 161354 537738
rect 161492 537738 161558 537754
rect 161492 537737 161508 537738
rect 161288 537688 161354 537704
rect 161490 537704 161508 537737
rect 161542 537737 161558 537738
rect 161684 537738 161750 537754
rect 161684 537737 161700 537738
rect 161542 537704 161700 537737
rect 161734 537704 161750 537738
rect 161306 537657 161336 537688
rect 161490 537677 161750 537704
rect 161892 537747 161958 537754
rect 162084 537747 162150 537754
rect 161892 537738 162150 537747
rect 161892 537704 161908 537738
rect 161942 537704 162100 537738
rect 162134 537704 162150 537738
rect 161892 537688 162150 537704
rect 162308 537738 162374 537754
rect 162308 537704 162324 537738
rect 162358 537704 162374 537738
rect 162308 537688 162374 537704
rect 161910 537677 162140 537688
rect 161510 537657 161540 537677
rect 161606 537657 161636 537677
rect 161702 537657 161732 537677
rect 161910 537657 161940 537677
rect 162006 537657 162036 537677
rect 162102 537657 162132 537677
rect 162326 537657 162356 537688
rect 161306 537026 161336 537057
rect 161510 537031 161540 537057
rect 161606 537026 161636 537057
rect 161702 537031 161732 537057
rect 161910 537031 161940 537057
rect 162006 537026 162036 537057
rect 162102 537031 162132 537057
rect 162326 537026 162356 537057
rect 161288 537010 161354 537026
rect 161288 536976 161304 537010
rect 161338 536976 161354 537010
rect 161288 536960 161354 536976
rect 161588 537010 161654 537026
rect 161588 536976 161604 537010
rect 161638 536976 161654 537010
rect 161588 536960 161654 536976
rect 161988 537010 162054 537026
rect 161988 536976 162004 537010
rect 162038 536976 162054 537010
rect 161988 536960 162054 536976
rect 162308 537010 162374 537026
rect 162308 536976 162324 537010
rect 162358 536976 162374 537010
rect 162308 536960 162374 536976
rect 157796 536718 157996 536734
rect 157796 536684 157812 536718
rect 157980 536684 157996 536718
rect 157796 536637 157996 536684
rect 158174 536718 158374 536734
rect 158174 536684 158190 536718
rect 158358 536684 158374 536718
rect 158174 536637 158374 536684
rect 158432 536718 158632 536734
rect 158432 536684 158448 536718
rect 158616 536684 158632 536718
rect 158432 536637 158632 536684
rect 158690 536718 158890 536734
rect 158690 536684 158706 536718
rect 158874 536684 158890 536718
rect 158690 536637 158890 536684
rect 158948 536718 159148 536734
rect 158948 536684 158964 536718
rect 159132 536684 159148 536718
rect 158948 536637 159148 536684
rect 159206 536718 159406 536734
rect 159206 536684 159222 536718
rect 159390 536684 159406 536718
rect 159206 536637 159406 536684
rect 159464 536718 159664 536734
rect 159464 536684 159480 536718
rect 159648 536684 159664 536718
rect 159464 536637 159664 536684
rect 159722 536718 159922 536734
rect 159722 536684 159738 536718
rect 159906 536684 159922 536718
rect 159722 536637 159922 536684
rect 159980 536718 160180 536734
rect 159980 536684 159996 536718
rect 160164 536684 160180 536718
rect 159980 536637 160180 536684
rect 160238 536718 160438 536734
rect 160238 536684 160254 536718
rect 160422 536684 160438 536718
rect 160238 536637 160438 536684
rect 160496 536718 160696 536734
rect 160496 536684 160512 536718
rect 160680 536684 160696 536718
rect 160496 536637 160696 536684
rect 160880 536718 161080 536734
rect 160880 536684 160896 536718
rect 161064 536684 161080 536718
rect 160880 536637 161080 536684
rect 161138 536718 161338 536734
rect 161138 536684 161154 536718
rect 161322 536684 161338 536718
rect 161138 536637 161338 536684
rect 161396 536718 161596 536734
rect 161396 536684 161412 536718
rect 161580 536684 161596 536718
rect 161396 536637 161596 536684
rect 161778 536718 161978 536734
rect 161778 536684 161794 536718
rect 161962 536684 161978 536718
rect 161778 536637 161978 536684
rect 162036 536718 162236 536734
rect 162036 536684 162052 536718
rect 162220 536684 162236 536718
rect 162036 536637 162236 536684
rect 162416 536718 162616 536734
rect 162416 536684 162432 536718
rect 162600 536684 162616 536718
rect 162416 536637 162616 536684
rect 157796 535990 157996 536037
rect 157796 535956 157812 535990
rect 157980 535956 157996 535990
rect 157796 535940 157996 535956
rect 158174 535990 158374 536037
rect 158174 535956 158190 535990
rect 158358 535956 158374 535990
rect 158174 535940 158374 535956
rect 158432 535990 158632 536037
rect 158432 535956 158448 535990
rect 158616 535956 158632 535990
rect 158432 535940 158632 535956
rect 158690 535990 158890 536037
rect 158690 535956 158706 535990
rect 158874 535956 158890 535990
rect 158690 535940 158890 535956
rect 158948 535990 159148 536037
rect 158948 535956 158964 535990
rect 159132 535956 159148 535990
rect 158948 535940 159148 535956
rect 159206 535990 159406 536037
rect 159206 535956 159222 535990
rect 159390 535956 159406 535990
rect 159206 535940 159406 535956
rect 159464 535990 159664 536037
rect 159464 535956 159480 535990
rect 159648 535956 159664 535990
rect 159464 535940 159664 535956
rect 159722 535990 159922 536037
rect 159722 535956 159738 535990
rect 159906 535956 159922 535990
rect 159722 535940 159922 535956
rect 159980 535990 160180 536037
rect 159980 535956 159996 535990
rect 160164 535956 160180 535990
rect 159980 535940 160180 535956
rect 160238 535990 160438 536037
rect 160238 535956 160254 535990
rect 160422 535956 160438 535990
rect 160238 535940 160438 535956
rect 160496 535990 160696 536037
rect 160496 535956 160512 535990
rect 160680 535956 160696 535990
rect 160496 535940 160696 535956
rect 160880 535990 161080 536037
rect 160880 535956 160896 535990
rect 161064 535956 161080 535990
rect 160880 535940 161080 535956
rect 161138 535990 161338 536037
rect 161138 535956 161154 535990
rect 161322 535956 161338 535990
rect 161138 535940 161338 535956
rect 161396 535990 161596 536037
rect 161396 535956 161412 535990
rect 161580 535956 161596 535990
rect 161396 535940 161596 535956
rect 161778 535990 161978 536037
rect 161778 535956 161794 535990
rect 161962 535956 161978 535990
rect 161778 535940 161978 535956
rect 162036 535990 162236 536037
rect 162036 535956 162052 535990
rect 162220 535956 162236 535990
rect 162036 535940 162236 535956
rect 162416 535990 162616 536037
rect 162416 535956 162432 535990
rect 162600 535956 162616 535990
rect 162416 535940 162616 535956
rect 172289 530564 172407 530590
rect 172573 530564 172603 530590
rect 172659 530564 172689 530590
rect 172745 530564 172775 530590
rect 172831 530564 172861 530590
rect 172928 530564 172958 530590
rect 173117 530564 174063 530590
rect 174221 530564 174615 530590
rect 174965 530564 174995 530590
rect 175051 530564 175081 530590
rect 175137 530564 175167 530590
rect 175223 530564 175253 530590
rect 175320 530564 175350 530590
rect 175601 530564 175631 530590
rect 175809 530564 175839 530590
rect 175900 530564 175930 530590
rect 176049 530564 176079 530590
rect 176145 530564 176175 530590
rect 176254 530564 176284 530590
rect 176353 530564 176383 530590
rect 176485 530564 176515 530590
rect 176557 530564 176587 530590
rect 176723 530564 176753 530590
rect 176819 530564 176849 530590
rect 176914 530564 176944 530590
rect 177169 530564 177199 530590
rect 177253 530564 177283 530590
rect 177736 530564 177766 530590
rect 177831 530564 177931 530590
rect 178089 530564 178189 530590
rect 178243 530564 178273 530590
rect 178453 530564 178483 530590
rect 178541 530564 178571 530590
rect 178737 530564 178767 530590
rect 178823 530564 178853 530590
rect 178909 530564 178939 530590
rect 178995 530564 179025 530590
rect 179092 530564 179122 530590
rect 179282 530564 179312 530590
rect 179379 530564 179409 530590
rect 179465 530564 179495 530590
rect 179551 530564 179581 530590
rect 179637 530564 179667 530590
rect 180293 530564 180323 530590
rect 180402 530564 180432 530590
rect 180498 530564 180528 530590
rect 180623 530564 180653 530590
rect 180719 530564 180749 530590
rect 180887 530564 180917 530590
rect 181259 530564 181289 530590
rect 181427 530564 181457 530590
rect 181523 530564 181553 530590
rect 181648 530564 181678 530590
rect 181744 530564 181774 530590
rect 181853 530564 181883 530590
rect 182042 530564 182072 530590
rect 182139 530564 182169 530590
rect 182225 530564 182255 530590
rect 182311 530564 182341 530590
rect 182397 530564 182427 530590
rect 182685 530564 182895 530590
rect 183146 530564 183176 530590
rect 183243 530564 183273 530590
rect 183329 530564 183359 530590
rect 183415 530564 183445 530590
rect 183501 530564 183531 530590
rect 183697 530564 184643 530590
rect 184801 530564 185011 530590
rect 185262 530564 185292 530590
rect 185359 530564 185389 530590
rect 185445 530564 185475 530590
rect 185531 530564 185561 530590
rect 185617 530564 185647 530590
rect 185813 530564 186759 530590
rect 172289 530428 172407 530454
rect 172369 530426 172407 530428
rect 172369 530410 172435 530426
rect 172261 530370 172327 530386
rect 172261 530336 172277 530370
rect 172311 530336 172327 530370
rect 172369 530376 172385 530410
rect 172419 530376 172435 530410
rect 172369 530360 172435 530376
rect 172573 530407 172603 530480
rect 172659 530407 172689 530480
rect 172745 530407 172775 530480
rect 172831 530407 172861 530480
rect 172928 530412 172958 530480
rect 173117 530428 174063 530454
rect 174221 530428 174615 530454
rect 172573 530401 172861 530407
rect 172573 530396 172862 530401
rect 172573 530374 172637 530396
rect 172574 530362 172637 530374
rect 172671 530362 172705 530396
rect 172739 530362 172773 530396
rect 172807 530362 172862 530396
rect 172261 530320 172327 530336
rect 172289 530318 172327 530320
rect 172574 530352 172862 530362
rect 172289 530288 172407 530318
rect 172574 530314 172604 530352
rect 172660 530314 172690 530352
rect 172746 530314 172776 530352
rect 172832 530314 172862 530352
rect 172909 530396 172969 530412
rect 172909 530362 172919 530396
rect 172953 530362 172969 530396
rect 173609 530406 174063 530428
rect 172909 530346 172969 530362
rect 173117 530370 173567 530386
rect 172928 530314 172958 530346
rect 173117 530336 173389 530370
rect 173423 530336 173567 530370
rect 173609 530372 173753 530406
rect 173787 530372 174063 530406
rect 174439 530406 174615 530428
rect 173609 530356 174063 530372
rect 174221 530370 174397 530386
rect 173117 530314 173567 530336
rect 174221 530336 174237 530370
rect 174271 530336 174347 530370
rect 174381 530336 174397 530370
rect 174439 530372 174455 530406
rect 174489 530372 174565 530406
rect 174599 530372 174615 530406
rect 174965 530407 174995 530480
rect 175051 530407 175081 530480
rect 175137 530407 175167 530480
rect 175223 530407 175253 530480
rect 175320 530412 175350 530480
rect 175601 530412 175631 530434
rect 174965 530401 175253 530407
rect 174965 530396 175254 530401
rect 174965 530374 175029 530396
rect 174439 530356 174615 530372
rect 174966 530362 175029 530374
rect 175063 530362 175097 530396
rect 175131 530362 175165 530396
rect 175199 530362 175254 530396
rect 174221 530314 174397 530336
rect 174966 530352 175254 530362
rect 174966 530314 174996 530352
rect 175052 530314 175082 530352
rect 175138 530314 175168 530352
rect 175224 530314 175254 530352
rect 175301 530396 175361 530412
rect 175301 530362 175311 530396
rect 175345 530362 175361 530396
rect 175301 530346 175361 530362
rect 175601 530396 175660 530412
rect 175601 530362 175616 530396
rect 175650 530362 175660 530396
rect 175601 530346 175660 530362
rect 175320 530314 175350 530346
rect 175601 530314 175631 530346
rect 173117 530288 174063 530314
rect 174221 530288 174615 530314
rect 175809 530312 175839 530480
rect 175900 530420 175930 530480
rect 176049 530448 176079 530480
rect 175977 530432 176079 530448
rect 175881 530404 175935 530420
rect 175881 530370 175891 530404
rect 175925 530370 175935 530404
rect 175977 530398 175987 530432
rect 176021 530418 176079 530432
rect 176145 530422 176175 530492
rect 176254 530470 176284 530492
rect 176021 530398 176038 530418
rect 175977 530382 176038 530398
rect 175881 530354 175935 530370
rect 175804 530296 175858 530312
rect 175804 530262 175814 530296
rect 175848 530262 175858 530296
rect 175804 530246 175858 530262
rect 175816 530198 175846 530246
rect 175900 530198 175930 530354
rect 176008 530198 176038 530382
rect 176121 530406 176175 530422
rect 176121 530372 176131 530406
rect 176165 530374 176175 530406
rect 176217 530454 176284 530470
rect 176217 530420 176227 530454
rect 176261 530420 176284 530454
rect 176485 530458 176515 530480
rect 176461 530442 176515 530458
rect 176217 530404 176284 530420
rect 176353 530410 176383 530436
rect 176353 530394 176419 530410
rect 176165 530372 176187 530374
rect 176121 530362 176187 530372
rect 176121 530356 176208 530362
rect 176145 530344 176208 530356
rect 176158 530332 176208 530344
rect 176082 530280 176136 530296
rect 176082 530246 176092 530280
rect 176126 530246 176136 530280
rect 176082 530230 176136 530246
rect 176092 530198 176122 530230
rect 176178 530198 176208 530332
rect 176353 530360 176375 530394
rect 176409 530360 176419 530394
rect 176461 530408 176471 530442
rect 176505 530408 176515 530442
rect 176461 530392 176515 530408
rect 176353 530344 176419 530360
rect 176353 530327 176383 530344
rect 176277 530297 176383 530327
rect 176277 530282 176307 530297
rect 176474 530198 176504 530392
rect 176557 530322 176587 530480
rect 176723 530458 176753 530492
rect 176819 530458 176849 530492
rect 176710 530448 176776 530458
rect 176710 530414 176726 530448
rect 176760 530414 176776 530448
rect 176710 530404 176776 530414
rect 176818 530442 176872 530458
rect 176818 530408 176828 530442
rect 176862 530408 176872 530442
rect 176818 530392 176872 530408
rect 176818 530362 176849 530392
rect 176711 530332 176849 530362
rect 176914 530351 176944 530480
rect 177169 530391 177199 530480
rect 177253 530465 177283 530480
rect 177253 530435 177316 530465
rect 177286 530412 177316 530435
rect 177736 530412 177766 530434
rect 177831 530412 177931 530480
rect 177286 530396 177340 530412
rect 177169 530381 177244 530391
rect 176914 530335 177031 530351
rect 176546 530306 176601 530322
rect 176546 530272 176557 530306
rect 176591 530272 176601 530306
rect 176546 530256 176601 530272
rect 176571 530198 176601 530256
rect 176711 530198 176741 530332
rect 176914 530315 176987 530335
rect 176902 530301 176987 530315
rect 177021 530301 177031 530335
rect 176790 530280 176856 530290
rect 176790 530246 176806 530280
rect 176840 530246 176856 530280
rect 176790 530236 176856 530246
rect 176902 530285 177031 530301
rect 177169 530347 177194 530381
rect 177228 530347 177244 530381
rect 177169 530337 177244 530347
rect 177286 530362 177296 530396
rect 177330 530362 177340 530396
rect 177286 530346 177340 530362
rect 177735 530396 177789 530412
rect 177735 530362 177745 530396
rect 177779 530362 177789 530396
rect 177735 530346 177789 530362
rect 177831 530396 177985 530412
rect 177831 530362 177941 530396
rect 177975 530362 177985 530396
rect 177831 530346 177985 530362
rect 178089 530396 178189 530480
rect 178089 530362 178145 530396
rect 178179 530362 178189 530396
rect 176810 530198 176840 530236
rect 176902 530198 176932 530285
rect 177169 530248 177199 530337
rect 177286 530293 177316 530346
rect 177736 530314 177766 530346
rect 177253 530263 177316 530293
rect 177253 530248 177283 530263
rect 172289 530088 172407 530114
rect 172574 530088 172604 530114
rect 172660 530088 172690 530114
rect 172746 530088 172776 530114
rect 172832 530088 172862 530114
rect 172928 530088 172958 530114
rect 173117 530088 174063 530114
rect 174221 530088 174615 530114
rect 174966 530088 174996 530114
rect 175052 530088 175082 530114
rect 175138 530088 175168 530114
rect 175224 530088 175254 530114
rect 175320 530088 175350 530114
rect 175601 530088 175631 530114
rect 175816 530088 175846 530114
rect 175900 530088 175930 530114
rect 176008 530088 176038 530114
rect 176092 530088 176122 530114
rect 176178 530088 176208 530114
rect 176277 530088 176307 530114
rect 176474 530088 176504 530114
rect 176571 530088 176601 530114
rect 176711 530088 176741 530114
rect 176810 530088 176840 530114
rect 176902 530088 176932 530114
rect 177169 530094 177199 530120
rect 177253 530094 177283 530120
rect 177831 530198 177931 530346
rect 178089 530198 178189 530362
rect 178243 530412 178273 530480
rect 178243 530396 178303 530412
rect 178453 530399 178483 530460
rect 178541 530445 178571 530460
rect 178541 530421 178577 530445
rect 178547 530412 178577 530421
rect 178243 530362 178259 530396
rect 178293 530362 178303 530396
rect 178243 530346 178303 530362
rect 178449 530383 178503 530399
rect 178449 530349 178459 530383
rect 178493 530349 178503 530383
rect 178243 530198 178273 530346
rect 178449 530333 178503 530349
rect 178547 530396 178623 530412
rect 178547 530362 178579 530396
rect 178613 530362 178623 530396
rect 178737 530407 178767 530480
rect 178823 530407 178853 530480
rect 178909 530407 178939 530480
rect 178995 530407 179025 530480
rect 179092 530412 179122 530480
rect 179282 530412 179312 530480
rect 178737 530401 179025 530407
rect 178737 530396 179026 530401
rect 178737 530374 178801 530396
rect 178547 530346 178623 530362
rect 178738 530362 178801 530374
rect 178835 530362 178869 530396
rect 178903 530362 178937 530396
rect 178971 530362 179026 530396
rect 178738 530352 179026 530362
rect 178453 530272 178483 530333
rect 178547 530311 178577 530346
rect 178738 530314 178768 530352
rect 178824 530314 178854 530352
rect 178910 530314 178940 530352
rect 178996 530314 179026 530352
rect 179073 530396 179133 530412
rect 179073 530362 179083 530396
rect 179117 530362 179133 530396
rect 179073 530346 179133 530362
rect 179271 530396 179331 530412
rect 179379 530407 179409 530480
rect 179465 530407 179495 530480
rect 179551 530407 179581 530480
rect 179637 530407 179667 530480
rect 180293 530412 180323 530434
rect 180402 530412 180432 530480
rect 180498 530448 180528 530480
rect 180623 530448 180653 530480
rect 180498 530432 180581 530448
rect 179379 530401 179667 530407
rect 179271 530362 179287 530396
rect 179321 530362 179331 530396
rect 179271 530346 179331 530362
rect 179378 530396 179667 530401
rect 179378 530362 179433 530396
rect 179467 530362 179501 530396
rect 179535 530362 179569 530396
rect 179603 530374 179667 530396
rect 180290 530396 180344 530412
rect 179603 530362 179666 530374
rect 179378 530352 179666 530362
rect 179092 530314 179122 530346
rect 179282 530314 179312 530346
rect 179378 530314 179408 530352
rect 179464 530314 179494 530352
rect 179550 530314 179580 530352
rect 179636 530314 179666 530352
rect 180290 530362 180300 530396
rect 180334 530362 180344 530396
rect 180290 530346 180344 530362
rect 180386 530396 180440 530412
rect 180386 530362 180396 530396
rect 180430 530362 180440 530396
rect 180498 530398 180537 530432
rect 180571 530398 180581 530432
rect 180498 530382 180581 530398
rect 180623 530432 180677 530448
rect 180623 530398 180633 530432
rect 180667 530398 180677 530432
rect 180719 530442 180749 530480
rect 180719 530432 180845 530442
rect 180719 530412 180795 530432
rect 180623 530382 180677 530398
rect 180779 530398 180795 530412
rect 180829 530398 180845 530432
rect 180779 530388 180845 530398
rect 180386 530346 180440 530362
rect 180293 530314 180323 530346
rect 178541 530287 178577 530311
rect 178541 530272 178571 530287
rect 180402 530237 180432 530346
rect 180623 530282 180653 530382
rect 180505 530252 180653 530282
rect 180695 530319 180749 530335
rect 180695 530285 180705 530319
rect 180739 530285 180749 530319
rect 180695 530269 180749 530285
rect 180505 530237 180535 530252
rect 180719 530237 180749 530269
rect 180791 530237 180821 530388
rect 180887 530335 180917 530480
rect 180863 530319 180917 530335
rect 180863 530285 180873 530319
rect 180907 530285 180917 530319
rect 180863 530269 180917 530285
rect 180887 530237 180917 530269
rect 181259 530335 181289 530480
rect 181427 530442 181457 530480
rect 181523 530448 181553 530480
rect 181648 530448 181678 530480
rect 181331 530432 181457 530442
rect 181331 530398 181347 530432
rect 181381 530412 181457 530432
rect 181499 530432 181553 530448
rect 181381 530398 181397 530412
rect 181331 530388 181397 530398
rect 181499 530398 181509 530432
rect 181543 530398 181553 530432
rect 181259 530319 181313 530335
rect 181259 530285 181269 530319
rect 181303 530285 181313 530319
rect 181259 530269 181313 530285
rect 181259 530237 181289 530269
rect 181355 530237 181385 530388
rect 181499 530382 181553 530398
rect 181595 530432 181678 530448
rect 181595 530398 181605 530432
rect 181639 530398 181678 530432
rect 181744 530412 181774 530480
rect 181853 530412 181883 530434
rect 182042 530412 182072 530480
rect 181595 530382 181678 530398
rect 181736 530396 181790 530412
rect 181427 530319 181481 530335
rect 181427 530285 181437 530319
rect 181471 530285 181481 530319
rect 181427 530269 181481 530285
rect 181523 530282 181553 530382
rect 181736 530362 181746 530396
rect 181780 530362 181790 530396
rect 181736 530346 181790 530362
rect 181832 530396 181886 530412
rect 181832 530362 181842 530396
rect 181876 530362 181886 530396
rect 181832 530346 181886 530362
rect 182031 530396 182091 530412
rect 182139 530407 182169 530480
rect 182225 530407 182255 530480
rect 182311 530407 182341 530480
rect 182397 530407 182427 530480
rect 182685 530428 182895 530454
rect 182139 530401 182427 530407
rect 182031 530362 182047 530396
rect 182081 530362 182091 530396
rect 182031 530346 182091 530362
rect 182138 530396 182427 530401
rect 182138 530362 182193 530396
rect 182227 530362 182261 530396
rect 182295 530362 182329 530396
rect 182363 530374 182427 530396
rect 182811 530422 182895 530428
rect 182811 530406 182953 530422
rect 183146 530412 183176 530480
rect 182363 530362 182426 530374
rect 182138 530352 182426 530362
rect 181427 530237 181457 530269
rect 181523 530252 181671 530282
rect 181641 530237 181671 530252
rect 181744 530237 181774 530346
rect 181853 530314 181883 530346
rect 182042 530314 182072 530346
rect 182138 530314 182168 530352
rect 182224 530314 182254 530352
rect 182310 530314 182340 530352
rect 182396 530314 182426 530352
rect 182627 530370 182769 530386
rect 182627 530336 182643 530370
rect 182677 530336 182769 530370
rect 182811 530372 182903 530406
rect 182937 530372 182953 530406
rect 182811 530356 182953 530372
rect 183135 530396 183195 530412
rect 183243 530407 183273 530480
rect 183329 530407 183359 530480
rect 183415 530407 183445 530480
rect 183501 530407 183531 530480
rect 183697 530428 184643 530454
rect 184801 530428 185011 530454
rect 183243 530401 183531 530407
rect 183135 530362 183151 530396
rect 183185 530362 183195 530396
rect 183135 530346 183195 530362
rect 183242 530396 183531 530401
rect 183242 530362 183297 530396
rect 183331 530362 183365 530396
rect 183399 530362 183433 530396
rect 183467 530374 183531 530396
rect 184189 530406 184643 530428
rect 183467 530362 183530 530374
rect 183242 530352 183530 530362
rect 182627 530320 182769 530336
rect 182685 530314 182769 530320
rect 183146 530314 183176 530346
rect 183242 530314 183272 530352
rect 183328 530314 183358 530352
rect 183414 530314 183444 530352
rect 183500 530314 183530 530352
rect 183697 530370 184147 530386
rect 183697 530336 183969 530370
rect 184003 530336 184147 530370
rect 184189 530372 184333 530406
rect 184367 530372 184643 530406
rect 184927 530422 185011 530428
rect 184927 530406 185069 530422
rect 185262 530412 185292 530480
rect 184189 530356 184643 530372
rect 184743 530370 184885 530386
rect 183697 530314 184147 530336
rect 184743 530336 184759 530370
rect 184793 530336 184885 530370
rect 184927 530372 185019 530406
rect 185053 530372 185069 530406
rect 184927 530356 185069 530372
rect 185251 530396 185311 530412
rect 185359 530407 185389 530480
rect 185445 530407 185475 530480
rect 185531 530407 185561 530480
rect 185617 530407 185647 530480
rect 186951 530560 187047 530590
rect 186951 530526 187001 530560
rect 187035 530526 187047 530560
rect 186951 530492 187047 530526
rect 186951 530458 187001 530492
rect 187035 530458 187047 530492
rect 185813 530428 186759 530454
rect 185359 530401 185647 530407
rect 185251 530362 185267 530396
rect 185301 530362 185311 530396
rect 185251 530346 185311 530362
rect 185358 530396 185647 530401
rect 185358 530362 185413 530396
rect 185447 530362 185481 530396
rect 185515 530362 185549 530396
rect 185583 530374 185647 530396
rect 186305 530406 186759 530428
rect 185583 530362 185646 530374
rect 185358 530352 185646 530362
rect 184743 530320 184885 530336
rect 184801 530314 184885 530320
rect 185262 530314 185292 530346
rect 185358 530314 185388 530352
rect 185444 530314 185474 530352
rect 185530 530314 185560 530352
rect 185616 530314 185646 530352
rect 185813 530370 186263 530386
rect 185813 530336 186085 530370
rect 186119 530336 186263 530370
rect 186305 530372 186449 530406
rect 186483 530372 186759 530406
rect 186305 530356 186759 530372
rect 186951 530379 187047 530458
rect 185813 530314 186263 530336
rect 180402 530127 180432 530153
rect 180505 530127 180535 530153
rect 180719 530127 180749 530153
rect 180791 530127 180821 530153
rect 180887 530127 180917 530153
rect 181259 530127 181289 530153
rect 181355 530127 181385 530153
rect 181427 530127 181457 530153
rect 181641 530127 181671 530153
rect 181744 530127 181774 530153
rect 182685 530288 182895 530314
rect 183697 530288 184643 530314
rect 184801 530288 185011 530314
rect 185813 530288 186759 530314
rect 186951 530229 187047 530370
rect 186951 530195 187001 530229
rect 187035 530195 187047 530229
rect 186951 530161 187047 530195
rect 186951 530127 187001 530161
rect 187035 530127 187047 530161
rect 177736 530088 177766 530114
rect 177831 530088 177931 530114
rect 178089 530088 178189 530114
rect 178243 530088 178273 530114
rect 178453 530088 178483 530114
rect 178541 530088 178571 530114
rect 178738 530088 178768 530114
rect 178824 530088 178854 530114
rect 178910 530088 178940 530114
rect 178996 530088 179026 530114
rect 179092 530088 179122 530114
rect 179282 530088 179312 530114
rect 179378 530088 179408 530114
rect 179464 530088 179494 530114
rect 179550 530088 179580 530114
rect 179636 530088 179666 530114
rect 180293 530088 180323 530114
rect 181853 530088 181883 530114
rect 182042 530088 182072 530114
rect 182138 530088 182168 530114
rect 182224 530088 182254 530114
rect 182310 530088 182340 530114
rect 182396 530088 182426 530114
rect 182685 530088 182895 530114
rect 183146 530088 183176 530114
rect 183242 530088 183272 530114
rect 183328 530088 183358 530114
rect 183414 530088 183444 530114
rect 183500 530088 183530 530114
rect 183697 530088 184643 530114
rect 184801 530088 185011 530114
rect 185262 530088 185292 530114
rect 185358 530088 185388 530114
rect 185444 530088 185474 530114
rect 185530 530088 185560 530114
rect 185616 530088 185646 530114
rect 185813 530088 186759 530114
rect 186951 530088 187047 530127
rect 187089 530564 187185 530590
rect 187285 530564 187403 530590
rect 187089 530530 187101 530564
rect 187135 530530 187185 530564
rect 187089 530496 187185 530530
rect 187089 530462 187101 530496
rect 187135 530462 187185 530496
rect 187089 530379 187185 530462
rect 187285 530428 187403 530454
rect 187285 530426 187323 530428
rect 187089 530229 187185 530370
rect 187257 530410 187323 530426
rect 187257 530376 187273 530410
rect 187307 530376 187323 530410
rect 187257 530360 187323 530376
rect 187365 530370 187431 530386
rect 187365 530336 187381 530370
rect 187415 530336 187431 530370
rect 187365 530320 187431 530336
rect 187365 530318 187403 530320
rect 187285 530288 187403 530318
rect 187089 530195 187101 530229
rect 187135 530195 187185 530229
rect 187089 530161 187185 530195
rect 187089 530127 187101 530161
rect 187135 530127 187185 530161
rect 187089 530088 187185 530127
rect 187285 530088 187403 530114
rect 172289 530020 172407 530046
rect 172565 530020 173511 530046
rect 173669 530020 174615 530046
rect 174887 530020 174917 530046
rect 174971 530020 175071 530046
rect 175229 530020 175329 530046
rect 175394 530020 175424 530046
rect 172289 529816 172407 529846
rect 172565 529820 173511 529846
rect 173669 529820 174615 529846
rect 172289 529814 172327 529816
rect 172261 529798 172327 529814
rect 172261 529764 172277 529798
rect 172311 529764 172327 529798
rect 172565 529798 173015 529820
rect 172261 529748 172327 529764
rect 172369 529758 172435 529774
rect 172369 529724 172385 529758
rect 172419 529724 172435 529758
rect 172565 529764 172837 529798
rect 172871 529764 173015 529798
rect 173669 529798 174119 529820
rect 172565 529748 173015 529764
rect 173057 529762 173511 529778
rect 172369 529708 172435 529724
rect 173057 529728 173201 529762
rect 173235 529728 173511 529762
rect 173669 529764 173941 529798
rect 173975 529764 174119 529798
rect 174887 529788 174917 529936
rect 173669 529748 174119 529764
rect 174161 529762 174615 529778
rect 172369 529706 172407 529708
rect 173057 529706 173511 529728
rect 174161 529728 174305 529762
rect 174339 529728 174615 529762
rect 174161 529706 174615 529728
rect 174857 529772 174917 529788
rect 174857 529738 174867 529772
rect 174901 529738 174917 529772
rect 174857 529722 174917 529738
rect 172289 529680 172407 529706
rect 172565 529680 173511 529706
rect 173669 529680 174615 529706
rect 174887 529654 174917 529722
rect 174971 529772 175071 529936
rect 175229 529788 175329 529936
rect 175601 530014 175631 530040
rect 175685 530014 175715 530040
rect 175952 530020 175982 530046
rect 176044 530020 176074 530046
rect 176143 530020 176173 530046
rect 176283 530020 176313 530046
rect 176380 530020 176410 530046
rect 176577 530020 176607 530046
rect 176676 530020 176706 530046
rect 176762 530020 176792 530046
rect 176846 530020 176876 530046
rect 176954 530020 176984 530046
rect 177038 530020 177068 530046
rect 177253 530020 177283 530046
rect 178265 530020 178295 530046
rect 178453 530020 178483 530046
rect 178668 530020 178698 530046
rect 178752 530020 178782 530046
rect 178860 530020 178890 530046
rect 178944 530020 178974 530046
rect 179030 530020 179060 530046
rect 179129 530020 179159 530046
rect 179326 530020 179356 530046
rect 179423 530020 179453 530046
rect 179563 530020 179593 530046
rect 179662 530020 179692 530046
rect 179754 530020 179784 530046
rect 175601 529871 175631 529886
rect 175568 529841 175631 529871
rect 175394 529788 175424 529820
rect 175568 529788 175598 529841
rect 175685 529797 175715 529886
rect 175952 529849 175982 529936
rect 176044 529898 176074 529936
rect 174971 529738 174981 529772
rect 175015 529738 175071 529772
rect 174971 529654 175071 529738
rect 175175 529772 175329 529788
rect 175175 529738 175185 529772
rect 175219 529738 175329 529772
rect 175175 529722 175329 529738
rect 175371 529772 175425 529788
rect 175371 529738 175381 529772
rect 175415 529738 175425 529772
rect 175371 529722 175425 529738
rect 175544 529772 175598 529788
rect 175544 529738 175554 529772
rect 175588 529738 175598 529772
rect 175640 529787 175715 529797
rect 175640 529753 175656 529787
rect 175690 529753 175715 529787
rect 175853 529833 175982 529849
rect 176028 529888 176094 529898
rect 176028 529854 176044 529888
rect 176078 529854 176094 529888
rect 176028 529844 176094 529854
rect 175853 529799 175863 529833
rect 175897 529819 175982 529833
rect 175897 529799 175970 529819
rect 176143 529802 176173 529936
rect 176283 529878 176313 529936
rect 176283 529862 176338 529878
rect 176283 529828 176293 529862
rect 176327 529828 176338 529862
rect 176283 529812 176338 529828
rect 175853 529783 175970 529799
rect 175640 529743 175715 529753
rect 175544 529722 175598 529738
rect 175229 529654 175329 529722
rect 175394 529700 175424 529722
rect 175568 529699 175598 529722
rect 175568 529669 175631 529699
rect 175601 529654 175631 529669
rect 175685 529654 175715 529743
rect 175940 529654 175970 529783
rect 176035 529772 176173 529802
rect 176035 529742 176066 529772
rect 176012 529726 176066 529742
rect 176012 529692 176022 529726
rect 176056 529692 176066 529726
rect 176012 529676 176066 529692
rect 176108 529720 176174 529730
rect 176108 529686 176124 529720
rect 176158 529686 176174 529720
rect 176108 529676 176174 529686
rect 176035 529642 176065 529676
rect 176131 529642 176161 529676
rect 176297 529654 176327 529812
rect 176380 529742 176410 529936
rect 176577 529837 176607 529852
rect 176501 529807 176607 529837
rect 176501 529790 176531 529807
rect 176465 529774 176531 529790
rect 176369 529726 176423 529742
rect 176369 529692 176379 529726
rect 176413 529692 176423 529726
rect 176465 529740 176475 529774
rect 176509 529740 176531 529774
rect 176676 529802 176706 529936
rect 176762 529904 176792 529936
rect 176748 529888 176802 529904
rect 176748 529854 176758 529888
rect 176792 529854 176802 529888
rect 176748 529838 176802 529854
rect 176676 529790 176726 529802
rect 176676 529778 176739 529790
rect 176676 529772 176763 529778
rect 176697 529762 176763 529772
rect 176697 529760 176719 529762
rect 176465 529724 176531 529740
rect 176501 529698 176531 529724
rect 176600 529714 176667 529730
rect 176369 529676 176423 529692
rect 176369 529654 176399 529676
rect 176600 529680 176623 529714
rect 176657 529680 176667 529714
rect 176600 529664 176667 529680
rect 176709 529728 176719 529760
rect 176753 529728 176763 529762
rect 176709 529712 176763 529728
rect 176846 529752 176876 529936
rect 176954 529780 176984 529936
rect 177038 529888 177068 529936
rect 177026 529872 177080 529888
rect 177026 529838 177036 529872
rect 177070 529838 177080 529872
rect 177026 529822 177080 529838
rect 176949 529764 177003 529780
rect 176846 529736 176907 529752
rect 176846 529716 176863 529736
rect 176600 529642 176630 529664
rect 176709 529642 176739 529712
rect 176805 529702 176863 529716
rect 176897 529702 176907 529736
rect 176949 529730 176959 529764
rect 176993 529730 177003 529764
rect 176949 529714 177003 529730
rect 176805 529686 176907 529702
rect 176805 529654 176835 529686
rect 176954 529654 176984 529714
rect 177045 529654 177075 529822
rect 177671 529981 177701 530007
rect 177767 529981 177797 530007
rect 177839 529981 177869 530007
rect 178053 529981 178083 530007
rect 178156 529981 178186 530007
rect 177671 529865 177701 529897
rect 177671 529849 177725 529865
rect 177253 529788 177283 529820
rect 177224 529772 177283 529788
rect 177224 529738 177234 529772
rect 177268 529738 177283 529772
rect 177224 529722 177283 529738
rect 177253 529700 177283 529722
rect 177671 529815 177681 529849
rect 177715 529815 177725 529849
rect 177671 529799 177725 529815
rect 177671 529654 177701 529799
rect 177767 529746 177797 529897
rect 177839 529865 177869 529897
rect 178053 529882 178083 529897
rect 177839 529849 177893 529865
rect 177839 529815 177849 529849
rect 177883 529815 177893 529849
rect 177839 529799 177893 529815
rect 177935 529852 178083 529882
rect 177935 529752 177965 529852
rect 178156 529788 178186 529897
rect 178668 529888 178698 529936
rect 178656 529872 178710 529888
rect 178656 529838 178666 529872
rect 178700 529838 178710 529872
rect 178656 529822 178710 529838
rect 178265 529788 178295 529820
rect 178453 529788 178483 529820
rect 178148 529772 178202 529788
rect 177743 529736 177809 529746
rect 177743 529702 177759 529736
rect 177793 529722 177809 529736
rect 177911 529736 177965 529752
rect 177793 529702 177869 529722
rect 177743 529692 177869 529702
rect 177839 529654 177869 529692
rect 177911 529702 177921 529736
rect 177955 529702 177965 529736
rect 177911 529686 177965 529702
rect 178007 529736 178090 529752
rect 178007 529702 178017 529736
rect 178051 529702 178090 529736
rect 178148 529738 178158 529772
rect 178192 529738 178202 529772
rect 178148 529722 178202 529738
rect 178244 529772 178298 529788
rect 178244 529738 178254 529772
rect 178288 529738 178298 529772
rect 178244 529722 178298 529738
rect 178453 529772 178512 529788
rect 178453 529738 178468 529772
rect 178502 529738 178512 529772
rect 178453 529722 178512 529738
rect 178007 529686 178090 529702
rect 177935 529654 177965 529686
rect 178060 529654 178090 529686
rect 178156 529654 178186 529722
rect 178265 529700 178295 529722
rect 178453 529700 178483 529722
rect 178661 529654 178691 529822
rect 178752 529780 178782 529936
rect 178733 529764 178787 529780
rect 178733 529730 178743 529764
rect 178777 529730 178787 529764
rect 178860 529752 178890 529936
rect 178944 529904 178974 529936
rect 178934 529888 178988 529904
rect 178934 529854 178944 529888
rect 178978 529854 178988 529888
rect 178934 529838 178988 529854
rect 179030 529802 179060 529936
rect 180021 530014 180051 530040
rect 180105 530014 180135 530040
rect 180293 530014 180323 530040
rect 180377 530014 180407 530040
rect 180644 530020 180674 530046
rect 180736 530020 180766 530046
rect 180835 530020 180865 530046
rect 180975 530020 181005 530046
rect 181072 530020 181102 530046
rect 181269 530020 181299 530046
rect 181368 530020 181398 530046
rect 181454 530020 181484 530046
rect 181538 530020 181568 530046
rect 181646 530020 181676 530046
rect 181730 530020 181760 530046
rect 181945 530020 181975 530046
rect 182133 530020 182343 530046
rect 182704 530020 182734 530046
rect 182799 530020 182899 530046
rect 183057 530020 183157 530046
rect 183211 530020 183241 530046
rect 183421 530020 184367 530046
rect 184525 530020 185471 530046
rect 185629 530020 186575 530046
rect 186733 530020 187127 530046
rect 187285 530020 187403 530046
rect 179129 529837 179159 529852
rect 179129 529807 179235 529837
rect 179010 529790 179060 529802
rect 178997 529778 179060 529790
rect 178733 529714 178787 529730
rect 178829 529736 178890 529752
rect 178752 529654 178782 529714
rect 178829 529702 178839 529736
rect 178873 529716 178890 529736
rect 178973 529772 179060 529778
rect 179205 529790 179235 529807
rect 179205 529774 179271 529790
rect 178973 529762 179039 529772
rect 178973 529728 178983 529762
rect 179017 529760 179039 529762
rect 179017 529728 179027 529760
rect 179205 529740 179227 529774
rect 179261 529740 179271 529774
rect 179326 529742 179356 529936
rect 179423 529878 179453 529936
rect 179398 529862 179453 529878
rect 179398 529828 179409 529862
rect 179443 529828 179453 529862
rect 179398 529812 179453 529828
rect 178873 529702 178931 529716
rect 178973 529712 179027 529728
rect 178829 529686 178931 529702
rect 178901 529654 178931 529686
rect 178997 529642 179027 529712
rect 179069 529714 179136 529730
rect 179069 529680 179079 529714
rect 179113 529680 179136 529714
rect 179205 529724 179271 529740
rect 179313 529726 179367 529742
rect 179205 529698 179235 529724
rect 179069 529664 179136 529680
rect 179106 529642 179136 529664
rect 179313 529692 179323 529726
rect 179357 529692 179367 529726
rect 179313 529676 179367 529692
rect 179337 529654 179367 529676
rect 179409 529654 179439 529812
rect 179563 529802 179593 529936
rect 179662 529898 179692 529936
rect 179642 529888 179708 529898
rect 179642 529854 179658 529888
rect 179692 529854 179708 529888
rect 179642 529844 179708 529854
rect 179754 529849 179784 529936
rect 179754 529833 179883 529849
rect 179754 529819 179839 529833
rect 179563 529772 179701 529802
rect 179670 529742 179701 529772
rect 179766 529799 179839 529819
rect 179873 529799 179883 529833
rect 179766 529783 179883 529799
rect 180021 529797 180051 529886
rect 180105 529871 180135 529886
rect 180293 529871 180323 529886
rect 180105 529841 180168 529871
rect 180021 529787 180096 529797
rect 179562 529720 179628 529730
rect 179562 529686 179578 529720
rect 179612 529686 179628 529720
rect 179562 529676 179628 529686
rect 179670 529726 179724 529742
rect 179670 529692 179680 529726
rect 179714 529692 179724 529726
rect 179670 529676 179724 529692
rect 179575 529642 179605 529676
rect 179671 529642 179701 529676
rect 179766 529654 179796 529783
rect 180021 529753 180046 529787
rect 180080 529753 180096 529787
rect 180021 529743 180096 529753
rect 180138 529788 180168 529841
rect 180260 529841 180323 529871
rect 180260 529788 180290 529841
rect 180377 529797 180407 529886
rect 180644 529849 180674 529936
rect 180736 529898 180766 529936
rect 180138 529772 180192 529788
rect 180021 529654 180051 529743
rect 180138 529738 180148 529772
rect 180182 529738 180192 529772
rect 180138 529722 180192 529738
rect 180236 529772 180290 529788
rect 180236 529738 180246 529772
rect 180280 529738 180290 529772
rect 180332 529787 180407 529797
rect 180332 529753 180348 529787
rect 180382 529753 180407 529787
rect 180545 529833 180674 529849
rect 180720 529888 180786 529898
rect 180720 529854 180736 529888
rect 180770 529854 180786 529888
rect 180720 529844 180786 529854
rect 180545 529799 180555 529833
rect 180589 529819 180674 529833
rect 180589 529799 180662 529819
rect 180835 529802 180865 529936
rect 180975 529878 181005 529936
rect 180975 529862 181030 529878
rect 180975 529828 180985 529862
rect 181019 529828 181030 529862
rect 180975 529812 181030 529828
rect 180545 529783 180662 529799
rect 180332 529743 180407 529753
rect 180236 529722 180290 529738
rect 180138 529699 180168 529722
rect 180105 529669 180168 529699
rect 180260 529699 180290 529722
rect 180260 529669 180323 529699
rect 180105 529654 180135 529669
rect 180293 529654 180323 529669
rect 180377 529654 180407 529743
rect 180632 529654 180662 529783
rect 180727 529772 180865 529802
rect 180727 529742 180758 529772
rect 180704 529726 180758 529742
rect 180704 529692 180714 529726
rect 180748 529692 180758 529726
rect 180704 529676 180758 529692
rect 180800 529720 180866 529730
rect 180800 529686 180816 529720
rect 180850 529686 180866 529720
rect 180800 529676 180866 529686
rect 180727 529642 180757 529676
rect 180823 529642 180853 529676
rect 180989 529654 181019 529812
rect 181072 529742 181102 529936
rect 181269 529837 181299 529852
rect 181193 529807 181299 529837
rect 181193 529790 181223 529807
rect 181157 529774 181223 529790
rect 181061 529726 181115 529742
rect 181061 529692 181071 529726
rect 181105 529692 181115 529726
rect 181157 529740 181167 529774
rect 181201 529740 181223 529774
rect 181368 529802 181398 529936
rect 181454 529904 181484 529936
rect 181440 529888 181494 529904
rect 181440 529854 181450 529888
rect 181484 529854 181494 529888
rect 181440 529838 181494 529854
rect 181368 529790 181418 529802
rect 181368 529778 181431 529790
rect 181368 529772 181455 529778
rect 181389 529762 181455 529772
rect 181389 529760 181411 529762
rect 181157 529724 181223 529740
rect 181193 529698 181223 529724
rect 181292 529714 181359 529730
rect 181061 529676 181115 529692
rect 181061 529654 181091 529676
rect 181292 529680 181315 529714
rect 181349 529680 181359 529714
rect 181292 529664 181359 529680
rect 181401 529728 181411 529760
rect 181445 529728 181455 529762
rect 181401 529712 181455 529728
rect 181538 529752 181568 529936
rect 181646 529780 181676 529936
rect 181730 529888 181760 529936
rect 181718 529872 181772 529888
rect 181718 529838 181728 529872
rect 181762 529838 181772 529872
rect 181718 529822 181772 529838
rect 181641 529764 181695 529780
rect 181538 529736 181599 529752
rect 181538 529716 181555 529736
rect 181292 529642 181322 529664
rect 181401 529642 181431 529712
rect 181497 529702 181555 529716
rect 181589 529702 181599 529736
rect 181641 529730 181651 529764
rect 181685 529730 181695 529764
rect 181641 529714 181695 529730
rect 181497 529686 181599 529702
rect 181497 529654 181527 529686
rect 181646 529654 181676 529714
rect 181737 529654 181767 529822
rect 182133 529820 182343 529846
rect 181945 529788 181975 529820
rect 182133 529814 182217 529820
rect 181916 529772 181975 529788
rect 181916 529738 181926 529772
rect 181960 529738 181975 529772
rect 182075 529798 182217 529814
rect 182075 529764 182091 529798
rect 182125 529764 182217 529798
rect 182704 529788 182734 529820
rect 182799 529788 182899 529936
rect 182075 529748 182217 529764
rect 182259 529762 182401 529778
rect 181916 529722 181975 529738
rect 181945 529700 181975 529722
rect 182259 529728 182351 529762
rect 182385 529728 182401 529762
rect 182259 529712 182401 529728
rect 182703 529772 182757 529788
rect 182703 529738 182713 529772
rect 182747 529738 182757 529772
rect 182703 529722 182757 529738
rect 182799 529772 182953 529788
rect 182799 529738 182909 529772
rect 182943 529738 182953 529772
rect 182799 529722 182953 529738
rect 183057 529772 183157 529936
rect 183057 529738 183113 529772
rect 183147 529738 183157 529772
rect 182259 529706 182343 529712
rect 182133 529680 182343 529706
rect 182704 529700 182734 529722
rect 182799 529654 182899 529722
rect 183057 529654 183157 529738
rect 183211 529788 183241 529936
rect 183421 529820 184367 529846
rect 184525 529820 185471 529846
rect 185629 529820 186575 529846
rect 186733 529820 187127 529846
rect 183421 529798 183871 529820
rect 183211 529772 183271 529788
rect 183211 529738 183227 529772
rect 183261 529738 183271 529772
rect 183421 529764 183693 529798
rect 183727 529764 183871 529798
rect 184525 529798 184975 529820
rect 183421 529748 183871 529764
rect 183913 529762 184367 529778
rect 183211 529722 183271 529738
rect 183913 529728 184057 529762
rect 184091 529728 184367 529762
rect 184525 529764 184797 529798
rect 184831 529764 184975 529798
rect 185629 529798 186079 529820
rect 184525 529748 184975 529764
rect 185017 529762 185471 529778
rect 183211 529654 183241 529722
rect 183913 529706 184367 529728
rect 185017 529728 185161 529762
rect 185195 529728 185471 529762
rect 185629 529764 185901 529798
rect 185935 529764 186079 529798
rect 186733 529798 186909 529820
rect 187285 529816 187403 529846
rect 185629 529748 186079 529764
rect 186121 529762 186575 529778
rect 185017 529706 185471 529728
rect 186121 529728 186265 529762
rect 186299 529728 186575 529762
rect 186733 529764 186749 529798
rect 186783 529764 186859 529798
rect 186893 529764 186909 529798
rect 187365 529814 187403 529816
rect 187365 529798 187431 529814
rect 186733 529748 186909 529764
rect 186951 529762 187127 529778
rect 186121 529706 186575 529728
rect 186951 529728 186967 529762
rect 187001 529728 187077 529762
rect 187111 529728 187127 529762
rect 186951 529706 187127 529728
rect 187257 529758 187323 529774
rect 187257 529724 187273 529758
rect 187307 529724 187323 529758
rect 187365 529764 187381 529798
rect 187415 529764 187431 529798
rect 187365 529748 187431 529764
rect 187257 529708 187323 529724
rect 183421 529680 184367 529706
rect 184525 529680 185471 529706
rect 185629 529680 186575 529706
rect 186733 529680 187127 529706
rect 187285 529706 187323 529708
rect 187285 529680 187403 529706
rect 172289 529544 172407 529570
rect 172565 529544 173511 529570
rect 173669 529544 174615 529570
rect 174887 529544 174917 529570
rect 174971 529544 175071 529570
rect 175229 529544 175329 529570
rect 175394 529544 175424 529570
rect 175601 529544 175631 529570
rect 175685 529544 175715 529570
rect 175940 529544 175970 529570
rect 176035 529544 176065 529570
rect 176131 529544 176161 529570
rect 176297 529544 176327 529570
rect 176369 529544 176399 529570
rect 176501 529544 176531 529570
rect 176600 529544 176630 529570
rect 176709 529544 176739 529570
rect 176805 529544 176835 529570
rect 176954 529544 176984 529570
rect 177045 529544 177075 529570
rect 177253 529544 177283 529570
rect 177671 529544 177701 529570
rect 177839 529544 177869 529570
rect 177935 529544 177965 529570
rect 178060 529544 178090 529570
rect 178156 529544 178186 529570
rect 178265 529544 178295 529570
rect 178453 529544 178483 529570
rect 178661 529544 178691 529570
rect 178752 529544 178782 529570
rect 178901 529544 178931 529570
rect 178997 529544 179027 529570
rect 179106 529544 179136 529570
rect 179205 529544 179235 529570
rect 179337 529544 179367 529570
rect 179409 529544 179439 529570
rect 179575 529544 179605 529570
rect 179671 529544 179701 529570
rect 179766 529544 179796 529570
rect 180021 529544 180051 529570
rect 180105 529544 180135 529570
rect 180293 529544 180323 529570
rect 180377 529544 180407 529570
rect 180632 529544 180662 529570
rect 180727 529544 180757 529570
rect 180823 529544 180853 529570
rect 180989 529544 181019 529570
rect 181061 529544 181091 529570
rect 181193 529544 181223 529570
rect 181292 529544 181322 529570
rect 181401 529544 181431 529570
rect 181497 529544 181527 529570
rect 181646 529544 181676 529570
rect 181737 529544 181767 529570
rect 181945 529544 181975 529570
rect 182133 529544 182343 529570
rect 182704 529544 182734 529570
rect 182799 529544 182899 529570
rect 183057 529544 183157 529570
rect 183211 529544 183241 529570
rect 183421 529544 184367 529570
rect 184525 529544 185471 529570
rect 185629 529544 186575 529570
rect 186733 529544 187127 529570
rect 187285 529544 187403 529570
rect 172289 529476 172407 529502
rect 172565 529476 173511 529502
rect 173669 529476 174615 529502
rect 175187 529476 175217 529502
rect 175355 529476 175385 529502
rect 175451 529476 175481 529502
rect 175576 529476 175606 529502
rect 175672 529476 175702 529502
rect 175781 529476 175811 529502
rect 175987 529476 176017 529502
rect 176073 529476 176103 529502
rect 176159 529476 176189 529502
rect 176245 529476 176275 529502
rect 176331 529476 176361 529502
rect 176417 529476 176447 529502
rect 176503 529476 176533 529502
rect 176589 529476 176619 529502
rect 176674 529476 176704 529502
rect 176760 529476 176790 529502
rect 176846 529476 176876 529502
rect 176932 529476 176962 529502
rect 177018 529476 177048 529502
rect 177104 529476 177134 529502
rect 177190 529476 177220 529502
rect 177276 529476 177306 529502
rect 177362 529476 177392 529502
rect 177448 529476 177478 529502
rect 177534 529476 177564 529502
rect 177620 529476 177650 529502
rect 177809 529476 177839 529502
rect 177893 529476 177923 529502
rect 178148 529476 178178 529502
rect 178243 529476 178273 529502
rect 178339 529476 178369 529502
rect 178505 529476 178535 529502
rect 178577 529476 178607 529502
rect 178709 529476 178739 529502
rect 178808 529476 178838 529502
rect 178917 529476 178947 529502
rect 179013 529476 179043 529502
rect 179162 529476 179192 529502
rect 179253 529476 179283 529502
rect 179461 529476 179491 529502
rect 179741 529476 179771 529502
rect 179829 529476 179859 529502
rect 180109 529476 180503 529502
rect 180754 529476 180784 529502
rect 180840 529476 180870 529502
rect 180926 529476 180956 529502
rect 181012 529476 181042 529502
rect 181098 529476 181128 529502
rect 181184 529476 181214 529502
rect 181270 529476 181300 529502
rect 181356 529476 181386 529502
rect 181442 529476 181472 529502
rect 181528 529476 181558 529502
rect 181614 529476 181644 529502
rect 181700 529476 181730 529502
rect 181785 529476 181815 529502
rect 181871 529476 181901 529502
rect 181957 529476 181987 529502
rect 182043 529476 182073 529502
rect 182129 529476 182159 529502
rect 182215 529476 182245 529502
rect 182301 529476 182331 529502
rect 182387 529476 182417 529502
rect 182593 529476 182623 529502
rect 182681 529476 182711 529502
rect 182869 529476 183815 529502
rect 183973 529476 184919 529502
rect 185261 529476 186207 529502
rect 186365 529476 186943 529502
rect 187285 529476 187403 529502
rect 172289 529340 172407 529366
rect 172565 529340 173511 529366
rect 173669 529340 174615 529366
rect 172369 529338 172407 529340
rect 172369 529322 172435 529338
rect 172261 529282 172327 529298
rect 172261 529248 172277 529282
rect 172311 529248 172327 529282
rect 172369 529288 172385 529322
rect 172419 529288 172435 529322
rect 173057 529318 173511 529340
rect 172369 529272 172435 529288
rect 172565 529282 173015 529298
rect 172261 529232 172327 529248
rect 172289 529230 172327 529232
rect 172565 529248 172837 529282
rect 172871 529248 173015 529282
rect 173057 529284 173201 529318
rect 173235 529284 173511 529318
rect 174161 529318 174615 529340
rect 173057 529268 173511 529284
rect 173669 529282 174119 529298
rect 172289 529200 172407 529230
rect 172565 529226 173015 529248
rect 173669 529248 173941 529282
rect 173975 529248 174119 529282
rect 174161 529284 174305 529318
rect 174339 529284 174615 529318
rect 174161 529268 174615 529284
rect 173669 529226 174119 529248
rect 175187 529247 175217 529392
rect 175355 529354 175385 529392
rect 175451 529360 175481 529392
rect 175576 529360 175606 529392
rect 175259 529344 175385 529354
rect 175259 529310 175275 529344
rect 175309 529324 175385 529344
rect 175427 529344 175481 529360
rect 175309 529310 175325 529324
rect 175259 529300 175325 529310
rect 175427 529310 175437 529344
rect 175471 529310 175481 529344
rect 175187 529231 175241 529247
rect 172565 529200 173511 529226
rect 173669 529200 174615 529226
rect 175187 529197 175197 529231
rect 175231 529197 175241 529231
rect 175187 529181 175241 529197
rect 175187 529149 175217 529181
rect 175283 529149 175313 529300
rect 175427 529294 175481 529310
rect 175523 529344 175606 529360
rect 175523 529310 175533 529344
rect 175567 529310 175606 529344
rect 175672 529324 175702 529392
rect 175781 529324 175811 529346
rect 175987 529333 176017 529392
rect 176073 529333 176103 529392
rect 176159 529333 176189 529392
rect 176245 529333 176275 529392
rect 176331 529333 176361 529392
rect 176417 529333 176447 529392
rect 176503 529333 176533 529392
rect 176589 529333 176619 529392
rect 176674 529333 176704 529392
rect 176760 529333 176790 529392
rect 176846 529333 176876 529392
rect 176932 529333 176962 529392
rect 177018 529333 177048 529392
rect 177104 529333 177134 529392
rect 177190 529333 177220 529392
rect 177276 529333 177306 529392
rect 175523 529294 175606 529310
rect 175664 529308 175718 529324
rect 175355 529231 175409 529247
rect 175355 529197 175365 529231
rect 175399 529197 175409 529231
rect 175355 529181 175409 529197
rect 175451 529194 175481 529294
rect 175664 529274 175674 529308
rect 175708 529274 175718 529308
rect 175664 529258 175718 529274
rect 175760 529308 175814 529324
rect 175760 529274 175770 529308
rect 175804 529274 175814 529308
rect 175760 529258 175814 529274
rect 175987 529308 177306 529333
rect 175987 529274 176212 529308
rect 176246 529274 176280 529308
rect 176314 529274 176348 529308
rect 176382 529274 176416 529308
rect 176450 529274 176484 529308
rect 176518 529274 176552 529308
rect 176586 529274 176620 529308
rect 176654 529274 176688 529308
rect 176722 529274 176756 529308
rect 176790 529274 176824 529308
rect 176858 529274 176892 529308
rect 176926 529274 176960 529308
rect 176994 529274 177028 529308
rect 177062 529274 177096 529308
rect 177130 529274 177164 529308
rect 177198 529274 177232 529308
rect 177266 529274 177306 529308
rect 175987 529258 177306 529274
rect 175355 529149 175385 529181
rect 175451 529164 175599 529194
rect 175569 529149 175599 529164
rect 175672 529149 175702 529258
rect 175781 529226 175811 529258
rect 175987 529226 176017 529258
rect 176073 529226 176103 529258
rect 176159 529226 176189 529258
rect 176245 529226 176275 529258
rect 176331 529226 176361 529258
rect 176417 529226 176447 529258
rect 176503 529226 176533 529258
rect 176589 529226 176619 529258
rect 176674 529226 176704 529258
rect 176760 529226 176790 529258
rect 176846 529226 176876 529258
rect 176932 529226 176962 529258
rect 177018 529226 177048 529258
rect 177104 529226 177134 529258
rect 177190 529226 177220 529258
rect 177276 529226 177306 529258
rect 177362 529343 177392 529392
rect 177448 529343 177478 529392
rect 177534 529343 177564 529392
rect 177620 529343 177650 529392
rect 177809 529377 177839 529392
rect 177776 529347 177839 529377
rect 177362 529308 177709 529343
rect 177776 529324 177806 529347
rect 177362 529274 177659 529308
rect 177693 529274 177709 529308
rect 177362 529241 177709 529274
rect 177752 529308 177806 529324
rect 177752 529274 177762 529308
rect 177796 529274 177806 529308
rect 177893 529303 177923 529392
rect 177752 529258 177806 529274
rect 177362 529226 177392 529241
rect 177448 529226 177478 529241
rect 177534 529226 177564 529241
rect 177620 529226 177650 529241
rect 175187 529039 175217 529065
rect 175283 529039 175313 529065
rect 175355 529039 175385 529065
rect 175569 529039 175599 529065
rect 175672 529039 175702 529065
rect 177776 529205 177806 529258
rect 177848 529293 177923 529303
rect 177848 529259 177864 529293
rect 177898 529259 177923 529293
rect 178148 529263 178178 529392
rect 178243 529370 178273 529404
rect 178339 529370 178369 529404
rect 178220 529354 178274 529370
rect 178220 529320 178230 529354
rect 178264 529320 178274 529354
rect 178220 529304 178274 529320
rect 178316 529360 178382 529370
rect 178316 529326 178332 529360
rect 178366 529326 178382 529360
rect 178316 529316 178382 529326
rect 177848 529249 177923 529259
rect 177776 529175 177839 529205
rect 177809 529160 177839 529175
rect 177893 529160 177923 529249
rect 178061 529247 178178 529263
rect 178061 529213 178071 529247
rect 178105 529227 178178 529247
rect 178243 529274 178274 529304
rect 178243 529244 178381 529274
rect 178105 529213 178190 529227
rect 178061 529197 178190 529213
rect 178160 529110 178190 529197
rect 178236 529192 178302 529202
rect 178236 529158 178252 529192
rect 178286 529158 178302 529192
rect 178236 529148 178302 529158
rect 178252 529110 178282 529148
rect 178351 529110 178381 529244
rect 178505 529234 178535 529392
rect 178577 529370 178607 529392
rect 178577 529354 178631 529370
rect 178577 529320 178587 529354
rect 178621 529320 178631 529354
rect 178808 529382 178838 529404
rect 178808 529366 178875 529382
rect 178709 529322 178739 529348
rect 178577 529304 178631 529320
rect 178673 529306 178739 529322
rect 178808 529332 178831 529366
rect 178865 529332 178875 529366
rect 178808 529316 178875 529332
rect 178917 529334 178947 529404
rect 179013 529360 179043 529392
rect 179013 529344 179115 529360
rect 178917 529318 178971 529334
rect 179013 529330 179071 529344
rect 178491 529218 178546 529234
rect 178491 529184 178501 529218
rect 178535 529184 178546 529218
rect 178491 529168 178546 529184
rect 178491 529110 178521 529168
rect 178588 529110 178618 529304
rect 178673 529272 178683 529306
rect 178717 529272 178739 529306
rect 178917 529286 178927 529318
rect 178905 529284 178927 529286
rect 178961 529284 178971 529318
rect 178905 529274 178971 529284
rect 178673 529256 178739 529272
rect 178709 529239 178739 529256
rect 178884 529268 178971 529274
rect 179054 529310 179071 529330
rect 179105 529310 179115 529344
rect 179162 529332 179192 529392
rect 179054 529294 179115 529310
rect 179157 529316 179211 529332
rect 178884 529256 178947 529268
rect 178884 529244 178934 529256
rect 178709 529209 178815 529239
rect 178785 529194 178815 529209
rect 172289 529000 172407 529026
rect 172565 529000 173511 529026
rect 173669 529000 174615 529026
rect 175781 529000 175811 529026
rect 175987 529000 176017 529026
rect 176073 529000 176103 529026
rect 176159 529000 176189 529026
rect 176245 529000 176275 529026
rect 176331 529000 176361 529026
rect 176417 529000 176447 529026
rect 176503 529000 176533 529026
rect 176589 529000 176619 529026
rect 176674 529000 176704 529026
rect 176760 529000 176790 529026
rect 176846 529000 176876 529026
rect 176932 529000 176962 529026
rect 177018 529000 177048 529026
rect 177104 529000 177134 529026
rect 177190 529000 177220 529026
rect 177276 529000 177306 529026
rect 177362 529000 177392 529026
rect 177448 529000 177478 529026
rect 177534 529000 177564 529026
rect 177620 529000 177650 529026
rect 177809 529006 177839 529032
rect 177893 529006 177923 529032
rect 178884 529110 178914 529244
rect 178956 529192 179010 529208
rect 178956 529158 178966 529192
rect 179000 529158 179010 529192
rect 178956 529142 179010 529158
rect 178970 529110 179000 529142
rect 179054 529110 179084 529294
rect 179157 529282 179167 529316
rect 179201 529282 179211 529316
rect 179157 529266 179211 529282
rect 179162 529110 179192 529266
rect 179253 529224 179283 529392
rect 179741 529357 179771 529372
rect 179461 529324 179491 529346
rect 179735 529333 179771 529357
rect 179735 529324 179765 529333
rect 179432 529308 179491 529324
rect 179432 529274 179442 529308
rect 179476 529274 179491 529308
rect 179432 529258 179491 529274
rect 179689 529308 179765 529324
rect 179829 529311 179859 529372
rect 180109 529340 180503 529366
rect 180754 529343 180784 529392
rect 180840 529343 180870 529392
rect 180926 529343 180956 529392
rect 181012 529343 181042 529392
rect 180327 529318 180503 529340
rect 179689 529274 179699 529308
rect 179733 529274 179765 529308
rect 179689 529258 179765 529274
rect 179461 529226 179491 529258
rect 179234 529208 179288 529224
rect 179234 529174 179244 529208
rect 179278 529174 179288 529208
rect 179234 529158 179288 529174
rect 179246 529110 179276 529158
rect 179735 529223 179765 529258
rect 179809 529295 179863 529311
rect 179809 529261 179819 529295
rect 179853 529261 179863 529295
rect 179809 529245 179863 529261
rect 180109 529282 180285 529298
rect 180109 529248 180125 529282
rect 180159 529248 180235 529282
rect 180269 529248 180285 529282
rect 180327 529284 180343 529318
rect 180377 529284 180453 529318
rect 180487 529284 180503 529318
rect 180327 529268 180503 529284
rect 180695 529308 181042 529343
rect 180695 529274 180711 529308
rect 180745 529274 181042 529308
rect 179735 529199 179771 529223
rect 179741 529184 179771 529199
rect 179829 529184 179859 529245
rect 180109 529226 180285 529248
rect 180695 529241 181042 529274
rect 180754 529226 180784 529241
rect 180840 529226 180870 529241
rect 180926 529226 180956 529241
rect 181012 529226 181042 529241
rect 181098 529333 181128 529392
rect 181184 529333 181214 529392
rect 181270 529333 181300 529392
rect 181356 529333 181386 529392
rect 181442 529333 181472 529392
rect 181528 529333 181558 529392
rect 181614 529333 181644 529392
rect 181700 529333 181730 529392
rect 181785 529333 181815 529392
rect 181871 529333 181901 529392
rect 181957 529333 181987 529392
rect 182043 529333 182073 529392
rect 182129 529333 182159 529392
rect 182215 529333 182245 529392
rect 182301 529333 182331 529392
rect 182387 529333 182417 529392
rect 181098 529308 182417 529333
rect 182593 529311 182623 529372
rect 182681 529357 182711 529372
rect 182681 529333 182717 529357
rect 182869 529340 183815 529366
rect 183973 529340 184919 529366
rect 185261 529340 186207 529366
rect 186365 529340 186943 529366
rect 182687 529324 182717 529333
rect 181098 529274 181138 529308
rect 181172 529274 181206 529308
rect 181240 529274 181274 529308
rect 181308 529274 181342 529308
rect 181376 529274 181410 529308
rect 181444 529274 181478 529308
rect 181512 529274 181546 529308
rect 181580 529274 181614 529308
rect 181648 529274 181682 529308
rect 181716 529274 181750 529308
rect 181784 529274 181818 529308
rect 181852 529274 181886 529308
rect 181920 529274 181954 529308
rect 181988 529274 182022 529308
rect 182056 529274 182090 529308
rect 182124 529274 182158 529308
rect 182192 529274 182417 529308
rect 181098 529258 182417 529274
rect 181098 529226 181128 529258
rect 181184 529226 181214 529258
rect 181270 529226 181300 529258
rect 181356 529226 181386 529258
rect 181442 529226 181472 529258
rect 181528 529226 181558 529258
rect 181614 529226 181644 529258
rect 181700 529226 181730 529258
rect 181785 529226 181815 529258
rect 181871 529226 181901 529258
rect 181957 529226 181987 529258
rect 182043 529226 182073 529258
rect 182129 529226 182159 529258
rect 182215 529226 182245 529258
rect 182301 529226 182331 529258
rect 182387 529226 182417 529258
rect 182589 529295 182643 529311
rect 182589 529261 182599 529295
rect 182633 529261 182643 529295
rect 182589 529245 182643 529261
rect 182687 529308 182763 529324
rect 182687 529274 182719 529308
rect 182753 529274 182763 529308
rect 183361 529318 183815 529340
rect 182687 529258 182763 529274
rect 182869 529282 183319 529298
rect 180109 529200 180503 529226
rect 182593 529184 182623 529245
rect 182687 529223 182717 529258
rect 182681 529199 182717 529223
rect 182869 529248 183141 529282
rect 183175 529248 183319 529282
rect 183361 529284 183505 529318
rect 183539 529284 183815 529318
rect 184465 529318 184919 529340
rect 183361 529268 183815 529284
rect 183973 529282 184423 529298
rect 182869 529226 183319 529248
rect 183973 529248 184245 529282
rect 184279 529248 184423 529282
rect 184465 529284 184609 529318
rect 184643 529284 184919 529318
rect 185753 529318 186207 529340
rect 184465 529268 184919 529284
rect 185261 529282 185711 529298
rect 183973 529226 184423 529248
rect 185261 529248 185533 529282
rect 185567 529248 185711 529282
rect 185753 529284 185897 529318
rect 185931 529284 186207 529318
rect 186671 529318 186943 529340
rect 187285 529340 187403 529366
rect 187285 529338 187323 529340
rect 185753 529268 186207 529284
rect 186365 529282 186629 529298
rect 185261 529226 185711 529248
rect 186365 529248 186381 529282
rect 186415 529248 186480 529282
rect 186514 529248 186579 529282
rect 186613 529248 186629 529282
rect 186671 529284 186687 529318
rect 186721 529284 186790 529318
rect 186824 529284 186893 529318
rect 186927 529284 186943 529318
rect 186671 529268 186943 529284
rect 187257 529322 187323 529338
rect 187257 529288 187273 529322
rect 187307 529288 187323 529322
rect 187257 529272 187323 529288
rect 187365 529282 187431 529298
rect 186365 529226 186629 529248
rect 187365 529248 187381 529282
rect 187415 529248 187431 529282
rect 187365 529232 187431 529248
rect 187365 529230 187403 529232
rect 182869 529200 183815 529226
rect 183973 529200 184919 529226
rect 182681 529184 182711 529199
rect 185261 529200 186207 529226
rect 186365 529200 186943 529226
rect 187285 529200 187403 529230
rect 178160 529000 178190 529026
rect 178252 529000 178282 529026
rect 178351 529000 178381 529026
rect 178491 529000 178521 529026
rect 178588 529000 178618 529026
rect 178785 529000 178815 529026
rect 178884 529000 178914 529026
rect 178970 529000 179000 529026
rect 179054 529000 179084 529026
rect 179162 529000 179192 529026
rect 179246 529000 179276 529026
rect 179461 529000 179491 529026
rect 179741 529000 179771 529026
rect 179829 529000 179859 529026
rect 180109 529000 180503 529026
rect 180754 529000 180784 529026
rect 180840 529000 180870 529026
rect 180926 529000 180956 529026
rect 181012 529000 181042 529026
rect 181098 529000 181128 529026
rect 181184 529000 181214 529026
rect 181270 529000 181300 529026
rect 181356 529000 181386 529026
rect 181442 529000 181472 529026
rect 181528 529000 181558 529026
rect 181614 529000 181644 529026
rect 181700 529000 181730 529026
rect 181785 529000 181815 529026
rect 181871 529000 181901 529026
rect 181957 529000 181987 529026
rect 182043 529000 182073 529026
rect 182129 529000 182159 529026
rect 182215 529000 182245 529026
rect 182301 529000 182331 529026
rect 182387 529000 182417 529026
rect 182593 529000 182623 529026
rect 182681 529000 182711 529026
rect 182869 529000 183815 529026
rect 183973 529000 184919 529026
rect 185261 529000 186207 529026
rect 186365 529000 186943 529026
rect 187285 529000 187403 529026
rect 172289 528932 172407 528958
rect 172565 528932 173511 528958
rect 173669 528932 174615 528958
rect 174773 528932 175719 528958
rect 175969 528932 175999 528958
rect 176057 528932 176087 528958
rect 176245 528932 176275 528958
rect 176333 528932 176363 528958
rect 177161 528932 177191 528958
rect 177552 528932 177582 528958
rect 177647 528932 177747 528958
rect 177905 528932 178005 528958
rect 178059 528932 178089 528958
rect 178454 528932 178484 528958
rect 178540 528932 178570 528958
rect 178626 528932 178656 528958
rect 178712 528932 178742 528958
rect 178798 528932 178828 528958
rect 178884 528932 178914 528958
rect 178970 528932 179000 528958
rect 179056 528932 179086 528958
rect 179142 528932 179172 528958
rect 179228 528932 179258 528958
rect 179314 528932 179344 528958
rect 179400 528932 179430 528958
rect 179485 528932 179515 528958
rect 179571 528932 179601 528958
rect 179657 528932 179687 528958
rect 179743 528932 179773 528958
rect 179829 528932 179859 528958
rect 179915 528932 179945 528958
rect 180001 528932 180031 528958
rect 180087 528932 180117 528958
rect 180293 528932 180323 528958
rect 180381 528932 180411 528958
rect 176567 528893 176597 528919
rect 176663 528893 176693 528919
rect 176735 528893 176765 528919
rect 176949 528893 176979 528919
rect 177052 528893 177082 528919
rect 176567 528777 176597 528809
rect 175969 528759 175999 528774
rect 172289 528728 172407 528758
rect 172565 528732 173511 528758
rect 173669 528732 174615 528758
rect 174773 528732 175719 528758
rect 175963 528735 175999 528759
rect 172289 528726 172327 528728
rect 172261 528710 172327 528726
rect 172261 528676 172277 528710
rect 172311 528676 172327 528710
rect 172565 528710 173015 528732
rect 172261 528660 172327 528676
rect 172369 528670 172435 528686
rect 172369 528636 172385 528670
rect 172419 528636 172435 528670
rect 172565 528676 172837 528710
rect 172871 528676 173015 528710
rect 173669 528710 174119 528732
rect 172565 528660 173015 528676
rect 173057 528674 173511 528690
rect 172369 528620 172435 528636
rect 173057 528640 173201 528674
rect 173235 528640 173511 528674
rect 173669 528676 173941 528710
rect 173975 528676 174119 528710
rect 174773 528710 175223 528732
rect 173669 528660 174119 528676
rect 174161 528674 174615 528690
rect 172369 528618 172407 528620
rect 173057 528618 173511 528640
rect 174161 528640 174305 528674
rect 174339 528640 174615 528674
rect 174773 528676 175045 528710
rect 175079 528676 175223 528710
rect 175963 528700 175993 528735
rect 176057 528713 176087 528774
rect 176245 528759 176275 528774
rect 176239 528735 176275 528759
rect 174773 528660 175223 528676
rect 175265 528674 175719 528690
rect 174161 528618 174615 528640
rect 175265 528640 175409 528674
rect 175443 528640 175719 528674
rect 175265 528618 175719 528640
rect 175917 528684 175993 528700
rect 175917 528650 175927 528684
rect 175961 528650 175993 528684
rect 175917 528634 175993 528650
rect 176037 528697 176091 528713
rect 176239 528700 176269 528735
rect 176333 528713 176363 528774
rect 176567 528761 176621 528777
rect 176567 528727 176577 528761
rect 176611 528727 176621 528761
rect 176037 528663 176047 528697
rect 176081 528663 176091 528697
rect 176037 528647 176091 528663
rect 176193 528684 176269 528700
rect 176193 528650 176203 528684
rect 176237 528650 176269 528684
rect 172289 528592 172407 528618
rect 172565 528592 173511 528618
rect 173669 528592 174615 528618
rect 174773 528592 175719 528618
rect 175963 528625 175993 528634
rect 175963 528601 175999 528625
rect 175969 528586 175999 528601
rect 176057 528586 176087 528647
rect 176193 528634 176269 528650
rect 176313 528697 176367 528713
rect 176313 528663 176323 528697
rect 176357 528663 176367 528697
rect 176313 528647 176367 528663
rect 176567 528711 176621 528727
rect 176239 528625 176269 528634
rect 176239 528601 176275 528625
rect 176245 528586 176275 528601
rect 176333 528586 176363 528647
rect 176567 528566 176597 528711
rect 176663 528658 176693 528809
rect 176735 528777 176765 528809
rect 176949 528794 176979 528809
rect 176735 528761 176789 528777
rect 176735 528727 176745 528761
rect 176779 528727 176789 528761
rect 176735 528711 176789 528727
rect 176831 528764 176979 528794
rect 176831 528664 176861 528764
rect 177052 528700 177082 528809
rect 177161 528700 177191 528732
rect 177552 528700 177582 528732
rect 177647 528700 177747 528848
rect 177044 528684 177098 528700
rect 176639 528648 176705 528658
rect 176639 528614 176655 528648
rect 176689 528634 176705 528648
rect 176807 528648 176861 528664
rect 176689 528614 176765 528634
rect 176639 528604 176765 528614
rect 176735 528566 176765 528604
rect 176807 528614 176817 528648
rect 176851 528614 176861 528648
rect 176807 528598 176861 528614
rect 176903 528648 176986 528664
rect 176903 528614 176913 528648
rect 176947 528614 176986 528648
rect 177044 528650 177054 528684
rect 177088 528650 177098 528684
rect 177044 528634 177098 528650
rect 177140 528684 177194 528700
rect 177140 528650 177150 528684
rect 177184 528650 177194 528684
rect 177140 528634 177194 528650
rect 177551 528684 177605 528700
rect 177551 528650 177561 528684
rect 177595 528650 177605 528684
rect 177551 528634 177605 528650
rect 177647 528684 177801 528700
rect 177647 528650 177757 528684
rect 177791 528650 177801 528684
rect 177647 528634 177801 528650
rect 177905 528684 178005 528848
rect 177905 528650 177961 528684
rect 177995 528650 178005 528684
rect 176903 528598 176986 528614
rect 176831 528566 176861 528598
rect 176956 528566 176986 528598
rect 177052 528566 177082 528634
rect 177161 528612 177191 528634
rect 177552 528612 177582 528634
rect 177647 528566 177747 528634
rect 177905 528566 178005 528650
rect 178059 528700 178089 528848
rect 180569 528926 180599 528952
rect 180653 528926 180683 528952
rect 180920 528932 180950 528958
rect 181012 528932 181042 528958
rect 181111 528932 181141 528958
rect 181251 528932 181281 528958
rect 181348 528932 181378 528958
rect 181545 528932 181575 528958
rect 181644 528932 181674 528958
rect 181730 528932 181760 528958
rect 181814 528932 181844 528958
rect 181922 528932 181952 528958
rect 182006 528932 182036 528958
rect 182221 528932 182251 528958
rect 182685 528932 183631 528958
rect 183789 528932 184735 528958
rect 184893 528932 185839 528958
rect 185997 528932 186943 528958
rect 187285 528932 187403 528958
rect 180569 528783 180599 528798
rect 180293 528759 180323 528774
rect 180287 528735 180323 528759
rect 178454 528717 178484 528732
rect 178540 528717 178570 528732
rect 178626 528717 178656 528732
rect 178712 528717 178742 528732
rect 178059 528684 178119 528700
rect 178059 528650 178075 528684
rect 178109 528650 178119 528684
rect 178059 528634 178119 528650
rect 178395 528684 178742 528717
rect 178395 528650 178411 528684
rect 178445 528650 178742 528684
rect 178059 528566 178089 528634
rect 178395 528615 178742 528650
rect 178454 528566 178484 528615
rect 178540 528566 178570 528615
rect 178626 528566 178656 528615
rect 178712 528566 178742 528615
rect 178798 528700 178828 528732
rect 178884 528700 178914 528732
rect 178970 528700 179000 528732
rect 179056 528700 179086 528732
rect 179142 528700 179172 528732
rect 179228 528700 179258 528732
rect 179314 528700 179344 528732
rect 179400 528700 179430 528732
rect 179485 528700 179515 528732
rect 179571 528700 179601 528732
rect 179657 528700 179687 528732
rect 179743 528700 179773 528732
rect 179829 528700 179859 528732
rect 179915 528700 179945 528732
rect 180001 528700 180031 528732
rect 180087 528700 180117 528732
rect 180287 528700 180317 528735
rect 180381 528713 180411 528774
rect 180536 528753 180599 528783
rect 178798 528684 180117 528700
rect 178798 528650 178838 528684
rect 178872 528650 178906 528684
rect 178940 528650 178974 528684
rect 179008 528650 179042 528684
rect 179076 528650 179110 528684
rect 179144 528650 179178 528684
rect 179212 528650 179246 528684
rect 179280 528650 179314 528684
rect 179348 528650 179382 528684
rect 179416 528650 179450 528684
rect 179484 528650 179518 528684
rect 179552 528650 179586 528684
rect 179620 528650 179654 528684
rect 179688 528650 179722 528684
rect 179756 528650 179790 528684
rect 179824 528650 179858 528684
rect 179892 528650 180117 528684
rect 178798 528625 180117 528650
rect 180241 528684 180317 528700
rect 180241 528650 180251 528684
rect 180285 528650 180317 528684
rect 180241 528634 180317 528650
rect 180361 528697 180415 528713
rect 180536 528700 180566 528753
rect 180653 528709 180683 528798
rect 180920 528761 180950 528848
rect 181012 528810 181042 528848
rect 180361 528663 180371 528697
rect 180405 528663 180415 528697
rect 180361 528647 180415 528663
rect 180512 528684 180566 528700
rect 180512 528650 180522 528684
rect 180556 528650 180566 528684
rect 180608 528699 180683 528709
rect 180608 528665 180624 528699
rect 180658 528665 180683 528699
rect 180821 528745 180950 528761
rect 180996 528800 181062 528810
rect 180996 528766 181012 528800
rect 181046 528766 181062 528800
rect 180996 528756 181062 528766
rect 180821 528711 180831 528745
rect 180865 528731 180950 528745
rect 180865 528711 180938 528731
rect 181111 528714 181141 528848
rect 181251 528790 181281 528848
rect 181251 528774 181306 528790
rect 181251 528740 181261 528774
rect 181295 528740 181306 528774
rect 181251 528724 181306 528740
rect 180821 528695 180938 528711
rect 180608 528655 180683 528665
rect 178798 528566 178828 528625
rect 178884 528566 178914 528625
rect 178970 528566 179000 528625
rect 179056 528566 179086 528625
rect 179142 528566 179172 528625
rect 179228 528566 179258 528625
rect 179314 528566 179344 528625
rect 179400 528566 179430 528625
rect 179485 528566 179515 528625
rect 179571 528566 179601 528625
rect 179657 528566 179687 528625
rect 179743 528566 179773 528625
rect 179829 528566 179859 528625
rect 179915 528566 179945 528625
rect 180001 528566 180031 528625
rect 180087 528566 180117 528625
rect 180287 528625 180317 528634
rect 180287 528601 180323 528625
rect 180293 528586 180323 528601
rect 180381 528586 180411 528647
rect 180512 528634 180566 528650
rect 180536 528611 180566 528634
rect 180536 528581 180599 528611
rect 180569 528566 180599 528581
rect 180653 528566 180683 528655
rect 180908 528566 180938 528695
rect 181003 528684 181141 528714
rect 181003 528654 181034 528684
rect 180980 528638 181034 528654
rect 180980 528604 180990 528638
rect 181024 528604 181034 528638
rect 180980 528588 181034 528604
rect 181076 528632 181142 528642
rect 181076 528598 181092 528632
rect 181126 528598 181142 528632
rect 181076 528588 181142 528598
rect 181003 528554 181033 528588
rect 181099 528554 181129 528588
rect 181265 528566 181295 528724
rect 181348 528654 181378 528848
rect 181545 528749 181575 528764
rect 181469 528719 181575 528749
rect 181469 528702 181499 528719
rect 181433 528686 181499 528702
rect 181337 528638 181391 528654
rect 181337 528604 181347 528638
rect 181381 528604 181391 528638
rect 181433 528652 181443 528686
rect 181477 528652 181499 528686
rect 181644 528714 181674 528848
rect 181730 528816 181760 528848
rect 181716 528800 181770 528816
rect 181716 528766 181726 528800
rect 181760 528766 181770 528800
rect 181716 528750 181770 528766
rect 181644 528702 181694 528714
rect 181644 528690 181707 528702
rect 181644 528684 181731 528690
rect 181665 528674 181731 528684
rect 181665 528672 181687 528674
rect 181433 528636 181499 528652
rect 181469 528610 181499 528636
rect 181568 528626 181635 528642
rect 181337 528588 181391 528604
rect 181337 528566 181367 528588
rect 181568 528592 181591 528626
rect 181625 528592 181635 528626
rect 181568 528576 181635 528592
rect 181677 528640 181687 528672
rect 181721 528640 181731 528674
rect 181677 528624 181731 528640
rect 181814 528664 181844 528848
rect 181922 528692 181952 528848
rect 182006 528800 182036 528848
rect 181994 528784 182048 528800
rect 181994 528750 182004 528784
rect 182038 528750 182048 528784
rect 181994 528734 182048 528750
rect 181917 528676 181971 528692
rect 181814 528648 181875 528664
rect 181814 528628 181831 528648
rect 181568 528554 181598 528576
rect 181677 528554 181707 528624
rect 181773 528614 181831 528628
rect 181865 528614 181875 528648
rect 181917 528642 181927 528676
rect 181961 528642 181971 528676
rect 181917 528626 181971 528642
rect 181773 528598 181875 528614
rect 181773 528566 181803 528598
rect 181922 528566 181952 528626
rect 182013 528566 182043 528734
rect 182685 528732 183631 528758
rect 183789 528732 184735 528758
rect 184893 528732 185839 528758
rect 185997 528732 186943 528758
rect 182221 528700 182251 528732
rect 182192 528684 182251 528700
rect 182192 528650 182202 528684
rect 182236 528650 182251 528684
rect 182685 528710 183135 528732
rect 182685 528676 182957 528710
rect 182991 528676 183135 528710
rect 183789 528710 184239 528732
rect 182685 528660 183135 528676
rect 183177 528674 183631 528690
rect 182192 528634 182251 528650
rect 182221 528612 182251 528634
rect 183177 528640 183321 528674
rect 183355 528640 183631 528674
rect 183789 528676 184061 528710
rect 184095 528676 184239 528710
rect 184893 528710 185343 528732
rect 183789 528660 184239 528676
rect 184281 528674 184735 528690
rect 183177 528618 183631 528640
rect 184281 528640 184425 528674
rect 184459 528640 184735 528674
rect 184893 528676 185165 528710
rect 185199 528676 185343 528710
rect 185997 528710 186447 528732
rect 187285 528728 187403 528758
rect 184893 528660 185343 528676
rect 185385 528674 185839 528690
rect 184281 528618 184735 528640
rect 185385 528640 185529 528674
rect 185563 528640 185839 528674
rect 185997 528676 186269 528710
rect 186303 528676 186447 528710
rect 187365 528726 187403 528728
rect 187365 528710 187431 528726
rect 185997 528660 186447 528676
rect 186489 528674 186943 528690
rect 185385 528618 185839 528640
rect 186489 528640 186633 528674
rect 186667 528640 186943 528674
rect 186489 528618 186943 528640
rect 187257 528670 187323 528686
rect 187257 528636 187273 528670
rect 187307 528636 187323 528670
rect 187365 528676 187381 528710
rect 187415 528676 187431 528710
rect 187365 528660 187431 528676
rect 187257 528620 187323 528636
rect 182685 528592 183631 528618
rect 183789 528592 184735 528618
rect 184893 528592 185839 528618
rect 185997 528592 186943 528618
rect 187285 528618 187323 528620
rect 187285 528592 187403 528618
rect 172289 528456 172407 528482
rect 172565 528456 173511 528482
rect 173669 528456 174615 528482
rect 174773 528456 175719 528482
rect 175969 528456 175999 528482
rect 176057 528456 176087 528482
rect 176245 528456 176275 528482
rect 176333 528456 176363 528482
rect 176567 528456 176597 528482
rect 176735 528456 176765 528482
rect 176831 528456 176861 528482
rect 176956 528456 176986 528482
rect 177052 528456 177082 528482
rect 177161 528456 177191 528482
rect 177552 528456 177582 528482
rect 177647 528456 177747 528482
rect 177905 528456 178005 528482
rect 178059 528456 178089 528482
rect 178454 528456 178484 528482
rect 178540 528456 178570 528482
rect 178626 528456 178656 528482
rect 178712 528456 178742 528482
rect 178798 528456 178828 528482
rect 178884 528456 178914 528482
rect 178970 528456 179000 528482
rect 179056 528456 179086 528482
rect 179142 528456 179172 528482
rect 179228 528456 179258 528482
rect 179314 528456 179344 528482
rect 179400 528456 179430 528482
rect 179485 528456 179515 528482
rect 179571 528456 179601 528482
rect 179657 528456 179687 528482
rect 179743 528456 179773 528482
rect 179829 528456 179859 528482
rect 179915 528456 179945 528482
rect 180001 528456 180031 528482
rect 180087 528456 180117 528482
rect 180293 528456 180323 528482
rect 180381 528456 180411 528482
rect 180569 528456 180599 528482
rect 180653 528456 180683 528482
rect 180908 528456 180938 528482
rect 181003 528456 181033 528482
rect 181099 528456 181129 528482
rect 181265 528456 181295 528482
rect 181337 528456 181367 528482
rect 181469 528456 181499 528482
rect 181568 528456 181598 528482
rect 181677 528456 181707 528482
rect 181773 528456 181803 528482
rect 181922 528456 181952 528482
rect 182013 528456 182043 528482
rect 182221 528456 182251 528482
rect 182685 528456 183631 528482
rect 183789 528456 184735 528482
rect 184893 528456 185839 528482
rect 185997 528456 186943 528482
rect 187285 528456 187403 528482
rect 172289 528388 172407 528414
rect 172565 528388 173511 528414
rect 173669 528388 174615 528414
rect 174957 528388 175903 528414
rect 176153 528388 176183 528414
rect 176237 528388 176267 528414
rect 176492 528388 176522 528414
rect 176587 528388 176617 528414
rect 176683 528388 176713 528414
rect 176849 528388 176879 528414
rect 176921 528388 176951 528414
rect 177053 528388 177083 528414
rect 177152 528388 177182 528414
rect 177261 528388 177291 528414
rect 177357 528388 177387 528414
rect 177506 528388 177536 528414
rect 177597 528388 177627 528414
rect 177805 528388 177835 528414
rect 177993 528388 178023 528414
rect 178081 528388 178111 528414
rect 178269 528388 178847 528414
rect 179005 528388 179035 528414
rect 179114 528388 179144 528414
rect 179210 528388 179240 528414
rect 179335 528388 179365 528414
rect 179431 528388 179461 528414
rect 179599 528388 179629 528414
rect 180109 528388 180687 528414
rect 181029 528388 181059 528414
rect 181138 528388 181168 528414
rect 181234 528388 181264 528414
rect 181359 528388 181389 528414
rect 181455 528388 181485 528414
rect 181623 528388 181653 528414
rect 181857 528388 182803 528414
rect 182961 528388 183907 528414
rect 184065 528388 185011 528414
rect 185261 528388 186207 528414
rect 186365 528388 186943 528414
rect 187285 528388 187403 528414
rect 172289 528252 172407 528278
rect 172565 528252 173511 528278
rect 173669 528252 174615 528278
rect 176153 528289 176183 528304
rect 174957 528252 175903 528278
rect 172369 528250 172407 528252
rect 172369 528234 172435 528250
rect 172261 528194 172327 528210
rect 172261 528160 172277 528194
rect 172311 528160 172327 528194
rect 172369 528200 172385 528234
rect 172419 528200 172435 528234
rect 173057 528230 173511 528252
rect 172369 528184 172435 528200
rect 172565 528194 173015 528210
rect 172261 528144 172327 528160
rect 172289 528142 172327 528144
rect 172565 528160 172837 528194
rect 172871 528160 173015 528194
rect 173057 528196 173201 528230
rect 173235 528196 173511 528230
rect 174161 528230 174615 528252
rect 173057 528180 173511 528196
rect 173669 528194 174119 528210
rect 172289 528112 172407 528142
rect 172565 528138 173015 528160
rect 173669 528160 173941 528194
rect 173975 528160 174119 528194
rect 174161 528196 174305 528230
rect 174339 528196 174615 528230
rect 175449 528230 175903 528252
rect 176120 528259 176183 528289
rect 176120 528236 176150 528259
rect 174161 528180 174615 528196
rect 174957 528194 175407 528210
rect 173669 528138 174119 528160
rect 174957 528160 175229 528194
rect 175263 528160 175407 528194
rect 175449 528196 175593 528230
rect 175627 528196 175903 528230
rect 175449 528180 175903 528196
rect 176096 528220 176150 528236
rect 176096 528186 176106 528220
rect 176140 528186 176150 528220
rect 176237 528215 176267 528304
rect 176096 528170 176150 528186
rect 174957 528138 175407 528160
rect 172565 528112 173511 528138
rect 173669 528112 174615 528138
rect 174957 528112 175903 528138
rect 176120 528117 176150 528170
rect 176192 528205 176267 528215
rect 176192 528171 176208 528205
rect 176242 528171 176267 528205
rect 176492 528175 176522 528304
rect 176587 528282 176617 528316
rect 176683 528282 176713 528316
rect 176564 528266 176618 528282
rect 176564 528232 176574 528266
rect 176608 528232 176618 528266
rect 176564 528216 176618 528232
rect 176660 528272 176726 528282
rect 176660 528238 176676 528272
rect 176710 528238 176726 528272
rect 176660 528228 176726 528238
rect 176192 528161 176267 528171
rect 176120 528087 176183 528117
rect 176153 528072 176183 528087
rect 176237 528072 176267 528161
rect 176405 528159 176522 528175
rect 176405 528125 176415 528159
rect 176449 528139 176522 528159
rect 176587 528186 176618 528216
rect 176587 528156 176725 528186
rect 176449 528125 176534 528139
rect 176405 528109 176534 528125
rect 176504 528022 176534 528109
rect 176580 528104 176646 528114
rect 176580 528070 176596 528104
rect 176630 528070 176646 528104
rect 176580 528060 176646 528070
rect 176596 528022 176626 528060
rect 176695 528022 176725 528156
rect 176849 528146 176879 528304
rect 176921 528282 176951 528304
rect 176921 528266 176975 528282
rect 176921 528232 176931 528266
rect 176965 528232 176975 528266
rect 177152 528294 177182 528316
rect 177152 528278 177219 528294
rect 177053 528234 177083 528260
rect 176921 528216 176975 528232
rect 177017 528218 177083 528234
rect 177152 528244 177175 528278
rect 177209 528244 177219 528278
rect 177152 528228 177219 528244
rect 177261 528246 177291 528316
rect 177357 528272 177387 528304
rect 177357 528256 177459 528272
rect 177261 528230 177315 528246
rect 177357 528242 177415 528256
rect 176835 528130 176890 528146
rect 176835 528096 176845 528130
rect 176879 528096 176890 528130
rect 176835 528080 176890 528096
rect 176835 528022 176865 528080
rect 176932 528022 176962 528216
rect 177017 528184 177027 528218
rect 177061 528184 177083 528218
rect 177261 528198 177271 528230
rect 177249 528196 177271 528198
rect 177305 528196 177315 528230
rect 177249 528186 177315 528196
rect 177017 528168 177083 528184
rect 177053 528151 177083 528168
rect 177228 528180 177315 528186
rect 177398 528222 177415 528242
rect 177449 528222 177459 528256
rect 177506 528244 177536 528304
rect 177398 528206 177459 528222
rect 177501 528228 177555 528244
rect 177228 528168 177291 528180
rect 177228 528156 177278 528168
rect 177053 528121 177159 528151
rect 177129 528106 177159 528121
rect 172289 527912 172407 527938
rect 172565 527912 173511 527938
rect 173669 527912 174615 527938
rect 174957 527912 175903 527938
rect 176153 527918 176183 527944
rect 176237 527918 176267 527944
rect 177228 528022 177258 528156
rect 177300 528104 177354 528120
rect 177300 528070 177310 528104
rect 177344 528070 177354 528104
rect 177300 528054 177354 528070
rect 177314 528022 177344 528054
rect 177398 528022 177428 528206
rect 177501 528194 177511 528228
rect 177545 528194 177555 528228
rect 177501 528178 177555 528194
rect 177506 528022 177536 528178
rect 177597 528136 177627 528304
rect 177805 528236 177835 528258
rect 177776 528220 177835 528236
rect 177993 528223 178023 528284
rect 178081 528269 178111 528284
rect 178081 528245 178117 528269
rect 178269 528252 178847 528278
rect 178087 528236 178117 528245
rect 177776 528186 177786 528220
rect 177820 528186 177835 528220
rect 177776 528170 177835 528186
rect 177805 528138 177835 528170
rect 177989 528207 178043 528223
rect 177989 528173 177999 528207
rect 178033 528173 178043 528207
rect 177989 528157 178043 528173
rect 178087 528220 178163 528236
rect 178087 528186 178119 528220
rect 178153 528186 178163 528220
rect 178575 528230 178847 528252
rect 179005 528236 179035 528258
rect 179114 528236 179144 528304
rect 179210 528272 179240 528304
rect 179335 528272 179365 528304
rect 179210 528256 179293 528272
rect 178087 528170 178163 528186
rect 178269 528194 178533 528210
rect 177578 528120 177632 528136
rect 177578 528086 177588 528120
rect 177622 528086 177632 528120
rect 177578 528070 177632 528086
rect 177590 528022 177620 528070
rect 177993 528096 178023 528157
rect 178087 528135 178117 528170
rect 178081 528111 178117 528135
rect 178269 528160 178285 528194
rect 178319 528160 178384 528194
rect 178418 528160 178483 528194
rect 178517 528160 178533 528194
rect 178575 528196 178591 528230
rect 178625 528196 178694 528230
rect 178728 528196 178797 528230
rect 178831 528196 178847 528230
rect 178575 528180 178847 528196
rect 179002 528220 179056 528236
rect 179002 528186 179012 528220
rect 179046 528186 179056 528220
rect 179002 528170 179056 528186
rect 179098 528220 179152 528236
rect 179098 528186 179108 528220
rect 179142 528186 179152 528220
rect 179210 528222 179249 528256
rect 179283 528222 179293 528256
rect 179210 528206 179293 528222
rect 179335 528256 179389 528272
rect 179335 528222 179345 528256
rect 179379 528222 179389 528256
rect 179431 528266 179461 528304
rect 179431 528256 179557 528266
rect 179431 528236 179507 528256
rect 179335 528206 179389 528222
rect 179491 528222 179507 528236
rect 179541 528222 179557 528256
rect 179491 528212 179557 528222
rect 179098 528170 179152 528186
rect 178269 528138 178533 528160
rect 179005 528138 179035 528170
rect 178269 528112 178847 528138
rect 178081 528096 178111 528111
rect 179114 528061 179144 528170
rect 179335 528106 179365 528206
rect 179217 528076 179365 528106
rect 179407 528143 179461 528159
rect 179407 528109 179417 528143
rect 179451 528109 179461 528143
rect 179407 528093 179461 528109
rect 179217 528061 179247 528076
rect 179431 528061 179461 528093
rect 179503 528061 179533 528212
rect 179599 528159 179629 528304
rect 180109 528252 180687 528278
rect 180415 528230 180687 528252
rect 181029 528236 181059 528258
rect 181138 528236 181168 528304
rect 181234 528272 181264 528304
rect 181359 528272 181389 528304
rect 181234 528256 181317 528272
rect 179575 528143 179629 528159
rect 179575 528109 179585 528143
rect 179619 528109 179629 528143
rect 180109 528194 180373 528210
rect 180109 528160 180125 528194
rect 180159 528160 180224 528194
rect 180258 528160 180323 528194
rect 180357 528160 180373 528194
rect 180415 528196 180431 528230
rect 180465 528196 180534 528230
rect 180568 528196 180637 528230
rect 180671 528196 180687 528230
rect 180415 528180 180687 528196
rect 181026 528220 181080 528236
rect 181026 528186 181036 528220
rect 181070 528186 181080 528220
rect 181026 528170 181080 528186
rect 181122 528220 181176 528236
rect 181122 528186 181132 528220
rect 181166 528186 181176 528220
rect 181234 528222 181273 528256
rect 181307 528222 181317 528256
rect 181234 528206 181317 528222
rect 181359 528256 181413 528272
rect 181359 528222 181369 528256
rect 181403 528222 181413 528256
rect 181455 528266 181485 528304
rect 181455 528256 181581 528266
rect 181455 528236 181531 528256
rect 181359 528206 181413 528222
rect 181515 528222 181531 528236
rect 181565 528222 181581 528256
rect 181515 528212 181581 528222
rect 181122 528170 181176 528186
rect 180109 528138 180373 528160
rect 181029 528138 181059 528170
rect 179575 528093 179629 528109
rect 179599 528061 179629 528093
rect 180109 528112 180687 528138
rect 179114 527951 179144 527977
rect 179217 527951 179247 527977
rect 179431 527951 179461 527977
rect 179503 527951 179533 527977
rect 179599 527951 179629 527977
rect 181138 528061 181168 528170
rect 181359 528106 181389 528206
rect 181241 528076 181389 528106
rect 181431 528143 181485 528159
rect 181431 528109 181441 528143
rect 181475 528109 181485 528143
rect 181431 528093 181485 528109
rect 181241 528061 181271 528076
rect 181455 528061 181485 528093
rect 181527 528061 181557 528212
rect 181623 528159 181653 528304
rect 181857 528252 182803 528278
rect 182961 528252 183907 528278
rect 184065 528252 185011 528278
rect 185261 528252 186207 528278
rect 186365 528252 186943 528278
rect 182349 528230 182803 528252
rect 181599 528143 181653 528159
rect 181599 528109 181609 528143
rect 181643 528109 181653 528143
rect 181857 528194 182307 528210
rect 181857 528160 182129 528194
rect 182163 528160 182307 528194
rect 182349 528196 182493 528230
rect 182527 528196 182803 528230
rect 183453 528230 183907 528252
rect 182349 528180 182803 528196
rect 182961 528194 183411 528210
rect 181857 528138 182307 528160
rect 182961 528160 183233 528194
rect 183267 528160 183411 528194
rect 183453 528196 183597 528230
rect 183631 528196 183907 528230
rect 184557 528230 185011 528252
rect 183453 528180 183907 528196
rect 184065 528194 184515 528210
rect 182961 528138 183411 528160
rect 184065 528160 184337 528194
rect 184371 528160 184515 528194
rect 184557 528196 184701 528230
rect 184735 528196 185011 528230
rect 185753 528230 186207 528252
rect 184557 528180 185011 528196
rect 185261 528194 185711 528210
rect 184065 528138 184515 528160
rect 185261 528160 185533 528194
rect 185567 528160 185711 528194
rect 185753 528196 185897 528230
rect 185931 528196 186207 528230
rect 186671 528230 186943 528252
rect 187285 528252 187403 528278
rect 187285 528250 187323 528252
rect 185753 528180 186207 528196
rect 186365 528194 186629 528210
rect 185261 528138 185711 528160
rect 186365 528160 186381 528194
rect 186415 528160 186480 528194
rect 186514 528160 186579 528194
rect 186613 528160 186629 528194
rect 186671 528196 186687 528230
rect 186721 528196 186790 528230
rect 186824 528196 186893 528230
rect 186927 528196 186943 528230
rect 186671 528180 186943 528196
rect 187257 528234 187323 528250
rect 187257 528200 187273 528234
rect 187307 528200 187323 528234
rect 187257 528184 187323 528200
rect 187365 528194 187431 528210
rect 186365 528138 186629 528160
rect 187365 528160 187381 528194
rect 187415 528160 187431 528194
rect 187365 528144 187431 528160
rect 187365 528142 187403 528144
rect 181857 528112 182803 528138
rect 182961 528112 183907 528138
rect 184065 528112 185011 528138
rect 181599 528093 181653 528109
rect 181623 528061 181653 528093
rect 181138 527951 181168 527977
rect 181241 527951 181271 527977
rect 181455 527951 181485 527977
rect 181527 527951 181557 527977
rect 181623 527951 181653 527977
rect 185261 528112 186207 528138
rect 186365 528112 186943 528138
rect 187285 528112 187403 528142
rect 176504 527912 176534 527938
rect 176596 527912 176626 527938
rect 176695 527912 176725 527938
rect 176835 527912 176865 527938
rect 176932 527912 176962 527938
rect 177129 527912 177159 527938
rect 177228 527912 177258 527938
rect 177314 527912 177344 527938
rect 177398 527912 177428 527938
rect 177506 527912 177536 527938
rect 177590 527912 177620 527938
rect 177805 527912 177835 527938
rect 177993 527912 178023 527938
rect 178081 527912 178111 527938
rect 178269 527912 178847 527938
rect 179005 527912 179035 527938
rect 180109 527912 180687 527938
rect 181029 527912 181059 527938
rect 181857 527912 182803 527938
rect 182961 527912 183907 527938
rect 184065 527912 185011 527938
rect 185261 527912 186207 527938
rect 186365 527912 186943 527938
rect 187285 527912 187403 527938
rect 172289 527844 172407 527870
rect 172565 527844 173511 527870
rect 173669 527844 174615 527870
rect 174773 527844 175719 527870
rect 175877 527844 176271 527870
rect 176448 527844 176478 527870
rect 176543 527844 176643 527870
rect 176801 527844 176901 527870
rect 176955 527844 176985 527870
rect 177165 527844 177283 527870
rect 177533 527844 178479 527870
rect 178637 527844 178847 527870
rect 179024 527844 179054 527870
rect 179119 527844 179219 527870
rect 179377 527844 179477 527870
rect 179531 527844 179561 527870
rect 179741 527844 180687 527870
rect 180845 527844 181791 527870
rect 181949 527844 182343 527870
rect 182685 527844 183631 527870
rect 183789 527844 184735 527870
rect 184893 527844 185839 527870
rect 185997 527844 186943 527870
rect 187285 527844 187403 527870
rect 172289 527640 172407 527670
rect 172565 527644 173511 527670
rect 173669 527644 174615 527670
rect 174773 527644 175719 527670
rect 175877 527644 176271 527670
rect 172289 527638 172327 527640
rect 172261 527622 172327 527638
rect 172261 527588 172277 527622
rect 172311 527588 172327 527622
rect 172565 527622 173015 527644
rect 172261 527572 172327 527588
rect 172369 527582 172435 527598
rect 172369 527548 172385 527582
rect 172419 527548 172435 527582
rect 172565 527588 172837 527622
rect 172871 527588 173015 527622
rect 173669 527622 174119 527644
rect 172565 527572 173015 527588
rect 173057 527586 173511 527602
rect 172369 527532 172435 527548
rect 173057 527552 173201 527586
rect 173235 527552 173511 527586
rect 173669 527588 173941 527622
rect 173975 527588 174119 527622
rect 174773 527622 175223 527644
rect 173669 527572 174119 527588
rect 174161 527586 174615 527602
rect 172369 527530 172407 527532
rect 173057 527530 173511 527552
rect 174161 527552 174305 527586
rect 174339 527552 174615 527586
rect 174773 527588 175045 527622
rect 175079 527588 175223 527622
rect 175877 527622 176053 527644
rect 174773 527572 175223 527588
rect 175265 527586 175719 527602
rect 174161 527530 174615 527552
rect 175265 527552 175409 527586
rect 175443 527552 175719 527586
rect 175877 527588 175893 527622
rect 175927 527588 176003 527622
rect 176037 527588 176053 527622
rect 176448 527612 176478 527644
rect 176543 527612 176643 527760
rect 175877 527572 176053 527588
rect 176095 527586 176271 527602
rect 175265 527530 175719 527552
rect 176095 527552 176111 527586
rect 176145 527552 176221 527586
rect 176255 527552 176271 527586
rect 176095 527530 176271 527552
rect 176447 527596 176501 527612
rect 176447 527562 176457 527596
rect 176491 527562 176501 527596
rect 176447 527546 176501 527562
rect 176543 527596 176697 527612
rect 176543 527562 176653 527596
rect 176687 527562 176697 527596
rect 176543 527546 176697 527562
rect 176801 527596 176901 527760
rect 176801 527562 176857 527596
rect 176891 527562 176901 527596
rect 172289 527504 172407 527530
rect 172565 527504 173511 527530
rect 173669 527504 174615 527530
rect 174773 527504 175719 527530
rect 175877 527504 176271 527530
rect 176448 527524 176478 527546
rect 176543 527478 176643 527546
rect 176801 527478 176901 527562
rect 176955 527612 176985 527760
rect 177165 527640 177283 527670
rect 177533 527644 178479 527670
rect 178637 527644 178847 527670
rect 177165 527638 177203 527640
rect 177137 527622 177203 527638
rect 176955 527596 177015 527612
rect 176955 527562 176971 527596
rect 177005 527562 177015 527596
rect 177137 527588 177153 527622
rect 177187 527588 177203 527622
rect 177533 527622 177983 527644
rect 178637 527638 178721 527644
rect 177137 527572 177203 527588
rect 177245 527582 177311 527598
rect 176955 527546 177015 527562
rect 177245 527548 177261 527582
rect 177295 527548 177311 527582
rect 177533 527588 177805 527622
rect 177839 527588 177983 527622
rect 178579 527622 178721 527638
rect 177533 527572 177983 527588
rect 178025 527586 178479 527602
rect 176955 527478 176985 527546
rect 177245 527532 177311 527548
rect 178025 527552 178169 527586
rect 178203 527552 178479 527586
rect 178579 527588 178595 527622
rect 178629 527588 178721 527622
rect 179024 527612 179054 527644
rect 179119 527612 179219 527760
rect 178579 527572 178721 527588
rect 178763 527586 178905 527602
rect 177245 527530 177283 527532
rect 178025 527530 178479 527552
rect 178763 527552 178855 527586
rect 178889 527552 178905 527586
rect 178763 527536 178905 527552
rect 179023 527596 179077 527612
rect 179023 527562 179033 527596
rect 179067 527562 179077 527596
rect 179023 527546 179077 527562
rect 179119 527596 179273 527612
rect 179119 527562 179229 527596
rect 179263 527562 179273 527596
rect 179119 527546 179273 527562
rect 179377 527596 179477 527760
rect 179377 527562 179433 527596
rect 179467 527562 179477 527596
rect 178763 527530 178847 527536
rect 177165 527504 177283 527530
rect 177533 527504 178479 527530
rect 178637 527504 178847 527530
rect 179024 527524 179054 527546
rect 179119 527478 179219 527546
rect 179377 527478 179477 527562
rect 179531 527612 179561 527760
rect 179741 527644 180687 527670
rect 180845 527644 181791 527670
rect 181949 527644 182343 527670
rect 182685 527644 183631 527670
rect 183789 527644 184735 527670
rect 184893 527644 185839 527670
rect 185997 527644 186943 527670
rect 179741 527622 180191 527644
rect 179531 527596 179591 527612
rect 179531 527562 179547 527596
rect 179581 527562 179591 527596
rect 179741 527588 180013 527622
rect 180047 527588 180191 527622
rect 180845 527622 181295 527644
rect 179741 527572 180191 527588
rect 180233 527586 180687 527602
rect 179531 527546 179591 527562
rect 180233 527552 180377 527586
rect 180411 527552 180687 527586
rect 180845 527588 181117 527622
rect 181151 527588 181295 527622
rect 181949 527622 182125 527644
rect 180845 527572 181295 527588
rect 181337 527586 181791 527602
rect 179531 527478 179561 527546
rect 180233 527530 180687 527552
rect 181337 527552 181481 527586
rect 181515 527552 181791 527586
rect 181949 527588 181965 527622
rect 181999 527588 182075 527622
rect 182109 527588 182125 527622
rect 182685 527622 183135 527644
rect 181949 527572 182125 527588
rect 182167 527586 182343 527602
rect 181337 527530 181791 527552
rect 182167 527552 182183 527586
rect 182217 527552 182293 527586
rect 182327 527552 182343 527586
rect 182685 527588 182957 527622
rect 182991 527588 183135 527622
rect 183789 527622 184239 527644
rect 182685 527572 183135 527588
rect 183177 527586 183631 527602
rect 182167 527530 182343 527552
rect 183177 527552 183321 527586
rect 183355 527552 183631 527586
rect 183789 527588 184061 527622
rect 184095 527588 184239 527622
rect 184893 527622 185343 527644
rect 183789 527572 184239 527588
rect 184281 527586 184735 527602
rect 183177 527530 183631 527552
rect 184281 527552 184425 527586
rect 184459 527552 184735 527586
rect 184893 527588 185165 527622
rect 185199 527588 185343 527622
rect 185997 527622 186447 527644
rect 187285 527640 187403 527670
rect 184893 527572 185343 527588
rect 185385 527586 185839 527602
rect 184281 527530 184735 527552
rect 185385 527552 185529 527586
rect 185563 527552 185839 527586
rect 185997 527588 186269 527622
rect 186303 527588 186447 527622
rect 187365 527638 187403 527640
rect 187365 527622 187431 527638
rect 185997 527572 186447 527588
rect 186489 527586 186943 527602
rect 185385 527530 185839 527552
rect 186489 527552 186633 527586
rect 186667 527552 186943 527586
rect 186489 527530 186943 527552
rect 187257 527582 187323 527598
rect 187257 527548 187273 527582
rect 187307 527548 187323 527582
rect 187365 527588 187381 527622
rect 187415 527588 187431 527622
rect 187365 527572 187431 527588
rect 187257 527532 187323 527548
rect 179741 527504 180687 527530
rect 180845 527504 181791 527530
rect 181949 527504 182343 527530
rect 182685 527504 183631 527530
rect 183789 527504 184735 527530
rect 184893 527504 185839 527530
rect 185997 527504 186943 527530
rect 187285 527530 187323 527532
rect 187285 527504 187403 527530
rect 172289 527368 172407 527394
rect 172565 527368 173511 527394
rect 173669 527368 174615 527394
rect 174773 527368 175719 527394
rect 175877 527368 176271 527394
rect 176448 527368 176478 527394
rect 176543 527368 176643 527394
rect 176801 527368 176901 527394
rect 176955 527368 176985 527394
rect 177165 527368 177283 527394
rect 177533 527368 178479 527394
rect 178637 527368 178847 527394
rect 179024 527368 179054 527394
rect 179119 527368 179219 527394
rect 179377 527368 179477 527394
rect 179531 527368 179561 527394
rect 179741 527368 180687 527394
rect 180845 527368 181791 527394
rect 181949 527368 182343 527394
rect 182685 527368 183631 527394
rect 183789 527368 184735 527394
rect 184893 527368 185839 527394
rect 185997 527368 186943 527394
rect 187285 527368 187403 527394
rect 172289 527300 172407 527326
rect 172565 527300 173511 527326
rect 173669 527300 174615 527326
rect 174957 527300 175903 527326
rect 176061 527300 177007 527326
rect 177165 527300 178111 527326
rect 178269 527300 179215 527326
rect 179373 527300 179767 527326
rect 180109 527300 181055 527326
rect 181213 527300 182159 527326
rect 182317 527300 183263 527326
rect 183421 527300 184367 527326
rect 184525 527300 184919 527326
rect 185261 527300 186207 527326
rect 186365 527300 186943 527326
rect 187285 527300 187403 527326
rect 172289 527164 172407 527190
rect 172565 527164 173511 527190
rect 173669 527164 174615 527190
rect 174957 527164 175903 527190
rect 176061 527164 177007 527190
rect 177165 527164 178111 527190
rect 178269 527164 179215 527190
rect 179373 527164 179767 527190
rect 180109 527164 181055 527190
rect 181213 527164 182159 527190
rect 182317 527164 183263 527190
rect 183421 527164 184367 527190
rect 184525 527164 184919 527190
rect 185261 527164 186207 527190
rect 186365 527164 186943 527190
rect 172369 527162 172407 527164
rect 172369 527146 172435 527162
rect 172261 527106 172327 527122
rect 172261 527072 172277 527106
rect 172311 527072 172327 527106
rect 172369 527112 172385 527146
rect 172419 527112 172435 527146
rect 173057 527142 173511 527164
rect 172369 527096 172435 527112
rect 172565 527106 173015 527122
rect 172261 527056 172327 527072
rect 172289 527054 172327 527056
rect 172565 527072 172837 527106
rect 172871 527072 173015 527106
rect 173057 527108 173201 527142
rect 173235 527108 173511 527142
rect 174161 527142 174615 527164
rect 173057 527092 173511 527108
rect 173669 527106 174119 527122
rect 172289 527024 172407 527054
rect 172565 527050 173015 527072
rect 173669 527072 173941 527106
rect 173975 527072 174119 527106
rect 174161 527108 174305 527142
rect 174339 527108 174615 527142
rect 175449 527142 175903 527164
rect 174161 527092 174615 527108
rect 174957 527106 175407 527122
rect 173669 527050 174119 527072
rect 174957 527072 175229 527106
rect 175263 527072 175407 527106
rect 175449 527108 175593 527142
rect 175627 527108 175903 527142
rect 176553 527142 177007 527164
rect 175449 527092 175903 527108
rect 176061 527106 176511 527122
rect 174957 527050 175407 527072
rect 176061 527072 176333 527106
rect 176367 527072 176511 527106
rect 176553 527108 176697 527142
rect 176731 527108 177007 527142
rect 177657 527142 178111 527164
rect 176553 527092 177007 527108
rect 177165 527106 177615 527122
rect 176061 527050 176511 527072
rect 177165 527072 177437 527106
rect 177471 527072 177615 527106
rect 177657 527108 177801 527142
rect 177835 527108 178111 527142
rect 178761 527142 179215 527164
rect 177657 527092 178111 527108
rect 178269 527106 178719 527122
rect 177165 527050 177615 527072
rect 178269 527072 178541 527106
rect 178575 527072 178719 527106
rect 178761 527108 178905 527142
rect 178939 527108 179215 527142
rect 179591 527142 179767 527164
rect 178761 527092 179215 527108
rect 179373 527106 179549 527122
rect 178269 527050 178719 527072
rect 179373 527072 179389 527106
rect 179423 527072 179499 527106
rect 179533 527072 179549 527106
rect 179591 527108 179607 527142
rect 179641 527108 179717 527142
rect 179751 527108 179767 527142
rect 180601 527142 181055 527164
rect 179591 527092 179767 527108
rect 180109 527106 180559 527122
rect 179373 527050 179549 527072
rect 180109 527072 180381 527106
rect 180415 527072 180559 527106
rect 180601 527108 180745 527142
rect 180779 527108 181055 527142
rect 181705 527142 182159 527164
rect 180601 527092 181055 527108
rect 181213 527106 181663 527122
rect 180109 527050 180559 527072
rect 181213 527072 181485 527106
rect 181519 527072 181663 527106
rect 181705 527108 181849 527142
rect 181883 527108 182159 527142
rect 182809 527142 183263 527164
rect 181705 527092 182159 527108
rect 182317 527106 182767 527122
rect 181213 527050 181663 527072
rect 182317 527072 182589 527106
rect 182623 527072 182767 527106
rect 182809 527108 182953 527142
rect 182987 527108 183263 527142
rect 183913 527142 184367 527164
rect 182809 527092 183263 527108
rect 183421 527106 183871 527122
rect 182317 527050 182767 527072
rect 183421 527072 183693 527106
rect 183727 527072 183871 527106
rect 183913 527108 184057 527142
rect 184091 527108 184367 527142
rect 184743 527142 184919 527164
rect 183913 527092 184367 527108
rect 184525 527106 184701 527122
rect 183421 527050 183871 527072
rect 184525 527072 184541 527106
rect 184575 527072 184651 527106
rect 184685 527072 184701 527106
rect 184743 527108 184759 527142
rect 184793 527108 184869 527142
rect 184903 527108 184919 527142
rect 185753 527142 186207 527164
rect 184743 527092 184919 527108
rect 185261 527106 185711 527122
rect 184525 527050 184701 527072
rect 185261 527072 185533 527106
rect 185567 527072 185711 527106
rect 185753 527108 185897 527142
rect 185931 527108 186207 527142
rect 186671 527142 186943 527164
rect 187285 527164 187403 527190
rect 187285 527162 187323 527164
rect 185753 527092 186207 527108
rect 186365 527106 186629 527122
rect 185261 527050 185711 527072
rect 186365 527072 186381 527106
rect 186415 527072 186480 527106
rect 186514 527072 186579 527106
rect 186613 527072 186629 527106
rect 186671 527108 186687 527142
rect 186721 527108 186790 527142
rect 186824 527108 186893 527142
rect 186927 527108 186943 527142
rect 186671 527092 186943 527108
rect 187257 527146 187323 527162
rect 187257 527112 187273 527146
rect 187307 527112 187323 527146
rect 187257 527096 187323 527112
rect 187365 527106 187431 527122
rect 186365 527050 186629 527072
rect 187365 527072 187381 527106
rect 187415 527072 187431 527106
rect 187365 527056 187431 527072
rect 187365 527054 187403 527056
rect 172565 527024 173511 527050
rect 173669 527024 174615 527050
rect 174957 527024 175903 527050
rect 176061 527024 177007 527050
rect 177165 527024 178111 527050
rect 178269 527024 179215 527050
rect 179373 527024 179767 527050
rect 180109 527024 181055 527050
rect 181213 527024 182159 527050
rect 182317 527024 183263 527050
rect 183421 527024 184367 527050
rect 184525 527024 184919 527050
rect 185261 527024 186207 527050
rect 186365 527024 186943 527050
rect 187285 527024 187403 527054
rect 172289 526824 172407 526850
rect 172565 526824 173511 526850
rect 173669 526824 174615 526850
rect 174957 526824 175903 526850
rect 176061 526824 177007 526850
rect 177165 526824 178111 526850
rect 178269 526824 179215 526850
rect 179373 526824 179767 526850
rect 180109 526824 181055 526850
rect 181213 526824 182159 526850
rect 182317 526824 183263 526850
rect 183421 526824 184367 526850
rect 184525 526824 184919 526850
rect 185261 526824 186207 526850
rect 186365 526824 186943 526850
rect 187285 526824 187403 526850
rect 172289 526756 172407 526782
rect 172565 526756 173511 526782
rect 173669 526756 174615 526782
rect 174773 526756 175719 526782
rect 175877 526756 176823 526782
rect 176981 526756 177191 526782
rect 177533 526756 178479 526782
rect 178637 526756 179583 526782
rect 179741 526756 180687 526782
rect 180845 526756 181791 526782
rect 181949 526756 182343 526782
rect 182685 526756 183631 526782
rect 183789 526756 184735 526782
rect 184893 526756 185839 526782
rect 185997 526756 186943 526782
rect 187285 526756 187403 526782
rect 172289 526552 172407 526582
rect 172565 526556 173511 526582
rect 173669 526556 174615 526582
rect 174773 526556 175719 526582
rect 175877 526556 176823 526582
rect 176981 526556 177191 526582
rect 177533 526556 178479 526582
rect 178637 526556 179583 526582
rect 179741 526556 180687 526582
rect 180845 526556 181791 526582
rect 181949 526556 182343 526582
rect 182685 526556 183631 526582
rect 183789 526556 184735 526582
rect 184893 526556 185839 526582
rect 185997 526556 186943 526582
rect 172289 526550 172327 526552
rect 172261 526534 172327 526550
rect 172261 526500 172277 526534
rect 172311 526500 172327 526534
rect 172565 526534 173015 526556
rect 172261 526484 172327 526500
rect 172369 526494 172435 526510
rect 172369 526460 172385 526494
rect 172419 526460 172435 526494
rect 172565 526500 172837 526534
rect 172871 526500 173015 526534
rect 173669 526534 174119 526556
rect 172565 526484 173015 526500
rect 173057 526498 173511 526514
rect 172369 526444 172435 526460
rect 173057 526464 173201 526498
rect 173235 526464 173511 526498
rect 173669 526500 173941 526534
rect 173975 526500 174119 526534
rect 174773 526534 175223 526556
rect 173669 526484 174119 526500
rect 174161 526498 174615 526514
rect 172369 526442 172407 526444
rect 173057 526442 173511 526464
rect 174161 526464 174305 526498
rect 174339 526464 174615 526498
rect 174773 526500 175045 526534
rect 175079 526500 175223 526534
rect 175877 526534 176327 526556
rect 176981 526550 177065 526556
rect 174773 526484 175223 526500
rect 175265 526498 175719 526514
rect 174161 526442 174615 526464
rect 175265 526464 175409 526498
rect 175443 526464 175719 526498
rect 175877 526500 176149 526534
rect 176183 526500 176327 526534
rect 176923 526534 177065 526550
rect 175877 526484 176327 526500
rect 176369 526498 176823 526514
rect 175265 526442 175719 526464
rect 176369 526464 176513 526498
rect 176547 526464 176823 526498
rect 176923 526500 176939 526534
rect 176973 526500 177065 526534
rect 177533 526534 177983 526556
rect 176923 526484 177065 526500
rect 177107 526498 177249 526514
rect 176369 526442 176823 526464
rect 177107 526464 177199 526498
rect 177233 526464 177249 526498
rect 177533 526500 177805 526534
rect 177839 526500 177983 526534
rect 178637 526534 179087 526556
rect 177533 526484 177983 526500
rect 178025 526498 178479 526514
rect 177107 526448 177249 526464
rect 178025 526464 178169 526498
rect 178203 526464 178479 526498
rect 178637 526500 178909 526534
rect 178943 526500 179087 526534
rect 179741 526534 180191 526556
rect 178637 526484 179087 526500
rect 179129 526498 179583 526514
rect 177107 526442 177191 526448
rect 178025 526442 178479 526464
rect 179129 526464 179273 526498
rect 179307 526464 179583 526498
rect 179741 526500 180013 526534
rect 180047 526500 180191 526534
rect 180845 526534 181295 526556
rect 179741 526484 180191 526500
rect 180233 526498 180687 526514
rect 179129 526442 179583 526464
rect 180233 526464 180377 526498
rect 180411 526464 180687 526498
rect 180845 526500 181117 526534
rect 181151 526500 181295 526534
rect 181949 526534 182125 526556
rect 180845 526484 181295 526500
rect 181337 526498 181791 526514
rect 180233 526442 180687 526464
rect 181337 526464 181481 526498
rect 181515 526464 181791 526498
rect 181949 526500 181965 526534
rect 181999 526500 182075 526534
rect 182109 526500 182125 526534
rect 182685 526534 183135 526556
rect 181949 526484 182125 526500
rect 182167 526498 182343 526514
rect 181337 526442 181791 526464
rect 182167 526464 182183 526498
rect 182217 526464 182293 526498
rect 182327 526464 182343 526498
rect 182685 526500 182957 526534
rect 182991 526500 183135 526534
rect 183789 526534 184239 526556
rect 182685 526484 183135 526500
rect 183177 526498 183631 526514
rect 182167 526442 182343 526464
rect 183177 526464 183321 526498
rect 183355 526464 183631 526498
rect 183789 526500 184061 526534
rect 184095 526500 184239 526534
rect 184893 526534 185343 526556
rect 183789 526484 184239 526500
rect 184281 526498 184735 526514
rect 183177 526442 183631 526464
rect 184281 526464 184425 526498
rect 184459 526464 184735 526498
rect 184893 526500 185165 526534
rect 185199 526500 185343 526534
rect 185997 526534 186447 526556
rect 187285 526552 187403 526582
rect 184893 526484 185343 526500
rect 185385 526498 185839 526514
rect 184281 526442 184735 526464
rect 185385 526464 185529 526498
rect 185563 526464 185839 526498
rect 185997 526500 186269 526534
rect 186303 526500 186447 526534
rect 187365 526550 187403 526552
rect 187365 526534 187431 526550
rect 185997 526484 186447 526500
rect 186489 526498 186943 526514
rect 185385 526442 185839 526464
rect 186489 526464 186633 526498
rect 186667 526464 186943 526498
rect 186489 526442 186943 526464
rect 187257 526494 187323 526510
rect 187257 526460 187273 526494
rect 187307 526460 187323 526494
rect 187365 526500 187381 526534
rect 187415 526500 187431 526534
rect 187365 526484 187431 526500
rect 187257 526444 187323 526460
rect 172289 526416 172407 526442
rect 172565 526416 173511 526442
rect 173669 526416 174615 526442
rect 174773 526416 175719 526442
rect 175877 526416 176823 526442
rect 176981 526416 177191 526442
rect 177533 526416 178479 526442
rect 178637 526416 179583 526442
rect 179741 526416 180687 526442
rect 180845 526416 181791 526442
rect 181949 526416 182343 526442
rect 182685 526416 183631 526442
rect 183789 526416 184735 526442
rect 184893 526416 185839 526442
rect 185997 526416 186943 526442
rect 187285 526442 187323 526444
rect 187285 526416 187403 526442
rect 172289 526280 172407 526306
rect 172565 526280 173511 526306
rect 173669 526280 174615 526306
rect 174773 526280 175719 526306
rect 175877 526280 176823 526306
rect 176981 526280 177191 526306
rect 177533 526280 178479 526306
rect 178637 526280 179583 526306
rect 179741 526280 180687 526306
rect 180845 526280 181791 526306
rect 181949 526280 182343 526306
rect 182685 526280 183631 526306
rect 183789 526280 184735 526306
rect 184893 526280 185839 526306
rect 185997 526280 186943 526306
rect 187285 526280 187403 526306
rect 172289 526212 172407 526238
rect 172565 526212 173511 526238
rect 173669 526212 174615 526238
rect 174957 526212 175903 526238
rect 176061 526212 177007 526238
rect 177165 526212 178111 526238
rect 178269 526212 179215 526238
rect 179373 526212 179767 526238
rect 180109 526212 181055 526238
rect 181213 526212 182159 526238
rect 182317 526212 183263 526238
rect 183421 526212 184367 526238
rect 184525 526212 184919 526238
rect 185261 526212 186207 526238
rect 186365 526212 186943 526238
rect 187285 526212 187403 526238
rect 172289 526076 172407 526102
rect 172565 526076 173511 526102
rect 173669 526076 174615 526102
rect 174957 526076 175903 526102
rect 176061 526076 177007 526102
rect 177165 526076 178111 526102
rect 178269 526076 179215 526102
rect 179373 526076 179767 526102
rect 180109 526076 181055 526102
rect 181213 526076 182159 526102
rect 182317 526076 183263 526102
rect 183421 526076 184367 526102
rect 184525 526076 184919 526102
rect 185261 526076 186207 526102
rect 186365 526076 186943 526102
rect 172369 526074 172407 526076
rect 172369 526058 172435 526074
rect 172261 526018 172327 526034
rect 172261 525984 172277 526018
rect 172311 525984 172327 526018
rect 172369 526024 172385 526058
rect 172419 526024 172435 526058
rect 173057 526054 173511 526076
rect 172369 526008 172435 526024
rect 172565 526018 173015 526034
rect 172261 525968 172327 525984
rect 172289 525966 172327 525968
rect 172565 525984 172837 526018
rect 172871 525984 173015 526018
rect 173057 526020 173201 526054
rect 173235 526020 173511 526054
rect 174161 526054 174615 526076
rect 173057 526004 173511 526020
rect 173669 526018 174119 526034
rect 172289 525936 172407 525966
rect 172565 525962 173015 525984
rect 173669 525984 173941 526018
rect 173975 525984 174119 526018
rect 174161 526020 174305 526054
rect 174339 526020 174615 526054
rect 175449 526054 175903 526076
rect 174161 526004 174615 526020
rect 174957 526018 175407 526034
rect 173669 525962 174119 525984
rect 174957 525984 175229 526018
rect 175263 525984 175407 526018
rect 175449 526020 175593 526054
rect 175627 526020 175903 526054
rect 176553 526054 177007 526076
rect 175449 526004 175903 526020
rect 176061 526018 176511 526034
rect 174957 525962 175407 525984
rect 176061 525984 176333 526018
rect 176367 525984 176511 526018
rect 176553 526020 176697 526054
rect 176731 526020 177007 526054
rect 177657 526054 178111 526076
rect 176553 526004 177007 526020
rect 177165 526018 177615 526034
rect 176061 525962 176511 525984
rect 177165 525984 177437 526018
rect 177471 525984 177615 526018
rect 177657 526020 177801 526054
rect 177835 526020 178111 526054
rect 178761 526054 179215 526076
rect 177657 526004 178111 526020
rect 178269 526018 178719 526034
rect 177165 525962 177615 525984
rect 178269 525984 178541 526018
rect 178575 525984 178719 526018
rect 178761 526020 178905 526054
rect 178939 526020 179215 526054
rect 179591 526054 179767 526076
rect 178761 526004 179215 526020
rect 179373 526018 179549 526034
rect 178269 525962 178719 525984
rect 179373 525984 179389 526018
rect 179423 525984 179499 526018
rect 179533 525984 179549 526018
rect 179591 526020 179607 526054
rect 179641 526020 179717 526054
rect 179751 526020 179767 526054
rect 180601 526054 181055 526076
rect 179591 526004 179767 526020
rect 180109 526018 180559 526034
rect 179373 525962 179549 525984
rect 180109 525984 180381 526018
rect 180415 525984 180559 526018
rect 180601 526020 180745 526054
rect 180779 526020 181055 526054
rect 181705 526054 182159 526076
rect 180601 526004 181055 526020
rect 181213 526018 181663 526034
rect 180109 525962 180559 525984
rect 181213 525984 181485 526018
rect 181519 525984 181663 526018
rect 181705 526020 181849 526054
rect 181883 526020 182159 526054
rect 182809 526054 183263 526076
rect 181705 526004 182159 526020
rect 182317 526018 182767 526034
rect 181213 525962 181663 525984
rect 182317 525984 182589 526018
rect 182623 525984 182767 526018
rect 182809 526020 182953 526054
rect 182987 526020 183263 526054
rect 183913 526054 184367 526076
rect 182809 526004 183263 526020
rect 183421 526018 183871 526034
rect 182317 525962 182767 525984
rect 183421 525984 183693 526018
rect 183727 525984 183871 526018
rect 183913 526020 184057 526054
rect 184091 526020 184367 526054
rect 184743 526054 184919 526076
rect 183913 526004 184367 526020
rect 184525 526018 184701 526034
rect 183421 525962 183871 525984
rect 184525 525984 184541 526018
rect 184575 525984 184651 526018
rect 184685 525984 184701 526018
rect 184743 526020 184759 526054
rect 184793 526020 184869 526054
rect 184903 526020 184919 526054
rect 185753 526054 186207 526076
rect 184743 526004 184919 526020
rect 185261 526018 185711 526034
rect 184525 525962 184701 525984
rect 185261 525984 185533 526018
rect 185567 525984 185711 526018
rect 185753 526020 185897 526054
rect 185931 526020 186207 526054
rect 186671 526054 186943 526076
rect 187285 526076 187403 526102
rect 187285 526074 187323 526076
rect 185753 526004 186207 526020
rect 186365 526018 186629 526034
rect 185261 525962 185711 525984
rect 186365 525984 186381 526018
rect 186415 525984 186480 526018
rect 186514 525984 186579 526018
rect 186613 525984 186629 526018
rect 186671 526020 186687 526054
rect 186721 526020 186790 526054
rect 186824 526020 186893 526054
rect 186927 526020 186943 526054
rect 186671 526004 186943 526020
rect 187257 526058 187323 526074
rect 187257 526024 187273 526058
rect 187307 526024 187323 526058
rect 187257 526008 187323 526024
rect 187365 526018 187431 526034
rect 186365 525962 186629 525984
rect 187365 525984 187381 526018
rect 187415 525984 187431 526018
rect 187365 525968 187431 525984
rect 187365 525966 187403 525968
rect 172565 525936 173511 525962
rect 173669 525936 174615 525962
rect 174957 525936 175903 525962
rect 176061 525936 177007 525962
rect 177165 525936 178111 525962
rect 178269 525936 179215 525962
rect 179373 525936 179767 525962
rect 180109 525936 181055 525962
rect 181213 525936 182159 525962
rect 182317 525936 183263 525962
rect 183421 525936 184367 525962
rect 184525 525936 184919 525962
rect 185261 525936 186207 525962
rect 186365 525936 186943 525962
rect 187285 525936 187403 525966
rect 172289 525736 172407 525762
rect 172565 525736 173511 525762
rect 173669 525736 174615 525762
rect 174957 525736 175903 525762
rect 176061 525736 177007 525762
rect 177165 525736 178111 525762
rect 178269 525736 179215 525762
rect 179373 525736 179767 525762
rect 180109 525736 181055 525762
rect 181213 525736 182159 525762
rect 182317 525736 183263 525762
rect 183421 525736 184367 525762
rect 184525 525736 184919 525762
rect 185261 525736 186207 525762
rect 186365 525736 186943 525762
rect 187285 525736 187403 525762
rect 172289 525668 172407 525694
rect 172565 525668 173511 525694
rect 173669 525668 174615 525694
rect 174773 525668 175719 525694
rect 175877 525668 176823 525694
rect 176981 525668 177191 525694
rect 177533 525668 178479 525694
rect 178637 525668 179583 525694
rect 179741 525668 180687 525694
rect 180845 525668 181791 525694
rect 181949 525668 182343 525694
rect 182685 525668 183631 525694
rect 183789 525668 184735 525694
rect 184893 525668 185839 525694
rect 185997 525668 186943 525694
rect 187285 525668 187403 525694
rect 172289 525464 172407 525494
rect 172565 525468 173511 525494
rect 173669 525468 174615 525494
rect 174773 525468 175719 525494
rect 175877 525468 176823 525494
rect 176981 525468 177191 525494
rect 177533 525468 178479 525494
rect 178637 525468 179583 525494
rect 179741 525468 180687 525494
rect 180845 525468 181791 525494
rect 181949 525468 182343 525494
rect 182685 525468 183631 525494
rect 183789 525468 184735 525494
rect 184893 525468 185839 525494
rect 185997 525468 186943 525494
rect 172289 525462 172327 525464
rect 172261 525446 172327 525462
rect 172261 525412 172277 525446
rect 172311 525412 172327 525446
rect 172565 525446 173015 525468
rect 172261 525396 172327 525412
rect 172369 525406 172435 525422
rect 172369 525372 172385 525406
rect 172419 525372 172435 525406
rect 172565 525412 172837 525446
rect 172871 525412 173015 525446
rect 173669 525446 174119 525468
rect 172565 525396 173015 525412
rect 173057 525410 173511 525426
rect 172369 525356 172435 525372
rect 173057 525376 173201 525410
rect 173235 525376 173511 525410
rect 173669 525412 173941 525446
rect 173975 525412 174119 525446
rect 174773 525446 175223 525468
rect 173669 525396 174119 525412
rect 174161 525410 174615 525426
rect 172369 525354 172407 525356
rect 173057 525354 173511 525376
rect 174161 525376 174305 525410
rect 174339 525376 174615 525410
rect 174773 525412 175045 525446
rect 175079 525412 175223 525446
rect 175877 525446 176327 525468
rect 176981 525462 177065 525468
rect 174773 525396 175223 525412
rect 175265 525410 175719 525426
rect 174161 525354 174615 525376
rect 175265 525376 175409 525410
rect 175443 525376 175719 525410
rect 175877 525412 176149 525446
rect 176183 525412 176327 525446
rect 176923 525446 177065 525462
rect 175877 525396 176327 525412
rect 176369 525410 176823 525426
rect 175265 525354 175719 525376
rect 176369 525376 176513 525410
rect 176547 525376 176823 525410
rect 176923 525412 176939 525446
rect 176973 525412 177065 525446
rect 177533 525446 177983 525468
rect 176923 525396 177065 525412
rect 177107 525410 177249 525426
rect 176369 525354 176823 525376
rect 177107 525376 177199 525410
rect 177233 525376 177249 525410
rect 177533 525412 177805 525446
rect 177839 525412 177983 525446
rect 178637 525446 179087 525468
rect 177533 525396 177983 525412
rect 178025 525410 178479 525426
rect 177107 525360 177249 525376
rect 178025 525376 178169 525410
rect 178203 525376 178479 525410
rect 178637 525412 178909 525446
rect 178943 525412 179087 525446
rect 179741 525446 180191 525468
rect 178637 525396 179087 525412
rect 179129 525410 179583 525426
rect 177107 525354 177191 525360
rect 178025 525354 178479 525376
rect 179129 525376 179273 525410
rect 179307 525376 179583 525410
rect 179741 525412 180013 525446
rect 180047 525412 180191 525446
rect 180845 525446 181295 525468
rect 179741 525396 180191 525412
rect 180233 525410 180687 525426
rect 179129 525354 179583 525376
rect 180233 525376 180377 525410
rect 180411 525376 180687 525410
rect 180845 525412 181117 525446
rect 181151 525412 181295 525446
rect 181949 525446 182125 525468
rect 180845 525396 181295 525412
rect 181337 525410 181791 525426
rect 180233 525354 180687 525376
rect 181337 525376 181481 525410
rect 181515 525376 181791 525410
rect 181949 525412 181965 525446
rect 181999 525412 182075 525446
rect 182109 525412 182125 525446
rect 182685 525446 183135 525468
rect 181949 525396 182125 525412
rect 182167 525410 182343 525426
rect 181337 525354 181791 525376
rect 182167 525376 182183 525410
rect 182217 525376 182293 525410
rect 182327 525376 182343 525410
rect 182685 525412 182957 525446
rect 182991 525412 183135 525446
rect 183789 525446 184239 525468
rect 182685 525396 183135 525412
rect 183177 525410 183631 525426
rect 182167 525354 182343 525376
rect 183177 525376 183321 525410
rect 183355 525376 183631 525410
rect 183789 525412 184061 525446
rect 184095 525412 184239 525446
rect 184893 525446 185343 525468
rect 183789 525396 184239 525412
rect 184281 525410 184735 525426
rect 183177 525354 183631 525376
rect 184281 525376 184425 525410
rect 184459 525376 184735 525410
rect 184893 525412 185165 525446
rect 185199 525412 185343 525446
rect 185997 525446 186447 525468
rect 187285 525464 187403 525494
rect 184893 525396 185343 525412
rect 185385 525410 185839 525426
rect 184281 525354 184735 525376
rect 185385 525376 185529 525410
rect 185563 525376 185839 525410
rect 185997 525412 186269 525446
rect 186303 525412 186447 525446
rect 187365 525462 187403 525464
rect 187365 525446 187431 525462
rect 185997 525396 186447 525412
rect 186489 525410 186943 525426
rect 185385 525354 185839 525376
rect 186489 525376 186633 525410
rect 186667 525376 186943 525410
rect 186489 525354 186943 525376
rect 187257 525406 187323 525422
rect 187257 525372 187273 525406
rect 187307 525372 187323 525406
rect 187365 525412 187381 525446
rect 187415 525412 187431 525446
rect 187365 525396 187431 525412
rect 187257 525356 187323 525372
rect 172289 525328 172407 525354
rect 172565 525328 173511 525354
rect 173669 525328 174615 525354
rect 174773 525328 175719 525354
rect 175877 525328 176823 525354
rect 176981 525328 177191 525354
rect 177533 525328 178479 525354
rect 178637 525328 179583 525354
rect 179741 525328 180687 525354
rect 180845 525328 181791 525354
rect 181949 525328 182343 525354
rect 182685 525328 183631 525354
rect 183789 525328 184735 525354
rect 184893 525328 185839 525354
rect 185997 525328 186943 525354
rect 187285 525354 187323 525356
rect 187285 525328 187403 525354
rect 172289 525192 172407 525218
rect 172565 525192 173511 525218
rect 173669 525192 174615 525218
rect 174773 525192 175719 525218
rect 175877 525192 176823 525218
rect 176981 525192 177191 525218
rect 177533 525192 178479 525218
rect 178637 525192 179583 525218
rect 179741 525192 180687 525218
rect 180845 525192 181791 525218
rect 181949 525192 182343 525218
rect 182685 525192 183631 525218
rect 183789 525192 184735 525218
rect 184893 525192 185839 525218
rect 185997 525192 186943 525218
rect 187285 525192 187403 525218
rect 172289 525124 172407 525150
rect 172565 525124 173511 525150
rect 173669 525124 174615 525150
rect 174957 525124 175903 525150
rect 176061 525124 177007 525150
rect 177165 525124 178111 525150
rect 178269 525124 179215 525150
rect 179373 525124 179767 525150
rect 180109 525124 181055 525150
rect 181213 525124 182159 525150
rect 182317 525124 183263 525150
rect 183421 525124 184367 525150
rect 184525 525124 184919 525150
rect 185261 525124 186207 525150
rect 186365 525124 186943 525150
rect 187285 525124 187403 525150
rect 172289 524988 172407 525014
rect 172565 524988 173511 525014
rect 173669 524988 174615 525014
rect 174957 524988 175903 525014
rect 176061 524988 177007 525014
rect 177165 524988 178111 525014
rect 178269 524988 179215 525014
rect 179373 524988 179767 525014
rect 180109 524988 181055 525014
rect 181213 524988 182159 525014
rect 182317 524988 183263 525014
rect 183421 524988 184367 525014
rect 184525 524988 184919 525014
rect 185261 524988 186207 525014
rect 186365 524988 186943 525014
rect 172369 524986 172407 524988
rect 172369 524970 172435 524986
rect 172261 524930 172327 524946
rect 172261 524896 172277 524930
rect 172311 524896 172327 524930
rect 172369 524936 172385 524970
rect 172419 524936 172435 524970
rect 173057 524966 173511 524988
rect 172369 524920 172435 524936
rect 172565 524930 173015 524946
rect 172261 524880 172327 524896
rect 172289 524878 172327 524880
rect 172565 524896 172837 524930
rect 172871 524896 173015 524930
rect 173057 524932 173201 524966
rect 173235 524932 173511 524966
rect 174161 524966 174615 524988
rect 173057 524916 173511 524932
rect 173669 524930 174119 524946
rect 172289 524848 172407 524878
rect 172565 524874 173015 524896
rect 173669 524896 173941 524930
rect 173975 524896 174119 524930
rect 174161 524932 174305 524966
rect 174339 524932 174615 524966
rect 175449 524966 175903 524988
rect 174161 524916 174615 524932
rect 174957 524930 175407 524946
rect 173669 524874 174119 524896
rect 174957 524896 175229 524930
rect 175263 524896 175407 524930
rect 175449 524932 175593 524966
rect 175627 524932 175903 524966
rect 176553 524966 177007 524988
rect 175449 524916 175903 524932
rect 176061 524930 176511 524946
rect 174957 524874 175407 524896
rect 176061 524896 176333 524930
rect 176367 524896 176511 524930
rect 176553 524932 176697 524966
rect 176731 524932 177007 524966
rect 177657 524966 178111 524988
rect 176553 524916 177007 524932
rect 177165 524930 177615 524946
rect 176061 524874 176511 524896
rect 177165 524896 177437 524930
rect 177471 524896 177615 524930
rect 177657 524932 177801 524966
rect 177835 524932 178111 524966
rect 178761 524966 179215 524988
rect 177657 524916 178111 524932
rect 178269 524930 178719 524946
rect 177165 524874 177615 524896
rect 178269 524896 178541 524930
rect 178575 524896 178719 524930
rect 178761 524932 178905 524966
rect 178939 524932 179215 524966
rect 179591 524966 179767 524988
rect 178761 524916 179215 524932
rect 179373 524930 179549 524946
rect 178269 524874 178719 524896
rect 179373 524896 179389 524930
rect 179423 524896 179499 524930
rect 179533 524896 179549 524930
rect 179591 524932 179607 524966
rect 179641 524932 179717 524966
rect 179751 524932 179767 524966
rect 180601 524966 181055 524988
rect 179591 524916 179767 524932
rect 180109 524930 180559 524946
rect 179373 524874 179549 524896
rect 180109 524896 180381 524930
rect 180415 524896 180559 524930
rect 180601 524932 180745 524966
rect 180779 524932 181055 524966
rect 181705 524966 182159 524988
rect 180601 524916 181055 524932
rect 181213 524930 181663 524946
rect 180109 524874 180559 524896
rect 181213 524896 181485 524930
rect 181519 524896 181663 524930
rect 181705 524932 181849 524966
rect 181883 524932 182159 524966
rect 182809 524966 183263 524988
rect 181705 524916 182159 524932
rect 182317 524930 182767 524946
rect 181213 524874 181663 524896
rect 182317 524896 182589 524930
rect 182623 524896 182767 524930
rect 182809 524932 182953 524966
rect 182987 524932 183263 524966
rect 183913 524966 184367 524988
rect 182809 524916 183263 524932
rect 183421 524930 183871 524946
rect 182317 524874 182767 524896
rect 183421 524896 183693 524930
rect 183727 524896 183871 524930
rect 183913 524932 184057 524966
rect 184091 524932 184367 524966
rect 184743 524966 184919 524988
rect 183913 524916 184367 524932
rect 184525 524930 184701 524946
rect 183421 524874 183871 524896
rect 184525 524896 184541 524930
rect 184575 524896 184651 524930
rect 184685 524896 184701 524930
rect 184743 524932 184759 524966
rect 184793 524932 184869 524966
rect 184903 524932 184919 524966
rect 185753 524966 186207 524988
rect 184743 524916 184919 524932
rect 185261 524930 185711 524946
rect 184525 524874 184701 524896
rect 185261 524896 185533 524930
rect 185567 524896 185711 524930
rect 185753 524932 185897 524966
rect 185931 524932 186207 524966
rect 186671 524966 186943 524988
rect 187285 524988 187403 525014
rect 187285 524986 187323 524988
rect 185753 524916 186207 524932
rect 186365 524930 186629 524946
rect 185261 524874 185711 524896
rect 186365 524896 186381 524930
rect 186415 524896 186480 524930
rect 186514 524896 186579 524930
rect 186613 524896 186629 524930
rect 186671 524932 186687 524966
rect 186721 524932 186790 524966
rect 186824 524932 186893 524966
rect 186927 524932 186943 524966
rect 186671 524916 186943 524932
rect 187257 524970 187323 524986
rect 187257 524936 187273 524970
rect 187307 524936 187323 524970
rect 187257 524920 187323 524936
rect 187365 524930 187431 524946
rect 186365 524874 186629 524896
rect 187365 524896 187381 524930
rect 187415 524896 187431 524930
rect 187365 524880 187431 524896
rect 187365 524878 187403 524880
rect 172565 524848 173511 524874
rect 173669 524848 174615 524874
rect 174957 524848 175903 524874
rect 176061 524848 177007 524874
rect 177165 524848 178111 524874
rect 178269 524848 179215 524874
rect 179373 524848 179767 524874
rect 180109 524848 181055 524874
rect 181213 524848 182159 524874
rect 182317 524848 183263 524874
rect 183421 524848 184367 524874
rect 184525 524848 184919 524874
rect 185261 524848 186207 524874
rect 186365 524848 186943 524874
rect 187285 524848 187403 524878
rect 172289 524648 172407 524674
rect 172565 524648 173511 524674
rect 173669 524648 174615 524674
rect 174957 524648 175903 524674
rect 176061 524648 177007 524674
rect 177165 524648 178111 524674
rect 178269 524648 179215 524674
rect 179373 524648 179767 524674
rect 180109 524648 181055 524674
rect 181213 524648 182159 524674
rect 182317 524648 183263 524674
rect 183421 524648 184367 524674
rect 184525 524648 184919 524674
rect 185261 524648 186207 524674
rect 186365 524648 186943 524674
rect 187285 524648 187403 524674
rect 172289 524580 172407 524606
rect 172565 524580 173511 524606
rect 173669 524580 174615 524606
rect 174773 524580 175719 524606
rect 175877 524580 176823 524606
rect 176981 524580 177191 524606
rect 177533 524580 178479 524606
rect 178637 524580 179583 524606
rect 179741 524580 180687 524606
rect 180845 524580 181791 524606
rect 181949 524580 182343 524606
rect 182685 524580 183631 524606
rect 183789 524580 184735 524606
rect 184893 524580 185839 524606
rect 185997 524580 186943 524606
rect 187285 524580 187403 524606
rect 172289 524376 172407 524406
rect 172565 524380 173511 524406
rect 173669 524380 174615 524406
rect 174773 524380 175719 524406
rect 175877 524380 176823 524406
rect 176981 524380 177191 524406
rect 177533 524380 178479 524406
rect 178637 524380 179583 524406
rect 179741 524380 180687 524406
rect 180845 524380 181791 524406
rect 181949 524380 182343 524406
rect 182685 524380 183631 524406
rect 183789 524380 184735 524406
rect 184893 524380 185839 524406
rect 185997 524380 186943 524406
rect 172289 524374 172327 524376
rect 172261 524358 172327 524374
rect 172261 524324 172277 524358
rect 172311 524324 172327 524358
rect 172565 524358 173015 524380
rect 172261 524308 172327 524324
rect 172369 524318 172435 524334
rect 172369 524284 172385 524318
rect 172419 524284 172435 524318
rect 172565 524324 172837 524358
rect 172871 524324 173015 524358
rect 173669 524358 174119 524380
rect 172565 524308 173015 524324
rect 173057 524322 173511 524338
rect 172369 524268 172435 524284
rect 173057 524288 173201 524322
rect 173235 524288 173511 524322
rect 173669 524324 173941 524358
rect 173975 524324 174119 524358
rect 174773 524358 175223 524380
rect 173669 524308 174119 524324
rect 174161 524322 174615 524338
rect 172369 524266 172407 524268
rect 173057 524266 173511 524288
rect 174161 524288 174305 524322
rect 174339 524288 174615 524322
rect 174773 524324 175045 524358
rect 175079 524324 175223 524358
rect 175877 524358 176327 524380
rect 176981 524374 177065 524380
rect 174773 524308 175223 524324
rect 175265 524322 175719 524338
rect 174161 524266 174615 524288
rect 175265 524288 175409 524322
rect 175443 524288 175719 524322
rect 175877 524324 176149 524358
rect 176183 524324 176327 524358
rect 176923 524358 177065 524374
rect 175877 524308 176327 524324
rect 176369 524322 176823 524338
rect 175265 524266 175719 524288
rect 176369 524288 176513 524322
rect 176547 524288 176823 524322
rect 176923 524324 176939 524358
rect 176973 524324 177065 524358
rect 177533 524358 177983 524380
rect 176923 524308 177065 524324
rect 177107 524322 177249 524338
rect 176369 524266 176823 524288
rect 177107 524288 177199 524322
rect 177233 524288 177249 524322
rect 177533 524324 177805 524358
rect 177839 524324 177983 524358
rect 178637 524358 179087 524380
rect 177533 524308 177983 524324
rect 178025 524322 178479 524338
rect 177107 524272 177249 524288
rect 178025 524288 178169 524322
rect 178203 524288 178479 524322
rect 178637 524324 178909 524358
rect 178943 524324 179087 524358
rect 179741 524358 180191 524380
rect 178637 524308 179087 524324
rect 179129 524322 179583 524338
rect 177107 524266 177191 524272
rect 178025 524266 178479 524288
rect 179129 524288 179273 524322
rect 179307 524288 179583 524322
rect 179741 524324 180013 524358
rect 180047 524324 180191 524358
rect 180845 524358 181295 524380
rect 179741 524308 180191 524324
rect 180233 524322 180687 524338
rect 179129 524266 179583 524288
rect 180233 524288 180377 524322
rect 180411 524288 180687 524322
rect 180845 524324 181117 524358
rect 181151 524324 181295 524358
rect 181949 524358 182125 524380
rect 180845 524308 181295 524324
rect 181337 524322 181791 524338
rect 180233 524266 180687 524288
rect 181337 524288 181481 524322
rect 181515 524288 181791 524322
rect 181949 524324 181965 524358
rect 181999 524324 182075 524358
rect 182109 524324 182125 524358
rect 182685 524358 183135 524380
rect 181949 524308 182125 524324
rect 182167 524322 182343 524338
rect 181337 524266 181791 524288
rect 182167 524288 182183 524322
rect 182217 524288 182293 524322
rect 182327 524288 182343 524322
rect 182685 524324 182957 524358
rect 182991 524324 183135 524358
rect 183789 524358 184239 524380
rect 182685 524308 183135 524324
rect 183177 524322 183631 524338
rect 182167 524266 182343 524288
rect 183177 524288 183321 524322
rect 183355 524288 183631 524322
rect 183789 524324 184061 524358
rect 184095 524324 184239 524358
rect 184893 524358 185343 524380
rect 183789 524308 184239 524324
rect 184281 524322 184735 524338
rect 183177 524266 183631 524288
rect 184281 524288 184425 524322
rect 184459 524288 184735 524322
rect 184893 524324 185165 524358
rect 185199 524324 185343 524358
rect 185997 524358 186447 524380
rect 187285 524376 187403 524406
rect 184893 524308 185343 524324
rect 185385 524322 185839 524338
rect 184281 524266 184735 524288
rect 185385 524288 185529 524322
rect 185563 524288 185839 524322
rect 185997 524324 186269 524358
rect 186303 524324 186447 524358
rect 187365 524374 187403 524376
rect 187365 524358 187431 524374
rect 185997 524308 186447 524324
rect 186489 524322 186943 524338
rect 185385 524266 185839 524288
rect 186489 524288 186633 524322
rect 186667 524288 186943 524322
rect 186489 524266 186943 524288
rect 187257 524318 187323 524334
rect 187257 524284 187273 524318
rect 187307 524284 187323 524318
rect 187365 524324 187381 524358
rect 187415 524324 187431 524358
rect 187365 524308 187431 524324
rect 187257 524268 187323 524284
rect 172289 524240 172407 524266
rect 172565 524240 173511 524266
rect 173669 524240 174615 524266
rect 174773 524240 175719 524266
rect 175877 524240 176823 524266
rect 176981 524240 177191 524266
rect 177533 524240 178479 524266
rect 178637 524240 179583 524266
rect 179741 524240 180687 524266
rect 180845 524240 181791 524266
rect 181949 524240 182343 524266
rect 182685 524240 183631 524266
rect 183789 524240 184735 524266
rect 184893 524240 185839 524266
rect 185997 524240 186943 524266
rect 187285 524266 187323 524268
rect 187285 524240 187403 524266
rect 172289 524104 172407 524130
rect 172565 524104 173511 524130
rect 173669 524104 174615 524130
rect 174773 524104 175719 524130
rect 175877 524104 176823 524130
rect 176981 524104 177191 524130
rect 177533 524104 178479 524130
rect 178637 524104 179583 524130
rect 179741 524104 180687 524130
rect 180845 524104 181791 524130
rect 181949 524104 182343 524130
rect 182685 524104 183631 524130
rect 183789 524104 184735 524130
rect 184893 524104 185839 524130
rect 185997 524104 186943 524130
rect 187285 524104 187403 524130
rect 172289 524036 172407 524062
rect 172565 524036 173511 524062
rect 173669 524036 174615 524062
rect 174957 524036 175903 524062
rect 176061 524036 177007 524062
rect 177165 524036 178111 524062
rect 178269 524036 179215 524062
rect 179373 524036 179767 524062
rect 180109 524036 181055 524062
rect 181213 524036 182159 524062
rect 182317 524036 183263 524062
rect 183421 524036 184367 524062
rect 184525 524036 184919 524062
rect 185261 524036 186207 524062
rect 186365 524036 186943 524062
rect 187285 524036 187403 524062
rect 172289 523900 172407 523926
rect 172565 523900 173511 523926
rect 173669 523900 174615 523926
rect 174957 523900 175903 523926
rect 176061 523900 177007 523926
rect 177165 523900 178111 523926
rect 178269 523900 179215 523926
rect 179373 523900 179767 523926
rect 180109 523900 181055 523926
rect 181213 523900 182159 523926
rect 182317 523900 183263 523926
rect 183421 523900 184367 523926
rect 184525 523900 184919 523926
rect 185261 523900 186207 523926
rect 186365 523900 186943 523926
rect 172369 523898 172407 523900
rect 172369 523882 172435 523898
rect 172261 523842 172327 523858
rect 172261 523808 172277 523842
rect 172311 523808 172327 523842
rect 172369 523848 172385 523882
rect 172419 523848 172435 523882
rect 173057 523878 173511 523900
rect 172369 523832 172435 523848
rect 172565 523842 173015 523858
rect 172261 523792 172327 523808
rect 172289 523790 172327 523792
rect 172565 523808 172837 523842
rect 172871 523808 173015 523842
rect 173057 523844 173201 523878
rect 173235 523844 173511 523878
rect 174161 523878 174615 523900
rect 173057 523828 173511 523844
rect 173669 523842 174119 523858
rect 172289 523760 172407 523790
rect 172565 523786 173015 523808
rect 173669 523808 173941 523842
rect 173975 523808 174119 523842
rect 174161 523844 174305 523878
rect 174339 523844 174615 523878
rect 175449 523878 175903 523900
rect 174161 523828 174615 523844
rect 174957 523842 175407 523858
rect 173669 523786 174119 523808
rect 174957 523808 175229 523842
rect 175263 523808 175407 523842
rect 175449 523844 175593 523878
rect 175627 523844 175903 523878
rect 176553 523878 177007 523900
rect 175449 523828 175903 523844
rect 176061 523842 176511 523858
rect 174957 523786 175407 523808
rect 176061 523808 176333 523842
rect 176367 523808 176511 523842
rect 176553 523844 176697 523878
rect 176731 523844 177007 523878
rect 177657 523878 178111 523900
rect 176553 523828 177007 523844
rect 177165 523842 177615 523858
rect 176061 523786 176511 523808
rect 177165 523808 177437 523842
rect 177471 523808 177615 523842
rect 177657 523844 177801 523878
rect 177835 523844 178111 523878
rect 178761 523878 179215 523900
rect 177657 523828 178111 523844
rect 178269 523842 178719 523858
rect 177165 523786 177615 523808
rect 178269 523808 178541 523842
rect 178575 523808 178719 523842
rect 178761 523844 178905 523878
rect 178939 523844 179215 523878
rect 179591 523878 179767 523900
rect 178761 523828 179215 523844
rect 179373 523842 179549 523858
rect 178269 523786 178719 523808
rect 179373 523808 179389 523842
rect 179423 523808 179499 523842
rect 179533 523808 179549 523842
rect 179591 523844 179607 523878
rect 179641 523844 179717 523878
rect 179751 523844 179767 523878
rect 180601 523878 181055 523900
rect 179591 523828 179767 523844
rect 180109 523842 180559 523858
rect 179373 523786 179549 523808
rect 180109 523808 180381 523842
rect 180415 523808 180559 523842
rect 180601 523844 180745 523878
rect 180779 523844 181055 523878
rect 181705 523878 182159 523900
rect 180601 523828 181055 523844
rect 181213 523842 181663 523858
rect 180109 523786 180559 523808
rect 181213 523808 181485 523842
rect 181519 523808 181663 523842
rect 181705 523844 181849 523878
rect 181883 523844 182159 523878
rect 182809 523878 183263 523900
rect 181705 523828 182159 523844
rect 182317 523842 182767 523858
rect 181213 523786 181663 523808
rect 182317 523808 182589 523842
rect 182623 523808 182767 523842
rect 182809 523844 182953 523878
rect 182987 523844 183263 523878
rect 183913 523878 184367 523900
rect 182809 523828 183263 523844
rect 183421 523842 183871 523858
rect 182317 523786 182767 523808
rect 183421 523808 183693 523842
rect 183727 523808 183871 523842
rect 183913 523844 184057 523878
rect 184091 523844 184367 523878
rect 184743 523878 184919 523900
rect 183913 523828 184367 523844
rect 184525 523842 184701 523858
rect 183421 523786 183871 523808
rect 184525 523808 184541 523842
rect 184575 523808 184651 523842
rect 184685 523808 184701 523842
rect 184743 523844 184759 523878
rect 184793 523844 184869 523878
rect 184903 523844 184919 523878
rect 185753 523878 186207 523900
rect 184743 523828 184919 523844
rect 185261 523842 185711 523858
rect 184525 523786 184701 523808
rect 185261 523808 185533 523842
rect 185567 523808 185711 523842
rect 185753 523844 185897 523878
rect 185931 523844 186207 523878
rect 186671 523878 186943 523900
rect 187285 523900 187403 523926
rect 187285 523898 187323 523900
rect 185753 523828 186207 523844
rect 186365 523842 186629 523858
rect 185261 523786 185711 523808
rect 186365 523808 186381 523842
rect 186415 523808 186480 523842
rect 186514 523808 186579 523842
rect 186613 523808 186629 523842
rect 186671 523844 186687 523878
rect 186721 523844 186790 523878
rect 186824 523844 186893 523878
rect 186927 523844 186943 523878
rect 186671 523828 186943 523844
rect 187257 523882 187323 523898
rect 187257 523848 187273 523882
rect 187307 523848 187323 523882
rect 187257 523832 187323 523848
rect 187365 523842 187431 523858
rect 186365 523786 186629 523808
rect 187365 523808 187381 523842
rect 187415 523808 187431 523842
rect 187365 523792 187431 523808
rect 187365 523790 187403 523792
rect 172565 523760 173511 523786
rect 173669 523760 174615 523786
rect 174957 523760 175903 523786
rect 176061 523760 177007 523786
rect 177165 523760 178111 523786
rect 178269 523760 179215 523786
rect 179373 523760 179767 523786
rect 180109 523760 181055 523786
rect 181213 523760 182159 523786
rect 182317 523760 183263 523786
rect 183421 523760 184367 523786
rect 184525 523760 184919 523786
rect 185261 523760 186207 523786
rect 186365 523760 186943 523786
rect 187285 523760 187403 523790
rect 172289 523560 172407 523586
rect 172565 523560 173511 523586
rect 173669 523560 174615 523586
rect 174957 523560 175903 523586
rect 176061 523560 177007 523586
rect 177165 523560 178111 523586
rect 178269 523560 179215 523586
rect 179373 523560 179767 523586
rect 180109 523560 181055 523586
rect 181213 523560 182159 523586
rect 182317 523560 183263 523586
rect 183421 523560 184367 523586
rect 184525 523560 184919 523586
rect 185261 523560 186207 523586
rect 186365 523560 186943 523586
rect 187285 523560 187403 523586
rect 172289 523492 172407 523518
rect 172565 523492 173511 523518
rect 173669 523492 174615 523518
rect 174773 523492 175719 523518
rect 175877 523492 176823 523518
rect 176981 523492 177191 523518
rect 177533 523492 178479 523518
rect 178637 523492 179583 523518
rect 179741 523492 180687 523518
rect 180845 523492 181791 523518
rect 181949 523492 182343 523518
rect 182685 523492 183631 523518
rect 183789 523492 184735 523518
rect 184893 523492 185839 523518
rect 185997 523492 186943 523518
rect 187285 523492 187403 523518
rect 172289 523288 172407 523318
rect 172565 523292 173511 523318
rect 173669 523292 174615 523318
rect 174773 523292 175719 523318
rect 175877 523292 176823 523318
rect 176981 523292 177191 523318
rect 177533 523292 178479 523318
rect 178637 523292 179583 523318
rect 179741 523292 180687 523318
rect 180845 523292 181791 523318
rect 181949 523292 182343 523318
rect 182685 523292 183631 523318
rect 183789 523292 184735 523318
rect 184893 523292 185839 523318
rect 185997 523292 186943 523318
rect 172289 523286 172327 523288
rect 172261 523270 172327 523286
rect 172261 523236 172277 523270
rect 172311 523236 172327 523270
rect 172565 523270 173015 523292
rect 172261 523220 172327 523236
rect 172369 523230 172435 523246
rect 172369 523196 172385 523230
rect 172419 523196 172435 523230
rect 172565 523236 172837 523270
rect 172871 523236 173015 523270
rect 173669 523270 174119 523292
rect 172565 523220 173015 523236
rect 173057 523234 173511 523250
rect 172369 523180 172435 523196
rect 173057 523200 173201 523234
rect 173235 523200 173511 523234
rect 173669 523236 173941 523270
rect 173975 523236 174119 523270
rect 174773 523270 175223 523292
rect 173669 523220 174119 523236
rect 174161 523234 174615 523250
rect 172369 523178 172407 523180
rect 173057 523178 173511 523200
rect 174161 523200 174305 523234
rect 174339 523200 174615 523234
rect 174773 523236 175045 523270
rect 175079 523236 175223 523270
rect 175877 523270 176327 523292
rect 176981 523286 177065 523292
rect 174773 523220 175223 523236
rect 175265 523234 175719 523250
rect 174161 523178 174615 523200
rect 175265 523200 175409 523234
rect 175443 523200 175719 523234
rect 175877 523236 176149 523270
rect 176183 523236 176327 523270
rect 176923 523270 177065 523286
rect 175877 523220 176327 523236
rect 176369 523234 176823 523250
rect 175265 523178 175719 523200
rect 176369 523200 176513 523234
rect 176547 523200 176823 523234
rect 176923 523236 176939 523270
rect 176973 523236 177065 523270
rect 177533 523270 177983 523292
rect 176923 523220 177065 523236
rect 177107 523234 177249 523250
rect 176369 523178 176823 523200
rect 177107 523200 177199 523234
rect 177233 523200 177249 523234
rect 177533 523236 177805 523270
rect 177839 523236 177983 523270
rect 178637 523270 179087 523292
rect 177533 523220 177983 523236
rect 178025 523234 178479 523250
rect 177107 523184 177249 523200
rect 178025 523200 178169 523234
rect 178203 523200 178479 523234
rect 178637 523236 178909 523270
rect 178943 523236 179087 523270
rect 179741 523270 180191 523292
rect 178637 523220 179087 523236
rect 179129 523234 179583 523250
rect 177107 523178 177191 523184
rect 178025 523178 178479 523200
rect 179129 523200 179273 523234
rect 179307 523200 179583 523234
rect 179741 523236 180013 523270
rect 180047 523236 180191 523270
rect 180845 523270 181295 523292
rect 179741 523220 180191 523236
rect 180233 523234 180687 523250
rect 179129 523178 179583 523200
rect 180233 523200 180377 523234
rect 180411 523200 180687 523234
rect 180845 523236 181117 523270
rect 181151 523236 181295 523270
rect 181949 523270 182125 523292
rect 180845 523220 181295 523236
rect 181337 523234 181791 523250
rect 180233 523178 180687 523200
rect 181337 523200 181481 523234
rect 181515 523200 181791 523234
rect 181949 523236 181965 523270
rect 181999 523236 182075 523270
rect 182109 523236 182125 523270
rect 182685 523270 183135 523292
rect 181949 523220 182125 523236
rect 182167 523234 182343 523250
rect 181337 523178 181791 523200
rect 182167 523200 182183 523234
rect 182217 523200 182293 523234
rect 182327 523200 182343 523234
rect 182685 523236 182957 523270
rect 182991 523236 183135 523270
rect 183789 523270 184239 523292
rect 182685 523220 183135 523236
rect 183177 523234 183631 523250
rect 182167 523178 182343 523200
rect 183177 523200 183321 523234
rect 183355 523200 183631 523234
rect 183789 523236 184061 523270
rect 184095 523236 184239 523270
rect 184893 523270 185343 523292
rect 183789 523220 184239 523236
rect 184281 523234 184735 523250
rect 183177 523178 183631 523200
rect 184281 523200 184425 523234
rect 184459 523200 184735 523234
rect 184893 523236 185165 523270
rect 185199 523236 185343 523270
rect 185997 523270 186447 523292
rect 187285 523288 187403 523318
rect 184893 523220 185343 523236
rect 185385 523234 185839 523250
rect 184281 523178 184735 523200
rect 185385 523200 185529 523234
rect 185563 523200 185839 523234
rect 185997 523236 186269 523270
rect 186303 523236 186447 523270
rect 187365 523286 187403 523288
rect 187365 523270 187431 523286
rect 185997 523220 186447 523236
rect 186489 523234 186943 523250
rect 185385 523178 185839 523200
rect 186489 523200 186633 523234
rect 186667 523200 186943 523234
rect 186489 523178 186943 523200
rect 187257 523230 187323 523246
rect 187257 523196 187273 523230
rect 187307 523196 187323 523230
rect 187365 523236 187381 523270
rect 187415 523236 187431 523270
rect 187365 523220 187431 523236
rect 187257 523180 187323 523196
rect 172289 523152 172407 523178
rect 172565 523152 173511 523178
rect 173669 523152 174615 523178
rect 174773 523152 175719 523178
rect 175877 523152 176823 523178
rect 176981 523152 177191 523178
rect 177533 523152 178479 523178
rect 178637 523152 179583 523178
rect 179741 523152 180687 523178
rect 180845 523152 181791 523178
rect 181949 523152 182343 523178
rect 182685 523152 183631 523178
rect 183789 523152 184735 523178
rect 184893 523152 185839 523178
rect 185997 523152 186943 523178
rect 187285 523178 187323 523180
rect 187285 523152 187403 523178
rect 172289 523016 172407 523042
rect 172565 523016 173511 523042
rect 173669 523016 174615 523042
rect 174773 523016 175719 523042
rect 175877 523016 176823 523042
rect 176981 523016 177191 523042
rect 177533 523016 178479 523042
rect 178637 523016 179583 523042
rect 179741 523016 180687 523042
rect 180845 523016 181791 523042
rect 181949 523016 182343 523042
rect 182685 523016 183631 523042
rect 183789 523016 184735 523042
rect 184893 523016 185839 523042
rect 185997 523016 186943 523042
rect 187285 523016 187403 523042
rect 172289 522948 172407 522974
rect 172565 522948 173511 522974
rect 173669 522948 174615 522974
rect 174957 522948 175903 522974
rect 176061 522948 177007 522974
rect 177165 522948 178111 522974
rect 178269 522948 179215 522974
rect 179373 522948 179767 522974
rect 180109 522948 181055 522974
rect 181213 522948 182159 522974
rect 182317 522948 183263 522974
rect 183421 522948 184367 522974
rect 184525 522948 184919 522974
rect 185261 522948 186207 522974
rect 186365 522948 186943 522974
rect 187285 522948 187403 522974
rect 172289 522812 172407 522838
rect 172565 522812 173511 522838
rect 173669 522812 174615 522838
rect 174957 522812 175903 522838
rect 176061 522812 177007 522838
rect 177165 522812 178111 522838
rect 178269 522812 179215 522838
rect 179373 522812 179767 522838
rect 180109 522812 181055 522838
rect 181213 522812 182159 522838
rect 182317 522812 183263 522838
rect 183421 522812 184367 522838
rect 184525 522812 184919 522838
rect 185261 522812 186207 522838
rect 186365 522812 186943 522838
rect 172369 522810 172407 522812
rect 172369 522794 172435 522810
rect 172261 522754 172327 522770
rect 172261 522720 172277 522754
rect 172311 522720 172327 522754
rect 172369 522760 172385 522794
rect 172419 522760 172435 522794
rect 173057 522790 173511 522812
rect 172369 522744 172435 522760
rect 172565 522754 173015 522770
rect 172261 522704 172327 522720
rect 172289 522702 172327 522704
rect 172565 522720 172837 522754
rect 172871 522720 173015 522754
rect 173057 522756 173201 522790
rect 173235 522756 173511 522790
rect 174161 522790 174615 522812
rect 173057 522740 173511 522756
rect 173669 522754 174119 522770
rect 172289 522672 172407 522702
rect 172565 522698 173015 522720
rect 173669 522720 173941 522754
rect 173975 522720 174119 522754
rect 174161 522756 174305 522790
rect 174339 522756 174615 522790
rect 175449 522790 175903 522812
rect 174161 522740 174615 522756
rect 174957 522754 175407 522770
rect 173669 522698 174119 522720
rect 174957 522720 175229 522754
rect 175263 522720 175407 522754
rect 175449 522756 175593 522790
rect 175627 522756 175903 522790
rect 176553 522790 177007 522812
rect 175449 522740 175903 522756
rect 176061 522754 176511 522770
rect 174957 522698 175407 522720
rect 176061 522720 176333 522754
rect 176367 522720 176511 522754
rect 176553 522756 176697 522790
rect 176731 522756 177007 522790
rect 177657 522790 178111 522812
rect 176553 522740 177007 522756
rect 177165 522754 177615 522770
rect 176061 522698 176511 522720
rect 177165 522720 177437 522754
rect 177471 522720 177615 522754
rect 177657 522756 177801 522790
rect 177835 522756 178111 522790
rect 178761 522790 179215 522812
rect 177657 522740 178111 522756
rect 178269 522754 178719 522770
rect 177165 522698 177615 522720
rect 178269 522720 178541 522754
rect 178575 522720 178719 522754
rect 178761 522756 178905 522790
rect 178939 522756 179215 522790
rect 179591 522790 179767 522812
rect 178761 522740 179215 522756
rect 179373 522754 179549 522770
rect 178269 522698 178719 522720
rect 179373 522720 179389 522754
rect 179423 522720 179499 522754
rect 179533 522720 179549 522754
rect 179591 522756 179607 522790
rect 179641 522756 179717 522790
rect 179751 522756 179767 522790
rect 180601 522790 181055 522812
rect 179591 522740 179767 522756
rect 180109 522754 180559 522770
rect 179373 522698 179549 522720
rect 180109 522720 180381 522754
rect 180415 522720 180559 522754
rect 180601 522756 180745 522790
rect 180779 522756 181055 522790
rect 181705 522790 182159 522812
rect 180601 522740 181055 522756
rect 181213 522754 181663 522770
rect 180109 522698 180559 522720
rect 181213 522720 181485 522754
rect 181519 522720 181663 522754
rect 181705 522756 181849 522790
rect 181883 522756 182159 522790
rect 182809 522790 183263 522812
rect 181705 522740 182159 522756
rect 182317 522754 182767 522770
rect 181213 522698 181663 522720
rect 182317 522720 182589 522754
rect 182623 522720 182767 522754
rect 182809 522756 182953 522790
rect 182987 522756 183263 522790
rect 183913 522790 184367 522812
rect 182809 522740 183263 522756
rect 183421 522754 183871 522770
rect 182317 522698 182767 522720
rect 183421 522720 183693 522754
rect 183727 522720 183871 522754
rect 183913 522756 184057 522790
rect 184091 522756 184367 522790
rect 184743 522790 184919 522812
rect 183913 522740 184367 522756
rect 184525 522754 184701 522770
rect 183421 522698 183871 522720
rect 184525 522720 184541 522754
rect 184575 522720 184651 522754
rect 184685 522720 184701 522754
rect 184743 522756 184759 522790
rect 184793 522756 184869 522790
rect 184903 522756 184919 522790
rect 185753 522790 186207 522812
rect 184743 522740 184919 522756
rect 185261 522754 185711 522770
rect 184525 522698 184701 522720
rect 185261 522720 185533 522754
rect 185567 522720 185711 522754
rect 185753 522756 185897 522790
rect 185931 522756 186207 522790
rect 186671 522790 186943 522812
rect 187285 522812 187403 522838
rect 187285 522810 187323 522812
rect 185753 522740 186207 522756
rect 186365 522754 186629 522770
rect 185261 522698 185711 522720
rect 186365 522720 186381 522754
rect 186415 522720 186480 522754
rect 186514 522720 186579 522754
rect 186613 522720 186629 522754
rect 186671 522756 186687 522790
rect 186721 522756 186790 522790
rect 186824 522756 186893 522790
rect 186927 522756 186943 522790
rect 186671 522740 186943 522756
rect 187257 522794 187323 522810
rect 187257 522760 187273 522794
rect 187307 522760 187323 522794
rect 187257 522744 187323 522760
rect 187365 522754 187431 522770
rect 186365 522698 186629 522720
rect 187365 522720 187381 522754
rect 187415 522720 187431 522754
rect 187365 522704 187431 522720
rect 187365 522702 187403 522704
rect 172565 522672 173511 522698
rect 173669 522672 174615 522698
rect 174957 522672 175903 522698
rect 176061 522672 177007 522698
rect 177165 522672 178111 522698
rect 178269 522672 179215 522698
rect 179373 522672 179767 522698
rect 180109 522672 181055 522698
rect 181213 522672 182159 522698
rect 182317 522672 183263 522698
rect 183421 522672 184367 522698
rect 184525 522672 184919 522698
rect 185261 522672 186207 522698
rect 186365 522672 186943 522698
rect 187285 522672 187403 522702
rect 172289 522472 172407 522498
rect 172565 522472 173511 522498
rect 173669 522472 174615 522498
rect 174957 522472 175903 522498
rect 176061 522472 177007 522498
rect 177165 522472 178111 522498
rect 178269 522472 179215 522498
rect 179373 522472 179767 522498
rect 180109 522472 181055 522498
rect 181213 522472 182159 522498
rect 182317 522472 183263 522498
rect 183421 522472 184367 522498
rect 184525 522472 184919 522498
rect 185261 522472 186207 522498
rect 186365 522472 186943 522498
rect 187285 522472 187403 522498
rect 172289 522404 172407 522430
rect 172565 522404 173511 522430
rect 173669 522404 174615 522430
rect 174773 522404 175719 522430
rect 175877 522404 176823 522430
rect 176981 522404 177191 522430
rect 177533 522404 178479 522430
rect 178637 522404 179583 522430
rect 179741 522404 180687 522430
rect 180845 522404 181791 522430
rect 181949 522404 182343 522430
rect 182685 522404 183631 522430
rect 183789 522404 184735 522430
rect 184893 522404 185839 522430
rect 185997 522404 186943 522430
rect 187285 522404 187403 522430
rect 172289 522200 172407 522230
rect 172565 522204 173511 522230
rect 173669 522204 174615 522230
rect 174773 522204 175719 522230
rect 175877 522204 176823 522230
rect 176981 522204 177191 522230
rect 177533 522204 178479 522230
rect 178637 522204 179583 522230
rect 179741 522204 180687 522230
rect 180845 522204 181791 522230
rect 181949 522204 182343 522230
rect 182685 522204 183631 522230
rect 183789 522204 184735 522230
rect 184893 522204 185839 522230
rect 185997 522204 186943 522230
rect 172289 522198 172327 522200
rect 172261 522182 172327 522198
rect 172261 522148 172277 522182
rect 172311 522148 172327 522182
rect 172565 522182 173015 522204
rect 172261 522132 172327 522148
rect 172369 522142 172435 522158
rect 172369 522108 172385 522142
rect 172419 522108 172435 522142
rect 172565 522148 172837 522182
rect 172871 522148 173015 522182
rect 173669 522182 174119 522204
rect 172565 522132 173015 522148
rect 173057 522146 173511 522162
rect 172369 522092 172435 522108
rect 173057 522112 173201 522146
rect 173235 522112 173511 522146
rect 173669 522148 173941 522182
rect 173975 522148 174119 522182
rect 174773 522182 175223 522204
rect 173669 522132 174119 522148
rect 174161 522146 174615 522162
rect 172369 522090 172407 522092
rect 173057 522090 173511 522112
rect 174161 522112 174305 522146
rect 174339 522112 174615 522146
rect 174773 522148 175045 522182
rect 175079 522148 175223 522182
rect 175877 522182 176327 522204
rect 176981 522198 177065 522204
rect 174773 522132 175223 522148
rect 175265 522146 175719 522162
rect 174161 522090 174615 522112
rect 175265 522112 175409 522146
rect 175443 522112 175719 522146
rect 175877 522148 176149 522182
rect 176183 522148 176327 522182
rect 176923 522182 177065 522198
rect 175877 522132 176327 522148
rect 176369 522146 176823 522162
rect 175265 522090 175719 522112
rect 176369 522112 176513 522146
rect 176547 522112 176823 522146
rect 176923 522148 176939 522182
rect 176973 522148 177065 522182
rect 177533 522182 177983 522204
rect 176923 522132 177065 522148
rect 177107 522146 177249 522162
rect 176369 522090 176823 522112
rect 177107 522112 177199 522146
rect 177233 522112 177249 522146
rect 177533 522148 177805 522182
rect 177839 522148 177983 522182
rect 178637 522182 179087 522204
rect 177533 522132 177983 522148
rect 178025 522146 178479 522162
rect 177107 522096 177249 522112
rect 178025 522112 178169 522146
rect 178203 522112 178479 522146
rect 178637 522148 178909 522182
rect 178943 522148 179087 522182
rect 179741 522182 180191 522204
rect 178637 522132 179087 522148
rect 179129 522146 179583 522162
rect 177107 522090 177191 522096
rect 178025 522090 178479 522112
rect 179129 522112 179273 522146
rect 179307 522112 179583 522146
rect 179741 522148 180013 522182
rect 180047 522148 180191 522182
rect 180845 522182 181295 522204
rect 179741 522132 180191 522148
rect 180233 522146 180687 522162
rect 179129 522090 179583 522112
rect 180233 522112 180377 522146
rect 180411 522112 180687 522146
rect 180845 522148 181117 522182
rect 181151 522148 181295 522182
rect 181949 522182 182125 522204
rect 180845 522132 181295 522148
rect 181337 522146 181791 522162
rect 180233 522090 180687 522112
rect 181337 522112 181481 522146
rect 181515 522112 181791 522146
rect 181949 522148 181965 522182
rect 181999 522148 182075 522182
rect 182109 522148 182125 522182
rect 182685 522182 183135 522204
rect 181949 522132 182125 522148
rect 182167 522146 182343 522162
rect 181337 522090 181791 522112
rect 182167 522112 182183 522146
rect 182217 522112 182293 522146
rect 182327 522112 182343 522146
rect 182685 522148 182957 522182
rect 182991 522148 183135 522182
rect 183789 522182 184239 522204
rect 182685 522132 183135 522148
rect 183177 522146 183631 522162
rect 182167 522090 182343 522112
rect 183177 522112 183321 522146
rect 183355 522112 183631 522146
rect 183789 522148 184061 522182
rect 184095 522148 184239 522182
rect 184893 522182 185343 522204
rect 183789 522132 184239 522148
rect 184281 522146 184735 522162
rect 183177 522090 183631 522112
rect 184281 522112 184425 522146
rect 184459 522112 184735 522146
rect 184893 522148 185165 522182
rect 185199 522148 185343 522182
rect 185997 522182 186447 522204
rect 187285 522200 187403 522230
rect 184893 522132 185343 522148
rect 185385 522146 185839 522162
rect 184281 522090 184735 522112
rect 185385 522112 185529 522146
rect 185563 522112 185839 522146
rect 185997 522148 186269 522182
rect 186303 522148 186447 522182
rect 187365 522198 187403 522200
rect 187365 522182 187431 522198
rect 185997 522132 186447 522148
rect 186489 522146 186943 522162
rect 185385 522090 185839 522112
rect 186489 522112 186633 522146
rect 186667 522112 186943 522146
rect 186489 522090 186943 522112
rect 187257 522142 187323 522158
rect 187257 522108 187273 522142
rect 187307 522108 187323 522142
rect 187365 522148 187381 522182
rect 187415 522148 187431 522182
rect 187365 522132 187431 522148
rect 187257 522092 187323 522108
rect 172289 522064 172407 522090
rect 172565 522064 173511 522090
rect 173669 522064 174615 522090
rect 174773 522064 175719 522090
rect 175877 522064 176823 522090
rect 176981 522064 177191 522090
rect 177533 522064 178479 522090
rect 178637 522064 179583 522090
rect 179741 522064 180687 522090
rect 180845 522064 181791 522090
rect 181949 522064 182343 522090
rect 182685 522064 183631 522090
rect 183789 522064 184735 522090
rect 184893 522064 185839 522090
rect 185997 522064 186943 522090
rect 187285 522090 187323 522092
rect 187285 522064 187403 522090
rect 172289 521928 172407 521954
rect 172565 521928 173511 521954
rect 173669 521928 174615 521954
rect 174773 521928 175719 521954
rect 175877 521928 176823 521954
rect 176981 521928 177191 521954
rect 177533 521928 178479 521954
rect 178637 521928 179583 521954
rect 179741 521928 180687 521954
rect 180845 521928 181791 521954
rect 181949 521928 182343 521954
rect 182685 521928 183631 521954
rect 183789 521928 184735 521954
rect 184893 521928 185839 521954
rect 185997 521928 186943 521954
rect 187285 521928 187403 521954
rect 172289 521860 172407 521886
rect 172565 521860 173511 521886
rect 173669 521860 174615 521886
rect 174957 521860 175903 521886
rect 176061 521860 177007 521886
rect 177165 521860 178111 521886
rect 178269 521860 179215 521886
rect 179373 521860 179767 521886
rect 180109 521860 181055 521886
rect 181213 521860 182159 521886
rect 182317 521860 183263 521886
rect 183421 521860 184367 521886
rect 184525 521860 184919 521886
rect 185261 521860 186207 521886
rect 186365 521860 186943 521886
rect 187285 521860 187403 521886
rect 172289 521724 172407 521750
rect 172565 521724 173511 521750
rect 173669 521724 174615 521750
rect 174957 521724 175903 521750
rect 176061 521724 177007 521750
rect 177165 521724 178111 521750
rect 178269 521724 179215 521750
rect 179373 521724 179767 521750
rect 180109 521724 181055 521750
rect 181213 521724 182159 521750
rect 182317 521724 183263 521750
rect 183421 521724 184367 521750
rect 184525 521724 184919 521750
rect 185261 521724 186207 521750
rect 186365 521724 186943 521750
rect 172369 521722 172407 521724
rect 172369 521706 172435 521722
rect 172261 521666 172327 521682
rect 172261 521632 172277 521666
rect 172311 521632 172327 521666
rect 172369 521672 172385 521706
rect 172419 521672 172435 521706
rect 173057 521702 173511 521724
rect 172369 521656 172435 521672
rect 172565 521666 173015 521682
rect 172261 521616 172327 521632
rect 172289 521614 172327 521616
rect 172565 521632 172837 521666
rect 172871 521632 173015 521666
rect 173057 521668 173201 521702
rect 173235 521668 173511 521702
rect 174161 521702 174615 521724
rect 173057 521652 173511 521668
rect 173669 521666 174119 521682
rect 172289 521584 172407 521614
rect 172565 521610 173015 521632
rect 173669 521632 173941 521666
rect 173975 521632 174119 521666
rect 174161 521668 174305 521702
rect 174339 521668 174615 521702
rect 175449 521702 175903 521724
rect 174161 521652 174615 521668
rect 174957 521666 175407 521682
rect 173669 521610 174119 521632
rect 174957 521632 175229 521666
rect 175263 521632 175407 521666
rect 175449 521668 175593 521702
rect 175627 521668 175903 521702
rect 176553 521702 177007 521724
rect 175449 521652 175903 521668
rect 176061 521666 176511 521682
rect 174957 521610 175407 521632
rect 176061 521632 176333 521666
rect 176367 521632 176511 521666
rect 176553 521668 176697 521702
rect 176731 521668 177007 521702
rect 177657 521702 178111 521724
rect 176553 521652 177007 521668
rect 177165 521666 177615 521682
rect 176061 521610 176511 521632
rect 177165 521632 177437 521666
rect 177471 521632 177615 521666
rect 177657 521668 177801 521702
rect 177835 521668 178111 521702
rect 178761 521702 179215 521724
rect 177657 521652 178111 521668
rect 178269 521666 178719 521682
rect 177165 521610 177615 521632
rect 178269 521632 178541 521666
rect 178575 521632 178719 521666
rect 178761 521668 178905 521702
rect 178939 521668 179215 521702
rect 179591 521702 179767 521724
rect 178761 521652 179215 521668
rect 179373 521666 179549 521682
rect 178269 521610 178719 521632
rect 179373 521632 179389 521666
rect 179423 521632 179499 521666
rect 179533 521632 179549 521666
rect 179591 521668 179607 521702
rect 179641 521668 179717 521702
rect 179751 521668 179767 521702
rect 180601 521702 181055 521724
rect 179591 521652 179767 521668
rect 180109 521666 180559 521682
rect 179373 521610 179549 521632
rect 180109 521632 180381 521666
rect 180415 521632 180559 521666
rect 180601 521668 180745 521702
rect 180779 521668 181055 521702
rect 181705 521702 182159 521724
rect 180601 521652 181055 521668
rect 181213 521666 181663 521682
rect 180109 521610 180559 521632
rect 181213 521632 181485 521666
rect 181519 521632 181663 521666
rect 181705 521668 181849 521702
rect 181883 521668 182159 521702
rect 182809 521702 183263 521724
rect 181705 521652 182159 521668
rect 182317 521666 182767 521682
rect 181213 521610 181663 521632
rect 182317 521632 182589 521666
rect 182623 521632 182767 521666
rect 182809 521668 182953 521702
rect 182987 521668 183263 521702
rect 183913 521702 184367 521724
rect 182809 521652 183263 521668
rect 183421 521666 183871 521682
rect 182317 521610 182767 521632
rect 183421 521632 183693 521666
rect 183727 521632 183871 521666
rect 183913 521668 184057 521702
rect 184091 521668 184367 521702
rect 184743 521702 184919 521724
rect 183913 521652 184367 521668
rect 184525 521666 184701 521682
rect 183421 521610 183871 521632
rect 184525 521632 184541 521666
rect 184575 521632 184651 521666
rect 184685 521632 184701 521666
rect 184743 521668 184759 521702
rect 184793 521668 184869 521702
rect 184903 521668 184919 521702
rect 185753 521702 186207 521724
rect 184743 521652 184919 521668
rect 185261 521666 185711 521682
rect 184525 521610 184701 521632
rect 185261 521632 185533 521666
rect 185567 521632 185711 521666
rect 185753 521668 185897 521702
rect 185931 521668 186207 521702
rect 186671 521702 186943 521724
rect 187285 521724 187403 521750
rect 187285 521722 187323 521724
rect 185753 521652 186207 521668
rect 186365 521666 186629 521682
rect 185261 521610 185711 521632
rect 186365 521632 186381 521666
rect 186415 521632 186480 521666
rect 186514 521632 186579 521666
rect 186613 521632 186629 521666
rect 186671 521668 186687 521702
rect 186721 521668 186790 521702
rect 186824 521668 186893 521702
rect 186927 521668 186943 521702
rect 186671 521652 186943 521668
rect 187257 521706 187323 521722
rect 187257 521672 187273 521706
rect 187307 521672 187323 521706
rect 187257 521656 187323 521672
rect 187365 521666 187431 521682
rect 186365 521610 186629 521632
rect 187365 521632 187381 521666
rect 187415 521632 187431 521666
rect 187365 521616 187431 521632
rect 187365 521614 187403 521616
rect 172565 521584 173511 521610
rect 173669 521584 174615 521610
rect 174957 521584 175903 521610
rect 176061 521584 177007 521610
rect 177165 521584 178111 521610
rect 178269 521584 179215 521610
rect 179373 521584 179767 521610
rect 180109 521584 181055 521610
rect 181213 521584 182159 521610
rect 182317 521584 183263 521610
rect 183421 521584 184367 521610
rect 184525 521584 184919 521610
rect 185261 521584 186207 521610
rect 186365 521584 186943 521610
rect 187285 521584 187403 521614
rect 172289 521384 172407 521410
rect 172565 521384 173511 521410
rect 173669 521384 174615 521410
rect 174957 521384 175903 521410
rect 176061 521384 177007 521410
rect 177165 521384 178111 521410
rect 178269 521384 179215 521410
rect 179373 521384 179767 521410
rect 180109 521384 181055 521410
rect 181213 521384 182159 521410
rect 182317 521384 183263 521410
rect 183421 521384 184367 521410
rect 184525 521384 184919 521410
rect 185261 521384 186207 521410
rect 186365 521384 186943 521410
rect 187285 521384 187403 521410
rect 172289 521316 172407 521342
rect 172565 521316 173511 521342
rect 173669 521316 174615 521342
rect 174773 521316 175719 521342
rect 175877 521316 176823 521342
rect 176981 521316 177191 521342
rect 177533 521316 178479 521342
rect 178637 521316 179583 521342
rect 179741 521316 180687 521342
rect 180845 521316 181791 521342
rect 181949 521316 182343 521342
rect 182685 521316 183631 521342
rect 183789 521316 184735 521342
rect 184893 521316 185839 521342
rect 185997 521316 186943 521342
rect 187285 521316 187403 521342
rect 172289 521112 172407 521142
rect 172565 521116 173511 521142
rect 173669 521116 174615 521142
rect 174773 521116 175719 521142
rect 175877 521116 176823 521142
rect 176981 521116 177191 521142
rect 177533 521116 178479 521142
rect 178637 521116 179583 521142
rect 179741 521116 180687 521142
rect 180845 521116 181791 521142
rect 181949 521116 182343 521142
rect 182685 521116 183631 521142
rect 183789 521116 184735 521142
rect 184893 521116 185839 521142
rect 185997 521116 186943 521142
rect 172289 521110 172327 521112
rect 172261 521094 172327 521110
rect 172261 521060 172277 521094
rect 172311 521060 172327 521094
rect 172565 521094 173015 521116
rect 172261 521044 172327 521060
rect 172369 521054 172435 521070
rect 172369 521020 172385 521054
rect 172419 521020 172435 521054
rect 172565 521060 172837 521094
rect 172871 521060 173015 521094
rect 173669 521094 174119 521116
rect 172565 521044 173015 521060
rect 173057 521058 173511 521074
rect 172369 521004 172435 521020
rect 173057 521024 173201 521058
rect 173235 521024 173511 521058
rect 173669 521060 173941 521094
rect 173975 521060 174119 521094
rect 174773 521094 175223 521116
rect 173669 521044 174119 521060
rect 174161 521058 174615 521074
rect 172369 521002 172407 521004
rect 173057 521002 173511 521024
rect 174161 521024 174305 521058
rect 174339 521024 174615 521058
rect 174773 521060 175045 521094
rect 175079 521060 175223 521094
rect 175877 521094 176327 521116
rect 176981 521110 177065 521116
rect 174773 521044 175223 521060
rect 175265 521058 175719 521074
rect 174161 521002 174615 521024
rect 175265 521024 175409 521058
rect 175443 521024 175719 521058
rect 175877 521060 176149 521094
rect 176183 521060 176327 521094
rect 176923 521094 177065 521110
rect 175877 521044 176327 521060
rect 176369 521058 176823 521074
rect 175265 521002 175719 521024
rect 176369 521024 176513 521058
rect 176547 521024 176823 521058
rect 176923 521060 176939 521094
rect 176973 521060 177065 521094
rect 177533 521094 177983 521116
rect 176923 521044 177065 521060
rect 177107 521058 177249 521074
rect 176369 521002 176823 521024
rect 177107 521024 177199 521058
rect 177233 521024 177249 521058
rect 177533 521060 177805 521094
rect 177839 521060 177983 521094
rect 178637 521094 179087 521116
rect 177533 521044 177983 521060
rect 178025 521058 178479 521074
rect 177107 521008 177249 521024
rect 178025 521024 178169 521058
rect 178203 521024 178479 521058
rect 178637 521060 178909 521094
rect 178943 521060 179087 521094
rect 179741 521094 180191 521116
rect 178637 521044 179087 521060
rect 179129 521058 179583 521074
rect 177107 521002 177191 521008
rect 178025 521002 178479 521024
rect 179129 521024 179273 521058
rect 179307 521024 179583 521058
rect 179741 521060 180013 521094
rect 180047 521060 180191 521094
rect 180845 521094 181295 521116
rect 179741 521044 180191 521060
rect 180233 521058 180687 521074
rect 179129 521002 179583 521024
rect 180233 521024 180377 521058
rect 180411 521024 180687 521058
rect 180845 521060 181117 521094
rect 181151 521060 181295 521094
rect 181949 521094 182125 521116
rect 180845 521044 181295 521060
rect 181337 521058 181791 521074
rect 180233 521002 180687 521024
rect 181337 521024 181481 521058
rect 181515 521024 181791 521058
rect 181949 521060 181965 521094
rect 181999 521060 182075 521094
rect 182109 521060 182125 521094
rect 182685 521094 183135 521116
rect 181949 521044 182125 521060
rect 182167 521058 182343 521074
rect 181337 521002 181791 521024
rect 182167 521024 182183 521058
rect 182217 521024 182293 521058
rect 182327 521024 182343 521058
rect 182685 521060 182957 521094
rect 182991 521060 183135 521094
rect 183789 521094 184239 521116
rect 182685 521044 183135 521060
rect 183177 521058 183631 521074
rect 182167 521002 182343 521024
rect 183177 521024 183321 521058
rect 183355 521024 183631 521058
rect 183789 521060 184061 521094
rect 184095 521060 184239 521094
rect 184893 521094 185343 521116
rect 183789 521044 184239 521060
rect 184281 521058 184735 521074
rect 183177 521002 183631 521024
rect 184281 521024 184425 521058
rect 184459 521024 184735 521058
rect 184893 521060 185165 521094
rect 185199 521060 185343 521094
rect 185997 521094 186447 521116
rect 187285 521112 187403 521142
rect 184893 521044 185343 521060
rect 185385 521058 185839 521074
rect 184281 521002 184735 521024
rect 185385 521024 185529 521058
rect 185563 521024 185839 521058
rect 185997 521060 186269 521094
rect 186303 521060 186447 521094
rect 187365 521110 187403 521112
rect 187365 521094 187431 521110
rect 185997 521044 186447 521060
rect 186489 521058 186943 521074
rect 185385 521002 185839 521024
rect 186489 521024 186633 521058
rect 186667 521024 186943 521058
rect 186489 521002 186943 521024
rect 187257 521054 187323 521070
rect 187257 521020 187273 521054
rect 187307 521020 187323 521054
rect 187365 521060 187381 521094
rect 187415 521060 187431 521094
rect 187365 521044 187431 521060
rect 187257 521004 187323 521020
rect 172289 520976 172407 521002
rect 172565 520976 173511 521002
rect 173669 520976 174615 521002
rect 174773 520976 175719 521002
rect 175877 520976 176823 521002
rect 176981 520976 177191 521002
rect 177533 520976 178479 521002
rect 178637 520976 179583 521002
rect 179741 520976 180687 521002
rect 180845 520976 181791 521002
rect 181949 520976 182343 521002
rect 182685 520976 183631 521002
rect 183789 520976 184735 521002
rect 184893 520976 185839 521002
rect 185997 520976 186943 521002
rect 187285 521002 187323 521004
rect 187285 520976 187403 521002
rect 172289 520840 172407 520866
rect 172565 520840 173511 520866
rect 173669 520840 174615 520866
rect 174773 520840 175719 520866
rect 175877 520840 176823 520866
rect 176981 520840 177191 520866
rect 177533 520840 178479 520866
rect 178637 520840 179583 520866
rect 179741 520840 180687 520866
rect 180845 520840 181791 520866
rect 181949 520840 182343 520866
rect 182685 520840 183631 520866
rect 183789 520840 184735 520866
rect 184893 520840 185839 520866
rect 185997 520840 186943 520866
rect 187285 520840 187403 520866
rect 172289 520772 172407 520798
rect 172565 520772 173511 520798
rect 173669 520772 174615 520798
rect 174957 520772 175903 520798
rect 176061 520772 177007 520798
rect 177165 520772 178111 520798
rect 178269 520772 179215 520798
rect 179373 520772 179767 520798
rect 180109 520772 181055 520798
rect 181213 520772 182159 520798
rect 182317 520772 183263 520798
rect 183421 520772 184367 520798
rect 184525 520772 184919 520798
rect 185261 520772 186207 520798
rect 186365 520772 186943 520798
rect 187285 520772 187403 520798
rect 172289 520636 172407 520662
rect 172565 520636 173511 520662
rect 173669 520636 174615 520662
rect 174957 520636 175903 520662
rect 176061 520636 177007 520662
rect 177165 520636 178111 520662
rect 178269 520636 179215 520662
rect 179373 520636 179767 520662
rect 180109 520636 181055 520662
rect 181213 520636 182159 520662
rect 182317 520636 183263 520662
rect 183421 520636 184367 520662
rect 184525 520636 184919 520662
rect 185261 520636 186207 520662
rect 186365 520636 186943 520662
rect 172369 520634 172407 520636
rect 172369 520618 172435 520634
rect 172261 520578 172327 520594
rect 172261 520544 172277 520578
rect 172311 520544 172327 520578
rect 172369 520584 172385 520618
rect 172419 520584 172435 520618
rect 173057 520614 173511 520636
rect 172369 520568 172435 520584
rect 172565 520578 173015 520594
rect 172261 520528 172327 520544
rect 172289 520526 172327 520528
rect 172565 520544 172837 520578
rect 172871 520544 173015 520578
rect 173057 520580 173201 520614
rect 173235 520580 173511 520614
rect 174161 520614 174615 520636
rect 173057 520564 173511 520580
rect 173669 520578 174119 520594
rect 172289 520496 172407 520526
rect 172565 520522 173015 520544
rect 173669 520544 173941 520578
rect 173975 520544 174119 520578
rect 174161 520580 174305 520614
rect 174339 520580 174615 520614
rect 175449 520614 175903 520636
rect 174161 520564 174615 520580
rect 174957 520578 175407 520594
rect 173669 520522 174119 520544
rect 174957 520544 175229 520578
rect 175263 520544 175407 520578
rect 175449 520580 175593 520614
rect 175627 520580 175903 520614
rect 176553 520614 177007 520636
rect 175449 520564 175903 520580
rect 176061 520578 176511 520594
rect 174957 520522 175407 520544
rect 176061 520544 176333 520578
rect 176367 520544 176511 520578
rect 176553 520580 176697 520614
rect 176731 520580 177007 520614
rect 177657 520614 178111 520636
rect 176553 520564 177007 520580
rect 177165 520578 177615 520594
rect 176061 520522 176511 520544
rect 177165 520544 177437 520578
rect 177471 520544 177615 520578
rect 177657 520580 177801 520614
rect 177835 520580 178111 520614
rect 178761 520614 179215 520636
rect 177657 520564 178111 520580
rect 178269 520578 178719 520594
rect 177165 520522 177615 520544
rect 178269 520544 178541 520578
rect 178575 520544 178719 520578
rect 178761 520580 178905 520614
rect 178939 520580 179215 520614
rect 179591 520614 179767 520636
rect 178761 520564 179215 520580
rect 179373 520578 179549 520594
rect 178269 520522 178719 520544
rect 179373 520544 179389 520578
rect 179423 520544 179499 520578
rect 179533 520544 179549 520578
rect 179591 520580 179607 520614
rect 179641 520580 179717 520614
rect 179751 520580 179767 520614
rect 180601 520614 181055 520636
rect 179591 520564 179767 520580
rect 180109 520578 180559 520594
rect 179373 520522 179549 520544
rect 180109 520544 180381 520578
rect 180415 520544 180559 520578
rect 180601 520580 180745 520614
rect 180779 520580 181055 520614
rect 181705 520614 182159 520636
rect 180601 520564 181055 520580
rect 181213 520578 181663 520594
rect 180109 520522 180559 520544
rect 181213 520544 181485 520578
rect 181519 520544 181663 520578
rect 181705 520580 181849 520614
rect 181883 520580 182159 520614
rect 182809 520614 183263 520636
rect 181705 520564 182159 520580
rect 182317 520578 182767 520594
rect 181213 520522 181663 520544
rect 182317 520544 182589 520578
rect 182623 520544 182767 520578
rect 182809 520580 182953 520614
rect 182987 520580 183263 520614
rect 183913 520614 184367 520636
rect 182809 520564 183263 520580
rect 183421 520578 183871 520594
rect 182317 520522 182767 520544
rect 183421 520544 183693 520578
rect 183727 520544 183871 520578
rect 183913 520580 184057 520614
rect 184091 520580 184367 520614
rect 184743 520614 184919 520636
rect 183913 520564 184367 520580
rect 184525 520578 184701 520594
rect 183421 520522 183871 520544
rect 184525 520544 184541 520578
rect 184575 520544 184651 520578
rect 184685 520544 184701 520578
rect 184743 520580 184759 520614
rect 184793 520580 184869 520614
rect 184903 520580 184919 520614
rect 185753 520614 186207 520636
rect 184743 520564 184919 520580
rect 185261 520578 185711 520594
rect 184525 520522 184701 520544
rect 185261 520544 185533 520578
rect 185567 520544 185711 520578
rect 185753 520580 185897 520614
rect 185931 520580 186207 520614
rect 186671 520614 186943 520636
rect 187285 520636 187403 520662
rect 187285 520634 187323 520636
rect 185753 520564 186207 520580
rect 186365 520578 186629 520594
rect 185261 520522 185711 520544
rect 186365 520544 186381 520578
rect 186415 520544 186480 520578
rect 186514 520544 186579 520578
rect 186613 520544 186629 520578
rect 186671 520580 186687 520614
rect 186721 520580 186790 520614
rect 186824 520580 186893 520614
rect 186927 520580 186943 520614
rect 186671 520564 186943 520580
rect 187257 520618 187323 520634
rect 187257 520584 187273 520618
rect 187307 520584 187323 520618
rect 187257 520568 187323 520584
rect 187365 520578 187431 520594
rect 186365 520522 186629 520544
rect 187365 520544 187381 520578
rect 187415 520544 187431 520578
rect 187365 520528 187431 520544
rect 187365 520526 187403 520528
rect 172565 520496 173511 520522
rect 173669 520496 174615 520522
rect 174957 520496 175903 520522
rect 176061 520496 177007 520522
rect 177165 520496 178111 520522
rect 178269 520496 179215 520522
rect 179373 520496 179767 520522
rect 180109 520496 181055 520522
rect 181213 520496 182159 520522
rect 182317 520496 183263 520522
rect 183421 520496 184367 520522
rect 184525 520496 184919 520522
rect 185261 520496 186207 520522
rect 186365 520496 186943 520522
rect 187285 520496 187403 520526
rect 172289 520296 172407 520322
rect 172565 520296 173511 520322
rect 173669 520296 174615 520322
rect 174957 520296 175903 520322
rect 176061 520296 177007 520322
rect 177165 520296 178111 520322
rect 178269 520296 179215 520322
rect 179373 520296 179767 520322
rect 180109 520296 181055 520322
rect 181213 520296 182159 520322
rect 182317 520296 183263 520322
rect 183421 520296 184367 520322
rect 184525 520296 184919 520322
rect 185261 520296 186207 520322
rect 186365 520296 186943 520322
rect 187285 520296 187403 520322
rect 172289 520228 172407 520254
rect 172565 520228 173511 520254
rect 173669 520228 174615 520254
rect 174773 520228 175719 520254
rect 175877 520228 176823 520254
rect 176981 520228 177191 520254
rect 177533 520228 178479 520254
rect 178637 520228 179583 520254
rect 179741 520228 180687 520254
rect 180845 520228 181791 520254
rect 181949 520228 182343 520254
rect 182685 520228 183631 520254
rect 183789 520228 184735 520254
rect 184893 520228 185839 520254
rect 185997 520228 186943 520254
rect 187285 520228 187403 520254
rect 172289 520024 172407 520054
rect 172565 520028 173511 520054
rect 173669 520028 174615 520054
rect 174773 520028 175719 520054
rect 175877 520028 176823 520054
rect 176981 520028 177191 520054
rect 177533 520028 178479 520054
rect 178637 520028 179583 520054
rect 179741 520028 180687 520054
rect 180845 520028 181791 520054
rect 181949 520028 182343 520054
rect 182685 520028 183631 520054
rect 183789 520028 184735 520054
rect 184893 520028 185839 520054
rect 185997 520028 186943 520054
rect 172289 520022 172327 520024
rect 172261 520006 172327 520022
rect 172261 519972 172277 520006
rect 172311 519972 172327 520006
rect 172565 520006 173015 520028
rect 172261 519956 172327 519972
rect 172369 519966 172435 519982
rect 172369 519932 172385 519966
rect 172419 519932 172435 519966
rect 172565 519972 172837 520006
rect 172871 519972 173015 520006
rect 173669 520006 174119 520028
rect 172565 519956 173015 519972
rect 173057 519970 173511 519986
rect 172369 519916 172435 519932
rect 173057 519936 173201 519970
rect 173235 519936 173511 519970
rect 173669 519972 173941 520006
rect 173975 519972 174119 520006
rect 174773 520006 175223 520028
rect 173669 519956 174119 519972
rect 174161 519970 174615 519986
rect 172369 519914 172407 519916
rect 173057 519914 173511 519936
rect 174161 519936 174305 519970
rect 174339 519936 174615 519970
rect 174773 519972 175045 520006
rect 175079 519972 175223 520006
rect 175877 520006 176327 520028
rect 176981 520022 177065 520028
rect 174773 519956 175223 519972
rect 175265 519970 175719 519986
rect 174161 519914 174615 519936
rect 175265 519936 175409 519970
rect 175443 519936 175719 519970
rect 175877 519972 176149 520006
rect 176183 519972 176327 520006
rect 176923 520006 177065 520022
rect 175877 519956 176327 519972
rect 176369 519970 176823 519986
rect 175265 519914 175719 519936
rect 176369 519936 176513 519970
rect 176547 519936 176823 519970
rect 176923 519972 176939 520006
rect 176973 519972 177065 520006
rect 177533 520006 177983 520028
rect 176923 519956 177065 519972
rect 177107 519970 177249 519986
rect 176369 519914 176823 519936
rect 177107 519936 177199 519970
rect 177233 519936 177249 519970
rect 177533 519972 177805 520006
rect 177839 519972 177983 520006
rect 178637 520006 179087 520028
rect 177533 519956 177983 519972
rect 178025 519970 178479 519986
rect 177107 519920 177249 519936
rect 178025 519936 178169 519970
rect 178203 519936 178479 519970
rect 178637 519972 178909 520006
rect 178943 519972 179087 520006
rect 179741 520006 180191 520028
rect 178637 519956 179087 519972
rect 179129 519970 179583 519986
rect 177107 519914 177191 519920
rect 178025 519914 178479 519936
rect 179129 519936 179273 519970
rect 179307 519936 179583 519970
rect 179741 519972 180013 520006
rect 180047 519972 180191 520006
rect 180845 520006 181295 520028
rect 179741 519956 180191 519972
rect 180233 519970 180687 519986
rect 179129 519914 179583 519936
rect 180233 519936 180377 519970
rect 180411 519936 180687 519970
rect 180845 519972 181117 520006
rect 181151 519972 181295 520006
rect 181949 520006 182125 520028
rect 180845 519956 181295 519972
rect 181337 519970 181791 519986
rect 180233 519914 180687 519936
rect 181337 519936 181481 519970
rect 181515 519936 181791 519970
rect 181949 519972 181965 520006
rect 181999 519972 182075 520006
rect 182109 519972 182125 520006
rect 182685 520006 183135 520028
rect 181949 519956 182125 519972
rect 182167 519970 182343 519986
rect 181337 519914 181791 519936
rect 182167 519936 182183 519970
rect 182217 519936 182293 519970
rect 182327 519936 182343 519970
rect 182685 519972 182957 520006
rect 182991 519972 183135 520006
rect 183789 520006 184239 520028
rect 182685 519956 183135 519972
rect 183177 519970 183631 519986
rect 182167 519914 182343 519936
rect 183177 519936 183321 519970
rect 183355 519936 183631 519970
rect 183789 519972 184061 520006
rect 184095 519972 184239 520006
rect 184893 520006 185343 520028
rect 183789 519956 184239 519972
rect 184281 519970 184735 519986
rect 183177 519914 183631 519936
rect 184281 519936 184425 519970
rect 184459 519936 184735 519970
rect 184893 519972 185165 520006
rect 185199 519972 185343 520006
rect 185997 520006 186447 520028
rect 187285 520024 187403 520054
rect 184893 519956 185343 519972
rect 185385 519970 185839 519986
rect 184281 519914 184735 519936
rect 185385 519936 185529 519970
rect 185563 519936 185839 519970
rect 185997 519972 186269 520006
rect 186303 519972 186447 520006
rect 187365 520022 187403 520024
rect 187365 520006 187431 520022
rect 185997 519956 186447 519972
rect 186489 519970 186943 519986
rect 185385 519914 185839 519936
rect 186489 519936 186633 519970
rect 186667 519936 186943 519970
rect 186489 519914 186943 519936
rect 187257 519966 187323 519982
rect 187257 519932 187273 519966
rect 187307 519932 187323 519966
rect 187365 519972 187381 520006
rect 187415 519972 187431 520006
rect 187365 519956 187431 519972
rect 187257 519916 187323 519932
rect 172289 519888 172407 519914
rect 172565 519888 173511 519914
rect 173669 519888 174615 519914
rect 174773 519888 175719 519914
rect 175877 519888 176823 519914
rect 176981 519888 177191 519914
rect 177533 519888 178479 519914
rect 178637 519888 179583 519914
rect 179741 519888 180687 519914
rect 180845 519888 181791 519914
rect 181949 519888 182343 519914
rect 182685 519888 183631 519914
rect 183789 519888 184735 519914
rect 184893 519888 185839 519914
rect 185997 519888 186943 519914
rect 187285 519914 187323 519916
rect 187285 519888 187403 519914
rect 172289 519752 172407 519778
rect 172565 519752 173511 519778
rect 173669 519752 174615 519778
rect 174773 519752 175719 519778
rect 175877 519752 176823 519778
rect 176981 519752 177191 519778
rect 177533 519752 178479 519778
rect 178637 519752 179583 519778
rect 179741 519752 180687 519778
rect 180845 519752 181791 519778
rect 181949 519752 182343 519778
rect 182685 519752 183631 519778
rect 183789 519752 184735 519778
rect 184893 519752 185839 519778
rect 185997 519752 186943 519778
rect 187285 519752 187403 519778
rect 172289 519684 172407 519710
rect 172565 519684 173511 519710
rect 173669 519684 174615 519710
rect 174957 519684 175903 519710
rect 176061 519684 177007 519710
rect 177165 519684 178111 519710
rect 178269 519684 179215 519710
rect 179373 519684 179767 519710
rect 180109 519684 181055 519710
rect 181213 519684 182159 519710
rect 182317 519684 183263 519710
rect 183421 519684 184367 519710
rect 184525 519684 184919 519710
rect 185261 519684 186207 519710
rect 186365 519684 186943 519710
rect 187285 519684 187403 519710
rect 172289 519548 172407 519574
rect 172565 519548 173511 519574
rect 173669 519548 174615 519574
rect 174957 519548 175903 519574
rect 176061 519548 177007 519574
rect 177165 519548 178111 519574
rect 178269 519548 179215 519574
rect 179373 519548 179767 519574
rect 180109 519548 181055 519574
rect 181213 519548 182159 519574
rect 182317 519548 183263 519574
rect 183421 519548 184367 519574
rect 184525 519548 184919 519574
rect 185261 519548 186207 519574
rect 186365 519548 186943 519574
rect 172369 519546 172407 519548
rect 172369 519530 172435 519546
rect 172261 519490 172327 519506
rect 172261 519456 172277 519490
rect 172311 519456 172327 519490
rect 172369 519496 172385 519530
rect 172419 519496 172435 519530
rect 173057 519526 173511 519548
rect 172369 519480 172435 519496
rect 172565 519490 173015 519506
rect 172261 519440 172327 519456
rect 172289 519438 172327 519440
rect 172565 519456 172837 519490
rect 172871 519456 173015 519490
rect 173057 519492 173201 519526
rect 173235 519492 173511 519526
rect 174161 519526 174615 519548
rect 173057 519476 173511 519492
rect 173669 519490 174119 519506
rect 172289 519408 172407 519438
rect 172565 519434 173015 519456
rect 173669 519456 173941 519490
rect 173975 519456 174119 519490
rect 174161 519492 174305 519526
rect 174339 519492 174615 519526
rect 175449 519526 175903 519548
rect 174161 519476 174615 519492
rect 174957 519490 175407 519506
rect 173669 519434 174119 519456
rect 174957 519456 175229 519490
rect 175263 519456 175407 519490
rect 175449 519492 175593 519526
rect 175627 519492 175903 519526
rect 176553 519526 177007 519548
rect 175449 519476 175903 519492
rect 176061 519490 176511 519506
rect 174957 519434 175407 519456
rect 176061 519456 176333 519490
rect 176367 519456 176511 519490
rect 176553 519492 176697 519526
rect 176731 519492 177007 519526
rect 177657 519526 178111 519548
rect 176553 519476 177007 519492
rect 177165 519490 177615 519506
rect 176061 519434 176511 519456
rect 177165 519456 177437 519490
rect 177471 519456 177615 519490
rect 177657 519492 177801 519526
rect 177835 519492 178111 519526
rect 178761 519526 179215 519548
rect 177657 519476 178111 519492
rect 178269 519490 178719 519506
rect 177165 519434 177615 519456
rect 178269 519456 178541 519490
rect 178575 519456 178719 519490
rect 178761 519492 178905 519526
rect 178939 519492 179215 519526
rect 179591 519526 179767 519548
rect 178761 519476 179215 519492
rect 179373 519490 179549 519506
rect 178269 519434 178719 519456
rect 179373 519456 179389 519490
rect 179423 519456 179499 519490
rect 179533 519456 179549 519490
rect 179591 519492 179607 519526
rect 179641 519492 179717 519526
rect 179751 519492 179767 519526
rect 180601 519526 181055 519548
rect 179591 519476 179767 519492
rect 180109 519490 180559 519506
rect 179373 519434 179549 519456
rect 180109 519456 180381 519490
rect 180415 519456 180559 519490
rect 180601 519492 180745 519526
rect 180779 519492 181055 519526
rect 181705 519526 182159 519548
rect 180601 519476 181055 519492
rect 181213 519490 181663 519506
rect 180109 519434 180559 519456
rect 181213 519456 181485 519490
rect 181519 519456 181663 519490
rect 181705 519492 181849 519526
rect 181883 519492 182159 519526
rect 182809 519526 183263 519548
rect 181705 519476 182159 519492
rect 182317 519490 182767 519506
rect 181213 519434 181663 519456
rect 182317 519456 182589 519490
rect 182623 519456 182767 519490
rect 182809 519492 182953 519526
rect 182987 519492 183263 519526
rect 183913 519526 184367 519548
rect 182809 519476 183263 519492
rect 183421 519490 183871 519506
rect 182317 519434 182767 519456
rect 183421 519456 183693 519490
rect 183727 519456 183871 519490
rect 183913 519492 184057 519526
rect 184091 519492 184367 519526
rect 184743 519526 184919 519548
rect 183913 519476 184367 519492
rect 184525 519490 184701 519506
rect 183421 519434 183871 519456
rect 184525 519456 184541 519490
rect 184575 519456 184651 519490
rect 184685 519456 184701 519490
rect 184743 519492 184759 519526
rect 184793 519492 184869 519526
rect 184903 519492 184919 519526
rect 185753 519526 186207 519548
rect 184743 519476 184919 519492
rect 185261 519490 185711 519506
rect 184525 519434 184701 519456
rect 185261 519456 185533 519490
rect 185567 519456 185711 519490
rect 185753 519492 185897 519526
rect 185931 519492 186207 519526
rect 186671 519526 186943 519548
rect 187285 519548 187403 519574
rect 187285 519546 187323 519548
rect 185753 519476 186207 519492
rect 186365 519490 186629 519506
rect 185261 519434 185711 519456
rect 186365 519456 186381 519490
rect 186415 519456 186480 519490
rect 186514 519456 186579 519490
rect 186613 519456 186629 519490
rect 186671 519492 186687 519526
rect 186721 519492 186790 519526
rect 186824 519492 186893 519526
rect 186927 519492 186943 519526
rect 186671 519476 186943 519492
rect 187257 519530 187323 519546
rect 187257 519496 187273 519530
rect 187307 519496 187323 519530
rect 187257 519480 187323 519496
rect 187365 519490 187431 519506
rect 186365 519434 186629 519456
rect 187365 519456 187381 519490
rect 187415 519456 187431 519490
rect 187365 519440 187431 519456
rect 187365 519438 187403 519440
rect 172565 519408 173511 519434
rect 173669 519408 174615 519434
rect 174957 519408 175903 519434
rect 176061 519408 177007 519434
rect 177165 519408 178111 519434
rect 178269 519408 179215 519434
rect 179373 519408 179767 519434
rect 180109 519408 181055 519434
rect 181213 519408 182159 519434
rect 182317 519408 183263 519434
rect 183421 519408 184367 519434
rect 184525 519408 184919 519434
rect 185261 519408 186207 519434
rect 186365 519408 186943 519434
rect 187285 519408 187403 519438
rect 172289 519208 172407 519234
rect 172565 519208 173511 519234
rect 173669 519208 174615 519234
rect 174957 519208 175903 519234
rect 176061 519208 177007 519234
rect 177165 519208 178111 519234
rect 178269 519208 179215 519234
rect 179373 519208 179767 519234
rect 180109 519208 181055 519234
rect 181213 519208 182159 519234
rect 182317 519208 183263 519234
rect 183421 519208 184367 519234
rect 184525 519208 184919 519234
rect 185261 519208 186207 519234
rect 186365 519208 186943 519234
rect 187285 519208 187403 519234
rect 172289 519140 172407 519166
rect 172565 519140 173511 519166
rect 173669 519140 174615 519166
rect 174773 519140 175719 519166
rect 175877 519140 176823 519166
rect 176981 519140 177191 519166
rect 177533 519140 178479 519166
rect 178637 519140 179583 519166
rect 179741 519140 180687 519166
rect 180845 519140 181791 519166
rect 181949 519140 182343 519166
rect 182685 519140 183631 519166
rect 183789 519140 184735 519166
rect 184893 519140 185839 519166
rect 185997 519140 186943 519166
rect 187285 519140 187403 519166
rect 172289 518936 172407 518966
rect 172565 518940 173511 518966
rect 173669 518940 174615 518966
rect 174773 518940 175719 518966
rect 175877 518940 176823 518966
rect 176981 518940 177191 518966
rect 177533 518940 178479 518966
rect 178637 518940 179583 518966
rect 179741 518940 180687 518966
rect 180845 518940 181791 518966
rect 181949 518940 182343 518966
rect 182685 518940 183631 518966
rect 183789 518940 184735 518966
rect 184893 518940 185839 518966
rect 185997 518940 186943 518966
rect 172289 518934 172327 518936
rect 172261 518918 172327 518934
rect 172261 518884 172277 518918
rect 172311 518884 172327 518918
rect 172565 518918 173015 518940
rect 172261 518868 172327 518884
rect 172369 518878 172435 518894
rect 172369 518844 172385 518878
rect 172419 518844 172435 518878
rect 172565 518884 172837 518918
rect 172871 518884 173015 518918
rect 173669 518918 174119 518940
rect 172565 518868 173015 518884
rect 173057 518882 173511 518898
rect 172369 518828 172435 518844
rect 173057 518848 173201 518882
rect 173235 518848 173511 518882
rect 173669 518884 173941 518918
rect 173975 518884 174119 518918
rect 174773 518918 175223 518940
rect 173669 518868 174119 518884
rect 174161 518882 174615 518898
rect 172369 518826 172407 518828
rect 173057 518826 173511 518848
rect 174161 518848 174305 518882
rect 174339 518848 174615 518882
rect 174773 518884 175045 518918
rect 175079 518884 175223 518918
rect 175877 518918 176327 518940
rect 176981 518934 177065 518940
rect 174773 518868 175223 518884
rect 175265 518882 175719 518898
rect 174161 518826 174615 518848
rect 175265 518848 175409 518882
rect 175443 518848 175719 518882
rect 175877 518884 176149 518918
rect 176183 518884 176327 518918
rect 176923 518918 177065 518934
rect 175877 518868 176327 518884
rect 176369 518882 176823 518898
rect 175265 518826 175719 518848
rect 176369 518848 176513 518882
rect 176547 518848 176823 518882
rect 176923 518884 176939 518918
rect 176973 518884 177065 518918
rect 177533 518918 177983 518940
rect 176923 518868 177065 518884
rect 177107 518882 177249 518898
rect 176369 518826 176823 518848
rect 177107 518848 177199 518882
rect 177233 518848 177249 518882
rect 177533 518884 177805 518918
rect 177839 518884 177983 518918
rect 178637 518918 179087 518940
rect 177533 518868 177983 518884
rect 178025 518882 178479 518898
rect 177107 518832 177249 518848
rect 178025 518848 178169 518882
rect 178203 518848 178479 518882
rect 178637 518884 178909 518918
rect 178943 518884 179087 518918
rect 179741 518918 180191 518940
rect 178637 518868 179087 518884
rect 179129 518882 179583 518898
rect 177107 518826 177191 518832
rect 178025 518826 178479 518848
rect 179129 518848 179273 518882
rect 179307 518848 179583 518882
rect 179741 518884 180013 518918
rect 180047 518884 180191 518918
rect 180845 518918 181295 518940
rect 179741 518868 180191 518884
rect 180233 518882 180687 518898
rect 179129 518826 179583 518848
rect 180233 518848 180377 518882
rect 180411 518848 180687 518882
rect 180845 518884 181117 518918
rect 181151 518884 181295 518918
rect 181949 518918 182125 518940
rect 180845 518868 181295 518884
rect 181337 518882 181791 518898
rect 180233 518826 180687 518848
rect 181337 518848 181481 518882
rect 181515 518848 181791 518882
rect 181949 518884 181965 518918
rect 181999 518884 182075 518918
rect 182109 518884 182125 518918
rect 182685 518918 183135 518940
rect 181949 518868 182125 518884
rect 182167 518882 182343 518898
rect 181337 518826 181791 518848
rect 182167 518848 182183 518882
rect 182217 518848 182293 518882
rect 182327 518848 182343 518882
rect 182685 518884 182957 518918
rect 182991 518884 183135 518918
rect 183789 518918 184239 518940
rect 182685 518868 183135 518884
rect 183177 518882 183631 518898
rect 182167 518826 182343 518848
rect 183177 518848 183321 518882
rect 183355 518848 183631 518882
rect 183789 518884 184061 518918
rect 184095 518884 184239 518918
rect 184893 518918 185343 518940
rect 183789 518868 184239 518884
rect 184281 518882 184735 518898
rect 183177 518826 183631 518848
rect 184281 518848 184425 518882
rect 184459 518848 184735 518882
rect 184893 518884 185165 518918
rect 185199 518884 185343 518918
rect 185997 518918 186447 518940
rect 187285 518936 187403 518966
rect 184893 518868 185343 518884
rect 185385 518882 185839 518898
rect 184281 518826 184735 518848
rect 185385 518848 185529 518882
rect 185563 518848 185839 518882
rect 185997 518884 186269 518918
rect 186303 518884 186447 518918
rect 187365 518934 187403 518936
rect 187365 518918 187431 518934
rect 185997 518868 186447 518884
rect 186489 518882 186943 518898
rect 185385 518826 185839 518848
rect 186489 518848 186633 518882
rect 186667 518848 186943 518882
rect 186489 518826 186943 518848
rect 187257 518878 187323 518894
rect 187257 518844 187273 518878
rect 187307 518844 187323 518878
rect 187365 518884 187381 518918
rect 187415 518884 187431 518918
rect 187365 518868 187431 518884
rect 187257 518828 187323 518844
rect 172289 518800 172407 518826
rect 172565 518800 173511 518826
rect 173669 518800 174615 518826
rect 174773 518800 175719 518826
rect 175877 518800 176823 518826
rect 176981 518800 177191 518826
rect 177533 518800 178479 518826
rect 178637 518800 179583 518826
rect 179741 518800 180687 518826
rect 180845 518800 181791 518826
rect 181949 518800 182343 518826
rect 182685 518800 183631 518826
rect 183789 518800 184735 518826
rect 184893 518800 185839 518826
rect 185997 518800 186943 518826
rect 187285 518826 187323 518828
rect 187285 518800 187403 518826
rect 172289 518664 172407 518690
rect 172565 518664 173511 518690
rect 173669 518664 174615 518690
rect 174773 518664 175719 518690
rect 175877 518664 176823 518690
rect 176981 518664 177191 518690
rect 177533 518664 178479 518690
rect 178637 518664 179583 518690
rect 179741 518664 180687 518690
rect 180845 518664 181791 518690
rect 181949 518664 182343 518690
rect 182685 518664 183631 518690
rect 183789 518664 184735 518690
rect 184893 518664 185839 518690
rect 185997 518664 186943 518690
rect 187285 518664 187403 518690
rect 172289 518596 172407 518622
rect 172565 518596 173511 518622
rect 173669 518596 174615 518622
rect 174957 518596 175903 518622
rect 176061 518596 177007 518622
rect 177165 518596 178111 518622
rect 178269 518596 179215 518622
rect 179373 518596 179767 518622
rect 180109 518596 181055 518622
rect 181213 518596 182159 518622
rect 182317 518596 183263 518622
rect 183421 518596 184367 518622
rect 184525 518596 184919 518622
rect 185261 518596 186207 518622
rect 186365 518596 186943 518622
rect 187285 518596 187403 518622
rect 172289 518460 172407 518486
rect 172565 518460 173511 518486
rect 173669 518460 174615 518486
rect 174957 518460 175903 518486
rect 176061 518460 177007 518486
rect 177165 518460 178111 518486
rect 178269 518460 179215 518486
rect 179373 518460 179767 518486
rect 180109 518460 181055 518486
rect 181213 518460 182159 518486
rect 182317 518460 183263 518486
rect 183421 518460 184367 518486
rect 184525 518460 184919 518486
rect 185261 518460 186207 518486
rect 186365 518460 186943 518486
rect 172369 518458 172407 518460
rect 172369 518442 172435 518458
rect 172261 518402 172327 518418
rect 172261 518368 172277 518402
rect 172311 518368 172327 518402
rect 172369 518408 172385 518442
rect 172419 518408 172435 518442
rect 173057 518438 173511 518460
rect 172369 518392 172435 518408
rect 172565 518402 173015 518418
rect 172261 518352 172327 518368
rect 172289 518350 172327 518352
rect 172565 518368 172837 518402
rect 172871 518368 173015 518402
rect 173057 518404 173201 518438
rect 173235 518404 173511 518438
rect 174161 518438 174615 518460
rect 173057 518388 173511 518404
rect 173669 518402 174119 518418
rect 172289 518320 172407 518350
rect 172565 518346 173015 518368
rect 173669 518368 173941 518402
rect 173975 518368 174119 518402
rect 174161 518404 174305 518438
rect 174339 518404 174615 518438
rect 175449 518438 175903 518460
rect 174161 518388 174615 518404
rect 174957 518402 175407 518418
rect 173669 518346 174119 518368
rect 174957 518368 175229 518402
rect 175263 518368 175407 518402
rect 175449 518404 175593 518438
rect 175627 518404 175903 518438
rect 176553 518438 177007 518460
rect 175449 518388 175903 518404
rect 176061 518402 176511 518418
rect 174957 518346 175407 518368
rect 176061 518368 176333 518402
rect 176367 518368 176511 518402
rect 176553 518404 176697 518438
rect 176731 518404 177007 518438
rect 177657 518438 178111 518460
rect 176553 518388 177007 518404
rect 177165 518402 177615 518418
rect 176061 518346 176511 518368
rect 177165 518368 177437 518402
rect 177471 518368 177615 518402
rect 177657 518404 177801 518438
rect 177835 518404 178111 518438
rect 178761 518438 179215 518460
rect 177657 518388 178111 518404
rect 178269 518402 178719 518418
rect 177165 518346 177615 518368
rect 178269 518368 178541 518402
rect 178575 518368 178719 518402
rect 178761 518404 178905 518438
rect 178939 518404 179215 518438
rect 179591 518438 179767 518460
rect 178761 518388 179215 518404
rect 179373 518402 179549 518418
rect 178269 518346 178719 518368
rect 179373 518368 179389 518402
rect 179423 518368 179499 518402
rect 179533 518368 179549 518402
rect 179591 518404 179607 518438
rect 179641 518404 179717 518438
rect 179751 518404 179767 518438
rect 180601 518438 181055 518460
rect 179591 518388 179767 518404
rect 180109 518402 180559 518418
rect 179373 518346 179549 518368
rect 180109 518368 180381 518402
rect 180415 518368 180559 518402
rect 180601 518404 180745 518438
rect 180779 518404 181055 518438
rect 181705 518438 182159 518460
rect 180601 518388 181055 518404
rect 181213 518402 181663 518418
rect 180109 518346 180559 518368
rect 181213 518368 181485 518402
rect 181519 518368 181663 518402
rect 181705 518404 181849 518438
rect 181883 518404 182159 518438
rect 182809 518438 183263 518460
rect 181705 518388 182159 518404
rect 182317 518402 182767 518418
rect 181213 518346 181663 518368
rect 182317 518368 182589 518402
rect 182623 518368 182767 518402
rect 182809 518404 182953 518438
rect 182987 518404 183263 518438
rect 183913 518438 184367 518460
rect 182809 518388 183263 518404
rect 183421 518402 183871 518418
rect 182317 518346 182767 518368
rect 183421 518368 183693 518402
rect 183727 518368 183871 518402
rect 183913 518404 184057 518438
rect 184091 518404 184367 518438
rect 184743 518438 184919 518460
rect 183913 518388 184367 518404
rect 184525 518402 184701 518418
rect 183421 518346 183871 518368
rect 184525 518368 184541 518402
rect 184575 518368 184651 518402
rect 184685 518368 184701 518402
rect 184743 518404 184759 518438
rect 184793 518404 184869 518438
rect 184903 518404 184919 518438
rect 185753 518438 186207 518460
rect 184743 518388 184919 518404
rect 185261 518402 185711 518418
rect 184525 518346 184701 518368
rect 185261 518368 185533 518402
rect 185567 518368 185711 518402
rect 185753 518404 185897 518438
rect 185931 518404 186207 518438
rect 186671 518438 186943 518460
rect 187285 518460 187403 518486
rect 187285 518458 187323 518460
rect 185753 518388 186207 518404
rect 186365 518402 186629 518418
rect 185261 518346 185711 518368
rect 186365 518368 186381 518402
rect 186415 518368 186480 518402
rect 186514 518368 186579 518402
rect 186613 518368 186629 518402
rect 186671 518404 186687 518438
rect 186721 518404 186790 518438
rect 186824 518404 186893 518438
rect 186927 518404 186943 518438
rect 186671 518388 186943 518404
rect 187257 518442 187323 518458
rect 187257 518408 187273 518442
rect 187307 518408 187323 518442
rect 187257 518392 187323 518408
rect 187365 518402 187431 518418
rect 186365 518346 186629 518368
rect 187365 518368 187381 518402
rect 187415 518368 187431 518402
rect 187365 518352 187431 518368
rect 187365 518350 187403 518352
rect 172565 518320 173511 518346
rect 173669 518320 174615 518346
rect 174957 518320 175903 518346
rect 176061 518320 177007 518346
rect 177165 518320 178111 518346
rect 178269 518320 179215 518346
rect 179373 518320 179767 518346
rect 180109 518320 181055 518346
rect 181213 518320 182159 518346
rect 182317 518320 183263 518346
rect 183421 518320 184367 518346
rect 184525 518320 184919 518346
rect 185261 518320 186207 518346
rect 186365 518320 186943 518346
rect 187285 518320 187403 518350
rect 172289 518120 172407 518146
rect 172565 518120 173511 518146
rect 173669 518120 174615 518146
rect 174957 518120 175903 518146
rect 176061 518120 177007 518146
rect 177165 518120 178111 518146
rect 178269 518120 179215 518146
rect 179373 518120 179767 518146
rect 180109 518120 181055 518146
rect 181213 518120 182159 518146
rect 182317 518120 183263 518146
rect 183421 518120 184367 518146
rect 184525 518120 184919 518146
rect 185261 518120 186207 518146
rect 186365 518120 186943 518146
rect 187285 518120 187403 518146
rect 172289 518052 172407 518078
rect 172565 518052 173511 518078
rect 173669 518052 174615 518078
rect 174773 518052 175719 518078
rect 175877 518052 176823 518078
rect 176981 518052 177191 518078
rect 177533 518052 178479 518078
rect 178637 518052 179583 518078
rect 179741 518052 180687 518078
rect 180845 518052 181791 518078
rect 181949 518052 182343 518078
rect 182685 518052 183631 518078
rect 183789 518052 184735 518078
rect 184893 518052 185839 518078
rect 185997 518052 186943 518078
rect 187285 518052 187403 518078
rect 172289 517848 172407 517878
rect 172565 517852 173511 517878
rect 173669 517852 174615 517878
rect 174773 517852 175719 517878
rect 175877 517852 176823 517878
rect 176981 517852 177191 517878
rect 177533 517852 178479 517878
rect 178637 517852 179583 517878
rect 179741 517852 180687 517878
rect 180845 517852 181791 517878
rect 181949 517852 182343 517878
rect 182685 517852 183631 517878
rect 183789 517852 184735 517878
rect 184893 517852 185839 517878
rect 185997 517852 186943 517878
rect 172289 517846 172327 517848
rect 172261 517830 172327 517846
rect 172261 517796 172277 517830
rect 172311 517796 172327 517830
rect 172565 517830 173015 517852
rect 172261 517780 172327 517796
rect 172369 517790 172435 517806
rect 172369 517756 172385 517790
rect 172419 517756 172435 517790
rect 172565 517796 172837 517830
rect 172871 517796 173015 517830
rect 173669 517830 174119 517852
rect 172565 517780 173015 517796
rect 173057 517794 173511 517810
rect 172369 517740 172435 517756
rect 173057 517760 173201 517794
rect 173235 517760 173511 517794
rect 173669 517796 173941 517830
rect 173975 517796 174119 517830
rect 174773 517830 175223 517852
rect 173669 517780 174119 517796
rect 174161 517794 174615 517810
rect 172369 517738 172407 517740
rect 173057 517738 173511 517760
rect 174161 517760 174305 517794
rect 174339 517760 174615 517794
rect 174773 517796 175045 517830
rect 175079 517796 175223 517830
rect 175877 517830 176327 517852
rect 176981 517846 177065 517852
rect 174773 517780 175223 517796
rect 175265 517794 175719 517810
rect 174161 517738 174615 517760
rect 175265 517760 175409 517794
rect 175443 517760 175719 517794
rect 175877 517796 176149 517830
rect 176183 517796 176327 517830
rect 176923 517830 177065 517846
rect 175877 517780 176327 517796
rect 176369 517794 176823 517810
rect 175265 517738 175719 517760
rect 176369 517760 176513 517794
rect 176547 517760 176823 517794
rect 176923 517796 176939 517830
rect 176973 517796 177065 517830
rect 177533 517830 177983 517852
rect 176923 517780 177065 517796
rect 177107 517794 177249 517810
rect 176369 517738 176823 517760
rect 177107 517760 177199 517794
rect 177233 517760 177249 517794
rect 177533 517796 177805 517830
rect 177839 517796 177983 517830
rect 178637 517830 179087 517852
rect 177533 517780 177983 517796
rect 178025 517794 178479 517810
rect 177107 517744 177249 517760
rect 178025 517760 178169 517794
rect 178203 517760 178479 517794
rect 178637 517796 178909 517830
rect 178943 517796 179087 517830
rect 179741 517830 180191 517852
rect 178637 517780 179087 517796
rect 179129 517794 179583 517810
rect 177107 517738 177191 517744
rect 178025 517738 178479 517760
rect 179129 517760 179273 517794
rect 179307 517760 179583 517794
rect 179741 517796 180013 517830
rect 180047 517796 180191 517830
rect 180845 517830 181295 517852
rect 179741 517780 180191 517796
rect 180233 517794 180687 517810
rect 179129 517738 179583 517760
rect 180233 517760 180377 517794
rect 180411 517760 180687 517794
rect 180845 517796 181117 517830
rect 181151 517796 181295 517830
rect 181949 517830 182125 517852
rect 180845 517780 181295 517796
rect 181337 517794 181791 517810
rect 180233 517738 180687 517760
rect 181337 517760 181481 517794
rect 181515 517760 181791 517794
rect 181949 517796 181965 517830
rect 181999 517796 182075 517830
rect 182109 517796 182125 517830
rect 182685 517830 183135 517852
rect 181949 517780 182125 517796
rect 182167 517794 182343 517810
rect 181337 517738 181791 517760
rect 182167 517760 182183 517794
rect 182217 517760 182293 517794
rect 182327 517760 182343 517794
rect 182685 517796 182957 517830
rect 182991 517796 183135 517830
rect 183789 517830 184239 517852
rect 182685 517780 183135 517796
rect 183177 517794 183631 517810
rect 182167 517738 182343 517760
rect 183177 517760 183321 517794
rect 183355 517760 183631 517794
rect 183789 517796 184061 517830
rect 184095 517796 184239 517830
rect 184893 517830 185343 517852
rect 183789 517780 184239 517796
rect 184281 517794 184735 517810
rect 183177 517738 183631 517760
rect 184281 517760 184425 517794
rect 184459 517760 184735 517794
rect 184893 517796 185165 517830
rect 185199 517796 185343 517830
rect 185997 517830 186447 517852
rect 187285 517848 187403 517878
rect 184893 517780 185343 517796
rect 185385 517794 185839 517810
rect 184281 517738 184735 517760
rect 185385 517760 185529 517794
rect 185563 517760 185839 517794
rect 185997 517796 186269 517830
rect 186303 517796 186447 517830
rect 187365 517846 187403 517848
rect 187365 517830 187431 517846
rect 185997 517780 186447 517796
rect 186489 517794 186943 517810
rect 185385 517738 185839 517760
rect 186489 517760 186633 517794
rect 186667 517760 186943 517794
rect 186489 517738 186943 517760
rect 187257 517790 187323 517806
rect 187257 517756 187273 517790
rect 187307 517756 187323 517790
rect 187365 517796 187381 517830
rect 187415 517796 187431 517830
rect 187365 517780 187431 517796
rect 187257 517740 187323 517756
rect 172289 517712 172407 517738
rect 172565 517712 173511 517738
rect 173669 517712 174615 517738
rect 174773 517712 175719 517738
rect 175877 517712 176823 517738
rect 176981 517712 177191 517738
rect 177533 517712 178479 517738
rect 178637 517712 179583 517738
rect 179741 517712 180687 517738
rect 180845 517712 181791 517738
rect 181949 517712 182343 517738
rect 182685 517712 183631 517738
rect 183789 517712 184735 517738
rect 184893 517712 185839 517738
rect 185997 517712 186943 517738
rect 187285 517738 187323 517740
rect 187285 517712 187403 517738
rect 172289 517576 172407 517602
rect 172565 517576 173511 517602
rect 173669 517576 174615 517602
rect 174773 517576 175719 517602
rect 175877 517576 176823 517602
rect 176981 517576 177191 517602
rect 177533 517576 178479 517602
rect 178637 517576 179583 517602
rect 179741 517576 180687 517602
rect 180845 517576 181791 517602
rect 181949 517576 182343 517602
rect 182685 517576 183631 517602
rect 183789 517576 184735 517602
rect 184893 517576 185839 517602
rect 185997 517576 186943 517602
rect 187285 517576 187403 517602
rect 172289 517508 172407 517534
rect 172565 517508 173511 517534
rect 173669 517508 174615 517534
rect 174957 517508 175903 517534
rect 176061 517508 177007 517534
rect 177165 517508 178111 517534
rect 178269 517508 179215 517534
rect 179373 517508 179767 517534
rect 180109 517508 181055 517534
rect 181213 517508 182159 517534
rect 182317 517508 183263 517534
rect 183421 517508 184367 517534
rect 184525 517508 184919 517534
rect 185261 517508 186207 517534
rect 186365 517508 186943 517534
rect 187285 517508 187403 517534
rect 172289 517372 172407 517398
rect 172565 517372 173511 517398
rect 173669 517372 174615 517398
rect 174957 517372 175903 517398
rect 176061 517372 177007 517398
rect 177165 517372 178111 517398
rect 178269 517372 179215 517398
rect 179373 517372 179767 517398
rect 180109 517372 181055 517398
rect 181213 517372 182159 517398
rect 182317 517372 183263 517398
rect 183421 517372 184367 517398
rect 184525 517372 184919 517398
rect 185261 517372 186207 517398
rect 186365 517372 186943 517398
rect 172369 517370 172407 517372
rect 172369 517354 172435 517370
rect 172261 517314 172327 517330
rect 172261 517280 172277 517314
rect 172311 517280 172327 517314
rect 172369 517320 172385 517354
rect 172419 517320 172435 517354
rect 173057 517350 173511 517372
rect 172369 517304 172435 517320
rect 172565 517314 173015 517330
rect 172261 517264 172327 517280
rect 172289 517262 172327 517264
rect 172565 517280 172837 517314
rect 172871 517280 173015 517314
rect 173057 517316 173201 517350
rect 173235 517316 173511 517350
rect 174161 517350 174615 517372
rect 173057 517300 173511 517316
rect 173669 517314 174119 517330
rect 172289 517232 172407 517262
rect 172565 517258 173015 517280
rect 173669 517280 173941 517314
rect 173975 517280 174119 517314
rect 174161 517316 174305 517350
rect 174339 517316 174615 517350
rect 175449 517350 175903 517372
rect 174161 517300 174615 517316
rect 174957 517314 175407 517330
rect 173669 517258 174119 517280
rect 174957 517280 175229 517314
rect 175263 517280 175407 517314
rect 175449 517316 175593 517350
rect 175627 517316 175903 517350
rect 176553 517350 177007 517372
rect 175449 517300 175903 517316
rect 176061 517314 176511 517330
rect 174957 517258 175407 517280
rect 176061 517280 176333 517314
rect 176367 517280 176511 517314
rect 176553 517316 176697 517350
rect 176731 517316 177007 517350
rect 177657 517350 178111 517372
rect 176553 517300 177007 517316
rect 177165 517314 177615 517330
rect 176061 517258 176511 517280
rect 177165 517280 177437 517314
rect 177471 517280 177615 517314
rect 177657 517316 177801 517350
rect 177835 517316 178111 517350
rect 178761 517350 179215 517372
rect 177657 517300 178111 517316
rect 178269 517314 178719 517330
rect 177165 517258 177615 517280
rect 178269 517280 178541 517314
rect 178575 517280 178719 517314
rect 178761 517316 178905 517350
rect 178939 517316 179215 517350
rect 179591 517350 179767 517372
rect 178761 517300 179215 517316
rect 179373 517314 179549 517330
rect 178269 517258 178719 517280
rect 179373 517280 179389 517314
rect 179423 517280 179499 517314
rect 179533 517280 179549 517314
rect 179591 517316 179607 517350
rect 179641 517316 179717 517350
rect 179751 517316 179767 517350
rect 180601 517350 181055 517372
rect 179591 517300 179767 517316
rect 180109 517314 180559 517330
rect 179373 517258 179549 517280
rect 180109 517280 180381 517314
rect 180415 517280 180559 517314
rect 180601 517316 180745 517350
rect 180779 517316 181055 517350
rect 181705 517350 182159 517372
rect 180601 517300 181055 517316
rect 181213 517314 181663 517330
rect 180109 517258 180559 517280
rect 181213 517280 181485 517314
rect 181519 517280 181663 517314
rect 181705 517316 181849 517350
rect 181883 517316 182159 517350
rect 182809 517350 183263 517372
rect 181705 517300 182159 517316
rect 182317 517314 182767 517330
rect 181213 517258 181663 517280
rect 182317 517280 182589 517314
rect 182623 517280 182767 517314
rect 182809 517316 182953 517350
rect 182987 517316 183263 517350
rect 183913 517350 184367 517372
rect 182809 517300 183263 517316
rect 183421 517314 183871 517330
rect 182317 517258 182767 517280
rect 183421 517280 183693 517314
rect 183727 517280 183871 517314
rect 183913 517316 184057 517350
rect 184091 517316 184367 517350
rect 184743 517350 184919 517372
rect 183913 517300 184367 517316
rect 184525 517314 184701 517330
rect 183421 517258 183871 517280
rect 184525 517280 184541 517314
rect 184575 517280 184651 517314
rect 184685 517280 184701 517314
rect 184743 517316 184759 517350
rect 184793 517316 184869 517350
rect 184903 517316 184919 517350
rect 185753 517350 186207 517372
rect 184743 517300 184919 517316
rect 185261 517314 185711 517330
rect 184525 517258 184701 517280
rect 185261 517280 185533 517314
rect 185567 517280 185711 517314
rect 185753 517316 185897 517350
rect 185931 517316 186207 517350
rect 186671 517350 186943 517372
rect 187285 517372 187403 517398
rect 187285 517370 187323 517372
rect 185753 517300 186207 517316
rect 186365 517314 186629 517330
rect 185261 517258 185711 517280
rect 186365 517280 186381 517314
rect 186415 517280 186480 517314
rect 186514 517280 186579 517314
rect 186613 517280 186629 517314
rect 186671 517316 186687 517350
rect 186721 517316 186790 517350
rect 186824 517316 186893 517350
rect 186927 517316 186943 517350
rect 186671 517300 186943 517316
rect 187257 517354 187323 517370
rect 187257 517320 187273 517354
rect 187307 517320 187323 517354
rect 187257 517304 187323 517320
rect 187365 517314 187431 517330
rect 186365 517258 186629 517280
rect 187365 517280 187381 517314
rect 187415 517280 187431 517314
rect 187365 517264 187431 517280
rect 187365 517262 187403 517264
rect 172565 517232 173511 517258
rect 173669 517232 174615 517258
rect 174957 517232 175903 517258
rect 176061 517232 177007 517258
rect 177165 517232 178111 517258
rect 178269 517232 179215 517258
rect 179373 517232 179767 517258
rect 180109 517232 181055 517258
rect 181213 517232 182159 517258
rect 182317 517232 183263 517258
rect 183421 517232 184367 517258
rect 184525 517232 184919 517258
rect 185261 517232 186207 517258
rect 186365 517232 186943 517258
rect 187285 517232 187403 517262
rect 172289 517032 172407 517058
rect 172565 517032 173511 517058
rect 173669 517032 174615 517058
rect 174957 517032 175903 517058
rect 176061 517032 177007 517058
rect 177165 517032 178111 517058
rect 178269 517032 179215 517058
rect 179373 517032 179767 517058
rect 180109 517032 181055 517058
rect 181213 517032 182159 517058
rect 182317 517032 183263 517058
rect 183421 517032 184367 517058
rect 184525 517032 184919 517058
rect 185261 517032 186207 517058
rect 186365 517032 186943 517058
rect 187285 517032 187403 517058
rect 172289 516964 172407 516990
rect 172565 516964 173511 516990
rect 173669 516964 174615 516990
rect 174773 516964 175719 516990
rect 175877 516964 176823 516990
rect 176981 516964 177191 516990
rect 177533 516964 178479 516990
rect 178637 516964 179583 516990
rect 179741 516964 180687 516990
rect 180845 516964 181791 516990
rect 181949 516964 182343 516990
rect 182685 516964 183631 516990
rect 183789 516964 184735 516990
rect 184893 516964 185839 516990
rect 185997 516964 186943 516990
rect 187285 516964 187403 516990
rect 172289 516760 172407 516790
rect 172565 516764 173511 516790
rect 173669 516764 174615 516790
rect 174773 516764 175719 516790
rect 175877 516764 176823 516790
rect 176981 516764 177191 516790
rect 177533 516764 178479 516790
rect 178637 516764 179583 516790
rect 179741 516764 180687 516790
rect 180845 516764 181791 516790
rect 181949 516764 182343 516790
rect 182685 516764 183631 516790
rect 183789 516764 184735 516790
rect 184893 516764 185839 516790
rect 185997 516764 186943 516790
rect 172289 516758 172327 516760
rect 172261 516742 172327 516758
rect 172261 516708 172277 516742
rect 172311 516708 172327 516742
rect 172565 516742 173015 516764
rect 172261 516692 172327 516708
rect 172369 516702 172435 516718
rect 172369 516668 172385 516702
rect 172419 516668 172435 516702
rect 172565 516708 172837 516742
rect 172871 516708 173015 516742
rect 173669 516742 174119 516764
rect 172565 516692 173015 516708
rect 173057 516706 173511 516722
rect 172369 516652 172435 516668
rect 173057 516672 173201 516706
rect 173235 516672 173511 516706
rect 173669 516708 173941 516742
rect 173975 516708 174119 516742
rect 174773 516742 175223 516764
rect 173669 516692 174119 516708
rect 174161 516706 174615 516722
rect 172369 516650 172407 516652
rect 173057 516650 173511 516672
rect 174161 516672 174305 516706
rect 174339 516672 174615 516706
rect 174773 516708 175045 516742
rect 175079 516708 175223 516742
rect 175877 516742 176327 516764
rect 176981 516758 177065 516764
rect 174773 516692 175223 516708
rect 175265 516706 175719 516722
rect 174161 516650 174615 516672
rect 175265 516672 175409 516706
rect 175443 516672 175719 516706
rect 175877 516708 176149 516742
rect 176183 516708 176327 516742
rect 176923 516742 177065 516758
rect 175877 516692 176327 516708
rect 176369 516706 176823 516722
rect 175265 516650 175719 516672
rect 176369 516672 176513 516706
rect 176547 516672 176823 516706
rect 176923 516708 176939 516742
rect 176973 516708 177065 516742
rect 177533 516742 177983 516764
rect 176923 516692 177065 516708
rect 177107 516706 177249 516722
rect 176369 516650 176823 516672
rect 177107 516672 177199 516706
rect 177233 516672 177249 516706
rect 177533 516708 177805 516742
rect 177839 516708 177983 516742
rect 178637 516742 179087 516764
rect 177533 516692 177983 516708
rect 178025 516706 178479 516722
rect 177107 516656 177249 516672
rect 178025 516672 178169 516706
rect 178203 516672 178479 516706
rect 178637 516708 178909 516742
rect 178943 516708 179087 516742
rect 179741 516742 180191 516764
rect 178637 516692 179087 516708
rect 179129 516706 179583 516722
rect 177107 516650 177191 516656
rect 178025 516650 178479 516672
rect 179129 516672 179273 516706
rect 179307 516672 179583 516706
rect 179741 516708 180013 516742
rect 180047 516708 180191 516742
rect 180845 516742 181295 516764
rect 179741 516692 180191 516708
rect 180233 516706 180687 516722
rect 179129 516650 179583 516672
rect 180233 516672 180377 516706
rect 180411 516672 180687 516706
rect 180845 516708 181117 516742
rect 181151 516708 181295 516742
rect 181949 516742 182125 516764
rect 180845 516692 181295 516708
rect 181337 516706 181791 516722
rect 180233 516650 180687 516672
rect 181337 516672 181481 516706
rect 181515 516672 181791 516706
rect 181949 516708 181965 516742
rect 181999 516708 182075 516742
rect 182109 516708 182125 516742
rect 182685 516742 183135 516764
rect 181949 516692 182125 516708
rect 182167 516706 182343 516722
rect 181337 516650 181791 516672
rect 182167 516672 182183 516706
rect 182217 516672 182293 516706
rect 182327 516672 182343 516706
rect 182685 516708 182957 516742
rect 182991 516708 183135 516742
rect 183789 516742 184239 516764
rect 182685 516692 183135 516708
rect 183177 516706 183631 516722
rect 182167 516650 182343 516672
rect 183177 516672 183321 516706
rect 183355 516672 183631 516706
rect 183789 516708 184061 516742
rect 184095 516708 184239 516742
rect 184893 516742 185343 516764
rect 183789 516692 184239 516708
rect 184281 516706 184735 516722
rect 183177 516650 183631 516672
rect 184281 516672 184425 516706
rect 184459 516672 184735 516706
rect 184893 516708 185165 516742
rect 185199 516708 185343 516742
rect 185997 516742 186447 516764
rect 187285 516760 187403 516790
rect 184893 516692 185343 516708
rect 185385 516706 185839 516722
rect 184281 516650 184735 516672
rect 185385 516672 185529 516706
rect 185563 516672 185839 516706
rect 185997 516708 186269 516742
rect 186303 516708 186447 516742
rect 187365 516758 187403 516760
rect 187365 516742 187431 516758
rect 185997 516692 186447 516708
rect 186489 516706 186943 516722
rect 185385 516650 185839 516672
rect 186489 516672 186633 516706
rect 186667 516672 186943 516706
rect 186489 516650 186943 516672
rect 187257 516702 187323 516718
rect 187257 516668 187273 516702
rect 187307 516668 187323 516702
rect 187365 516708 187381 516742
rect 187415 516708 187431 516742
rect 187365 516692 187431 516708
rect 187257 516652 187323 516668
rect 172289 516624 172407 516650
rect 172565 516624 173511 516650
rect 173669 516624 174615 516650
rect 174773 516624 175719 516650
rect 175877 516624 176823 516650
rect 176981 516624 177191 516650
rect 177533 516624 178479 516650
rect 178637 516624 179583 516650
rect 179741 516624 180687 516650
rect 180845 516624 181791 516650
rect 181949 516624 182343 516650
rect 182685 516624 183631 516650
rect 183789 516624 184735 516650
rect 184893 516624 185839 516650
rect 185997 516624 186943 516650
rect 187285 516650 187323 516652
rect 187285 516624 187403 516650
rect 172289 516488 172407 516514
rect 172565 516488 173511 516514
rect 173669 516488 174615 516514
rect 174773 516488 175719 516514
rect 175877 516488 176823 516514
rect 176981 516488 177191 516514
rect 177533 516488 178479 516514
rect 178637 516488 179583 516514
rect 179741 516488 180687 516514
rect 180845 516488 181791 516514
rect 181949 516488 182343 516514
rect 182685 516488 183631 516514
rect 183789 516488 184735 516514
rect 184893 516488 185839 516514
rect 185997 516488 186943 516514
rect 187285 516488 187403 516514
rect 172289 516420 172407 516446
rect 172565 516420 173511 516446
rect 173669 516420 174615 516446
rect 174957 516420 175903 516446
rect 176061 516420 177007 516446
rect 177165 516420 178111 516446
rect 178269 516420 179215 516446
rect 179373 516420 179767 516446
rect 180109 516420 181055 516446
rect 181213 516420 182159 516446
rect 182317 516420 183263 516446
rect 183421 516420 184367 516446
rect 184525 516420 184919 516446
rect 185261 516420 186207 516446
rect 186365 516420 186943 516446
rect 187285 516420 187403 516446
rect 172289 516284 172407 516310
rect 172565 516284 173511 516310
rect 173669 516284 174615 516310
rect 174957 516284 175903 516310
rect 176061 516284 177007 516310
rect 177165 516284 178111 516310
rect 178269 516284 179215 516310
rect 179373 516284 179767 516310
rect 180109 516284 181055 516310
rect 181213 516284 182159 516310
rect 182317 516284 183263 516310
rect 183421 516284 184367 516310
rect 184525 516284 184919 516310
rect 185261 516284 186207 516310
rect 186365 516284 186943 516310
rect 172369 516282 172407 516284
rect 172369 516266 172435 516282
rect 172261 516226 172327 516242
rect 172261 516192 172277 516226
rect 172311 516192 172327 516226
rect 172369 516232 172385 516266
rect 172419 516232 172435 516266
rect 173057 516262 173511 516284
rect 172369 516216 172435 516232
rect 172565 516226 173015 516242
rect 172261 516176 172327 516192
rect 172289 516174 172327 516176
rect 172565 516192 172837 516226
rect 172871 516192 173015 516226
rect 173057 516228 173201 516262
rect 173235 516228 173511 516262
rect 174161 516262 174615 516284
rect 173057 516212 173511 516228
rect 173669 516226 174119 516242
rect 172289 516144 172407 516174
rect 172565 516170 173015 516192
rect 173669 516192 173941 516226
rect 173975 516192 174119 516226
rect 174161 516228 174305 516262
rect 174339 516228 174615 516262
rect 175449 516262 175903 516284
rect 174161 516212 174615 516228
rect 174957 516226 175407 516242
rect 173669 516170 174119 516192
rect 174957 516192 175229 516226
rect 175263 516192 175407 516226
rect 175449 516228 175593 516262
rect 175627 516228 175903 516262
rect 176553 516262 177007 516284
rect 175449 516212 175903 516228
rect 176061 516226 176511 516242
rect 174957 516170 175407 516192
rect 176061 516192 176333 516226
rect 176367 516192 176511 516226
rect 176553 516228 176697 516262
rect 176731 516228 177007 516262
rect 177657 516262 178111 516284
rect 176553 516212 177007 516228
rect 177165 516226 177615 516242
rect 176061 516170 176511 516192
rect 177165 516192 177437 516226
rect 177471 516192 177615 516226
rect 177657 516228 177801 516262
rect 177835 516228 178111 516262
rect 178761 516262 179215 516284
rect 177657 516212 178111 516228
rect 178269 516226 178719 516242
rect 177165 516170 177615 516192
rect 178269 516192 178541 516226
rect 178575 516192 178719 516226
rect 178761 516228 178905 516262
rect 178939 516228 179215 516262
rect 179591 516262 179767 516284
rect 178761 516212 179215 516228
rect 179373 516226 179549 516242
rect 178269 516170 178719 516192
rect 179373 516192 179389 516226
rect 179423 516192 179499 516226
rect 179533 516192 179549 516226
rect 179591 516228 179607 516262
rect 179641 516228 179717 516262
rect 179751 516228 179767 516262
rect 180601 516262 181055 516284
rect 179591 516212 179767 516228
rect 180109 516226 180559 516242
rect 179373 516170 179549 516192
rect 180109 516192 180381 516226
rect 180415 516192 180559 516226
rect 180601 516228 180745 516262
rect 180779 516228 181055 516262
rect 181705 516262 182159 516284
rect 180601 516212 181055 516228
rect 181213 516226 181663 516242
rect 180109 516170 180559 516192
rect 181213 516192 181485 516226
rect 181519 516192 181663 516226
rect 181705 516228 181849 516262
rect 181883 516228 182159 516262
rect 182809 516262 183263 516284
rect 181705 516212 182159 516228
rect 182317 516226 182767 516242
rect 181213 516170 181663 516192
rect 182317 516192 182589 516226
rect 182623 516192 182767 516226
rect 182809 516228 182953 516262
rect 182987 516228 183263 516262
rect 183913 516262 184367 516284
rect 182809 516212 183263 516228
rect 183421 516226 183871 516242
rect 182317 516170 182767 516192
rect 183421 516192 183693 516226
rect 183727 516192 183871 516226
rect 183913 516228 184057 516262
rect 184091 516228 184367 516262
rect 184743 516262 184919 516284
rect 183913 516212 184367 516228
rect 184525 516226 184701 516242
rect 183421 516170 183871 516192
rect 184525 516192 184541 516226
rect 184575 516192 184651 516226
rect 184685 516192 184701 516226
rect 184743 516228 184759 516262
rect 184793 516228 184869 516262
rect 184903 516228 184919 516262
rect 185753 516262 186207 516284
rect 184743 516212 184919 516228
rect 185261 516226 185711 516242
rect 184525 516170 184701 516192
rect 185261 516192 185533 516226
rect 185567 516192 185711 516226
rect 185753 516228 185897 516262
rect 185931 516228 186207 516262
rect 186671 516262 186943 516284
rect 187285 516284 187403 516310
rect 187285 516282 187323 516284
rect 185753 516212 186207 516228
rect 186365 516226 186629 516242
rect 185261 516170 185711 516192
rect 186365 516192 186381 516226
rect 186415 516192 186480 516226
rect 186514 516192 186579 516226
rect 186613 516192 186629 516226
rect 186671 516228 186687 516262
rect 186721 516228 186790 516262
rect 186824 516228 186893 516262
rect 186927 516228 186943 516262
rect 186671 516212 186943 516228
rect 187257 516266 187323 516282
rect 187257 516232 187273 516266
rect 187307 516232 187323 516266
rect 187257 516216 187323 516232
rect 187365 516226 187431 516242
rect 186365 516170 186629 516192
rect 187365 516192 187381 516226
rect 187415 516192 187431 516226
rect 187365 516176 187431 516192
rect 187365 516174 187403 516176
rect 172565 516144 173511 516170
rect 173669 516144 174615 516170
rect 174957 516144 175903 516170
rect 176061 516144 177007 516170
rect 177165 516144 178111 516170
rect 178269 516144 179215 516170
rect 179373 516144 179767 516170
rect 180109 516144 181055 516170
rect 181213 516144 182159 516170
rect 182317 516144 183263 516170
rect 183421 516144 184367 516170
rect 184525 516144 184919 516170
rect 185261 516144 186207 516170
rect 186365 516144 186943 516170
rect 187285 516144 187403 516174
rect 172289 515944 172407 515970
rect 172565 515944 173511 515970
rect 173669 515944 174615 515970
rect 174957 515944 175903 515970
rect 176061 515944 177007 515970
rect 177165 515944 178111 515970
rect 178269 515944 179215 515970
rect 179373 515944 179767 515970
rect 180109 515944 181055 515970
rect 181213 515944 182159 515970
rect 182317 515944 183263 515970
rect 183421 515944 184367 515970
rect 184525 515944 184919 515970
rect 185261 515944 186207 515970
rect 186365 515944 186943 515970
rect 187285 515944 187403 515970
rect 172289 515876 172407 515902
rect 172565 515876 173143 515902
rect 173486 515876 173516 515902
rect 173582 515876 173612 515902
rect 173668 515876 173698 515902
rect 173754 515876 173784 515902
rect 173840 515876 173870 515902
rect 174037 515876 174615 515902
rect 174957 515876 175903 515902
rect 176061 515876 177007 515902
rect 177165 515876 177283 515902
rect 177533 515876 178479 515902
rect 178637 515876 179583 515902
rect 179741 515876 179859 515902
rect 180109 515876 181055 515902
rect 181213 515876 181791 515902
rect 182133 515876 182163 515902
rect 182221 515876 182251 515902
rect 182685 515876 183631 515902
rect 183789 515876 184735 515902
rect 184893 515876 185011 515902
rect 185261 515876 186207 515902
rect 186458 515876 186488 515902
rect 186554 515876 186584 515902
rect 186640 515876 186670 515902
rect 186726 515876 186756 515902
rect 186812 515876 186842 515902
rect 187009 515876 187127 515902
rect 187285 515876 187403 515902
rect 172289 515672 172407 515702
rect 172565 515676 173143 515702
rect 174037 515676 174615 515702
rect 174957 515676 175903 515702
rect 176061 515676 177007 515702
rect 172289 515670 172327 515672
rect 172261 515654 172327 515670
rect 172261 515620 172277 515654
rect 172311 515620 172327 515654
rect 172565 515654 172829 515676
rect 172261 515604 172327 515620
rect 172369 515614 172435 515630
rect 172369 515580 172385 515614
rect 172419 515580 172435 515614
rect 172565 515620 172581 515654
rect 172615 515620 172680 515654
rect 172714 515620 172779 515654
rect 172813 515620 172829 515654
rect 173486 515644 173516 515676
rect 172565 515604 172829 515620
rect 172871 515618 173143 515634
rect 172369 515564 172435 515580
rect 172871 515584 172887 515618
rect 172921 515584 172990 515618
rect 173024 515584 173093 515618
rect 173127 515584 173143 515618
rect 172369 515562 172407 515564
rect 172871 515562 173143 515584
rect 173475 515628 173535 515644
rect 173475 515594 173491 515628
rect 173525 515594 173535 515628
rect 173475 515578 173535 515594
rect 173582 515638 173612 515676
rect 173668 515638 173698 515676
rect 173754 515638 173784 515676
rect 173840 515638 173870 515676
rect 173582 515628 173870 515638
rect 173582 515594 173637 515628
rect 173671 515594 173705 515628
rect 173739 515594 173773 515628
rect 173807 515616 173870 515628
rect 174037 515654 174301 515676
rect 174037 515620 174053 515654
rect 174087 515620 174152 515654
rect 174186 515620 174251 515654
rect 174285 515620 174301 515654
rect 174957 515654 175407 515676
rect 173807 515594 173871 515616
rect 174037 515604 174301 515620
rect 174343 515618 174615 515634
rect 173582 515589 173871 515594
rect 173583 515583 173871 515589
rect 172289 515536 172407 515562
rect 172565 515536 173143 515562
rect 173486 515510 173516 515578
rect 173583 515510 173613 515583
rect 173669 515510 173699 515583
rect 173755 515510 173785 515583
rect 173841 515510 173871 515583
rect 174343 515584 174359 515618
rect 174393 515584 174462 515618
rect 174496 515584 174565 515618
rect 174599 515584 174615 515618
rect 174957 515620 175229 515654
rect 175263 515620 175407 515654
rect 176061 515654 176511 515676
rect 177165 515672 177283 515702
rect 177533 515676 178479 515702
rect 178637 515676 179583 515702
rect 177165 515670 177203 515672
rect 174957 515604 175407 515620
rect 175449 515618 175903 515634
rect 174343 515562 174615 515584
rect 175449 515584 175593 515618
rect 175627 515584 175903 515618
rect 176061 515620 176333 515654
rect 176367 515620 176511 515654
rect 177137 515654 177203 515670
rect 176061 515604 176511 515620
rect 176553 515618 177007 515634
rect 175449 515562 175903 515584
rect 176553 515584 176697 515618
rect 176731 515584 177007 515618
rect 177137 515620 177153 515654
rect 177187 515620 177203 515654
rect 177533 515654 177983 515676
rect 177137 515604 177203 515620
rect 177245 515614 177311 515630
rect 176553 515562 177007 515584
rect 177245 515580 177261 515614
rect 177295 515580 177311 515614
rect 177533 515620 177805 515654
rect 177839 515620 177983 515654
rect 178637 515654 179087 515676
rect 179741 515672 179859 515702
rect 180109 515676 181055 515702
rect 181213 515676 181791 515702
rect 179741 515670 179779 515672
rect 177533 515604 177983 515620
rect 178025 515618 178479 515634
rect 177245 515564 177311 515580
rect 178025 515584 178169 515618
rect 178203 515584 178479 515618
rect 178637 515620 178909 515654
rect 178943 515620 179087 515654
rect 179713 515654 179779 515670
rect 178637 515604 179087 515620
rect 179129 515618 179583 515634
rect 177245 515562 177283 515564
rect 178025 515562 178479 515584
rect 179129 515584 179273 515618
rect 179307 515584 179583 515618
rect 179713 515620 179729 515654
rect 179763 515620 179779 515654
rect 180109 515654 180559 515676
rect 179713 515604 179779 515620
rect 179821 515614 179887 515630
rect 179129 515562 179583 515584
rect 179821 515580 179837 515614
rect 179871 515580 179887 515614
rect 180109 515620 180381 515654
rect 180415 515620 180559 515654
rect 181213 515654 181477 515676
rect 182133 515657 182163 515718
rect 182221 515703 182251 515718
rect 182221 515679 182257 515703
rect 180109 515604 180559 515620
rect 180601 515618 181055 515634
rect 179821 515564 179887 515580
rect 180601 515584 180745 515618
rect 180779 515584 181055 515618
rect 181213 515620 181229 515654
rect 181263 515620 181328 515654
rect 181362 515620 181427 515654
rect 181461 515620 181477 515654
rect 182131 515641 182185 515657
rect 181213 515604 181477 515620
rect 181519 515618 181791 515634
rect 179821 515562 179859 515564
rect 180601 515562 181055 515584
rect 181519 515584 181535 515618
rect 181569 515584 181638 515618
rect 181672 515584 181741 515618
rect 181775 515584 181791 515618
rect 182131 515607 182141 515641
rect 182175 515607 182185 515641
rect 182131 515591 182185 515607
rect 182227 515644 182257 515679
rect 182685 515676 183631 515702
rect 183789 515676 184735 515702
rect 182685 515654 183135 515676
rect 182227 515628 182303 515644
rect 182227 515594 182259 515628
rect 182293 515594 182303 515628
rect 182685 515620 182957 515654
rect 182991 515620 183135 515654
rect 183789 515654 184239 515676
rect 184893 515672 185011 515702
rect 185261 515676 186207 515702
rect 184893 515670 184931 515672
rect 182685 515604 183135 515620
rect 183177 515618 183631 515634
rect 181519 515562 181791 515584
rect 174037 515536 174615 515562
rect 174957 515536 175903 515562
rect 176061 515536 177007 515562
rect 177165 515536 177283 515562
rect 177533 515536 178479 515562
rect 178637 515536 179583 515562
rect 179741 515536 179859 515562
rect 180109 515536 181055 515562
rect 181213 515536 181791 515562
rect 182133 515530 182163 515591
rect 182227 515578 182303 515594
rect 183177 515584 183321 515618
rect 183355 515584 183631 515618
rect 183789 515620 184061 515654
rect 184095 515620 184239 515654
rect 184865 515654 184931 515670
rect 183789 515604 184239 515620
rect 184281 515618 184735 515634
rect 182227 515569 182257 515578
rect 182221 515545 182257 515569
rect 183177 515562 183631 515584
rect 184281 515584 184425 515618
rect 184459 515584 184735 515618
rect 184865 515620 184881 515654
rect 184915 515620 184931 515654
rect 185261 515654 185711 515676
rect 184865 515604 184931 515620
rect 184973 515614 185039 515630
rect 184281 515562 184735 515584
rect 184973 515580 184989 515614
rect 185023 515580 185039 515614
rect 185261 515620 185533 515654
rect 185567 515620 185711 515654
rect 186458 515644 186488 515676
rect 185261 515604 185711 515620
rect 185753 515618 186207 515634
rect 184973 515564 185039 515580
rect 185753 515584 185897 515618
rect 185931 515584 186207 515618
rect 184973 515562 185011 515564
rect 185753 515562 186207 515584
rect 186447 515628 186507 515644
rect 186447 515594 186463 515628
rect 186497 515594 186507 515628
rect 186447 515578 186507 515594
rect 186554 515638 186584 515676
rect 186640 515638 186670 515676
rect 186726 515638 186756 515676
rect 186812 515638 186842 515676
rect 187009 515672 187127 515702
rect 187285 515672 187403 515702
rect 187009 515670 187047 515672
rect 186554 515628 186842 515638
rect 186554 515594 186609 515628
rect 186643 515594 186677 515628
rect 186711 515594 186745 515628
rect 186779 515616 186842 515628
rect 186981 515654 187047 515670
rect 186981 515620 186997 515654
rect 187031 515620 187047 515654
rect 187365 515670 187403 515672
rect 187365 515654 187431 515670
rect 186779 515594 186843 515616
rect 186981 515604 187047 515620
rect 187089 515614 187155 515630
rect 186554 515589 186843 515594
rect 186555 515583 186843 515589
rect 182221 515530 182251 515545
rect 182685 515536 183631 515562
rect 183789 515536 184735 515562
rect 184893 515536 185011 515562
rect 185261 515536 186207 515562
rect 186458 515510 186488 515578
rect 186555 515510 186585 515583
rect 186641 515510 186671 515583
rect 186727 515510 186757 515583
rect 186813 515510 186843 515583
rect 187089 515580 187105 515614
rect 187139 515580 187155 515614
rect 187089 515564 187155 515580
rect 187257 515614 187323 515630
rect 187257 515580 187273 515614
rect 187307 515580 187323 515614
rect 187365 515620 187381 515654
rect 187415 515620 187431 515654
rect 187365 515604 187431 515620
rect 187257 515564 187323 515580
rect 187089 515562 187127 515564
rect 187009 515536 187127 515562
rect 187285 515562 187323 515564
rect 187285 515536 187403 515562
rect 172289 515400 172407 515426
rect 172565 515400 173143 515426
rect 173486 515400 173516 515426
rect 173583 515400 173613 515426
rect 173669 515400 173699 515426
rect 173755 515400 173785 515426
rect 173841 515400 173871 515426
rect 174037 515400 174615 515426
rect 174957 515400 175903 515426
rect 176061 515400 177007 515426
rect 177165 515400 177283 515426
rect 177533 515400 178479 515426
rect 178637 515400 179583 515426
rect 179741 515400 179859 515426
rect 180109 515400 181055 515426
rect 181213 515400 181791 515426
rect 182133 515400 182163 515426
rect 182221 515400 182251 515426
rect 182685 515400 183631 515426
rect 183789 515400 184735 515426
rect 184893 515400 185011 515426
rect 185261 515400 186207 515426
rect 186458 515400 186488 515426
rect 186555 515400 186585 515426
rect 186641 515400 186671 515426
rect 186727 515400 186757 515426
rect 186813 515400 186843 515426
rect 187009 515400 187127 515426
rect 187285 515400 187403 515426
<< polycont >>
rect 164730 541117 164764 541151
rect 165033 541124 165067 541158
rect 165225 541124 165259 541158
rect 165417 541124 165451 541158
rect 165609 541124 165643 541158
rect 165801 541124 165835 541158
rect 165993 541124 166027 541158
rect 166410 541117 166444 541151
rect 166210 540317 166244 540351
rect 164730 540007 164764 540041
rect 164937 540014 164971 540048
rect 165129 540014 165163 540048
rect 165321 540014 165355 540048
rect 165513 540014 165547 540048
rect 165705 540014 165739 540048
rect 165897 540014 165931 540048
rect 166210 540007 166244 540041
rect 166410 540007 166444 540041
rect 168530 541117 168564 541151
rect 168833 541124 168867 541158
rect 169025 541124 169059 541158
rect 169217 541124 169251 541158
rect 169409 541124 169443 541158
rect 169601 541124 169635 541158
rect 169793 541124 169827 541158
rect 170210 541117 170244 541151
rect 170010 540317 170044 540351
rect 168530 540007 168564 540041
rect 168737 540014 168771 540048
rect 168929 540014 168963 540048
rect 169121 540014 169155 540048
rect 169313 540014 169347 540048
rect 169505 540014 169539 540048
rect 169697 540014 169731 540048
rect 170010 540007 170044 540041
rect 170210 540007 170244 540041
rect 172230 541117 172264 541151
rect 172533 541124 172567 541158
rect 172725 541124 172759 541158
rect 172917 541124 172951 541158
rect 173109 541124 173143 541158
rect 173301 541124 173335 541158
rect 173493 541124 173527 541158
rect 173910 541117 173944 541151
rect 173710 540317 173744 540351
rect 172230 540007 172264 540041
rect 172437 540014 172471 540048
rect 172629 540014 172663 540048
rect 172821 540014 172855 540048
rect 173013 540014 173047 540048
rect 173205 540014 173239 540048
rect 173397 540014 173431 540048
rect 173710 540007 173744 540041
rect 173910 540007 173944 540041
rect 175730 541117 175764 541151
rect 176033 541124 176067 541158
rect 176225 541124 176259 541158
rect 176417 541124 176451 541158
rect 176609 541124 176643 541158
rect 176801 541124 176835 541158
rect 176993 541124 177027 541158
rect 177410 541117 177444 541151
rect 177210 540317 177244 540351
rect 175730 540007 175764 540041
rect 175937 540014 175971 540048
rect 176129 540014 176163 540048
rect 176321 540014 176355 540048
rect 176513 540014 176547 540048
rect 176705 540014 176739 540048
rect 176897 540014 176931 540048
rect 177210 540007 177244 540041
rect 177410 540007 177444 540041
rect 179330 541117 179364 541151
rect 179633 541124 179667 541158
rect 179825 541124 179859 541158
rect 180017 541124 180051 541158
rect 180209 541124 180243 541158
rect 180401 541124 180435 541158
rect 180593 541124 180627 541158
rect 181010 541117 181044 541151
rect 180810 540317 180844 540351
rect 179330 540007 179364 540041
rect 179537 540014 179571 540048
rect 179729 540014 179763 540048
rect 179921 540014 179955 540048
rect 180113 540014 180147 540048
rect 180305 540014 180339 540048
rect 180497 540014 180531 540048
rect 180810 540007 180844 540041
rect 181010 540007 181044 540041
rect 182630 541117 182664 541151
rect 182933 541124 182967 541158
rect 183125 541124 183159 541158
rect 183317 541124 183351 541158
rect 183509 541124 183543 541158
rect 183701 541124 183735 541158
rect 183893 541124 183927 541158
rect 184310 541117 184344 541151
rect 184110 540317 184144 540351
rect 182630 540007 182664 540041
rect 182837 540014 182871 540048
rect 183029 540014 183063 540048
rect 183221 540014 183255 540048
rect 183413 540014 183447 540048
rect 183605 540014 183639 540048
rect 183797 540014 183831 540048
rect 184110 540007 184144 540041
rect 184310 540007 184344 540041
rect 185930 541117 185964 541151
rect 186233 541124 186267 541158
rect 186425 541124 186459 541158
rect 186617 541124 186651 541158
rect 186809 541124 186843 541158
rect 187001 541124 187035 541158
rect 187193 541124 187227 541158
rect 187610 541117 187644 541151
rect 187410 540317 187444 540351
rect 185930 540007 185964 540041
rect 186137 540014 186171 540048
rect 186329 540014 186363 540048
rect 186521 540014 186555 540048
rect 186713 540014 186747 540048
rect 186905 540014 186939 540048
rect 187097 540014 187131 540048
rect 187410 540007 187444 540041
rect 187610 540007 187644 540041
rect 189230 541117 189264 541151
rect 189533 541124 189567 541158
rect 189725 541124 189759 541158
rect 189917 541124 189951 541158
rect 190109 541124 190143 541158
rect 190301 541124 190335 541158
rect 190493 541124 190527 541158
rect 190910 541117 190944 541151
rect 190710 540317 190744 540351
rect 189230 540007 189264 540041
rect 189437 540014 189471 540048
rect 189629 540014 189663 540048
rect 189821 540014 189855 540048
rect 190013 540014 190047 540048
rect 190205 540014 190239 540048
rect 190397 540014 190431 540048
rect 190710 540007 190744 540041
rect 190910 540007 190944 540041
rect 158728 538467 158896 538501
rect 159104 538467 159272 538501
rect 159362 538467 159530 538501
rect 159620 538467 159788 538501
rect 159878 538467 160046 538501
rect 160136 538467 160304 538501
rect 160394 538467 160562 538501
rect 160652 538467 160820 538501
rect 160910 538467 161078 538501
rect 161168 538467 161336 538501
rect 161548 538467 161716 538501
rect 161948 538467 162116 538501
rect 162328 538467 162496 538501
rect 158728 538157 158896 538191
rect 159104 538157 159272 538191
rect 159362 538157 159530 538191
rect 159620 538157 159788 538191
rect 159878 538157 160046 538191
rect 160136 538157 160304 538191
rect 160394 538157 160562 538191
rect 160652 538157 160820 538191
rect 160910 538157 161078 538191
rect 161168 538157 161336 538191
rect 161548 538157 161716 538191
rect 161948 538157 162116 538191
rect 162328 538157 162496 538191
rect 164714 539604 164748 539638
rect 165037 539611 165071 539645
rect 165229 539611 165263 539645
rect 165421 539611 165455 539645
rect 165613 539611 165647 539645
rect 165805 539611 165839 539645
rect 165997 539611 166031 539645
rect 166214 539604 166248 539638
rect 166414 539604 166448 539638
rect 166214 538876 166248 538910
rect 164714 538476 164748 538510
rect 164941 538483 164975 538517
rect 165133 538483 165167 538517
rect 165325 538483 165359 538517
rect 165517 538483 165551 538517
rect 165709 538483 165743 538517
rect 165901 538483 165935 538517
rect 166414 538476 166448 538510
rect 168514 539604 168548 539638
rect 168837 539611 168871 539645
rect 169029 539611 169063 539645
rect 169221 539611 169255 539645
rect 169413 539611 169447 539645
rect 169605 539611 169639 539645
rect 169797 539611 169831 539645
rect 170014 539604 170048 539638
rect 170214 539604 170248 539638
rect 170014 538876 170048 538910
rect 168514 538476 168548 538510
rect 168741 538483 168775 538517
rect 168933 538483 168967 538517
rect 169125 538483 169159 538517
rect 169317 538483 169351 538517
rect 169509 538483 169543 538517
rect 169701 538483 169735 538517
rect 170214 538476 170248 538510
rect 172214 539604 172248 539638
rect 172537 539611 172571 539645
rect 172729 539611 172763 539645
rect 172921 539611 172955 539645
rect 173113 539611 173147 539645
rect 173305 539611 173339 539645
rect 173497 539611 173531 539645
rect 173714 539604 173748 539638
rect 173914 539604 173948 539638
rect 173714 538876 173748 538910
rect 172214 538476 172248 538510
rect 172441 538483 172475 538517
rect 172633 538483 172667 538517
rect 172825 538483 172859 538517
rect 173017 538483 173051 538517
rect 173209 538483 173243 538517
rect 173401 538483 173435 538517
rect 173914 538476 173948 538510
rect 175714 539604 175748 539638
rect 176037 539611 176071 539645
rect 176229 539611 176263 539645
rect 176421 539611 176455 539645
rect 176613 539611 176647 539645
rect 176805 539611 176839 539645
rect 176997 539611 177031 539645
rect 177214 539604 177248 539638
rect 177414 539604 177448 539638
rect 177214 538876 177248 538910
rect 175714 538476 175748 538510
rect 175941 538483 175975 538517
rect 176133 538483 176167 538517
rect 176325 538483 176359 538517
rect 176517 538483 176551 538517
rect 176709 538483 176743 538517
rect 176901 538483 176935 538517
rect 177414 538476 177448 538510
rect 179314 539604 179348 539638
rect 179637 539611 179671 539645
rect 179829 539611 179863 539645
rect 180021 539611 180055 539645
rect 180213 539611 180247 539645
rect 180405 539611 180439 539645
rect 180597 539611 180631 539645
rect 180814 539604 180848 539638
rect 181014 539604 181048 539638
rect 180814 538876 180848 538910
rect 179314 538476 179348 538510
rect 179541 538483 179575 538517
rect 179733 538483 179767 538517
rect 179925 538483 179959 538517
rect 180117 538483 180151 538517
rect 180309 538483 180343 538517
rect 180501 538483 180535 538517
rect 181014 538476 181048 538510
rect 182614 539604 182648 539638
rect 182937 539611 182971 539645
rect 183129 539611 183163 539645
rect 183321 539611 183355 539645
rect 183513 539611 183547 539645
rect 183705 539611 183739 539645
rect 183897 539611 183931 539645
rect 184114 539604 184148 539638
rect 184314 539604 184348 539638
rect 184114 538876 184148 538910
rect 182614 538476 182648 538510
rect 182841 538483 182875 538517
rect 183033 538483 183067 538517
rect 183225 538483 183259 538517
rect 183417 538483 183451 538517
rect 183609 538483 183643 538517
rect 183801 538483 183835 538517
rect 184314 538476 184348 538510
rect 185914 539604 185948 539638
rect 186237 539611 186271 539645
rect 186429 539611 186463 539645
rect 186621 539611 186655 539645
rect 186813 539611 186847 539645
rect 187005 539611 187039 539645
rect 187197 539611 187231 539645
rect 187414 539604 187448 539638
rect 187614 539604 187648 539638
rect 187414 538876 187448 538910
rect 185914 538476 185948 538510
rect 186141 538483 186175 538517
rect 186333 538483 186367 538517
rect 186525 538483 186559 538517
rect 186717 538483 186751 538517
rect 186909 538483 186943 538517
rect 187101 538483 187135 538517
rect 187614 538476 187648 538510
rect 189214 539604 189248 539638
rect 189537 539611 189571 539645
rect 189729 539611 189763 539645
rect 189921 539611 189955 539645
rect 190113 539611 190147 539645
rect 190305 539611 190339 539645
rect 190497 539611 190531 539645
rect 190714 539604 190748 539638
rect 190914 539604 190948 539638
rect 190714 538876 190748 538910
rect 189214 538476 189248 538510
rect 189441 538483 189475 538517
rect 189633 538483 189667 538517
rect 189825 538483 189859 538517
rect 190017 538483 190051 538517
rect 190209 538483 190243 538517
rect 190401 538483 190435 538517
rect 190914 538476 190948 538510
rect 161304 537704 161338 537738
rect 161508 537704 161542 537738
rect 161700 537704 161734 537738
rect 161908 537704 161942 537738
rect 162100 537704 162134 537738
rect 162324 537704 162358 537738
rect 161304 536976 161338 537010
rect 161604 536976 161638 537010
rect 162004 536976 162038 537010
rect 162324 536976 162358 537010
rect 157812 536684 157980 536718
rect 158190 536684 158358 536718
rect 158448 536684 158616 536718
rect 158706 536684 158874 536718
rect 158964 536684 159132 536718
rect 159222 536684 159390 536718
rect 159480 536684 159648 536718
rect 159738 536684 159906 536718
rect 159996 536684 160164 536718
rect 160254 536684 160422 536718
rect 160512 536684 160680 536718
rect 160896 536684 161064 536718
rect 161154 536684 161322 536718
rect 161412 536684 161580 536718
rect 161794 536684 161962 536718
rect 162052 536684 162220 536718
rect 162432 536684 162600 536718
rect 157812 535956 157980 535990
rect 158190 535956 158358 535990
rect 158448 535956 158616 535990
rect 158706 535956 158874 535990
rect 158964 535956 159132 535990
rect 159222 535956 159390 535990
rect 159480 535956 159648 535990
rect 159738 535956 159906 535990
rect 159996 535956 160164 535990
rect 160254 535956 160422 535990
rect 160512 535956 160680 535990
rect 160896 535956 161064 535990
rect 161154 535956 161322 535990
rect 161412 535956 161580 535990
rect 161794 535956 161962 535990
rect 162052 535956 162220 535990
rect 162432 535956 162600 535990
rect 172277 530336 172311 530370
rect 172385 530376 172419 530410
rect 172637 530362 172671 530396
rect 172705 530362 172739 530396
rect 172773 530362 172807 530396
rect 172919 530362 172953 530396
rect 173389 530336 173423 530370
rect 173753 530372 173787 530406
rect 174237 530336 174271 530370
rect 174347 530336 174381 530370
rect 174455 530372 174489 530406
rect 174565 530372 174599 530406
rect 175029 530362 175063 530396
rect 175097 530362 175131 530396
rect 175165 530362 175199 530396
rect 175311 530362 175345 530396
rect 175616 530362 175650 530396
rect 175891 530370 175925 530404
rect 175987 530398 176021 530432
rect 175814 530262 175848 530296
rect 176131 530372 176165 530406
rect 176227 530420 176261 530454
rect 176092 530246 176126 530280
rect 176375 530360 176409 530394
rect 176471 530408 176505 530442
rect 176726 530414 176760 530448
rect 176828 530408 176862 530442
rect 176557 530272 176591 530306
rect 176987 530301 177021 530335
rect 176806 530246 176840 530280
rect 177194 530347 177228 530381
rect 177296 530362 177330 530396
rect 177745 530362 177779 530396
rect 177941 530362 177975 530396
rect 178145 530362 178179 530396
rect 178259 530362 178293 530396
rect 178459 530349 178493 530383
rect 178579 530362 178613 530396
rect 178801 530362 178835 530396
rect 178869 530362 178903 530396
rect 178937 530362 178971 530396
rect 179083 530362 179117 530396
rect 179287 530362 179321 530396
rect 179433 530362 179467 530396
rect 179501 530362 179535 530396
rect 179569 530362 179603 530396
rect 180300 530362 180334 530396
rect 180396 530362 180430 530396
rect 180537 530398 180571 530432
rect 180633 530398 180667 530432
rect 180795 530398 180829 530432
rect 180705 530285 180739 530319
rect 180873 530285 180907 530319
rect 181347 530398 181381 530432
rect 181509 530398 181543 530432
rect 181269 530285 181303 530319
rect 181605 530398 181639 530432
rect 181437 530285 181471 530319
rect 181746 530362 181780 530396
rect 181842 530362 181876 530396
rect 182047 530362 182081 530396
rect 182193 530362 182227 530396
rect 182261 530362 182295 530396
rect 182329 530362 182363 530396
rect 182643 530336 182677 530370
rect 182903 530372 182937 530406
rect 183151 530362 183185 530396
rect 183297 530362 183331 530396
rect 183365 530362 183399 530396
rect 183433 530362 183467 530396
rect 183969 530336 184003 530370
rect 184333 530372 184367 530406
rect 184759 530336 184793 530370
rect 185019 530372 185053 530406
rect 187001 530526 187035 530560
rect 187001 530458 187035 530492
rect 185267 530362 185301 530396
rect 185413 530362 185447 530396
rect 185481 530362 185515 530396
rect 185549 530362 185583 530396
rect 186085 530336 186119 530370
rect 186449 530372 186483 530406
rect 187001 530195 187035 530229
rect 187001 530127 187035 530161
rect 187101 530530 187135 530564
rect 187101 530462 187135 530496
rect 187273 530376 187307 530410
rect 187381 530336 187415 530370
rect 187101 530195 187135 530229
rect 187101 530127 187135 530161
rect 172277 529764 172311 529798
rect 172385 529724 172419 529758
rect 172837 529764 172871 529798
rect 173201 529728 173235 529762
rect 173941 529764 173975 529798
rect 174305 529728 174339 529762
rect 174867 529738 174901 529772
rect 174981 529738 175015 529772
rect 175185 529738 175219 529772
rect 175381 529738 175415 529772
rect 175554 529738 175588 529772
rect 175656 529753 175690 529787
rect 176044 529854 176078 529888
rect 175863 529799 175897 529833
rect 176293 529828 176327 529862
rect 176022 529692 176056 529726
rect 176124 529686 176158 529720
rect 176379 529692 176413 529726
rect 176475 529740 176509 529774
rect 176758 529854 176792 529888
rect 176623 529680 176657 529714
rect 176719 529728 176753 529762
rect 177036 529838 177070 529872
rect 176863 529702 176897 529736
rect 176959 529730 176993 529764
rect 177234 529738 177268 529772
rect 177681 529815 177715 529849
rect 177849 529815 177883 529849
rect 178666 529838 178700 529872
rect 177759 529702 177793 529736
rect 177921 529702 177955 529736
rect 178017 529702 178051 529736
rect 178158 529738 178192 529772
rect 178254 529738 178288 529772
rect 178468 529738 178502 529772
rect 178743 529730 178777 529764
rect 178944 529854 178978 529888
rect 178839 529702 178873 529736
rect 178983 529728 179017 529762
rect 179227 529740 179261 529774
rect 179409 529828 179443 529862
rect 179079 529680 179113 529714
rect 179323 529692 179357 529726
rect 179658 529854 179692 529888
rect 179839 529799 179873 529833
rect 179578 529686 179612 529720
rect 179680 529692 179714 529726
rect 180046 529753 180080 529787
rect 180148 529738 180182 529772
rect 180246 529738 180280 529772
rect 180348 529753 180382 529787
rect 180736 529854 180770 529888
rect 180555 529799 180589 529833
rect 180985 529828 181019 529862
rect 180714 529692 180748 529726
rect 180816 529686 180850 529720
rect 181071 529692 181105 529726
rect 181167 529740 181201 529774
rect 181450 529854 181484 529888
rect 181315 529680 181349 529714
rect 181411 529728 181445 529762
rect 181728 529838 181762 529872
rect 181555 529702 181589 529736
rect 181651 529730 181685 529764
rect 181926 529738 181960 529772
rect 182091 529764 182125 529798
rect 182351 529728 182385 529762
rect 182713 529738 182747 529772
rect 182909 529738 182943 529772
rect 183113 529738 183147 529772
rect 183227 529738 183261 529772
rect 183693 529764 183727 529798
rect 184057 529728 184091 529762
rect 184797 529764 184831 529798
rect 185161 529728 185195 529762
rect 185901 529764 185935 529798
rect 186265 529728 186299 529762
rect 186749 529764 186783 529798
rect 186859 529764 186893 529798
rect 186967 529728 187001 529762
rect 187077 529728 187111 529762
rect 187273 529724 187307 529758
rect 187381 529764 187415 529798
rect 172277 529248 172311 529282
rect 172385 529288 172419 529322
rect 172837 529248 172871 529282
rect 173201 529284 173235 529318
rect 173941 529248 173975 529282
rect 174305 529284 174339 529318
rect 175275 529310 175309 529344
rect 175437 529310 175471 529344
rect 175197 529197 175231 529231
rect 175533 529310 175567 529344
rect 175365 529197 175399 529231
rect 175674 529274 175708 529308
rect 175770 529274 175804 529308
rect 176212 529274 176246 529308
rect 176280 529274 176314 529308
rect 176348 529274 176382 529308
rect 176416 529274 176450 529308
rect 176484 529274 176518 529308
rect 176552 529274 176586 529308
rect 176620 529274 176654 529308
rect 176688 529274 176722 529308
rect 176756 529274 176790 529308
rect 176824 529274 176858 529308
rect 176892 529274 176926 529308
rect 176960 529274 176994 529308
rect 177028 529274 177062 529308
rect 177096 529274 177130 529308
rect 177164 529274 177198 529308
rect 177232 529274 177266 529308
rect 177659 529274 177693 529308
rect 177762 529274 177796 529308
rect 177864 529259 177898 529293
rect 178230 529320 178264 529354
rect 178332 529326 178366 529360
rect 178071 529213 178105 529247
rect 178252 529158 178286 529192
rect 178587 529320 178621 529354
rect 178831 529332 178865 529366
rect 178501 529184 178535 529218
rect 178683 529272 178717 529306
rect 178927 529284 178961 529318
rect 179071 529310 179105 529344
rect 178966 529158 179000 529192
rect 179167 529282 179201 529316
rect 179442 529274 179476 529308
rect 179699 529274 179733 529308
rect 179244 529174 179278 529208
rect 179819 529261 179853 529295
rect 180125 529248 180159 529282
rect 180235 529248 180269 529282
rect 180343 529284 180377 529318
rect 180453 529284 180487 529318
rect 180711 529274 180745 529308
rect 181138 529274 181172 529308
rect 181206 529274 181240 529308
rect 181274 529274 181308 529308
rect 181342 529274 181376 529308
rect 181410 529274 181444 529308
rect 181478 529274 181512 529308
rect 181546 529274 181580 529308
rect 181614 529274 181648 529308
rect 181682 529274 181716 529308
rect 181750 529274 181784 529308
rect 181818 529274 181852 529308
rect 181886 529274 181920 529308
rect 181954 529274 181988 529308
rect 182022 529274 182056 529308
rect 182090 529274 182124 529308
rect 182158 529274 182192 529308
rect 182599 529261 182633 529295
rect 182719 529274 182753 529308
rect 183141 529248 183175 529282
rect 183505 529284 183539 529318
rect 184245 529248 184279 529282
rect 184609 529284 184643 529318
rect 185533 529248 185567 529282
rect 185897 529284 185931 529318
rect 186381 529248 186415 529282
rect 186480 529248 186514 529282
rect 186579 529248 186613 529282
rect 186687 529284 186721 529318
rect 186790 529284 186824 529318
rect 186893 529284 186927 529318
rect 187273 529288 187307 529322
rect 187381 529248 187415 529282
rect 172277 528676 172311 528710
rect 172385 528636 172419 528670
rect 172837 528676 172871 528710
rect 173201 528640 173235 528674
rect 173941 528676 173975 528710
rect 174305 528640 174339 528674
rect 175045 528676 175079 528710
rect 175409 528640 175443 528674
rect 175927 528650 175961 528684
rect 176577 528727 176611 528761
rect 176047 528663 176081 528697
rect 176203 528650 176237 528684
rect 176323 528663 176357 528697
rect 176745 528727 176779 528761
rect 176655 528614 176689 528648
rect 176817 528614 176851 528648
rect 176913 528614 176947 528648
rect 177054 528650 177088 528684
rect 177150 528650 177184 528684
rect 177561 528650 177595 528684
rect 177757 528650 177791 528684
rect 177961 528650 177995 528684
rect 178075 528650 178109 528684
rect 178411 528650 178445 528684
rect 178838 528650 178872 528684
rect 178906 528650 178940 528684
rect 178974 528650 179008 528684
rect 179042 528650 179076 528684
rect 179110 528650 179144 528684
rect 179178 528650 179212 528684
rect 179246 528650 179280 528684
rect 179314 528650 179348 528684
rect 179382 528650 179416 528684
rect 179450 528650 179484 528684
rect 179518 528650 179552 528684
rect 179586 528650 179620 528684
rect 179654 528650 179688 528684
rect 179722 528650 179756 528684
rect 179790 528650 179824 528684
rect 179858 528650 179892 528684
rect 180251 528650 180285 528684
rect 180371 528663 180405 528697
rect 180522 528650 180556 528684
rect 180624 528665 180658 528699
rect 181012 528766 181046 528800
rect 180831 528711 180865 528745
rect 181261 528740 181295 528774
rect 180990 528604 181024 528638
rect 181092 528598 181126 528632
rect 181347 528604 181381 528638
rect 181443 528652 181477 528686
rect 181726 528766 181760 528800
rect 181591 528592 181625 528626
rect 181687 528640 181721 528674
rect 182004 528750 182038 528784
rect 181831 528614 181865 528648
rect 181927 528642 181961 528676
rect 182202 528650 182236 528684
rect 182957 528676 182991 528710
rect 183321 528640 183355 528674
rect 184061 528676 184095 528710
rect 184425 528640 184459 528674
rect 185165 528676 185199 528710
rect 185529 528640 185563 528674
rect 186269 528676 186303 528710
rect 186633 528640 186667 528674
rect 187273 528636 187307 528670
rect 187381 528676 187415 528710
rect 172277 528160 172311 528194
rect 172385 528200 172419 528234
rect 172837 528160 172871 528194
rect 173201 528196 173235 528230
rect 173941 528160 173975 528194
rect 174305 528196 174339 528230
rect 175229 528160 175263 528194
rect 175593 528196 175627 528230
rect 176106 528186 176140 528220
rect 176208 528171 176242 528205
rect 176574 528232 176608 528266
rect 176676 528238 176710 528272
rect 176415 528125 176449 528159
rect 176596 528070 176630 528104
rect 176931 528232 176965 528266
rect 177175 528244 177209 528278
rect 176845 528096 176879 528130
rect 177027 528184 177061 528218
rect 177271 528196 177305 528230
rect 177415 528222 177449 528256
rect 177310 528070 177344 528104
rect 177511 528194 177545 528228
rect 177786 528186 177820 528220
rect 177999 528173 178033 528207
rect 178119 528186 178153 528220
rect 177588 528086 177622 528120
rect 178285 528160 178319 528194
rect 178384 528160 178418 528194
rect 178483 528160 178517 528194
rect 178591 528196 178625 528230
rect 178694 528196 178728 528230
rect 178797 528196 178831 528230
rect 179012 528186 179046 528220
rect 179108 528186 179142 528220
rect 179249 528222 179283 528256
rect 179345 528222 179379 528256
rect 179507 528222 179541 528256
rect 179417 528109 179451 528143
rect 179585 528109 179619 528143
rect 180125 528160 180159 528194
rect 180224 528160 180258 528194
rect 180323 528160 180357 528194
rect 180431 528196 180465 528230
rect 180534 528196 180568 528230
rect 180637 528196 180671 528230
rect 181036 528186 181070 528220
rect 181132 528186 181166 528220
rect 181273 528222 181307 528256
rect 181369 528222 181403 528256
rect 181531 528222 181565 528256
rect 181441 528109 181475 528143
rect 181609 528109 181643 528143
rect 182129 528160 182163 528194
rect 182493 528196 182527 528230
rect 183233 528160 183267 528194
rect 183597 528196 183631 528230
rect 184337 528160 184371 528194
rect 184701 528196 184735 528230
rect 185533 528160 185567 528194
rect 185897 528196 185931 528230
rect 186381 528160 186415 528194
rect 186480 528160 186514 528194
rect 186579 528160 186613 528194
rect 186687 528196 186721 528230
rect 186790 528196 186824 528230
rect 186893 528196 186927 528230
rect 187273 528200 187307 528234
rect 187381 528160 187415 528194
rect 172277 527588 172311 527622
rect 172385 527548 172419 527582
rect 172837 527588 172871 527622
rect 173201 527552 173235 527586
rect 173941 527588 173975 527622
rect 174305 527552 174339 527586
rect 175045 527588 175079 527622
rect 175409 527552 175443 527586
rect 175893 527588 175927 527622
rect 176003 527588 176037 527622
rect 176111 527552 176145 527586
rect 176221 527552 176255 527586
rect 176457 527562 176491 527596
rect 176653 527562 176687 527596
rect 176857 527562 176891 527596
rect 176971 527562 177005 527596
rect 177153 527588 177187 527622
rect 177261 527548 177295 527582
rect 177805 527588 177839 527622
rect 178169 527552 178203 527586
rect 178595 527588 178629 527622
rect 178855 527552 178889 527586
rect 179033 527562 179067 527596
rect 179229 527562 179263 527596
rect 179433 527562 179467 527596
rect 179547 527562 179581 527596
rect 180013 527588 180047 527622
rect 180377 527552 180411 527586
rect 181117 527588 181151 527622
rect 181481 527552 181515 527586
rect 181965 527588 181999 527622
rect 182075 527588 182109 527622
rect 182183 527552 182217 527586
rect 182293 527552 182327 527586
rect 182957 527588 182991 527622
rect 183321 527552 183355 527586
rect 184061 527588 184095 527622
rect 184425 527552 184459 527586
rect 185165 527588 185199 527622
rect 185529 527552 185563 527586
rect 186269 527588 186303 527622
rect 186633 527552 186667 527586
rect 187273 527548 187307 527582
rect 187381 527588 187415 527622
rect 172277 527072 172311 527106
rect 172385 527112 172419 527146
rect 172837 527072 172871 527106
rect 173201 527108 173235 527142
rect 173941 527072 173975 527106
rect 174305 527108 174339 527142
rect 175229 527072 175263 527106
rect 175593 527108 175627 527142
rect 176333 527072 176367 527106
rect 176697 527108 176731 527142
rect 177437 527072 177471 527106
rect 177801 527108 177835 527142
rect 178541 527072 178575 527106
rect 178905 527108 178939 527142
rect 179389 527072 179423 527106
rect 179499 527072 179533 527106
rect 179607 527108 179641 527142
rect 179717 527108 179751 527142
rect 180381 527072 180415 527106
rect 180745 527108 180779 527142
rect 181485 527072 181519 527106
rect 181849 527108 181883 527142
rect 182589 527072 182623 527106
rect 182953 527108 182987 527142
rect 183693 527072 183727 527106
rect 184057 527108 184091 527142
rect 184541 527072 184575 527106
rect 184651 527072 184685 527106
rect 184759 527108 184793 527142
rect 184869 527108 184903 527142
rect 185533 527072 185567 527106
rect 185897 527108 185931 527142
rect 186381 527072 186415 527106
rect 186480 527072 186514 527106
rect 186579 527072 186613 527106
rect 186687 527108 186721 527142
rect 186790 527108 186824 527142
rect 186893 527108 186927 527142
rect 187273 527112 187307 527146
rect 187381 527072 187415 527106
rect 172277 526500 172311 526534
rect 172385 526460 172419 526494
rect 172837 526500 172871 526534
rect 173201 526464 173235 526498
rect 173941 526500 173975 526534
rect 174305 526464 174339 526498
rect 175045 526500 175079 526534
rect 175409 526464 175443 526498
rect 176149 526500 176183 526534
rect 176513 526464 176547 526498
rect 176939 526500 176973 526534
rect 177199 526464 177233 526498
rect 177805 526500 177839 526534
rect 178169 526464 178203 526498
rect 178909 526500 178943 526534
rect 179273 526464 179307 526498
rect 180013 526500 180047 526534
rect 180377 526464 180411 526498
rect 181117 526500 181151 526534
rect 181481 526464 181515 526498
rect 181965 526500 181999 526534
rect 182075 526500 182109 526534
rect 182183 526464 182217 526498
rect 182293 526464 182327 526498
rect 182957 526500 182991 526534
rect 183321 526464 183355 526498
rect 184061 526500 184095 526534
rect 184425 526464 184459 526498
rect 185165 526500 185199 526534
rect 185529 526464 185563 526498
rect 186269 526500 186303 526534
rect 186633 526464 186667 526498
rect 187273 526460 187307 526494
rect 187381 526500 187415 526534
rect 172277 525984 172311 526018
rect 172385 526024 172419 526058
rect 172837 525984 172871 526018
rect 173201 526020 173235 526054
rect 173941 525984 173975 526018
rect 174305 526020 174339 526054
rect 175229 525984 175263 526018
rect 175593 526020 175627 526054
rect 176333 525984 176367 526018
rect 176697 526020 176731 526054
rect 177437 525984 177471 526018
rect 177801 526020 177835 526054
rect 178541 525984 178575 526018
rect 178905 526020 178939 526054
rect 179389 525984 179423 526018
rect 179499 525984 179533 526018
rect 179607 526020 179641 526054
rect 179717 526020 179751 526054
rect 180381 525984 180415 526018
rect 180745 526020 180779 526054
rect 181485 525984 181519 526018
rect 181849 526020 181883 526054
rect 182589 525984 182623 526018
rect 182953 526020 182987 526054
rect 183693 525984 183727 526018
rect 184057 526020 184091 526054
rect 184541 525984 184575 526018
rect 184651 525984 184685 526018
rect 184759 526020 184793 526054
rect 184869 526020 184903 526054
rect 185533 525984 185567 526018
rect 185897 526020 185931 526054
rect 186381 525984 186415 526018
rect 186480 525984 186514 526018
rect 186579 525984 186613 526018
rect 186687 526020 186721 526054
rect 186790 526020 186824 526054
rect 186893 526020 186927 526054
rect 187273 526024 187307 526058
rect 187381 525984 187415 526018
rect 172277 525412 172311 525446
rect 172385 525372 172419 525406
rect 172837 525412 172871 525446
rect 173201 525376 173235 525410
rect 173941 525412 173975 525446
rect 174305 525376 174339 525410
rect 175045 525412 175079 525446
rect 175409 525376 175443 525410
rect 176149 525412 176183 525446
rect 176513 525376 176547 525410
rect 176939 525412 176973 525446
rect 177199 525376 177233 525410
rect 177805 525412 177839 525446
rect 178169 525376 178203 525410
rect 178909 525412 178943 525446
rect 179273 525376 179307 525410
rect 180013 525412 180047 525446
rect 180377 525376 180411 525410
rect 181117 525412 181151 525446
rect 181481 525376 181515 525410
rect 181965 525412 181999 525446
rect 182075 525412 182109 525446
rect 182183 525376 182217 525410
rect 182293 525376 182327 525410
rect 182957 525412 182991 525446
rect 183321 525376 183355 525410
rect 184061 525412 184095 525446
rect 184425 525376 184459 525410
rect 185165 525412 185199 525446
rect 185529 525376 185563 525410
rect 186269 525412 186303 525446
rect 186633 525376 186667 525410
rect 187273 525372 187307 525406
rect 187381 525412 187415 525446
rect 172277 524896 172311 524930
rect 172385 524936 172419 524970
rect 172837 524896 172871 524930
rect 173201 524932 173235 524966
rect 173941 524896 173975 524930
rect 174305 524932 174339 524966
rect 175229 524896 175263 524930
rect 175593 524932 175627 524966
rect 176333 524896 176367 524930
rect 176697 524932 176731 524966
rect 177437 524896 177471 524930
rect 177801 524932 177835 524966
rect 178541 524896 178575 524930
rect 178905 524932 178939 524966
rect 179389 524896 179423 524930
rect 179499 524896 179533 524930
rect 179607 524932 179641 524966
rect 179717 524932 179751 524966
rect 180381 524896 180415 524930
rect 180745 524932 180779 524966
rect 181485 524896 181519 524930
rect 181849 524932 181883 524966
rect 182589 524896 182623 524930
rect 182953 524932 182987 524966
rect 183693 524896 183727 524930
rect 184057 524932 184091 524966
rect 184541 524896 184575 524930
rect 184651 524896 184685 524930
rect 184759 524932 184793 524966
rect 184869 524932 184903 524966
rect 185533 524896 185567 524930
rect 185897 524932 185931 524966
rect 186381 524896 186415 524930
rect 186480 524896 186514 524930
rect 186579 524896 186613 524930
rect 186687 524932 186721 524966
rect 186790 524932 186824 524966
rect 186893 524932 186927 524966
rect 187273 524936 187307 524970
rect 187381 524896 187415 524930
rect 172277 524324 172311 524358
rect 172385 524284 172419 524318
rect 172837 524324 172871 524358
rect 173201 524288 173235 524322
rect 173941 524324 173975 524358
rect 174305 524288 174339 524322
rect 175045 524324 175079 524358
rect 175409 524288 175443 524322
rect 176149 524324 176183 524358
rect 176513 524288 176547 524322
rect 176939 524324 176973 524358
rect 177199 524288 177233 524322
rect 177805 524324 177839 524358
rect 178169 524288 178203 524322
rect 178909 524324 178943 524358
rect 179273 524288 179307 524322
rect 180013 524324 180047 524358
rect 180377 524288 180411 524322
rect 181117 524324 181151 524358
rect 181481 524288 181515 524322
rect 181965 524324 181999 524358
rect 182075 524324 182109 524358
rect 182183 524288 182217 524322
rect 182293 524288 182327 524322
rect 182957 524324 182991 524358
rect 183321 524288 183355 524322
rect 184061 524324 184095 524358
rect 184425 524288 184459 524322
rect 185165 524324 185199 524358
rect 185529 524288 185563 524322
rect 186269 524324 186303 524358
rect 186633 524288 186667 524322
rect 187273 524284 187307 524318
rect 187381 524324 187415 524358
rect 172277 523808 172311 523842
rect 172385 523848 172419 523882
rect 172837 523808 172871 523842
rect 173201 523844 173235 523878
rect 173941 523808 173975 523842
rect 174305 523844 174339 523878
rect 175229 523808 175263 523842
rect 175593 523844 175627 523878
rect 176333 523808 176367 523842
rect 176697 523844 176731 523878
rect 177437 523808 177471 523842
rect 177801 523844 177835 523878
rect 178541 523808 178575 523842
rect 178905 523844 178939 523878
rect 179389 523808 179423 523842
rect 179499 523808 179533 523842
rect 179607 523844 179641 523878
rect 179717 523844 179751 523878
rect 180381 523808 180415 523842
rect 180745 523844 180779 523878
rect 181485 523808 181519 523842
rect 181849 523844 181883 523878
rect 182589 523808 182623 523842
rect 182953 523844 182987 523878
rect 183693 523808 183727 523842
rect 184057 523844 184091 523878
rect 184541 523808 184575 523842
rect 184651 523808 184685 523842
rect 184759 523844 184793 523878
rect 184869 523844 184903 523878
rect 185533 523808 185567 523842
rect 185897 523844 185931 523878
rect 186381 523808 186415 523842
rect 186480 523808 186514 523842
rect 186579 523808 186613 523842
rect 186687 523844 186721 523878
rect 186790 523844 186824 523878
rect 186893 523844 186927 523878
rect 187273 523848 187307 523882
rect 187381 523808 187415 523842
rect 172277 523236 172311 523270
rect 172385 523196 172419 523230
rect 172837 523236 172871 523270
rect 173201 523200 173235 523234
rect 173941 523236 173975 523270
rect 174305 523200 174339 523234
rect 175045 523236 175079 523270
rect 175409 523200 175443 523234
rect 176149 523236 176183 523270
rect 176513 523200 176547 523234
rect 176939 523236 176973 523270
rect 177199 523200 177233 523234
rect 177805 523236 177839 523270
rect 178169 523200 178203 523234
rect 178909 523236 178943 523270
rect 179273 523200 179307 523234
rect 180013 523236 180047 523270
rect 180377 523200 180411 523234
rect 181117 523236 181151 523270
rect 181481 523200 181515 523234
rect 181965 523236 181999 523270
rect 182075 523236 182109 523270
rect 182183 523200 182217 523234
rect 182293 523200 182327 523234
rect 182957 523236 182991 523270
rect 183321 523200 183355 523234
rect 184061 523236 184095 523270
rect 184425 523200 184459 523234
rect 185165 523236 185199 523270
rect 185529 523200 185563 523234
rect 186269 523236 186303 523270
rect 186633 523200 186667 523234
rect 187273 523196 187307 523230
rect 187381 523236 187415 523270
rect 172277 522720 172311 522754
rect 172385 522760 172419 522794
rect 172837 522720 172871 522754
rect 173201 522756 173235 522790
rect 173941 522720 173975 522754
rect 174305 522756 174339 522790
rect 175229 522720 175263 522754
rect 175593 522756 175627 522790
rect 176333 522720 176367 522754
rect 176697 522756 176731 522790
rect 177437 522720 177471 522754
rect 177801 522756 177835 522790
rect 178541 522720 178575 522754
rect 178905 522756 178939 522790
rect 179389 522720 179423 522754
rect 179499 522720 179533 522754
rect 179607 522756 179641 522790
rect 179717 522756 179751 522790
rect 180381 522720 180415 522754
rect 180745 522756 180779 522790
rect 181485 522720 181519 522754
rect 181849 522756 181883 522790
rect 182589 522720 182623 522754
rect 182953 522756 182987 522790
rect 183693 522720 183727 522754
rect 184057 522756 184091 522790
rect 184541 522720 184575 522754
rect 184651 522720 184685 522754
rect 184759 522756 184793 522790
rect 184869 522756 184903 522790
rect 185533 522720 185567 522754
rect 185897 522756 185931 522790
rect 186381 522720 186415 522754
rect 186480 522720 186514 522754
rect 186579 522720 186613 522754
rect 186687 522756 186721 522790
rect 186790 522756 186824 522790
rect 186893 522756 186927 522790
rect 187273 522760 187307 522794
rect 187381 522720 187415 522754
rect 172277 522148 172311 522182
rect 172385 522108 172419 522142
rect 172837 522148 172871 522182
rect 173201 522112 173235 522146
rect 173941 522148 173975 522182
rect 174305 522112 174339 522146
rect 175045 522148 175079 522182
rect 175409 522112 175443 522146
rect 176149 522148 176183 522182
rect 176513 522112 176547 522146
rect 176939 522148 176973 522182
rect 177199 522112 177233 522146
rect 177805 522148 177839 522182
rect 178169 522112 178203 522146
rect 178909 522148 178943 522182
rect 179273 522112 179307 522146
rect 180013 522148 180047 522182
rect 180377 522112 180411 522146
rect 181117 522148 181151 522182
rect 181481 522112 181515 522146
rect 181965 522148 181999 522182
rect 182075 522148 182109 522182
rect 182183 522112 182217 522146
rect 182293 522112 182327 522146
rect 182957 522148 182991 522182
rect 183321 522112 183355 522146
rect 184061 522148 184095 522182
rect 184425 522112 184459 522146
rect 185165 522148 185199 522182
rect 185529 522112 185563 522146
rect 186269 522148 186303 522182
rect 186633 522112 186667 522146
rect 187273 522108 187307 522142
rect 187381 522148 187415 522182
rect 172277 521632 172311 521666
rect 172385 521672 172419 521706
rect 172837 521632 172871 521666
rect 173201 521668 173235 521702
rect 173941 521632 173975 521666
rect 174305 521668 174339 521702
rect 175229 521632 175263 521666
rect 175593 521668 175627 521702
rect 176333 521632 176367 521666
rect 176697 521668 176731 521702
rect 177437 521632 177471 521666
rect 177801 521668 177835 521702
rect 178541 521632 178575 521666
rect 178905 521668 178939 521702
rect 179389 521632 179423 521666
rect 179499 521632 179533 521666
rect 179607 521668 179641 521702
rect 179717 521668 179751 521702
rect 180381 521632 180415 521666
rect 180745 521668 180779 521702
rect 181485 521632 181519 521666
rect 181849 521668 181883 521702
rect 182589 521632 182623 521666
rect 182953 521668 182987 521702
rect 183693 521632 183727 521666
rect 184057 521668 184091 521702
rect 184541 521632 184575 521666
rect 184651 521632 184685 521666
rect 184759 521668 184793 521702
rect 184869 521668 184903 521702
rect 185533 521632 185567 521666
rect 185897 521668 185931 521702
rect 186381 521632 186415 521666
rect 186480 521632 186514 521666
rect 186579 521632 186613 521666
rect 186687 521668 186721 521702
rect 186790 521668 186824 521702
rect 186893 521668 186927 521702
rect 187273 521672 187307 521706
rect 187381 521632 187415 521666
rect 172277 521060 172311 521094
rect 172385 521020 172419 521054
rect 172837 521060 172871 521094
rect 173201 521024 173235 521058
rect 173941 521060 173975 521094
rect 174305 521024 174339 521058
rect 175045 521060 175079 521094
rect 175409 521024 175443 521058
rect 176149 521060 176183 521094
rect 176513 521024 176547 521058
rect 176939 521060 176973 521094
rect 177199 521024 177233 521058
rect 177805 521060 177839 521094
rect 178169 521024 178203 521058
rect 178909 521060 178943 521094
rect 179273 521024 179307 521058
rect 180013 521060 180047 521094
rect 180377 521024 180411 521058
rect 181117 521060 181151 521094
rect 181481 521024 181515 521058
rect 181965 521060 181999 521094
rect 182075 521060 182109 521094
rect 182183 521024 182217 521058
rect 182293 521024 182327 521058
rect 182957 521060 182991 521094
rect 183321 521024 183355 521058
rect 184061 521060 184095 521094
rect 184425 521024 184459 521058
rect 185165 521060 185199 521094
rect 185529 521024 185563 521058
rect 186269 521060 186303 521094
rect 186633 521024 186667 521058
rect 187273 521020 187307 521054
rect 187381 521060 187415 521094
rect 172277 520544 172311 520578
rect 172385 520584 172419 520618
rect 172837 520544 172871 520578
rect 173201 520580 173235 520614
rect 173941 520544 173975 520578
rect 174305 520580 174339 520614
rect 175229 520544 175263 520578
rect 175593 520580 175627 520614
rect 176333 520544 176367 520578
rect 176697 520580 176731 520614
rect 177437 520544 177471 520578
rect 177801 520580 177835 520614
rect 178541 520544 178575 520578
rect 178905 520580 178939 520614
rect 179389 520544 179423 520578
rect 179499 520544 179533 520578
rect 179607 520580 179641 520614
rect 179717 520580 179751 520614
rect 180381 520544 180415 520578
rect 180745 520580 180779 520614
rect 181485 520544 181519 520578
rect 181849 520580 181883 520614
rect 182589 520544 182623 520578
rect 182953 520580 182987 520614
rect 183693 520544 183727 520578
rect 184057 520580 184091 520614
rect 184541 520544 184575 520578
rect 184651 520544 184685 520578
rect 184759 520580 184793 520614
rect 184869 520580 184903 520614
rect 185533 520544 185567 520578
rect 185897 520580 185931 520614
rect 186381 520544 186415 520578
rect 186480 520544 186514 520578
rect 186579 520544 186613 520578
rect 186687 520580 186721 520614
rect 186790 520580 186824 520614
rect 186893 520580 186927 520614
rect 187273 520584 187307 520618
rect 187381 520544 187415 520578
rect 172277 519972 172311 520006
rect 172385 519932 172419 519966
rect 172837 519972 172871 520006
rect 173201 519936 173235 519970
rect 173941 519972 173975 520006
rect 174305 519936 174339 519970
rect 175045 519972 175079 520006
rect 175409 519936 175443 519970
rect 176149 519972 176183 520006
rect 176513 519936 176547 519970
rect 176939 519972 176973 520006
rect 177199 519936 177233 519970
rect 177805 519972 177839 520006
rect 178169 519936 178203 519970
rect 178909 519972 178943 520006
rect 179273 519936 179307 519970
rect 180013 519972 180047 520006
rect 180377 519936 180411 519970
rect 181117 519972 181151 520006
rect 181481 519936 181515 519970
rect 181965 519972 181999 520006
rect 182075 519972 182109 520006
rect 182183 519936 182217 519970
rect 182293 519936 182327 519970
rect 182957 519972 182991 520006
rect 183321 519936 183355 519970
rect 184061 519972 184095 520006
rect 184425 519936 184459 519970
rect 185165 519972 185199 520006
rect 185529 519936 185563 519970
rect 186269 519972 186303 520006
rect 186633 519936 186667 519970
rect 187273 519932 187307 519966
rect 187381 519972 187415 520006
rect 172277 519456 172311 519490
rect 172385 519496 172419 519530
rect 172837 519456 172871 519490
rect 173201 519492 173235 519526
rect 173941 519456 173975 519490
rect 174305 519492 174339 519526
rect 175229 519456 175263 519490
rect 175593 519492 175627 519526
rect 176333 519456 176367 519490
rect 176697 519492 176731 519526
rect 177437 519456 177471 519490
rect 177801 519492 177835 519526
rect 178541 519456 178575 519490
rect 178905 519492 178939 519526
rect 179389 519456 179423 519490
rect 179499 519456 179533 519490
rect 179607 519492 179641 519526
rect 179717 519492 179751 519526
rect 180381 519456 180415 519490
rect 180745 519492 180779 519526
rect 181485 519456 181519 519490
rect 181849 519492 181883 519526
rect 182589 519456 182623 519490
rect 182953 519492 182987 519526
rect 183693 519456 183727 519490
rect 184057 519492 184091 519526
rect 184541 519456 184575 519490
rect 184651 519456 184685 519490
rect 184759 519492 184793 519526
rect 184869 519492 184903 519526
rect 185533 519456 185567 519490
rect 185897 519492 185931 519526
rect 186381 519456 186415 519490
rect 186480 519456 186514 519490
rect 186579 519456 186613 519490
rect 186687 519492 186721 519526
rect 186790 519492 186824 519526
rect 186893 519492 186927 519526
rect 187273 519496 187307 519530
rect 187381 519456 187415 519490
rect 172277 518884 172311 518918
rect 172385 518844 172419 518878
rect 172837 518884 172871 518918
rect 173201 518848 173235 518882
rect 173941 518884 173975 518918
rect 174305 518848 174339 518882
rect 175045 518884 175079 518918
rect 175409 518848 175443 518882
rect 176149 518884 176183 518918
rect 176513 518848 176547 518882
rect 176939 518884 176973 518918
rect 177199 518848 177233 518882
rect 177805 518884 177839 518918
rect 178169 518848 178203 518882
rect 178909 518884 178943 518918
rect 179273 518848 179307 518882
rect 180013 518884 180047 518918
rect 180377 518848 180411 518882
rect 181117 518884 181151 518918
rect 181481 518848 181515 518882
rect 181965 518884 181999 518918
rect 182075 518884 182109 518918
rect 182183 518848 182217 518882
rect 182293 518848 182327 518882
rect 182957 518884 182991 518918
rect 183321 518848 183355 518882
rect 184061 518884 184095 518918
rect 184425 518848 184459 518882
rect 185165 518884 185199 518918
rect 185529 518848 185563 518882
rect 186269 518884 186303 518918
rect 186633 518848 186667 518882
rect 187273 518844 187307 518878
rect 187381 518884 187415 518918
rect 172277 518368 172311 518402
rect 172385 518408 172419 518442
rect 172837 518368 172871 518402
rect 173201 518404 173235 518438
rect 173941 518368 173975 518402
rect 174305 518404 174339 518438
rect 175229 518368 175263 518402
rect 175593 518404 175627 518438
rect 176333 518368 176367 518402
rect 176697 518404 176731 518438
rect 177437 518368 177471 518402
rect 177801 518404 177835 518438
rect 178541 518368 178575 518402
rect 178905 518404 178939 518438
rect 179389 518368 179423 518402
rect 179499 518368 179533 518402
rect 179607 518404 179641 518438
rect 179717 518404 179751 518438
rect 180381 518368 180415 518402
rect 180745 518404 180779 518438
rect 181485 518368 181519 518402
rect 181849 518404 181883 518438
rect 182589 518368 182623 518402
rect 182953 518404 182987 518438
rect 183693 518368 183727 518402
rect 184057 518404 184091 518438
rect 184541 518368 184575 518402
rect 184651 518368 184685 518402
rect 184759 518404 184793 518438
rect 184869 518404 184903 518438
rect 185533 518368 185567 518402
rect 185897 518404 185931 518438
rect 186381 518368 186415 518402
rect 186480 518368 186514 518402
rect 186579 518368 186613 518402
rect 186687 518404 186721 518438
rect 186790 518404 186824 518438
rect 186893 518404 186927 518438
rect 187273 518408 187307 518442
rect 187381 518368 187415 518402
rect 172277 517796 172311 517830
rect 172385 517756 172419 517790
rect 172837 517796 172871 517830
rect 173201 517760 173235 517794
rect 173941 517796 173975 517830
rect 174305 517760 174339 517794
rect 175045 517796 175079 517830
rect 175409 517760 175443 517794
rect 176149 517796 176183 517830
rect 176513 517760 176547 517794
rect 176939 517796 176973 517830
rect 177199 517760 177233 517794
rect 177805 517796 177839 517830
rect 178169 517760 178203 517794
rect 178909 517796 178943 517830
rect 179273 517760 179307 517794
rect 180013 517796 180047 517830
rect 180377 517760 180411 517794
rect 181117 517796 181151 517830
rect 181481 517760 181515 517794
rect 181965 517796 181999 517830
rect 182075 517796 182109 517830
rect 182183 517760 182217 517794
rect 182293 517760 182327 517794
rect 182957 517796 182991 517830
rect 183321 517760 183355 517794
rect 184061 517796 184095 517830
rect 184425 517760 184459 517794
rect 185165 517796 185199 517830
rect 185529 517760 185563 517794
rect 186269 517796 186303 517830
rect 186633 517760 186667 517794
rect 187273 517756 187307 517790
rect 187381 517796 187415 517830
rect 172277 517280 172311 517314
rect 172385 517320 172419 517354
rect 172837 517280 172871 517314
rect 173201 517316 173235 517350
rect 173941 517280 173975 517314
rect 174305 517316 174339 517350
rect 175229 517280 175263 517314
rect 175593 517316 175627 517350
rect 176333 517280 176367 517314
rect 176697 517316 176731 517350
rect 177437 517280 177471 517314
rect 177801 517316 177835 517350
rect 178541 517280 178575 517314
rect 178905 517316 178939 517350
rect 179389 517280 179423 517314
rect 179499 517280 179533 517314
rect 179607 517316 179641 517350
rect 179717 517316 179751 517350
rect 180381 517280 180415 517314
rect 180745 517316 180779 517350
rect 181485 517280 181519 517314
rect 181849 517316 181883 517350
rect 182589 517280 182623 517314
rect 182953 517316 182987 517350
rect 183693 517280 183727 517314
rect 184057 517316 184091 517350
rect 184541 517280 184575 517314
rect 184651 517280 184685 517314
rect 184759 517316 184793 517350
rect 184869 517316 184903 517350
rect 185533 517280 185567 517314
rect 185897 517316 185931 517350
rect 186381 517280 186415 517314
rect 186480 517280 186514 517314
rect 186579 517280 186613 517314
rect 186687 517316 186721 517350
rect 186790 517316 186824 517350
rect 186893 517316 186927 517350
rect 187273 517320 187307 517354
rect 187381 517280 187415 517314
rect 172277 516708 172311 516742
rect 172385 516668 172419 516702
rect 172837 516708 172871 516742
rect 173201 516672 173235 516706
rect 173941 516708 173975 516742
rect 174305 516672 174339 516706
rect 175045 516708 175079 516742
rect 175409 516672 175443 516706
rect 176149 516708 176183 516742
rect 176513 516672 176547 516706
rect 176939 516708 176973 516742
rect 177199 516672 177233 516706
rect 177805 516708 177839 516742
rect 178169 516672 178203 516706
rect 178909 516708 178943 516742
rect 179273 516672 179307 516706
rect 180013 516708 180047 516742
rect 180377 516672 180411 516706
rect 181117 516708 181151 516742
rect 181481 516672 181515 516706
rect 181965 516708 181999 516742
rect 182075 516708 182109 516742
rect 182183 516672 182217 516706
rect 182293 516672 182327 516706
rect 182957 516708 182991 516742
rect 183321 516672 183355 516706
rect 184061 516708 184095 516742
rect 184425 516672 184459 516706
rect 185165 516708 185199 516742
rect 185529 516672 185563 516706
rect 186269 516708 186303 516742
rect 186633 516672 186667 516706
rect 187273 516668 187307 516702
rect 187381 516708 187415 516742
rect 172277 516192 172311 516226
rect 172385 516232 172419 516266
rect 172837 516192 172871 516226
rect 173201 516228 173235 516262
rect 173941 516192 173975 516226
rect 174305 516228 174339 516262
rect 175229 516192 175263 516226
rect 175593 516228 175627 516262
rect 176333 516192 176367 516226
rect 176697 516228 176731 516262
rect 177437 516192 177471 516226
rect 177801 516228 177835 516262
rect 178541 516192 178575 516226
rect 178905 516228 178939 516262
rect 179389 516192 179423 516226
rect 179499 516192 179533 516226
rect 179607 516228 179641 516262
rect 179717 516228 179751 516262
rect 180381 516192 180415 516226
rect 180745 516228 180779 516262
rect 181485 516192 181519 516226
rect 181849 516228 181883 516262
rect 182589 516192 182623 516226
rect 182953 516228 182987 516262
rect 183693 516192 183727 516226
rect 184057 516228 184091 516262
rect 184541 516192 184575 516226
rect 184651 516192 184685 516226
rect 184759 516228 184793 516262
rect 184869 516228 184903 516262
rect 185533 516192 185567 516226
rect 185897 516228 185931 516262
rect 186381 516192 186415 516226
rect 186480 516192 186514 516226
rect 186579 516192 186613 516226
rect 186687 516228 186721 516262
rect 186790 516228 186824 516262
rect 186893 516228 186927 516262
rect 187273 516232 187307 516266
rect 187381 516192 187415 516226
rect 172277 515620 172311 515654
rect 172385 515580 172419 515614
rect 172581 515620 172615 515654
rect 172680 515620 172714 515654
rect 172779 515620 172813 515654
rect 172887 515584 172921 515618
rect 172990 515584 173024 515618
rect 173093 515584 173127 515618
rect 173491 515594 173525 515628
rect 173637 515594 173671 515628
rect 173705 515594 173739 515628
rect 173773 515594 173807 515628
rect 174053 515620 174087 515654
rect 174152 515620 174186 515654
rect 174251 515620 174285 515654
rect 174359 515584 174393 515618
rect 174462 515584 174496 515618
rect 174565 515584 174599 515618
rect 175229 515620 175263 515654
rect 175593 515584 175627 515618
rect 176333 515620 176367 515654
rect 176697 515584 176731 515618
rect 177153 515620 177187 515654
rect 177261 515580 177295 515614
rect 177805 515620 177839 515654
rect 178169 515584 178203 515618
rect 178909 515620 178943 515654
rect 179273 515584 179307 515618
rect 179729 515620 179763 515654
rect 179837 515580 179871 515614
rect 180381 515620 180415 515654
rect 180745 515584 180779 515618
rect 181229 515620 181263 515654
rect 181328 515620 181362 515654
rect 181427 515620 181461 515654
rect 181535 515584 181569 515618
rect 181638 515584 181672 515618
rect 181741 515584 181775 515618
rect 182141 515607 182175 515641
rect 182259 515594 182293 515628
rect 182957 515620 182991 515654
rect 183321 515584 183355 515618
rect 184061 515620 184095 515654
rect 184425 515584 184459 515618
rect 184881 515620 184915 515654
rect 184989 515580 185023 515614
rect 185533 515620 185567 515654
rect 185897 515584 185931 515618
rect 186463 515594 186497 515628
rect 186609 515594 186643 515628
rect 186677 515594 186711 515628
rect 186745 515594 186779 515628
rect 186997 515620 187031 515654
rect 187105 515580 187139 515614
rect 187273 515580 187307 515614
rect 187381 515620 187415 515654
<< xpolycontact >>
rect 164318 537549 164388 537981
rect 164318 536033 164388 536465
rect 164636 537549 164706 537981
rect 164636 536033 164706 536465
rect 164954 537549 165024 537981
rect 164954 536033 165024 536465
rect 165272 537549 165342 537981
rect 165272 536033 165342 536465
rect 165590 537549 165660 537981
rect 165590 536033 165660 536465
rect 165908 537549 165978 537981
rect 165908 536033 165978 536465
rect 166226 537549 166296 537981
rect 166226 536033 166296 536465
rect 166544 537549 166614 537981
rect 166544 536033 166614 536465
rect 168090 537549 168160 537981
rect 168090 536033 168160 536465
rect 168408 537549 168478 537981
rect 168408 536033 168478 536465
rect 168726 537549 168796 537981
rect 168726 536033 168796 536465
rect 169044 537549 169114 537981
rect 169044 536033 169114 536465
rect 171826 537549 171896 537981
rect 171826 536033 171896 536465
rect 172144 537549 172214 537981
rect 172144 536033 172214 536465
rect 175344 537549 175414 537981
rect 175344 536033 175414 536465
rect 178944 537549 179014 537981
rect 178944 536593 179014 537025
rect 182244 537549 182314 537981
rect 182244 536873 182314 537305
rect 185544 537549 185614 537981
rect 185544 537013 185614 537445
rect 188844 537549 188914 537981
rect 188844 536917 188914 537349
rect 164288 535209 164358 535641
rect 164288 533693 164358 534125
rect 164606 535209 164676 535641
rect 164606 533693 164676 534125
rect 164924 535209 164994 535641
rect 164924 533693 164994 534125
rect 165242 535209 165312 535641
rect 165242 533693 165312 534125
rect 165560 535209 165630 535641
rect 165560 533693 165630 534125
rect 165878 535209 165948 535641
rect 165878 533693 165948 534125
rect 166196 535209 166266 535641
rect 166196 533693 166266 534125
rect 166514 535209 166584 535641
rect 166514 533693 166584 534125
<< ppolyres >>
rect 188844 537349 188914 537549
<< xpolyres >>
rect 164318 536465 164388 537549
rect 164636 536465 164706 537549
rect 164954 536465 165024 537549
rect 165272 536465 165342 537549
rect 165590 536465 165660 537549
rect 165908 536465 165978 537549
rect 166226 536465 166296 537549
rect 166544 536465 166614 537549
rect 168090 536465 168160 537549
rect 168408 536465 168478 537549
rect 168726 536465 168796 537549
rect 169044 536465 169114 537549
rect 171826 536465 171896 537549
rect 172144 536465 172214 537549
rect 175344 536465 175414 537549
rect 178944 537025 179014 537549
rect 182244 537305 182314 537549
rect 185544 537445 185614 537549
rect 164288 534125 164358 535209
rect 164606 534125 164676 535209
rect 164924 534125 164994 535209
rect 165242 534125 165312 535209
rect 165560 534125 165630 535209
rect 165878 534125 165948 535209
rect 166196 534125 166266 535209
rect 166514 534125 166584 535209
<< rmp >>
rect 186951 530370 187047 530379
rect 187089 530370 187185 530379
<< locali >>
rect 164520 541287 166650 541307
rect 164520 541277 164620 541287
rect 164520 539897 164540 541277
rect 164580 541247 164620 541277
rect 166540 541267 166650 541287
rect 166540 541247 166580 541267
rect 164580 541217 166580 541247
rect 164580 539947 164600 541217
rect 164714 541117 164730 541151
rect 164764 541117 164780 541151
rect 165017 541124 165033 541158
rect 165067 541124 165083 541158
rect 165209 541124 165225 541158
rect 165259 541124 165275 541158
rect 165401 541124 165417 541158
rect 165451 541124 165467 541158
rect 165593 541124 165609 541158
rect 165643 541124 165659 541158
rect 165785 541124 165801 541158
rect 165835 541124 165851 541158
rect 165977 541124 165993 541158
rect 166027 541124 166043 541158
rect 166394 541117 166410 541151
rect 166444 541117 166460 541151
rect 164686 541067 164720 541083
rect 164686 540075 164720 540091
rect 164774 541067 164808 541083
rect 164774 540075 164808 540091
rect 164889 541074 164923 541090
rect 164889 540082 164923 540098
rect 164985 541074 165019 541090
rect 164985 540082 165019 540098
rect 165081 541074 165115 541090
rect 165081 540082 165115 540098
rect 165177 541074 165211 541090
rect 165177 540082 165211 540098
rect 165273 541074 165307 541090
rect 165273 540082 165307 540098
rect 165369 541074 165403 541090
rect 165369 540082 165403 540098
rect 165465 541074 165499 541090
rect 165465 540082 165499 540098
rect 165561 541074 165595 541090
rect 165561 540082 165595 540098
rect 165657 541074 165691 541090
rect 165657 540082 165691 540098
rect 165753 541074 165787 541090
rect 165753 540082 165787 540098
rect 165849 541074 165883 541090
rect 165849 540082 165883 540098
rect 165945 541074 165979 541090
rect 165945 540082 165979 540098
rect 166041 541074 166075 541090
rect 166366 541067 166400 541083
rect 166194 540317 166210 540351
rect 166244 540317 166260 540351
rect 166041 540082 166075 540098
rect 166166 540267 166200 540283
rect 166166 540075 166200 540091
rect 166254 540267 166288 540283
rect 166254 540075 166288 540091
rect 166366 540075 166400 540091
rect 166454 541067 166488 541083
rect 166454 540075 166488 540091
rect 166560 540247 166580 541217
rect 166620 540247 166650 541267
rect 166560 540117 166570 540247
rect 166630 540117 166650 540247
rect 164714 540007 164730 540041
rect 164764 540007 164780 540041
rect 164921 540014 164937 540048
rect 164971 540014 164987 540048
rect 165113 540014 165129 540048
rect 165163 540014 165179 540048
rect 165305 540014 165321 540048
rect 165355 540014 165371 540048
rect 165497 540014 165513 540048
rect 165547 540014 165563 540048
rect 165689 540014 165705 540048
rect 165739 540014 165755 540048
rect 165881 540014 165897 540048
rect 165931 540014 165947 540048
rect 166194 540007 166210 540041
rect 166244 540007 166260 540041
rect 166394 540007 166410 540041
rect 166444 540007 166460 540041
rect 166560 539947 166580 540117
rect 164580 539927 166580 539947
rect 164580 539897 164620 539927
rect 164520 539887 164620 539897
rect 166540 539887 166580 539927
rect 166620 539887 166650 540117
rect 164520 539857 166650 539887
rect 168320 541287 170450 541307
rect 168320 541277 168420 541287
rect 168320 539897 168340 541277
rect 168380 541247 168420 541277
rect 170340 541267 170450 541287
rect 170340 541247 170380 541267
rect 168380 541217 170380 541247
rect 168380 539947 168400 541217
rect 168514 541117 168530 541151
rect 168564 541117 168580 541151
rect 168817 541124 168833 541158
rect 168867 541124 168883 541158
rect 169009 541124 169025 541158
rect 169059 541124 169075 541158
rect 169201 541124 169217 541158
rect 169251 541124 169267 541158
rect 169393 541124 169409 541158
rect 169443 541124 169459 541158
rect 169585 541124 169601 541158
rect 169635 541124 169651 541158
rect 169777 541124 169793 541158
rect 169827 541124 169843 541158
rect 170194 541117 170210 541151
rect 170244 541117 170260 541151
rect 168486 541067 168520 541083
rect 168486 540075 168520 540091
rect 168574 541067 168608 541083
rect 168574 540075 168608 540091
rect 168689 541074 168723 541090
rect 168689 540082 168723 540098
rect 168785 541074 168819 541090
rect 168785 540082 168819 540098
rect 168881 541074 168915 541090
rect 168881 540082 168915 540098
rect 168977 541074 169011 541090
rect 168977 540082 169011 540098
rect 169073 541074 169107 541090
rect 169073 540082 169107 540098
rect 169169 541074 169203 541090
rect 169169 540082 169203 540098
rect 169265 541074 169299 541090
rect 169265 540082 169299 540098
rect 169361 541074 169395 541090
rect 169361 540082 169395 540098
rect 169457 541074 169491 541090
rect 169457 540082 169491 540098
rect 169553 541074 169587 541090
rect 169553 540082 169587 540098
rect 169649 541074 169683 541090
rect 169649 540082 169683 540098
rect 169745 541074 169779 541090
rect 169745 540082 169779 540098
rect 169841 541074 169875 541090
rect 170166 541067 170200 541083
rect 169994 540317 170010 540351
rect 170044 540317 170060 540351
rect 169841 540082 169875 540098
rect 169966 540267 170000 540283
rect 169966 540075 170000 540091
rect 170054 540267 170088 540283
rect 170054 540075 170088 540091
rect 170166 540075 170200 540091
rect 170254 541067 170288 541083
rect 170254 540075 170288 540091
rect 170360 540247 170380 541217
rect 170420 540247 170450 541267
rect 170360 540117 170370 540247
rect 170430 540117 170450 540247
rect 168514 540007 168530 540041
rect 168564 540007 168580 540041
rect 168721 540014 168737 540048
rect 168771 540014 168787 540048
rect 168913 540014 168929 540048
rect 168963 540014 168979 540048
rect 169105 540014 169121 540048
rect 169155 540014 169171 540048
rect 169297 540014 169313 540048
rect 169347 540014 169363 540048
rect 169489 540014 169505 540048
rect 169539 540014 169555 540048
rect 169681 540014 169697 540048
rect 169731 540014 169747 540048
rect 169994 540007 170010 540041
rect 170044 540007 170060 540041
rect 170194 540007 170210 540041
rect 170244 540007 170260 540041
rect 170360 539947 170380 540117
rect 168380 539927 170380 539947
rect 168380 539897 168420 539927
rect 168320 539887 168420 539897
rect 170340 539887 170380 539927
rect 170420 539887 170450 540117
rect 168320 539857 170450 539887
rect 172020 541287 174150 541307
rect 172020 541277 172120 541287
rect 172020 539897 172040 541277
rect 172080 541247 172120 541277
rect 174040 541267 174150 541287
rect 174040 541247 174080 541267
rect 172080 541217 174080 541247
rect 172080 539947 172100 541217
rect 172214 541117 172230 541151
rect 172264 541117 172280 541151
rect 172517 541124 172533 541158
rect 172567 541124 172583 541158
rect 172709 541124 172725 541158
rect 172759 541124 172775 541158
rect 172901 541124 172917 541158
rect 172951 541124 172967 541158
rect 173093 541124 173109 541158
rect 173143 541124 173159 541158
rect 173285 541124 173301 541158
rect 173335 541124 173351 541158
rect 173477 541124 173493 541158
rect 173527 541124 173543 541158
rect 173894 541117 173910 541151
rect 173944 541117 173960 541151
rect 172186 541067 172220 541083
rect 172186 540075 172220 540091
rect 172274 541067 172308 541083
rect 172274 540075 172308 540091
rect 172389 541074 172423 541090
rect 172389 540082 172423 540098
rect 172485 541074 172519 541090
rect 172485 540082 172519 540098
rect 172581 541074 172615 541090
rect 172581 540082 172615 540098
rect 172677 541074 172711 541090
rect 172677 540082 172711 540098
rect 172773 541074 172807 541090
rect 172773 540082 172807 540098
rect 172869 541074 172903 541090
rect 172869 540082 172903 540098
rect 172965 541074 172999 541090
rect 172965 540082 172999 540098
rect 173061 541074 173095 541090
rect 173061 540082 173095 540098
rect 173157 541074 173191 541090
rect 173157 540082 173191 540098
rect 173253 541074 173287 541090
rect 173253 540082 173287 540098
rect 173349 541074 173383 541090
rect 173349 540082 173383 540098
rect 173445 541074 173479 541090
rect 173445 540082 173479 540098
rect 173541 541074 173575 541090
rect 173866 541067 173900 541083
rect 173694 540317 173710 540351
rect 173744 540317 173760 540351
rect 173541 540082 173575 540098
rect 173666 540267 173700 540283
rect 173666 540075 173700 540091
rect 173754 540267 173788 540283
rect 173754 540075 173788 540091
rect 173866 540075 173900 540091
rect 173954 541067 173988 541083
rect 173954 540075 173988 540091
rect 174060 540247 174080 541217
rect 174120 540247 174150 541267
rect 174060 540117 174070 540247
rect 174130 540117 174150 540247
rect 172214 540007 172230 540041
rect 172264 540007 172280 540041
rect 172421 540014 172437 540048
rect 172471 540014 172487 540048
rect 172613 540014 172629 540048
rect 172663 540014 172679 540048
rect 172805 540014 172821 540048
rect 172855 540014 172871 540048
rect 172997 540014 173013 540048
rect 173047 540014 173063 540048
rect 173189 540014 173205 540048
rect 173239 540014 173255 540048
rect 173381 540014 173397 540048
rect 173431 540014 173447 540048
rect 173694 540007 173710 540041
rect 173744 540007 173760 540041
rect 173894 540007 173910 540041
rect 173944 540007 173960 540041
rect 174060 539947 174080 540117
rect 172080 539927 174080 539947
rect 172080 539897 172120 539927
rect 172020 539887 172120 539897
rect 174040 539887 174080 539927
rect 174120 539887 174150 540117
rect 172020 539857 174150 539887
rect 175520 541287 177650 541307
rect 175520 541277 175620 541287
rect 175520 539897 175540 541277
rect 175580 541247 175620 541277
rect 177540 541267 177650 541287
rect 177540 541247 177580 541267
rect 175580 541217 177580 541247
rect 175580 539947 175600 541217
rect 175714 541117 175730 541151
rect 175764 541117 175780 541151
rect 176017 541124 176033 541158
rect 176067 541124 176083 541158
rect 176209 541124 176225 541158
rect 176259 541124 176275 541158
rect 176401 541124 176417 541158
rect 176451 541124 176467 541158
rect 176593 541124 176609 541158
rect 176643 541124 176659 541158
rect 176785 541124 176801 541158
rect 176835 541124 176851 541158
rect 176977 541124 176993 541158
rect 177027 541124 177043 541158
rect 177394 541117 177410 541151
rect 177444 541117 177460 541151
rect 175686 541067 175720 541083
rect 175686 540075 175720 540091
rect 175774 541067 175808 541083
rect 175774 540075 175808 540091
rect 175889 541074 175923 541090
rect 175889 540082 175923 540098
rect 175985 541074 176019 541090
rect 175985 540082 176019 540098
rect 176081 541074 176115 541090
rect 176081 540082 176115 540098
rect 176177 541074 176211 541090
rect 176177 540082 176211 540098
rect 176273 541074 176307 541090
rect 176273 540082 176307 540098
rect 176369 541074 176403 541090
rect 176369 540082 176403 540098
rect 176465 541074 176499 541090
rect 176465 540082 176499 540098
rect 176561 541074 176595 541090
rect 176561 540082 176595 540098
rect 176657 541074 176691 541090
rect 176657 540082 176691 540098
rect 176753 541074 176787 541090
rect 176753 540082 176787 540098
rect 176849 541074 176883 541090
rect 176849 540082 176883 540098
rect 176945 541074 176979 541090
rect 176945 540082 176979 540098
rect 177041 541074 177075 541090
rect 177366 541067 177400 541083
rect 177194 540317 177210 540351
rect 177244 540317 177260 540351
rect 177041 540082 177075 540098
rect 177166 540267 177200 540283
rect 177166 540075 177200 540091
rect 177254 540267 177288 540283
rect 177254 540075 177288 540091
rect 177366 540075 177400 540091
rect 177454 541067 177488 541083
rect 177454 540075 177488 540091
rect 177560 540247 177580 541217
rect 177620 540247 177650 541267
rect 177560 540117 177570 540247
rect 177630 540117 177650 540247
rect 175714 540007 175730 540041
rect 175764 540007 175780 540041
rect 175921 540014 175937 540048
rect 175971 540014 175987 540048
rect 176113 540014 176129 540048
rect 176163 540014 176179 540048
rect 176305 540014 176321 540048
rect 176355 540014 176371 540048
rect 176497 540014 176513 540048
rect 176547 540014 176563 540048
rect 176689 540014 176705 540048
rect 176739 540014 176755 540048
rect 176881 540014 176897 540048
rect 176931 540014 176947 540048
rect 177194 540007 177210 540041
rect 177244 540007 177260 540041
rect 177394 540007 177410 540041
rect 177444 540007 177460 540041
rect 177560 539947 177580 540117
rect 175580 539927 177580 539947
rect 175580 539897 175620 539927
rect 175520 539887 175620 539897
rect 177540 539887 177580 539927
rect 177620 539887 177650 540117
rect 175520 539857 177650 539887
rect 179120 541287 181250 541307
rect 179120 541277 179220 541287
rect 179120 539897 179140 541277
rect 179180 541247 179220 541277
rect 181140 541267 181250 541287
rect 181140 541247 181180 541267
rect 179180 541217 181180 541247
rect 179180 539947 179200 541217
rect 179314 541117 179330 541151
rect 179364 541117 179380 541151
rect 179617 541124 179633 541158
rect 179667 541124 179683 541158
rect 179809 541124 179825 541158
rect 179859 541124 179875 541158
rect 180001 541124 180017 541158
rect 180051 541124 180067 541158
rect 180193 541124 180209 541158
rect 180243 541124 180259 541158
rect 180385 541124 180401 541158
rect 180435 541124 180451 541158
rect 180577 541124 180593 541158
rect 180627 541124 180643 541158
rect 180994 541117 181010 541151
rect 181044 541117 181060 541151
rect 179286 541067 179320 541083
rect 179286 540075 179320 540091
rect 179374 541067 179408 541083
rect 179374 540075 179408 540091
rect 179489 541074 179523 541090
rect 179489 540082 179523 540098
rect 179585 541074 179619 541090
rect 179585 540082 179619 540098
rect 179681 541074 179715 541090
rect 179681 540082 179715 540098
rect 179777 541074 179811 541090
rect 179777 540082 179811 540098
rect 179873 541074 179907 541090
rect 179873 540082 179907 540098
rect 179969 541074 180003 541090
rect 179969 540082 180003 540098
rect 180065 541074 180099 541090
rect 180065 540082 180099 540098
rect 180161 541074 180195 541090
rect 180161 540082 180195 540098
rect 180257 541074 180291 541090
rect 180257 540082 180291 540098
rect 180353 541074 180387 541090
rect 180353 540082 180387 540098
rect 180449 541074 180483 541090
rect 180449 540082 180483 540098
rect 180545 541074 180579 541090
rect 180545 540082 180579 540098
rect 180641 541074 180675 541090
rect 180966 541067 181000 541083
rect 180794 540317 180810 540351
rect 180844 540317 180860 540351
rect 180641 540082 180675 540098
rect 180766 540267 180800 540283
rect 180766 540075 180800 540091
rect 180854 540267 180888 540283
rect 180854 540075 180888 540091
rect 180966 540075 181000 540091
rect 181054 541067 181088 541083
rect 181054 540075 181088 540091
rect 181160 540247 181180 541217
rect 181220 540247 181250 541267
rect 181160 540117 181170 540247
rect 181230 540117 181250 540247
rect 179314 540007 179330 540041
rect 179364 540007 179380 540041
rect 179521 540014 179537 540048
rect 179571 540014 179587 540048
rect 179713 540014 179729 540048
rect 179763 540014 179779 540048
rect 179905 540014 179921 540048
rect 179955 540014 179971 540048
rect 180097 540014 180113 540048
rect 180147 540014 180163 540048
rect 180289 540014 180305 540048
rect 180339 540014 180355 540048
rect 180481 540014 180497 540048
rect 180531 540014 180547 540048
rect 180794 540007 180810 540041
rect 180844 540007 180860 540041
rect 180994 540007 181010 540041
rect 181044 540007 181060 540041
rect 181160 539947 181180 540117
rect 179180 539927 181180 539947
rect 179180 539897 179220 539927
rect 179120 539887 179220 539897
rect 181140 539887 181180 539927
rect 181220 539887 181250 540117
rect 179120 539857 181250 539887
rect 182420 541287 184550 541307
rect 182420 541277 182520 541287
rect 182420 539897 182440 541277
rect 182480 541247 182520 541277
rect 184440 541267 184550 541287
rect 184440 541247 184480 541267
rect 182480 541217 184480 541247
rect 182480 539947 182500 541217
rect 182614 541117 182630 541151
rect 182664 541117 182680 541151
rect 182917 541124 182933 541158
rect 182967 541124 182983 541158
rect 183109 541124 183125 541158
rect 183159 541124 183175 541158
rect 183301 541124 183317 541158
rect 183351 541124 183367 541158
rect 183493 541124 183509 541158
rect 183543 541124 183559 541158
rect 183685 541124 183701 541158
rect 183735 541124 183751 541158
rect 183877 541124 183893 541158
rect 183927 541124 183943 541158
rect 184294 541117 184310 541151
rect 184344 541117 184360 541151
rect 182586 541067 182620 541083
rect 182586 540075 182620 540091
rect 182674 541067 182708 541083
rect 182674 540075 182708 540091
rect 182789 541074 182823 541090
rect 182789 540082 182823 540098
rect 182885 541074 182919 541090
rect 182885 540082 182919 540098
rect 182981 541074 183015 541090
rect 182981 540082 183015 540098
rect 183077 541074 183111 541090
rect 183077 540082 183111 540098
rect 183173 541074 183207 541090
rect 183173 540082 183207 540098
rect 183269 541074 183303 541090
rect 183269 540082 183303 540098
rect 183365 541074 183399 541090
rect 183365 540082 183399 540098
rect 183461 541074 183495 541090
rect 183461 540082 183495 540098
rect 183557 541074 183591 541090
rect 183557 540082 183591 540098
rect 183653 541074 183687 541090
rect 183653 540082 183687 540098
rect 183749 541074 183783 541090
rect 183749 540082 183783 540098
rect 183845 541074 183879 541090
rect 183845 540082 183879 540098
rect 183941 541074 183975 541090
rect 184266 541067 184300 541083
rect 184094 540317 184110 540351
rect 184144 540317 184160 540351
rect 183941 540082 183975 540098
rect 184066 540267 184100 540283
rect 184066 540075 184100 540091
rect 184154 540267 184188 540283
rect 184154 540075 184188 540091
rect 184266 540075 184300 540091
rect 184354 541067 184388 541083
rect 184354 540075 184388 540091
rect 184460 540247 184480 541217
rect 184520 540247 184550 541267
rect 184460 540117 184470 540247
rect 184530 540117 184550 540247
rect 182614 540007 182630 540041
rect 182664 540007 182680 540041
rect 182821 540014 182837 540048
rect 182871 540014 182887 540048
rect 183013 540014 183029 540048
rect 183063 540014 183079 540048
rect 183205 540014 183221 540048
rect 183255 540014 183271 540048
rect 183397 540014 183413 540048
rect 183447 540014 183463 540048
rect 183589 540014 183605 540048
rect 183639 540014 183655 540048
rect 183781 540014 183797 540048
rect 183831 540014 183847 540048
rect 184094 540007 184110 540041
rect 184144 540007 184160 540041
rect 184294 540007 184310 540041
rect 184344 540007 184360 540041
rect 184460 539947 184480 540117
rect 182480 539927 184480 539947
rect 182480 539897 182520 539927
rect 182420 539887 182520 539897
rect 184440 539887 184480 539927
rect 184520 539887 184550 540117
rect 182420 539857 184550 539887
rect 185720 541287 187850 541307
rect 185720 541277 185820 541287
rect 185720 539897 185740 541277
rect 185780 541247 185820 541277
rect 187740 541267 187850 541287
rect 187740 541247 187780 541267
rect 185780 541217 187780 541247
rect 185780 539947 185800 541217
rect 185914 541117 185930 541151
rect 185964 541117 185980 541151
rect 186217 541124 186233 541158
rect 186267 541124 186283 541158
rect 186409 541124 186425 541158
rect 186459 541124 186475 541158
rect 186601 541124 186617 541158
rect 186651 541124 186667 541158
rect 186793 541124 186809 541158
rect 186843 541124 186859 541158
rect 186985 541124 187001 541158
rect 187035 541124 187051 541158
rect 187177 541124 187193 541158
rect 187227 541124 187243 541158
rect 187594 541117 187610 541151
rect 187644 541117 187660 541151
rect 185886 541067 185920 541083
rect 185886 540075 185920 540091
rect 185974 541067 186008 541083
rect 185974 540075 186008 540091
rect 186089 541074 186123 541090
rect 186089 540082 186123 540098
rect 186185 541074 186219 541090
rect 186185 540082 186219 540098
rect 186281 541074 186315 541090
rect 186281 540082 186315 540098
rect 186377 541074 186411 541090
rect 186377 540082 186411 540098
rect 186473 541074 186507 541090
rect 186473 540082 186507 540098
rect 186569 541074 186603 541090
rect 186569 540082 186603 540098
rect 186665 541074 186699 541090
rect 186665 540082 186699 540098
rect 186761 541074 186795 541090
rect 186761 540082 186795 540098
rect 186857 541074 186891 541090
rect 186857 540082 186891 540098
rect 186953 541074 186987 541090
rect 186953 540082 186987 540098
rect 187049 541074 187083 541090
rect 187049 540082 187083 540098
rect 187145 541074 187179 541090
rect 187145 540082 187179 540098
rect 187241 541074 187275 541090
rect 187566 541067 187600 541083
rect 187394 540317 187410 540351
rect 187444 540317 187460 540351
rect 187241 540082 187275 540098
rect 187366 540267 187400 540283
rect 187366 540075 187400 540091
rect 187454 540267 187488 540283
rect 187454 540075 187488 540091
rect 187566 540075 187600 540091
rect 187654 541067 187688 541083
rect 187654 540075 187688 540091
rect 187760 540247 187780 541217
rect 187820 540247 187850 541267
rect 187760 540117 187770 540247
rect 187830 540117 187850 540247
rect 185914 540007 185930 540041
rect 185964 540007 185980 540041
rect 186121 540014 186137 540048
rect 186171 540014 186187 540048
rect 186313 540014 186329 540048
rect 186363 540014 186379 540048
rect 186505 540014 186521 540048
rect 186555 540014 186571 540048
rect 186697 540014 186713 540048
rect 186747 540014 186763 540048
rect 186889 540014 186905 540048
rect 186939 540014 186955 540048
rect 187081 540014 187097 540048
rect 187131 540014 187147 540048
rect 187394 540007 187410 540041
rect 187444 540007 187460 540041
rect 187594 540007 187610 540041
rect 187644 540007 187660 540041
rect 187760 539947 187780 540117
rect 185780 539927 187780 539947
rect 185780 539897 185820 539927
rect 185720 539887 185820 539897
rect 187740 539887 187780 539927
rect 187820 539887 187850 540117
rect 185720 539857 187850 539887
rect 189020 541287 191150 541307
rect 189020 541277 189120 541287
rect 189020 539897 189040 541277
rect 189080 541247 189120 541277
rect 191040 541267 191150 541287
rect 191040 541247 191080 541267
rect 189080 541217 191080 541247
rect 189080 539947 189100 541217
rect 189214 541117 189230 541151
rect 189264 541117 189280 541151
rect 189517 541124 189533 541158
rect 189567 541124 189583 541158
rect 189709 541124 189725 541158
rect 189759 541124 189775 541158
rect 189901 541124 189917 541158
rect 189951 541124 189967 541158
rect 190093 541124 190109 541158
rect 190143 541124 190159 541158
rect 190285 541124 190301 541158
rect 190335 541124 190351 541158
rect 190477 541124 190493 541158
rect 190527 541124 190543 541158
rect 190894 541117 190910 541151
rect 190944 541117 190960 541151
rect 189186 541067 189220 541083
rect 189186 540075 189220 540091
rect 189274 541067 189308 541083
rect 189274 540075 189308 540091
rect 189389 541074 189423 541090
rect 189389 540082 189423 540098
rect 189485 541074 189519 541090
rect 189485 540082 189519 540098
rect 189581 541074 189615 541090
rect 189581 540082 189615 540098
rect 189677 541074 189711 541090
rect 189677 540082 189711 540098
rect 189773 541074 189807 541090
rect 189773 540082 189807 540098
rect 189869 541074 189903 541090
rect 189869 540082 189903 540098
rect 189965 541074 189999 541090
rect 189965 540082 189999 540098
rect 190061 541074 190095 541090
rect 190061 540082 190095 540098
rect 190157 541074 190191 541090
rect 190157 540082 190191 540098
rect 190253 541074 190287 541090
rect 190253 540082 190287 540098
rect 190349 541074 190383 541090
rect 190349 540082 190383 540098
rect 190445 541074 190479 541090
rect 190445 540082 190479 540098
rect 190541 541074 190575 541090
rect 190866 541067 190900 541083
rect 190694 540317 190710 540351
rect 190744 540317 190760 540351
rect 190541 540082 190575 540098
rect 190666 540267 190700 540283
rect 190666 540075 190700 540091
rect 190754 540267 190788 540283
rect 190754 540075 190788 540091
rect 190866 540075 190900 540091
rect 190954 541067 190988 541083
rect 190954 540075 190988 540091
rect 191060 540247 191080 541217
rect 191120 540247 191150 541267
rect 191060 540117 191070 540247
rect 191130 540117 191150 540247
rect 189214 540007 189230 540041
rect 189264 540007 189280 540041
rect 189421 540014 189437 540048
rect 189471 540014 189487 540048
rect 189613 540014 189629 540048
rect 189663 540014 189679 540048
rect 189805 540014 189821 540048
rect 189855 540014 189871 540048
rect 189997 540014 190013 540048
rect 190047 540014 190063 540048
rect 190189 540014 190205 540048
rect 190239 540014 190255 540048
rect 190381 540014 190397 540048
rect 190431 540014 190447 540048
rect 190694 540007 190710 540041
rect 190744 540007 190760 540041
rect 190894 540007 190910 540041
rect 190944 540007 190960 540041
rect 191060 539947 191080 540117
rect 189080 539927 191080 539947
rect 189080 539897 189120 539927
rect 189020 539887 189120 539897
rect 191040 539887 191080 539927
rect 191120 539887 191150 540117
rect 191810 540277 191990 540293
rect 191810 540081 191990 540097
rect 189020 539857 191150 539887
rect 164520 539767 166640 539787
rect 164520 539747 164620 539767
rect 157630 538737 162870 538757
rect 157630 538697 157710 538737
rect 162770 538697 162870 538737
rect 157630 538677 162870 538697
rect 157630 538657 157710 538677
rect 157630 537997 157650 538657
rect 157690 538037 157710 538657
rect 158712 538467 158728 538501
rect 158896 538467 158912 538501
rect 159088 538467 159104 538501
rect 159272 538467 159288 538501
rect 159346 538467 159362 538501
rect 159530 538467 159546 538501
rect 159604 538467 159620 538501
rect 159788 538467 159804 538501
rect 159862 538467 159878 538501
rect 160046 538467 160062 538501
rect 160120 538467 160136 538501
rect 160304 538467 160320 538501
rect 160378 538467 160394 538501
rect 160562 538467 160578 538501
rect 160636 538467 160652 538501
rect 160820 538467 160836 538501
rect 160894 538467 160910 538501
rect 161078 538467 161094 538501
rect 161152 538467 161168 538501
rect 161336 538467 161352 538501
rect 161532 538467 161548 538501
rect 161716 538467 161732 538501
rect 161932 538467 161948 538501
rect 162116 538467 162132 538501
rect 162312 538467 162328 538501
rect 162496 538467 162512 538501
rect 158666 538417 158700 538433
rect 158666 538225 158700 538241
rect 158924 538417 158958 538433
rect 158924 538225 158958 538241
rect 159042 538417 159076 538433
rect 159042 538225 159076 538241
rect 159300 538417 159334 538433
rect 159300 538225 159334 538241
rect 159558 538417 159592 538433
rect 159558 538225 159592 538241
rect 159816 538417 159850 538433
rect 159816 538225 159850 538241
rect 160074 538417 160108 538433
rect 160074 538225 160108 538241
rect 160332 538417 160366 538433
rect 160332 538225 160366 538241
rect 160590 538417 160624 538433
rect 160590 538225 160624 538241
rect 160848 538417 160882 538433
rect 160848 538225 160882 538241
rect 161106 538417 161140 538433
rect 161106 538225 161140 538241
rect 161364 538417 161398 538433
rect 161364 538225 161398 538241
rect 161486 538417 161520 538433
rect 161486 538225 161520 538241
rect 161744 538417 161778 538433
rect 161744 538225 161778 538241
rect 161886 538417 161920 538433
rect 161886 538225 161920 538241
rect 162144 538417 162178 538433
rect 162144 538225 162178 538241
rect 162266 538417 162300 538433
rect 162266 538225 162300 538241
rect 162524 538417 162558 538433
rect 162524 538225 162558 538241
rect 158712 538157 158728 538191
rect 158896 538157 158912 538191
rect 159088 538157 159104 538191
rect 159272 538157 159288 538191
rect 159346 538157 159362 538191
rect 159530 538157 159546 538191
rect 159604 538157 159620 538191
rect 159788 538157 159804 538191
rect 159862 538157 159878 538191
rect 160046 538157 160062 538191
rect 160120 538157 160136 538191
rect 160304 538157 160320 538191
rect 160378 538157 160394 538191
rect 160562 538157 160578 538191
rect 160636 538157 160652 538191
rect 160820 538157 160836 538191
rect 160894 538157 160910 538191
rect 161078 538157 161094 538191
rect 161152 538157 161168 538191
rect 161336 538157 161352 538191
rect 161532 538157 161548 538191
rect 161716 538157 161732 538191
rect 161932 538157 161948 538191
rect 162116 538157 162132 538191
rect 162312 538157 162328 538191
rect 162496 538157 162512 538191
rect 162790 538037 162810 538677
rect 162850 538037 162870 538677
rect 164520 538347 164540 539747
rect 164580 539727 164620 539747
rect 166540 539747 166640 539767
rect 166540 539727 166580 539747
rect 164580 539707 166580 539727
rect 164580 538387 164600 539707
rect 166540 539687 166580 539707
rect 164698 539604 164714 539638
rect 164748 539604 164764 539638
rect 165021 539611 165037 539645
rect 165071 539611 165087 539645
rect 165213 539611 165229 539645
rect 165263 539611 165279 539645
rect 165405 539611 165421 539645
rect 165455 539611 165471 539645
rect 165597 539611 165613 539645
rect 165647 539611 165663 539645
rect 165789 539611 165805 539645
rect 165839 539611 165855 539645
rect 165981 539611 165997 539645
rect 166031 539611 166047 539645
rect 166198 539604 166214 539638
rect 166248 539604 166264 539638
rect 166398 539604 166414 539638
rect 166448 539604 166464 539638
rect 164670 539545 164704 539561
rect 164670 538553 164704 538569
rect 164758 539545 164792 539561
rect 164758 538553 164792 538569
rect 164893 539552 164927 539568
rect 164893 538560 164927 538576
rect 164989 539552 165023 539568
rect 164989 538560 165023 538576
rect 165085 539552 165119 539568
rect 165085 538560 165119 538576
rect 165181 539552 165215 539568
rect 165181 538560 165215 538576
rect 165277 539552 165311 539568
rect 165277 538560 165311 538576
rect 165373 539552 165407 539568
rect 165373 538560 165407 538576
rect 165469 539552 165503 539568
rect 165469 538560 165503 538576
rect 165565 539552 165599 539568
rect 165565 538560 165599 538576
rect 165661 539552 165695 539568
rect 165661 538560 165695 538576
rect 165757 539552 165791 539568
rect 165757 538560 165791 538576
rect 165853 539552 165887 539568
rect 165853 538560 165887 538576
rect 165949 539552 165983 539568
rect 165949 538560 165983 538576
rect 166045 539552 166079 539568
rect 166170 539545 166204 539561
rect 166170 538953 166204 538969
rect 166258 539545 166292 539561
rect 166258 538953 166292 538969
rect 166370 539545 166404 539561
rect 166198 538876 166214 538910
rect 166248 538876 166264 538910
rect 166045 538560 166079 538576
rect 166370 538553 166404 538569
rect 166458 539545 166492 539561
rect 166458 538553 166492 538569
rect 166560 539297 166580 539687
rect 166560 539207 166570 539297
rect 164698 538476 164714 538510
rect 164748 538476 164764 538510
rect 164925 538483 164941 538517
rect 164975 538483 164991 538517
rect 165117 538483 165133 538517
rect 165167 538483 165183 538517
rect 165309 538483 165325 538517
rect 165359 538483 165375 538517
rect 165501 538483 165517 538517
rect 165551 538483 165567 538517
rect 165693 538483 165709 538517
rect 165743 538483 165759 538517
rect 165885 538483 165901 538517
rect 165935 538483 165951 538517
rect 166398 538476 166414 538510
rect 166448 538476 166464 538510
rect 166560 538387 166580 539207
rect 164580 538367 166580 538387
rect 164580 538347 164620 538367
rect 164520 538327 164620 538347
rect 166540 538347 166580 538367
rect 166620 538347 166640 539747
rect 166540 538327 166640 538347
rect 164520 538307 166640 538327
rect 168320 539767 170440 539787
rect 168320 539747 168420 539767
rect 168320 538347 168340 539747
rect 168380 539727 168420 539747
rect 170340 539747 170440 539767
rect 170340 539727 170380 539747
rect 168380 539707 170380 539727
rect 168380 538387 168400 539707
rect 170340 539687 170380 539707
rect 168498 539604 168514 539638
rect 168548 539604 168564 539638
rect 168821 539611 168837 539645
rect 168871 539611 168887 539645
rect 169013 539611 169029 539645
rect 169063 539611 169079 539645
rect 169205 539611 169221 539645
rect 169255 539611 169271 539645
rect 169397 539611 169413 539645
rect 169447 539611 169463 539645
rect 169589 539611 169605 539645
rect 169639 539611 169655 539645
rect 169781 539611 169797 539645
rect 169831 539611 169847 539645
rect 169998 539604 170014 539638
rect 170048 539604 170064 539638
rect 170198 539604 170214 539638
rect 170248 539604 170264 539638
rect 168470 539545 168504 539561
rect 168470 538553 168504 538569
rect 168558 539545 168592 539561
rect 168558 538553 168592 538569
rect 168693 539552 168727 539568
rect 168693 538560 168727 538576
rect 168789 539552 168823 539568
rect 168789 538560 168823 538576
rect 168885 539552 168919 539568
rect 168885 538560 168919 538576
rect 168981 539552 169015 539568
rect 168981 538560 169015 538576
rect 169077 539552 169111 539568
rect 169077 538560 169111 538576
rect 169173 539552 169207 539568
rect 169173 538560 169207 538576
rect 169269 539552 169303 539568
rect 169269 538560 169303 538576
rect 169365 539552 169399 539568
rect 169365 538560 169399 538576
rect 169461 539552 169495 539568
rect 169461 538560 169495 538576
rect 169557 539552 169591 539568
rect 169557 538560 169591 538576
rect 169653 539552 169687 539568
rect 169653 538560 169687 538576
rect 169749 539552 169783 539568
rect 169749 538560 169783 538576
rect 169845 539552 169879 539568
rect 169970 539545 170004 539561
rect 169970 538953 170004 538969
rect 170058 539545 170092 539561
rect 170058 538953 170092 538969
rect 170170 539545 170204 539561
rect 169998 538876 170014 538910
rect 170048 538876 170064 538910
rect 169845 538560 169879 538576
rect 170170 538553 170204 538569
rect 170258 539545 170292 539561
rect 170258 538553 170292 538569
rect 170360 539297 170380 539687
rect 170360 539207 170370 539297
rect 168498 538476 168514 538510
rect 168548 538476 168564 538510
rect 168725 538483 168741 538517
rect 168775 538483 168791 538517
rect 168917 538483 168933 538517
rect 168967 538483 168983 538517
rect 169109 538483 169125 538517
rect 169159 538483 169175 538517
rect 169301 538483 169317 538517
rect 169351 538483 169367 538517
rect 169493 538483 169509 538517
rect 169543 538483 169559 538517
rect 169685 538483 169701 538517
rect 169735 538483 169751 538517
rect 170198 538476 170214 538510
rect 170248 538476 170264 538510
rect 170360 538387 170380 539207
rect 168380 538367 170380 538387
rect 168380 538347 168420 538367
rect 168320 538327 168420 538347
rect 170340 538347 170380 538367
rect 170420 538347 170440 539747
rect 170340 538327 170440 538347
rect 168320 538307 170440 538327
rect 172020 539767 174140 539787
rect 172020 539747 172120 539767
rect 172020 538347 172040 539747
rect 172080 539727 172120 539747
rect 174040 539747 174140 539767
rect 174040 539727 174080 539747
rect 172080 539707 174080 539727
rect 172080 538387 172100 539707
rect 174040 539687 174080 539707
rect 172198 539604 172214 539638
rect 172248 539604 172264 539638
rect 172521 539611 172537 539645
rect 172571 539611 172587 539645
rect 172713 539611 172729 539645
rect 172763 539611 172779 539645
rect 172905 539611 172921 539645
rect 172955 539611 172971 539645
rect 173097 539611 173113 539645
rect 173147 539611 173163 539645
rect 173289 539611 173305 539645
rect 173339 539611 173355 539645
rect 173481 539611 173497 539645
rect 173531 539611 173547 539645
rect 173698 539604 173714 539638
rect 173748 539604 173764 539638
rect 173898 539604 173914 539638
rect 173948 539604 173964 539638
rect 172170 539545 172204 539561
rect 172170 538553 172204 538569
rect 172258 539545 172292 539561
rect 172258 538553 172292 538569
rect 172393 539552 172427 539568
rect 172393 538560 172427 538576
rect 172489 539552 172523 539568
rect 172489 538560 172523 538576
rect 172585 539552 172619 539568
rect 172585 538560 172619 538576
rect 172681 539552 172715 539568
rect 172681 538560 172715 538576
rect 172777 539552 172811 539568
rect 172777 538560 172811 538576
rect 172873 539552 172907 539568
rect 172873 538560 172907 538576
rect 172969 539552 173003 539568
rect 172969 538560 173003 538576
rect 173065 539552 173099 539568
rect 173065 538560 173099 538576
rect 173161 539552 173195 539568
rect 173161 538560 173195 538576
rect 173257 539552 173291 539568
rect 173257 538560 173291 538576
rect 173353 539552 173387 539568
rect 173353 538560 173387 538576
rect 173449 539552 173483 539568
rect 173449 538560 173483 538576
rect 173545 539552 173579 539568
rect 173670 539545 173704 539561
rect 173670 538953 173704 538969
rect 173758 539545 173792 539561
rect 173758 538953 173792 538969
rect 173870 539545 173904 539561
rect 173698 538876 173714 538910
rect 173748 538876 173764 538910
rect 173545 538560 173579 538576
rect 173870 538553 173904 538569
rect 173958 539545 173992 539561
rect 173958 538553 173992 538569
rect 174060 539297 174080 539687
rect 174060 539207 174070 539297
rect 172198 538476 172214 538510
rect 172248 538476 172264 538510
rect 172425 538483 172441 538517
rect 172475 538483 172491 538517
rect 172617 538483 172633 538517
rect 172667 538483 172683 538517
rect 172809 538483 172825 538517
rect 172859 538483 172875 538517
rect 173001 538483 173017 538517
rect 173051 538483 173067 538517
rect 173193 538483 173209 538517
rect 173243 538483 173259 538517
rect 173385 538483 173401 538517
rect 173435 538483 173451 538517
rect 173898 538476 173914 538510
rect 173948 538476 173964 538510
rect 174060 538387 174080 539207
rect 172080 538367 174080 538387
rect 172080 538347 172120 538367
rect 172020 538327 172120 538347
rect 174040 538347 174080 538367
rect 174120 538347 174140 539747
rect 174040 538327 174140 538347
rect 172020 538307 174140 538327
rect 175520 539767 177640 539787
rect 175520 539747 175620 539767
rect 175520 538347 175540 539747
rect 175580 539727 175620 539747
rect 177540 539747 177640 539767
rect 177540 539727 177580 539747
rect 175580 539707 177580 539727
rect 175580 538387 175600 539707
rect 177540 539687 177580 539707
rect 175698 539604 175714 539638
rect 175748 539604 175764 539638
rect 176021 539611 176037 539645
rect 176071 539611 176087 539645
rect 176213 539611 176229 539645
rect 176263 539611 176279 539645
rect 176405 539611 176421 539645
rect 176455 539611 176471 539645
rect 176597 539611 176613 539645
rect 176647 539611 176663 539645
rect 176789 539611 176805 539645
rect 176839 539611 176855 539645
rect 176981 539611 176997 539645
rect 177031 539611 177047 539645
rect 177198 539604 177214 539638
rect 177248 539604 177264 539638
rect 177398 539604 177414 539638
rect 177448 539604 177464 539638
rect 175670 539545 175704 539561
rect 175670 538553 175704 538569
rect 175758 539545 175792 539561
rect 175758 538553 175792 538569
rect 175893 539552 175927 539568
rect 175893 538560 175927 538576
rect 175989 539552 176023 539568
rect 175989 538560 176023 538576
rect 176085 539552 176119 539568
rect 176085 538560 176119 538576
rect 176181 539552 176215 539568
rect 176181 538560 176215 538576
rect 176277 539552 176311 539568
rect 176277 538560 176311 538576
rect 176373 539552 176407 539568
rect 176373 538560 176407 538576
rect 176469 539552 176503 539568
rect 176469 538560 176503 538576
rect 176565 539552 176599 539568
rect 176565 538560 176599 538576
rect 176661 539552 176695 539568
rect 176661 538560 176695 538576
rect 176757 539552 176791 539568
rect 176757 538560 176791 538576
rect 176853 539552 176887 539568
rect 176853 538560 176887 538576
rect 176949 539552 176983 539568
rect 176949 538560 176983 538576
rect 177045 539552 177079 539568
rect 177170 539545 177204 539561
rect 177170 538953 177204 538969
rect 177258 539545 177292 539561
rect 177258 538953 177292 538969
rect 177370 539545 177404 539561
rect 177198 538876 177214 538910
rect 177248 538876 177264 538910
rect 177045 538560 177079 538576
rect 177370 538553 177404 538569
rect 177458 539545 177492 539561
rect 177458 538553 177492 538569
rect 177560 539297 177580 539687
rect 177560 539207 177570 539297
rect 175698 538476 175714 538510
rect 175748 538476 175764 538510
rect 175925 538483 175941 538517
rect 175975 538483 175991 538517
rect 176117 538483 176133 538517
rect 176167 538483 176183 538517
rect 176309 538483 176325 538517
rect 176359 538483 176375 538517
rect 176501 538483 176517 538517
rect 176551 538483 176567 538517
rect 176693 538483 176709 538517
rect 176743 538483 176759 538517
rect 176885 538483 176901 538517
rect 176935 538483 176951 538517
rect 177398 538476 177414 538510
rect 177448 538476 177464 538510
rect 177560 538387 177580 539207
rect 175580 538367 177580 538387
rect 175580 538347 175620 538367
rect 175520 538327 175620 538347
rect 177540 538347 177580 538367
rect 177620 538347 177640 539747
rect 177540 538327 177640 538347
rect 175520 538307 177640 538327
rect 179120 539767 181240 539787
rect 179120 539747 179220 539767
rect 179120 538347 179140 539747
rect 179180 539727 179220 539747
rect 181140 539747 181240 539767
rect 181140 539727 181180 539747
rect 179180 539707 181180 539727
rect 179180 538387 179200 539707
rect 181140 539687 181180 539707
rect 179298 539604 179314 539638
rect 179348 539604 179364 539638
rect 179621 539611 179637 539645
rect 179671 539611 179687 539645
rect 179813 539611 179829 539645
rect 179863 539611 179879 539645
rect 180005 539611 180021 539645
rect 180055 539611 180071 539645
rect 180197 539611 180213 539645
rect 180247 539611 180263 539645
rect 180389 539611 180405 539645
rect 180439 539611 180455 539645
rect 180581 539611 180597 539645
rect 180631 539611 180647 539645
rect 180798 539604 180814 539638
rect 180848 539604 180864 539638
rect 180998 539604 181014 539638
rect 181048 539604 181064 539638
rect 179270 539545 179304 539561
rect 179270 538553 179304 538569
rect 179358 539545 179392 539561
rect 179358 538553 179392 538569
rect 179493 539552 179527 539568
rect 179493 538560 179527 538576
rect 179589 539552 179623 539568
rect 179589 538560 179623 538576
rect 179685 539552 179719 539568
rect 179685 538560 179719 538576
rect 179781 539552 179815 539568
rect 179781 538560 179815 538576
rect 179877 539552 179911 539568
rect 179877 538560 179911 538576
rect 179973 539552 180007 539568
rect 179973 538560 180007 538576
rect 180069 539552 180103 539568
rect 180069 538560 180103 538576
rect 180165 539552 180199 539568
rect 180165 538560 180199 538576
rect 180261 539552 180295 539568
rect 180261 538560 180295 538576
rect 180357 539552 180391 539568
rect 180357 538560 180391 538576
rect 180453 539552 180487 539568
rect 180453 538560 180487 538576
rect 180549 539552 180583 539568
rect 180549 538560 180583 538576
rect 180645 539552 180679 539568
rect 180770 539545 180804 539561
rect 180770 538953 180804 538969
rect 180858 539545 180892 539561
rect 180858 538953 180892 538969
rect 180970 539545 181004 539561
rect 180798 538876 180814 538910
rect 180848 538876 180864 538910
rect 180645 538560 180679 538576
rect 180970 538553 181004 538569
rect 181058 539545 181092 539561
rect 181058 538553 181092 538569
rect 181160 539297 181180 539687
rect 181160 539207 181170 539297
rect 179298 538476 179314 538510
rect 179348 538476 179364 538510
rect 179525 538483 179541 538517
rect 179575 538483 179591 538517
rect 179717 538483 179733 538517
rect 179767 538483 179783 538517
rect 179909 538483 179925 538517
rect 179959 538483 179975 538517
rect 180101 538483 180117 538517
rect 180151 538483 180167 538517
rect 180293 538483 180309 538517
rect 180343 538483 180359 538517
rect 180485 538483 180501 538517
rect 180535 538483 180551 538517
rect 180998 538476 181014 538510
rect 181048 538476 181064 538510
rect 181160 538387 181180 539207
rect 179180 538367 181180 538387
rect 179180 538347 179220 538367
rect 179120 538327 179220 538347
rect 181140 538347 181180 538367
rect 181220 538347 181240 539747
rect 181140 538327 181240 538347
rect 179120 538307 181240 538327
rect 182420 539767 184540 539787
rect 182420 539747 182520 539767
rect 182420 538347 182440 539747
rect 182480 539727 182520 539747
rect 184440 539747 184540 539767
rect 184440 539727 184480 539747
rect 182480 539707 184480 539727
rect 182480 538387 182500 539707
rect 184440 539687 184480 539707
rect 182598 539604 182614 539638
rect 182648 539604 182664 539638
rect 182921 539611 182937 539645
rect 182971 539611 182987 539645
rect 183113 539611 183129 539645
rect 183163 539611 183179 539645
rect 183305 539611 183321 539645
rect 183355 539611 183371 539645
rect 183497 539611 183513 539645
rect 183547 539611 183563 539645
rect 183689 539611 183705 539645
rect 183739 539611 183755 539645
rect 183881 539611 183897 539645
rect 183931 539611 183947 539645
rect 184098 539604 184114 539638
rect 184148 539604 184164 539638
rect 184298 539604 184314 539638
rect 184348 539604 184364 539638
rect 182570 539545 182604 539561
rect 182570 538553 182604 538569
rect 182658 539545 182692 539561
rect 182658 538553 182692 538569
rect 182793 539552 182827 539568
rect 182793 538560 182827 538576
rect 182889 539552 182923 539568
rect 182889 538560 182923 538576
rect 182985 539552 183019 539568
rect 182985 538560 183019 538576
rect 183081 539552 183115 539568
rect 183081 538560 183115 538576
rect 183177 539552 183211 539568
rect 183177 538560 183211 538576
rect 183273 539552 183307 539568
rect 183273 538560 183307 538576
rect 183369 539552 183403 539568
rect 183369 538560 183403 538576
rect 183465 539552 183499 539568
rect 183465 538560 183499 538576
rect 183561 539552 183595 539568
rect 183561 538560 183595 538576
rect 183657 539552 183691 539568
rect 183657 538560 183691 538576
rect 183753 539552 183787 539568
rect 183753 538560 183787 538576
rect 183849 539552 183883 539568
rect 183849 538560 183883 538576
rect 183945 539552 183979 539568
rect 184070 539545 184104 539561
rect 184070 538953 184104 538969
rect 184158 539545 184192 539561
rect 184158 538953 184192 538969
rect 184270 539545 184304 539561
rect 184098 538876 184114 538910
rect 184148 538876 184164 538910
rect 183945 538560 183979 538576
rect 184270 538553 184304 538569
rect 184358 539545 184392 539561
rect 184358 538553 184392 538569
rect 184460 539297 184480 539687
rect 184460 539207 184470 539297
rect 182598 538476 182614 538510
rect 182648 538476 182664 538510
rect 182825 538483 182841 538517
rect 182875 538483 182891 538517
rect 183017 538483 183033 538517
rect 183067 538483 183083 538517
rect 183209 538483 183225 538517
rect 183259 538483 183275 538517
rect 183401 538483 183417 538517
rect 183451 538483 183467 538517
rect 183593 538483 183609 538517
rect 183643 538483 183659 538517
rect 183785 538483 183801 538517
rect 183835 538483 183851 538517
rect 184298 538476 184314 538510
rect 184348 538476 184364 538510
rect 184460 538387 184480 539207
rect 182480 538367 184480 538387
rect 182480 538347 182520 538367
rect 182420 538327 182520 538347
rect 184440 538347 184480 538367
rect 184520 538347 184540 539747
rect 184440 538327 184540 538347
rect 182420 538307 184540 538327
rect 185720 539767 187840 539787
rect 185720 539747 185820 539767
rect 185720 538347 185740 539747
rect 185780 539727 185820 539747
rect 187740 539747 187840 539767
rect 187740 539727 187780 539747
rect 185780 539707 187780 539727
rect 185780 538387 185800 539707
rect 187740 539687 187780 539707
rect 185898 539604 185914 539638
rect 185948 539604 185964 539638
rect 186221 539611 186237 539645
rect 186271 539611 186287 539645
rect 186413 539611 186429 539645
rect 186463 539611 186479 539645
rect 186605 539611 186621 539645
rect 186655 539611 186671 539645
rect 186797 539611 186813 539645
rect 186847 539611 186863 539645
rect 186989 539611 187005 539645
rect 187039 539611 187055 539645
rect 187181 539611 187197 539645
rect 187231 539611 187247 539645
rect 187398 539604 187414 539638
rect 187448 539604 187464 539638
rect 187598 539604 187614 539638
rect 187648 539604 187664 539638
rect 185870 539545 185904 539561
rect 185870 538553 185904 538569
rect 185958 539545 185992 539561
rect 185958 538553 185992 538569
rect 186093 539552 186127 539568
rect 186093 538560 186127 538576
rect 186189 539552 186223 539568
rect 186189 538560 186223 538576
rect 186285 539552 186319 539568
rect 186285 538560 186319 538576
rect 186381 539552 186415 539568
rect 186381 538560 186415 538576
rect 186477 539552 186511 539568
rect 186477 538560 186511 538576
rect 186573 539552 186607 539568
rect 186573 538560 186607 538576
rect 186669 539552 186703 539568
rect 186669 538560 186703 538576
rect 186765 539552 186799 539568
rect 186765 538560 186799 538576
rect 186861 539552 186895 539568
rect 186861 538560 186895 538576
rect 186957 539552 186991 539568
rect 186957 538560 186991 538576
rect 187053 539552 187087 539568
rect 187053 538560 187087 538576
rect 187149 539552 187183 539568
rect 187149 538560 187183 538576
rect 187245 539552 187279 539568
rect 187370 539545 187404 539561
rect 187370 538953 187404 538969
rect 187458 539545 187492 539561
rect 187458 538953 187492 538969
rect 187570 539545 187604 539561
rect 187398 538876 187414 538910
rect 187448 538876 187464 538910
rect 187245 538560 187279 538576
rect 187570 538553 187604 538569
rect 187658 539545 187692 539561
rect 187658 538553 187692 538569
rect 187760 539297 187780 539687
rect 187760 539207 187770 539297
rect 185898 538476 185914 538510
rect 185948 538476 185964 538510
rect 186125 538483 186141 538517
rect 186175 538483 186191 538517
rect 186317 538483 186333 538517
rect 186367 538483 186383 538517
rect 186509 538483 186525 538517
rect 186559 538483 186575 538517
rect 186701 538483 186717 538517
rect 186751 538483 186767 538517
rect 186893 538483 186909 538517
rect 186943 538483 186959 538517
rect 187085 538483 187101 538517
rect 187135 538483 187151 538517
rect 187598 538476 187614 538510
rect 187648 538476 187664 538510
rect 187760 538387 187780 539207
rect 185780 538367 187780 538387
rect 185780 538347 185820 538367
rect 185720 538327 185820 538347
rect 187740 538347 187780 538367
rect 187820 538347 187840 539747
rect 187740 538327 187840 538347
rect 185720 538307 187840 538327
rect 189020 539767 191140 539787
rect 189020 539747 189120 539767
rect 189020 538347 189040 539747
rect 189080 539727 189120 539747
rect 191040 539747 191140 539767
rect 191040 539727 191080 539747
rect 189080 539707 191080 539727
rect 189080 538387 189100 539707
rect 191040 539687 191080 539707
rect 189198 539604 189214 539638
rect 189248 539604 189264 539638
rect 189521 539611 189537 539645
rect 189571 539611 189587 539645
rect 189713 539611 189729 539645
rect 189763 539611 189779 539645
rect 189905 539611 189921 539645
rect 189955 539611 189971 539645
rect 190097 539611 190113 539645
rect 190147 539611 190163 539645
rect 190289 539611 190305 539645
rect 190339 539611 190355 539645
rect 190481 539611 190497 539645
rect 190531 539611 190547 539645
rect 190698 539604 190714 539638
rect 190748 539604 190764 539638
rect 190898 539604 190914 539638
rect 190948 539604 190964 539638
rect 189170 539545 189204 539561
rect 189170 538553 189204 538569
rect 189258 539545 189292 539561
rect 189258 538553 189292 538569
rect 189393 539552 189427 539568
rect 189393 538560 189427 538576
rect 189489 539552 189523 539568
rect 189489 538560 189523 538576
rect 189585 539552 189619 539568
rect 189585 538560 189619 538576
rect 189681 539552 189715 539568
rect 189681 538560 189715 538576
rect 189777 539552 189811 539568
rect 189777 538560 189811 538576
rect 189873 539552 189907 539568
rect 189873 538560 189907 538576
rect 189969 539552 190003 539568
rect 189969 538560 190003 538576
rect 190065 539552 190099 539568
rect 190065 538560 190099 538576
rect 190161 539552 190195 539568
rect 190161 538560 190195 538576
rect 190257 539552 190291 539568
rect 190257 538560 190291 538576
rect 190353 539552 190387 539568
rect 190353 538560 190387 538576
rect 190449 539552 190483 539568
rect 190449 538560 190483 538576
rect 190545 539552 190579 539568
rect 190670 539545 190704 539561
rect 190670 538953 190704 538969
rect 190758 539545 190792 539561
rect 190758 538953 190792 538969
rect 190870 539545 190904 539561
rect 190698 538876 190714 538910
rect 190748 538876 190764 538910
rect 190545 538560 190579 538576
rect 190870 538553 190904 538569
rect 190958 539545 190992 539561
rect 190958 538553 190992 538569
rect 191060 539297 191080 539687
rect 191060 539207 191070 539297
rect 189198 538476 189214 538510
rect 189248 538476 189264 538510
rect 189425 538483 189441 538517
rect 189475 538483 189491 538517
rect 189617 538483 189633 538517
rect 189667 538483 189683 538517
rect 189809 538483 189825 538517
rect 189859 538483 189875 538517
rect 190001 538483 190017 538517
rect 190051 538483 190067 538517
rect 190193 538483 190209 538517
rect 190243 538483 190259 538517
rect 190385 538483 190401 538517
rect 190435 538483 190451 538517
rect 190898 538476 190914 538510
rect 190948 538476 190964 538510
rect 191060 538387 191080 539207
rect 189080 538367 191080 538387
rect 189080 538347 189120 538367
rect 189020 538327 189120 538347
rect 191040 538347 191080 538367
rect 191120 538347 191140 539747
rect 191040 538327 191140 538347
rect 189020 538307 191140 538327
rect 157690 538017 162870 538037
rect 157690 537997 157730 538017
rect 157630 537977 157730 537997
rect 162770 537977 162870 538017
rect 157630 537957 162870 537977
rect 164188 538077 164284 538111
rect 166648 538077 166744 538111
rect 164188 538015 164222 538077
rect 157590 537857 162850 537877
rect 157590 537817 157650 537857
rect 162750 537817 162850 537857
rect 157590 537797 162790 537817
rect 157590 537757 157670 537797
rect 157590 535817 157610 537757
rect 157650 535817 157670 537757
rect 161288 537704 161304 537738
rect 161338 537704 161354 537738
rect 161492 537704 161508 537738
rect 161542 537704 161558 537738
rect 161684 537704 161700 537738
rect 161734 537704 161750 537738
rect 161892 537704 161908 537738
rect 161942 537704 161958 537738
rect 162084 537704 162100 537738
rect 162134 537704 162150 537738
rect 162308 537704 162324 537738
rect 162358 537704 162374 537738
rect 161260 537645 161294 537661
rect 161260 537053 161294 537069
rect 161348 537645 161382 537661
rect 161348 537053 161382 537069
rect 161460 537645 161494 537661
rect 161460 537053 161494 537069
rect 161556 537645 161590 537661
rect 161556 537053 161590 537069
rect 161652 537645 161686 537661
rect 161652 537053 161686 537069
rect 161748 537645 161782 537661
rect 161748 537053 161782 537069
rect 161860 537645 161894 537661
rect 161860 537053 161894 537069
rect 161956 537645 161990 537661
rect 161956 537053 161990 537069
rect 162052 537645 162086 537661
rect 162052 537053 162086 537069
rect 162148 537645 162182 537661
rect 162148 537053 162182 537069
rect 162280 537645 162314 537661
rect 162280 537053 162314 537069
rect 162368 537645 162402 537661
rect 162368 537053 162402 537069
rect 161288 536976 161304 537010
rect 161338 536976 161354 537010
rect 161588 536976 161604 537010
rect 161638 536976 161654 537010
rect 161988 536976 162004 537010
rect 162038 536976 162054 537010
rect 162308 536976 162324 537010
rect 162358 536976 162374 537010
rect 157796 536684 157812 536718
rect 157980 536684 157996 536718
rect 158174 536684 158190 536718
rect 158358 536684 158374 536718
rect 158432 536684 158448 536718
rect 158616 536684 158632 536718
rect 158690 536684 158706 536718
rect 158874 536684 158890 536718
rect 158948 536684 158964 536718
rect 159132 536684 159148 536718
rect 159206 536684 159222 536718
rect 159390 536684 159406 536718
rect 159464 536684 159480 536718
rect 159648 536684 159664 536718
rect 159722 536684 159738 536718
rect 159906 536684 159922 536718
rect 159980 536684 159996 536718
rect 160164 536684 160180 536718
rect 160238 536684 160254 536718
rect 160422 536684 160438 536718
rect 160496 536684 160512 536718
rect 160680 536684 160696 536718
rect 160880 536684 160896 536718
rect 161064 536684 161080 536718
rect 161138 536684 161154 536718
rect 161322 536684 161338 536718
rect 161396 536684 161412 536718
rect 161580 536684 161596 536718
rect 161778 536684 161794 536718
rect 161962 536684 161978 536718
rect 162036 536684 162052 536718
rect 162220 536684 162236 536718
rect 162416 536684 162432 536718
rect 162600 536684 162616 536718
rect 157750 536625 157784 536641
rect 157750 536033 157784 536049
rect 158008 536625 158042 536641
rect 158008 536033 158042 536049
rect 158128 536625 158162 536641
rect 158128 536033 158162 536049
rect 158386 536625 158420 536641
rect 158386 536033 158420 536049
rect 158644 536625 158678 536641
rect 158644 536033 158678 536049
rect 158902 536625 158936 536641
rect 158902 536033 158936 536049
rect 159160 536625 159194 536641
rect 159160 536033 159194 536049
rect 159418 536625 159452 536641
rect 159418 536033 159452 536049
rect 159676 536625 159710 536641
rect 159676 536033 159710 536049
rect 159934 536625 159968 536641
rect 159934 536033 159968 536049
rect 160192 536625 160226 536641
rect 160192 536033 160226 536049
rect 160450 536625 160484 536641
rect 160450 536033 160484 536049
rect 160708 536625 160742 536641
rect 160708 536033 160742 536049
rect 160834 536625 160868 536641
rect 160834 536033 160868 536049
rect 161092 536625 161126 536641
rect 161092 536033 161126 536049
rect 161350 536625 161384 536641
rect 161350 536033 161384 536049
rect 161608 536625 161642 536641
rect 161608 536033 161642 536049
rect 161732 536625 161766 536641
rect 161732 536033 161766 536049
rect 161990 536625 162024 536641
rect 161990 536033 162024 536049
rect 162248 536625 162282 536641
rect 162248 536033 162282 536049
rect 162370 536625 162404 536641
rect 162370 536033 162404 536049
rect 162628 536625 162662 536641
rect 162628 536033 162662 536049
rect 157796 535956 157812 535990
rect 157980 535956 157996 535990
rect 158174 535956 158190 535990
rect 158358 535956 158374 535990
rect 158432 535956 158448 535990
rect 158616 535956 158632 535990
rect 158690 535956 158706 535990
rect 158874 535956 158890 535990
rect 158948 535956 158964 535990
rect 159132 535956 159148 535990
rect 159206 535956 159222 535990
rect 159390 535956 159406 535990
rect 159464 535956 159480 535990
rect 159648 535956 159664 535990
rect 159722 535956 159738 535990
rect 159906 535956 159922 535990
rect 159980 535956 159996 535990
rect 160164 535956 160180 535990
rect 160238 535956 160254 535990
rect 160422 535956 160438 535990
rect 160496 535956 160512 535990
rect 160680 535956 160696 535990
rect 160880 535956 160896 535990
rect 161064 535956 161080 535990
rect 161138 535956 161154 535990
rect 161322 535956 161338 535990
rect 161396 535956 161412 535990
rect 161580 535956 161596 535990
rect 161778 535956 161794 535990
rect 161962 535956 161978 535990
rect 162036 535956 162052 535990
rect 162220 535956 162236 535990
rect 162416 535956 162432 535990
rect 162600 535956 162616 535990
rect 157590 535797 157670 535817
rect 162770 535797 162790 537797
rect 162830 535797 162850 537817
rect 166710 538015 166744 538077
rect 164188 535937 164222 535999
rect 166710 535937 166744 535999
rect 164188 535903 164284 535937
rect 166648 535903 166744 535937
rect 167960 538077 168056 538111
rect 169148 538077 169244 538111
rect 167960 538015 167994 538077
rect 169210 538015 169244 538077
rect 167960 535937 167994 535999
rect 169210 535937 169244 535999
rect 167960 535903 168056 535937
rect 169148 535903 169244 535937
rect 171696 538077 171792 538111
rect 172248 538077 172344 538111
rect 171696 538015 171730 538077
rect 172310 538015 172344 538077
rect 171696 535937 171730 535999
rect 172310 535937 172344 535999
rect 171696 535903 171792 535937
rect 172248 535903 172344 535937
rect 175214 538077 175310 538111
rect 175448 538077 175544 538111
rect 175214 538015 175248 538077
rect 175510 538015 175544 538077
rect 175214 535937 175248 535999
rect 178814 538077 178910 538111
rect 179048 538077 179144 538111
rect 178814 538015 178848 538077
rect 179110 538015 179144 538077
rect 178814 536497 178848 536559
rect 182114 538077 182210 538111
rect 182348 538077 182444 538111
rect 182114 538015 182148 538077
rect 182410 538015 182444 538077
rect 182114 536777 182148 536839
rect 185414 538077 185510 538111
rect 185648 538077 185744 538111
rect 185414 538015 185448 538077
rect 185710 538015 185744 538077
rect 185414 536917 185448 536979
rect 185710 536917 185744 536979
rect 185414 536883 185510 536917
rect 185648 536883 185744 536917
rect 188714 538077 188810 538111
rect 188948 538077 189044 538111
rect 188714 538015 188748 538077
rect 189010 538015 189044 538077
rect 182410 536777 182444 536839
rect 188714 536821 188748 536883
rect 189010 536821 189044 536883
rect 188714 536787 188810 536821
rect 188948 536787 189044 536821
rect 182114 536743 182210 536777
rect 182348 536743 182444 536777
rect 179110 536497 179144 536559
rect 178814 536463 178910 536497
rect 179048 536463 179144 536497
rect 175510 535937 175544 535999
rect 175214 535903 175310 535937
rect 175448 535903 175544 535937
rect 157590 535777 162850 535797
rect 157590 535737 157670 535777
rect 162750 535737 162850 535777
rect 157590 535717 162850 535737
rect 164158 535737 164254 535771
rect 166618 535737 166714 535771
rect 164158 535675 164192 535737
rect 166680 535675 166714 535737
rect 164158 533597 164192 533659
rect 166680 533597 166714 533659
rect 164158 533563 164254 533597
rect 166618 533563 166714 533597
rect 172210 530594 172239 530628
rect 172273 530594 172331 530628
rect 172365 530594 172423 530628
rect 172457 530594 172515 530628
rect 172549 530594 172607 530628
rect 172641 530594 172699 530628
rect 172733 530594 172791 530628
rect 172825 530594 172883 530628
rect 172917 530594 172975 530628
rect 173009 530594 173067 530628
rect 173101 530594 173159 530628
rect 173193 530594 173251 530628
rect 173285 530594 173343 530628
rect 173377 530594 173435 530628
rect 173469 530594 173527 530628
rect 173561 530594 173619 530628
rect 173653 530594 173711 530628
rect 173745 530594 173803 530628
rect 173837 530594 173895 530628
rect 173929 530594 173987 530628
rect 174021 530594 174079 530628
rect 174113 530594 174171 530628
rect 174205 530594 174263 530628
rect 174297 530594 174355 530628
rect 174389 530594 174447 530628
rect 174481 530594 174539 530628
rect 174573 530594 174631 530628
rect 174665 530594 174723 530628
rect 174757 530594 174815 530628
rect 174849 530594 174907 530628
rect 174941 530594 174999 530628
rect 175033 530594 175091 530628
rect 175125 530594 175183 530628
rect 175217 530594 175275 530628
rect 175309 530594 175367 530628
rect 175401 530594 175459 530628
rect 175493 530594 175551 530628
rect 175585 530594 175643 530628
rect 175677 530594 175735 530628
rect 175769 530594 175827 530628
rect 175861 530594 175919 530628
rect 175953 530594 176011 530628
rect 176045 530594 176103 530628
rect 176137 530594 176195 530628
rect 176229 530594 176287 530628
rect 176321 530594 176379 530628
rect 176413 530594 176471 530628
rect 176505 530594 176563 530628
rect 176597 530594 176655 530628
rect 176689 530594 176747 530628
rect 176781 530594 176839 530628
rect 176873 530594 176931 530628
rect 176965 530594 177023 530628
rect 177057 530594 177115 530628
rect 177149 530594 177207 530628
rect 177241 530594 177299 530628
rect 177333 530594 177391 530628
rect 177425 530594 177483 530628
rect 177517 530594 177575 530628
rect 177609 530594 177667 530628
rect 177701 530594 177759 530628
rect 177793 530594 177851 530628
rect 177885 530594 177943 530628
rect 177977 530594 178035 530628
rect 178069 530594 178127 530628
rect 178161 530594 178219 530628
rect 178253 530594 178311 530628
rect 178345 530594 178403 530628
rect 178437 530594 178495 530628
rect 178529 530594 178587 530628
rect 178621 530594 178679 530628
rect 178713 530594 178771 530628
rect 178805 530594 178863 530628
rect 178897 530594 178955 530628
rect 178989 530594 179047 530628
rect 179081 530594 179139 530628
rect 179173 530594 179231 530628
rect 179265 530594 179323 530628
rect 179357 530594 179415 530628
rect 179449 530594 179507 530628
rect 179541 530594 179599 530628
rect 179633 530594 179691 530628
rect 179725 530594 179783 530628
rect 179817 530594 179875 530628
rect 179909 530594 179967 530628
rect 180001 530594 180059 530628
rect 180093 530594 180151 530628
rect 180185 530594 180243 530628
rect 180277 530594 180335 530628
rect 180369 530594 180427 530628
rect 180461 530594 180519 530628
rect 180553 530594 180611 530628
rect 180645 530594 180703 530628
rect 180737 530594 180795 530628
rect 180829 530594 180887 530628
rect 180921 530594 180979 530628
rect 181013 530594 181071 530628
rect 181105 530594 181163 530628
rect 181197 530594 181255 530628
rect 181289 530594 181347 530628
rect 181381 530594 181439 530628
rect 181473 530594 181531 530628
rect 181565 530594 181623 530628
rect 181657 530594 181715 530628
rect 181749 530594 181807 530628
rect 181841 530594 181899 530628
rect 181933 530594 181991 530628
rect 182025 530594 182083 530628
rect 182117 530594 182175 530628
rect 182209 530594 182267 530628
rect 182301 530594 182359 530628
rect 182393 530594 182451 530628
rect 182485 530594 182543 530628
rect 182577 530594 182635 530628
rect 182669 530594 182727 530628
rect 182761 530594 182819 530628
rect 182853 530594 182911 530628
rect 182945 530594 183003 530628
rect 183037 530594 183095 530628
rect 183129 530594 183187 530628
rect 183221 530594 183279 530628
rect 183313 530594 183371 530628
rect 183405 530594 183463 530628
rect 183497 530594 183555 530628
rect 183589 530594 183647 530628
rect 183681 530594 183739 530628
rect 183773 530594 183831 530628
rect 183865 530594 183923 530628
rect 183957 530594 184015 530628
rect 184049 530594 184107 530628
rect 184141 530594 184199 530628
rect 184233 530594 184291 530628
rect 184325 530594 184383 530628
rect 184417 530594 184475 530628
rect 184509 530594 184567 530628
rect 184601 530594 184659 530628
rect 184693 530594 184751 530628
rect 184785 530594 184843 530628
rect 184877 530594 184935 530628
rect 184969 530594 185027 530628
rect 185061 530594 185119 530628
rect 185153 530594 185211 530628
rect 185245 530594 185303 530628
rect 185337 530594 185395 530628
rect 185429 530594 185487 530628
rect 185521 530594 185579 530628
rect 185613 530594 185671 530628
rect 185705 530594 185763 530628
rect 185797 530594 185855 530628
rect 185889 530594 185947 530628
rect 185981 530594 186039 530628
rect 186073 530594 186131 530628
rect 186165 530594 186223 530628
rect 186257 530594 186315 530628
rect 186349 530594 186407 530628
rect 186441 530594 186499 530628
rect 186533 530594 186591 530628
rect 186625 530594 186683 530628
rect 186717 530594 186775 530628
rect 186809 530594 186867 530628
rect 186901 530594 186959 530628
rect 186993 530594 187051 530628
rect 187085 530594 187143 530628
rect 187177 530594 187235 530628
rect 187269 530594 187327 530628
rect 187361 530594 187419 530628
rect 187453 530594 187482 530628
rect 172227 530531 172469 530594
rect 172227 530497 172245 530531
rect 172279 530497 172417 530531
rect 172451 530497 172469 530531
rect 172515 530548 172571 530594
rect 172515 530514 172528 530548
rect 172562 530514 172571 530548
rect 172692 530548 172743 530594
rect 172515 530498 172571 530514
rect 172605 530526 172657 530542
rect 172227 530444 172469 530497
rect 172605 530492 172614 530526
rect 172648 530492 172657 530526
rect 172692 530514 172700 530548
rect 172734 530514 172743 530548
rect 172872 530548 172927 530594
rect 172692 530498 172743 530514
rect 172777 530526 172836 530542
rect 172605 530464 172657 530492
rect 172777 530492 172786 530526
rect 172820 530492 172836 530526
rect 172872 530514 172883 530548
rect 172917 530514 172927 530548
rect 172872 530498 172927 530514
rect 172961 530544 173021 530560
rect 172961 530510 172969 530544
rect 173003 530510 173021 530544
rect 172961 530494 173021 530510
rect 172777 530464 172836 530492
rect 172506 530458 172836 530464
rect 172227 530370 172331 530444
rect 172506 530424 172515 530458
rect 172549 530430 172836 530458
rect 172549 530424 172587 530430
rect 172227 530336 172277 530370
rect 172311 530336 172331 530370
rect 172365 530376 172385 530410
rect 172419 530376 172469 530410
rect 172365 530302 172469 530376
rect 172227 530255 172469 530302
rect 172506 530328 172587 530424
rect 172883 530396 172953 530460
rect 172621 530362 172637 530396
rect 172671 530362 172705 530396
rect 172739 530362 172773 530396
rect 172807 530362 172849 530396
rect 172506 530304 172657 530328
rect 172506 530294 172615 530304
rect 172605 530270 172615 530294
rect 172649 530270 172657 530304
rect 172815 530312 172849 530362
rect 172883 530390 172919 530396
rect 172917 530362 172919 530390
rect 172917 530356 172953 530362
rect 172883 530346 172953 530356
rect 172987 530312 173021 530494
rect 173055 530533 174124 530594
rect 173055 530499 173073 530533
rect 173107 530499 174073 530533
rect 174107 530499 174124 530533
rect 173055 530485 174124 530499
rect 174159 530533 174677 530594
rect 174159 530499 174177 530533
rect 174211 530499 174625 530533
rect 174659 530499 174677 530533
rect 173372 530370 173440 530485
rect 174159 530440 174677 530499
rect 174803 530500 174861 530594
rect 174803 530466 174815 530500
rect 174849 530466 174861 530500
rect 174907 530548 174963 530594
rect 174907 530514 174920 530548
rect 174954 530514 174963 530548
rect 175084 530548 175135 530594
rect 174907 530498 174963 530514
rect 174997 530526 175049 530542
rect 174803 530449 174861 530466
rect 174997 530492 175006 530526
rect 175040 530492 175049 530526
rect 175084 530514 175092 530548
rect 175126 530514 175135 530548
rect 175264 530548 175319 530594
rect 175084 530498 175135 530514
rect 175169 530526 175228 530542
rect 174997 530464 175049 530492
rect 175169 530492 175178 530526
rect 175212 530492 175228 530526
rect 175264 530514 175275 530548
rect 175309 530514 175319 530548
rect 175264 530498 175319 530514
rect 175353 530544 175413 530560
rect 175353 530510 175361 530544
rect 175395 530510 175413 530544
rect 175353 530494 175413 530510
rect 175169 530464 175228 530492
rect 174898 530458 175228 530464
rect 173372 530336 173389 530370
rect 173423 530336 173440 530370
rect 173372 530319 173440 530336
rect 173736 530406 173806 530421
rect 173736 530372 173753 530406
rect 173787 530372 173806 530406
rect 172815 530290 173021 530312
rect 172815 530278 172969 530290
rect 172227 530221 172245 530255
rect 172279 530221 172417 530255
rect 172451 530221 172469 530255
rect 172227 530160 172469 530221
rect 172227 530126 172245 530160
rect 172279 530126 172417 530160
rect 172451 530126 172469 530160
rect 172227 530084 172469 530126
rect 172514 530242 172571 530258
rect 172514 530208 172529 530242
rect 172563 530208 172571 530242
rect 172514 530174 172571 530208
rect 172514 530140 172529 530174
rect 172563 530140 172571 530174
rect 172514 530084 172571 530140
rect 172605 530244 172657 530270
rect 172959 530256 172969 530278
rect 173003 530256 173021 530290
rect 172605 530236 172829 530244
rect 172605 530202 172615 530236
rect 172649 530210 172829 530236
rect 172649 530202 172657 530210
rect 172605 530168 172657 530202
rect 172777 530195 172829 530210
rect 172605 530134 172615 530168
rect 172649 530134 172657 530168
rect 172605 530118 172657 530134
rect 172692 530160 172743 530176
rect 172692 530126 172701 530160
rect 172735 530126 172743 530160
rect 172692 530084 172743 530126
rect 172777 530161 172787 530195
rect 172821 530161 172829 530195
rect 172777 530118 172829 530161
rect 172863 530228 172925 530244
rect 172863 530194 172883 530228
rect 172917 530194 172925 530228
rect 172863 530160 172925 530194
rect 172863 530126 172883 530160
rect 172917 530126 172925 530160
rect 172863 530084 172925 530126
rect 172959 530168 173021 530256
rect 173736 530171 173806 530372
rect 174159 530370 174401 530440
rect 174898 530424 174907 530458
rect 174941 530430 175228 530458
rect 174941 530424 174979 530430
rect 174159 530336 174237 530370
rect 174271 530336 174347 530370
rect 174381 530336 174401 530370
rect 174435 530372 174455 530406
rect 174489 530372 174565 530406
rect 174599 530372 174677 530406
rect 174435 530302 174677 530372
rect 174898 530328 174979 530424
rect 175275 530396 175345 530460
rect 175013 530362 175029 530396
rect 175063 530362 175097 530396
rect 175131 530362 175165 530396
rect 175199 530362 175241 530396
rect 174159 530262 174677 530302
rect 174159 530228 174177 530262
rect 174211 530228 174625 530262
rect 174659 530228 174677 530262
rect 172959 530134 172969 530168
rect 173003 530134 173021 530168
rect 172959 530118 173021 530134
rect 173055 530160 174124 530171
rect 173055 530126 173073 530160
rect 173107 530126 174073 530160
rect 174107 530126 174124 530160
rect 173055 530084 174124 530126
rect 174159 530160 174677 530228
rect 174159 530126 174177 530160
rect 174211 530126 174625 530160
rect 174659 530126 174677 530160
rect 174159 530084 174677 530126
rect 174803 530282 174861 530317
rect 174898 530304 175049 530328
rect 174898 530294 175007 530304
rect 174803 530248 174815 530282
rect 174849 530248 174861 530282
rect 174997 530270 175007 530294
rect 175041 530270 175049 530304
rect 175207 530312 175241 530362
rect 175275 530390 175311 530396
rect 175309 530362 175311 530390
rect 175309 530356 175345 530362
rect 175275 530346 175345 530356
rect 175379 530312 175413 530494
rect 175207 530290 175413 530312
rect 175207 530278 175361 530290
rect 174803 530189 174861 530248
rect 174803 530155 174815 530189
rect 174849 530155 174861 530189
rect 174803 530084 174861 530155
rect 174906 530242 174963 530258
rect 174906 530208 174921 530242
rect 174955 530208 174963 530242
rect 174906 530174 174963 530208
rect 174906 530140 174921 530174
rect 174955 530140 174963 530174
rect 174906 530084 174963 530140
rect 174997 530244 175049 530270
rect 175351 530256 175361 530278
rect 175395 530256 175413 530290
rect 174997 530236 175221 530244
rect 174997 530202 175007 530236
rect 175041 530210 175221 530236
rect 175041 530202 175049 530210
rect 174997 530168 175049 530202
rect 175169 530195 175221 530210
rect 174997 530134 175007 530168
rect 175041 530134 175049 530168
rect 174997 530118 175049 530134
rect 175084 530160 175135 530176
rect 175084 530126 175093 530160
rect 175127 530126 175135 530160
rect 175084 530084 175135 530126
rect 175169 530161 175179 530195
rect 175213 530161 175221 530195
rect 175169 530118 175221 530161
rect 175255 530228 175317 530244
rect 175255 530194 175275 530228
rect 175309 530194 175317 530228
rect 175255 530160 175317 530194
rect 175255 530126 175275 530160
rect 175309 530126 175317 530160
rect 175255 530084 175317 530126
rect 175351 530168 175413 530256
rect 175351 530134 175361 530168
rect 175395 530134 175413 530168
rect 175540 530502 175591 530558
rect 175625 530552 175686 530594
rect 175983 530556 176021 530594
rect 175625 530518 175641 530552
rect 175675 530518 175686 530552
rect 175625 530502 175686 530518
rect 175735 530536 175949 530552
rect 175735 530502 175765 530536
rect 175799 530518 175949 530536
rect 175540 530468 175557 530502
rect 175540 530452 175591 530468
rect 175540 530322 175582 530452
rect 175735 530447 175799 530502
rect 175734 530412 175799 530447
rect 175616 530396 175799 530412
rect 175650 530362 175799 530396
rect 175616 530352 175799 530362
rect 175833 530458 175881 530484
rect 175833 530424 175847 530458
rect 175915 530472 175949 530518
rect 176017 530522 176021 530556
rect 175983 530506 176021 530522
rect 176055 530552 176245 530560
rect 176055 530518 176195 530552
rect 176229 530518 176245 530552
rect 176289 530522 176305 530556
rect 176339 530522 176359 530556
rect 176055 530504 176245 530518
rect 175915 530438 176021 530472
rect 175833 530404 175881 530424
rect 175977 530432 176021 530438
rect 175833 530370 175891 530404
rect 175925 530395 175941 530404
rect 175977 530398 175987 530432
rect 175977 530382 176021 530398
rect 175833 530361 175907 530370
rect 175616 530346 175764 530352
rect 175540 530288 175551 530322
rect 175585 530288 175591 530322
rect 175540 530264 175591 530288
rect 175540 530230 175557 530264
rect 175540 530196 175591 530230
rect 175540 530162 175557 530196
rect 175540 530146 175591 530162
rect 175625 530228 175686 530312
rect 175625 530194 175641 530228
rect 175675 530194 175686 530228
rect 175730 530228 175764 530346
rect 175833 530330 175941 530361
rect 176055 530348 176089 530504
rect 176008 530314 176089 530348
rect 176123 530406 176193 530470
rect 176123 530390 176131 530406
rect 176165 530372 176193 530406
rect 176157 530356 176193 530372
rect 176123 530346 176193 530356
rect 176227 530454 176269 530470
rect 176261 530420 176269 530454
rect 176008 530296 176042 530314
rect 176227 530312 176269 530420
rect 175798 530262 175814 530296
rect 175848 530262 176042 530296
rect 176134 530280 176269 530312
rect 175730 530194 175890 530228
rect 175625 530160 175686 530194
rect 175856 530186 175890 530194
rect 175351 530118 175413 530134
rect 175625 530126 175641 530160
rect 175675 530126 175686 530160
rect 175625 530084 175686 530126
rect 175754 530126 175770 530160
rect 175804 530126 175820 530160
rect 176008 530186 176042 530262
rect 176076 530246 176092 530280
rect 176126 530278 176269 530280
rect 176307 530444 176359 530522
rect 176401 530552 176467 530594
rect 176401 530518 176417 530552
rect 176451 530518 176467 530552
rect 176987 530556 177053 530594
rect 176401 530502 176467 530518
rect 176642 530516 176763 530550
rect 176797 530516 176813 530550
rect 176854 530516 176870 530550
rect 176904 530516 176953 530550
rect 176987 530522 177003 530556
rect 177037 530522 177053 530556
rect 177193 530552 177259 530594
rect 177125 530526 177159 530542
rect 176307 530306 176341 530444
rect 176443 530442 176495 530458
rect 176375 530394 176409 530410
rect 176443 530408 176471 530442
rect 176529 530424 176567 530458
rect 176505 530408 176601 530424
rect 176642 530374 176676 530516
rect 176710 530448 176781 530458
rect 176710 530414 176726 530448
rect 176760 530414 176781 530448
rect 176409 530360 176713 530374
rect 176375 530340 176713 530360
rect 176126 530254 176168 530278
rect 176076 530220 176123 530246
rect 176157 530220 176168 530254
rect 176307 530272 176557 530306
rect 176591 530272 176607 530306
rect 176307 530244 176341 530272
rect 176229 530210 176341 530244
rect 175856 530136 175890 530152
rect 175924 530160 175974 530176
rect 175754 530084 175820 530126
rect 175924 530126 175940 530160
rect 175924 530084 175974 530126
rect 176008 530161 176182 530186
rect 176008 530127 176132 530161
rect 176166 530127 176182 530161
rect 176008 530118 176182 530127
rect 176229 530168 176263 530210
rect 176430 530204 176645 530238
rect 176430 530186 176464 530204
rect 176229 530118 176263 530134
rect 176297 530160 176371 530176
rect 176297 530126 176317 530160
rect 176351 530126 176371 530160
rect 176611 530186 176645 530204
rect 176430 530136 176464 530152
rect 176498 530136 176514 530170
rect 176548 530136 176564 530170
rect 176611 530136 176645 530152
rect 176679 530184 176713 530340
rect 176747 530296 176781 530414
rect 176815 530442 176885 530458
rect 176815 530408 176828 530442
rect 176862 530408 176885 530442
rect 176815 530390 176885 530408
rect 176815 530356 176839 530390
rect 176873 530356 176885 530390
rect 176815 530334 176885 530356
rect 176747 530280 176840 530296
rect 176747 530254 176806 530280
rect 176781 530246 176806 530254
rect 176781 530220 176840 530246
rect 176919 530244 176953 530516
rect 177193 530518 177209 530552
rect 177243 530518 177259 530552
rect 177293 530526 177344 530542
rect 176987 530335 177079 530488
rect 177021 530322 177079 530335
rect 177021 530301 177023 530322
rect 176987 530288 177023 530301
rect 177057 530288 177079 530322
rect 176987 530278 177079 530288
rect 176747 530218 176840 530220
rect 176874 530210 176953 530244
rect 176874 530184 176908 530210
rect 176679 530162 176815 530184
rect 176297 530084 176371 530126
rect 176498 530084 176564 530136
rect 176679 530128 176765 530162
rect 176799 530128 176815 530162
rect 176679 530118 176815 530128
rect 176858 530168 176908 530184
rect 176892 530134 176908 530168
rect 176858 530118 176908 530134
rect 176942 530160 176992 530176
rect 176976 530126 176992 530160
rect 176942 530084 176992 530126
rect 177026 530121 177091 530278
rect 177125 530254 177159 530492
rect 177327 530492 177344 530526
rect 177293 530484 177344 530492
rect 177194 530450 177344 530484
rect 177379 530500 177437 530594
rect 177379 530466 177391 530500
rect 177425 530466 177437 530500
rect 177194 530390 177240 530450
rect 177379 530449 177437 530466
rect 177655 530526 177732 530560
rect 177655 530492 177692 530526
rect 177726 530492 177732 530526
rect 177766 530552 177831 530594
rect 177766 530518 177782 530552
rect 177816 530518 177831 530552
rect 177766 530502 177831 530518
rect 177935 530526 177991 530560
rect 177655 530446 177732 530492
rect 177935 530492 177941 530526
rect 177975 530492 177991 530526
rect 177935 530468 177991 530492
rect 177194 530381 177206 530390
rect 177228 530347 177240 530356
rect 177194 530252 177240 530347
rect 177274 530396 177344 530416
rect 177274 530362 177296 530396
rect 177330 530362 177344 530396
rect 177274 530322 177344 530362
rect 177274 530288 177299 530322
rect 177333 530288 177344 530322
rect 177274 530286 177344 530288
rect 177379 530282 177437 530317
rect 177194 530236 177344 530252
rect 177194 530218 177293 530236
rect 177125 530168 177159 530202
rect 177327 530202 177344 530236
rect 177125 530118 177159 530134
rect 177193 530150 177209 530184
rect 177243 530150 177259 530184
rect 177193 530084 177259 530150
rect 177293 530168 177344 530202
rect 177327 530134 177344 530168
rect 177293 530118 177344 530134
rect 177379 530248 177391 530282
rect 177425 530248 177437 530282
rect 177379 530189 177437 530248
rect 177379 530155 177391 530189
rect 177425 530155 177437 530189
rect 177379 530084 177437 530155
rect 177655 530312 177711 530446
rect 177766 530434 177991 530468
rect 178029 530526 178109 530560
rect 178029 530492 178045 530526
rect 178079 530492 178109 530526
rect 178189 530552 178243 530594
rect 178189 530518 178199 530552
rect 178233 530518 178243 530552
rect 178189 530502 178243 530518
rect 178277 530526 178334 530560
rect 177766 530412 177856 530434
rect 177745 530396 177856 530412
rect 178029 530400 178109 530492
rect 178277 530492 178283 530526
rect 178317 530492 178334 530526
rect 178277 530468 178334 530492
rect 177779 530362 177856 530396
rect 177745 530346 177856 530362
rect 177655 530186 177732 530312
rect 177766 530254 177856 530346
rect 177890 530396 178109 530400
rect 177890 530362 177941 530396
rect 177975 530362 178109 530396
rect 177890 530288 178109 530362
rect 177766 530210 177991 530254
rect 177655 530152 177667 530186
rect 177726 530152 177732 530186
rect 177935 530186 177991 530210
rect 177655 530118 177732 530152
rect 177766 530160 177831 530176
rect 177766 530126 177782 530160
rect 177816 530126 177831 530160
rect 177766 530084 177831 530126
rect 177935 530152 177941 530186
rect 177975 530152 177991 530186
rect 177935 530118 177991 530152
rect 178029 530186 178109 530288
rect 178143 530434 178334 530468
rect 178391 530522 178443 530560
rect 178391 530488 178409 530522
rect 178479 530552 178545 530594
rect 178479 530518 178495 530552
rect 178529 530518 178545 530552
rect 178581 530539 178615 530560
rect 178391 530459 178443 530488
rect 178581 530484 178615 530505
rect 178679 530548 178735 530594
rect 178679 530514 178692 530548
rect 178726 530514 178735 530548
rect 178856 530548 178907 530594
rect 178679 530498 178735 530514
rect 178769 530526 178821 530542
rect 178143 530396 178185 530434
rect 178143 530362 178145 530396
rect 178179 530362 178185 530396
rect 178143 530254 178185 530362
rect 178219 530396 178357 530400
rect 178219 530362 178259 530396
rect 178293 530362 178357 530396
rect 178219 530322 178357 530362
rect 178253 530288 178357 530322
rect 178391 530299 178425 530459
rect 178482 530450 178615 530484
rect 178769 530492 178771 530526
rect 178812 530492 178821 530526
rect 178856 530514 178864 530548
rect 178898 530514 178907 530548
rect 179036 530548 179091 530594
rect 178856 530498 178907 530514
rect 178941 530526 179000 530542
rect 178769 530464 178821 530492
rect 178941 530492 178950 530526
rect 178984 530492 179000 530526
rect 179036 530514 179047 530548
rect 179081 530514 179091 530548
rect 179036 530498 179091 530514
rect 179125 530544 179185 530560
rect 179125 530510 179133 530544
rect 179167 530510 179185 530544
rect 179125 530494 179185 530510
rect 178941 530464 179000 530492
rect 178482 530399 178516 530450
rect 178670 530430 179000 530464
rect 178459 530383 178516 530399
rect 178493 530349 178516 530383
rect 178459 530333 178516 530349
rect 178563 530396 178629 530414
rect 178563 530362 178579 530396
rect 178613 530390 178629 530396
rect 178563 530356 178587 530362
rect 178621 530356 178629 530390
rect 178563 530340 178629 530356
rect 178482 530304 178516 530333
rect 178670 530328 178751 530430
rect 179047 530396 179117 530460
rect 178785 530362 178801 530396
rect 178835 530362 178869 530396
rect 178903 530362 178937 530396
rect 178971 530362 179013 530396
rect 178670 530304 178821 530328
rect 178143 530210 178334 530254
rect 178029 530152 178045 530186
rect 178079 530152 178109 530186
rect 178277 530186 178334 530210
rect 178029 530118 178109 530152
rect 178189 530160 178243 530176
rect 178189 530126 178199 530160
rect 178233 530126 178243 530160
rect 178189 530084 178243 530126
rect 178277 530152 178283 530186
rect 178317 530152 178334 530186
rect 178277 530118 178334 530152
rect 178391 530249 178445 530299
rect 178482 530270 178615 530304
rect 178670 530294 178779 530304
rect 178391 530215 178409 530249
rect 178443 530215 178445 530249
rect 178581 530236 178615 530270
rect 178769 530270 178779 530294
rect 178813 530270 178821 530304
rect 178979 530312 179013 530362
rect 179047 530390 179083 530396
rect 179081 530362 179083 530390
rect 179081 530356 179117 530362
rect 179047 530346 179117 530356
rect 179151 530312 179185 530494
rect 178979 530290 179185 530312
rect 178979 530278 179133 530290
rect 178391 530186 178445 530215
rect 178391 530152 178403 530186
rect 178437 530168 178445 530186
rect 178391 530134 178409 530152
rect 178443 530134 178445 530168
rect 178391 530118 178445 530134
rect 178479 530202 178495 530236
rect 178529 530202 178545 530236
rect 178479 530168 178545 530202
rect 178479 530134 178495 530168
rect 178529 530134 178545 530168
rect 178479 530084 178545 530134
rect 178581 530168 178615 530202
rect 178581 530118 178615 530134
rect 178678 530242 178735 530258
rect 178678 530208 178693 530242
rect 178727 530208 178735 530242
rect 178678 530174 178735 530208
rect 178678 530140 178693 530174
rect 178727 530140 178735 530174
rect 178678 530084 178735 530140
rect 178769 530244 178821 530270
rect 179123 530256 179133 530278
rect 179167 530256 179185 530290
rect 178769 530236 178993 530244
rect 178769 530202 178779 530236
rect 178813 530210 178993 530236
rect 178813 530202 178821 530210
rect 178769 530168 178821 530202
rect 178941 530195 178993 530210
rect 178769 530134 178779 530168
rect 178813 530134 178821 530168
rect 178769 530118 178821 530134
rect 178856 530160 178907 530176
rect 178856 530126 178865 530160
rect 178899 530126 178907 530160
rect 178856 530084 178907 530126
rect 178941 530161 178951 530195
rect 178985 530161 178993 530195
rect 178941 530118 178993 530161
rect 179027 530228 179089 530244
rect 179027 530194 179047 530228
rect 179081 530194 179089 530228
rect 179027 530160 179089 530194
rect 179027 530126 179047 530160
rect 179081 530126 179089 530160
rect 179027 530084 179089 530126
rect 179123 530168 179185 530256
rect 179123 530134 179133 530168
rect 179167 530134 179185 530168
rect 179123 530118 179185 530134
rect 179219 530544 179279 530560
rect 179219 530510 179237 530544
rect 179271 530510 179279 530544
rect 179219 530494 179279 530510
rect 179313 530548 179368 530594
rect 179313 530514 179323 530548
rect 179357 530514 179368 530548
rect 179497 530548 179548 530594
rect 179313 530498 179368 530514
rect 179404 530526 179463 530542
rect 179219 530312 179253 530494
rect 179404 530492 179415 530526
rect 179454 530492 179463 530526
rect 179497 530514 179506 530548
rect 179540 530514 179548 530548
rect 179669 530548 179725 530594
rect 179497 530498 179548 530514
rect 179583 530526 179635 530542
rect 179404 530464 179463 530492
rect 179583 530492 179592 530526
rect 179626 530492 179635 530526
rect 179669 530514 179678 530548
rect 179712 530514 179725 530548
rect 179669 530498 179725 530514
rect 179955 530500 180013 530594
rect 179583 530464 179635 530492
rect 179955 530466 179967 530500
rect 180001 530466 180013 530500
rect 179287 530396 179357 530460
rect 179404 530430 179734 530464
rect 179955 530449 180013 530466
rect 180232 530533 180283 530560
rect 180232 530499 180249 530533
rect 180317 530552 180383 530594
rect 180317 530518 180333 530552
rect 180367 530518 180383 530552
rect 180317 530514 180383 530518
rect 180468 530537 180574 530560
rect 179321 530390 179357 530396
rect 179321 530362 179323 530390
rect 179287 530356 179323 530362
rect 179287 530346 179357 530356
rect 179391 530362 179433 530396
rect 179467 530362 179501 530396
rect 179535 530362 179569 530396
rect 179603 530362 179619 530396
rect 179391 530312 179425 530362
rect 179653 530328 179734 530430
rect 179219 530290 179425 530312
rect 179219 530256 179237 530290
rect 179271 530278 179425 530290
rect 179583 530304 179734 530328
rect 180232 530446 180283 530499
rect 180468 530503 180540 530537
rect 180468 530487 180574 530503
rect 180468 530480 180503 530487
rect 180317 530446 180503 530480
rect 179271 530256 179281 530278
rect 179219 530168 179281 530256
rect 179583 530270 179591 530304
rect 179625 530294 179734 530304
rect 179625 530270 179635 530294
rect 179583 530244 179635 530270
rect 179955 530282 180013 530317
rect 179219 530134 179237 530168
rect 179271 530134 179281 530168
rect 179219 530118 179281 530134
rect 179315 530228 179377 530244
rect 179315 530194 179323 530228
rect 179357 530194 179377 530228
rect 179315 530160 179377 530194
rect 179315 530126 179323 530160
rect 179357 530126 179377 530160
rect 179315 530084 179377 530126
rect 179411 530236 179635 530244
rect 179411 530210 179591 530236
rect 179411 530195 179463 530210
rect 179411 530161 179419 530195
rect 179453 530161 179463 530195
rect 179583 530202 179591 530210
rect 179625 530202 179635 530236
rect 179411 530118 179463 530161
rect 179497 530160 179548 530176
rect 179497 530126 179505 530160
rect 179539 530126 179548 530160
rect 179497 530084 179548 530126
rect 179583 530168 179635 530202
rect 179583 530134 179591 530168
rect 179625 530134 179635 530168
rect 179583 530118 179635 530134
rect 179669 530242 179726 530258
rect 179669 530208 179677 530242
rect 179711 530208 179726 530242
rect 179669 530174 179726 530208
rect 179669 530140 179677 530174
rect 179711 530140 179726 530174
rect 179669 530084 179726 530140
rect 179955 530248 179967 530282
rect 180001 530248 180013 530282
rect 179955 530189 180013 530248
rect 179955 530155 179967 530189
rect 180001 530155 180013 530189
rect 179955 530084 180013 530155
rect 180232 530312 180266 530446
rect 180317 530412 180351 530446
rect 180300 530396 180351 530412
rect 180334 530362 180351 530396
rect 180300 530346 180351 530362
rect 180396 530396 180435 530412
rect 180430 530362 180435 530396
rect 180396 530346 180435 530362
rect 180232 530296 180299 530312
rect 180232 530262 180249 530296
rect 180283 530262 180299 530296
rect 180232 530228 180299 530262
rect 180232 530194 180249 530228
rect 180283 530194 180299 530228
rect 180232 530186 180299 530194
rect 180232 530152 180243 530186
rect 180277 530160 180299 530186
rect 180232 530126 180249 530152
rect 180283 530126 180299 530160
rect 180232 530118 180299 530126
rect 180333 530296 180367 530312
rect 180333 530228 180367 530262
rect 180333 530160 180367 530194
rect 180333 530084 180367 530126
rect 180401 530152 180435 530346
rect 180469 530220 180503 530446
rect 180537 530432 180571 530448
rect 180537 530288 180571 530398
rect 180612 530432 180667 530560
rect 180612 530398 180633 530432
rect 180612 530390 180667 530398
rect 180645 530356 180667 530390
rect 180612 530328 180667 530356
rect 180701 530526 180739 530560
rect 180701 530492 180703 530526
rect 180737 530492 180739 530526
rect 180701 530319 180739 530492
rect 180775 530537 180877 530594
rect 180809 530503 180843 530537
rect 180775 530487 180877 530503
rect 180921 530537 180970 530553
rect 180921 530503 180927 530537
rect 180961 530503 180970 530537
rect 180921 530432 180970 530503
rect 181206 530537 181255 530553
rect 181206 530503 181215 530537
rect 181249 530503 181255 530537
rect 181206 530432 181255 530503
rect 181299 530537 181401 530594
rect 181333 530503 181367 530537
rect 181299 530487 181401 530503
rect 180779 530398 180795 530432
rect 180829 530398 181025 530432
rect 180701 530288 180705 530319
rect 180537 530285 180705 530288
rect 180537 530254 180739 530285
rect 180773 530322 180923 530323
rect 180773 530288 180795 530322
rect 180829 530319 180923 530322
rect 180829 530288 180873 530319
rect 180773 530285 180873 530288
rect 180907 530285 180923 530319
rect 180469 530186 180569 530220
rect 180603 530186 180644 530220
rect 180678 530186 180694 530220
rect 180773 530152 180807 530285
rect 180957 530236 181025 530398
rect 180401 530118 180807 530152
rect 180841 530220 180875 530236
rect 180841 530084 180875 530186
rect 180922 530220 181025 530236
rect 180922 530186 180927 530220
rect 180961 530186 181025 530220
rect 180922 530154 181025 530186
rect 181151 530398 181347 530432
rect 181381 530398 181397 530432
rect 181151 530236 181219 530398
rect 181253 530322 181403 530323
rect 181253 530288 181255 530322
rect 181289 530319 181403 530322
rect 181253 530285 181269 530288
rect 181303 530285 181403 530319
rect 181151 530220 181254 530236
rect 181151 530186 181215 530220
rect 181249 530186 181254 530220
rect 181151 530154 181254 530186
rect 181301 530220 181335 530236
rect 181301 530084 181335 530186
rect 181369 530152 181403 530285
rect 181437 530322 181475 530560
rect 181509 530432 181564 530560
rect 181602 530537 181708 530560
rect 181636 530503 181708 530537
rect 181793 530552 181859 530594
rect 181793 530518 181809 530552
rect 181843 530518 181859 530552
rect 181793 530514 181859 530518
rect 181893 530533 181944 530560
rect 181602 530487 181708 530503
rect 181673 530480 181708 530487
rect 181927 530499 181944 530533
rect 181543 530398 181564 530432
rect 181509 530390 181564 530398
rect 181605 530432 181639 530448
rect 181509 530356 181531 530390
rect 181509 530328 181564 530356
rect 181437 530319 181439 530322
rect 181473 530288 181475 530322
rect 181605 530288 181639 530398
rect 181471 530285 181639 530288
rect 181437 530254 181639 530285
rect 181673 530446 181859 530480
rect 181893 530446 181944 530499
rect 181673 530220 181707 530446
rect 181825 530412 181859 530446
rect 181482 530186 181498 530220
rect 181532 530186 181573 530220
rect 181607 530186 181707 530220
rect 181741 530396 181780 530412
rect 181741 530362 181746 530396
rect 181741 530346 181780 530362
rect 181825 530396 181876 530412
rect 181825 530362 181842 530396
rect 181825 530346 181876 530362
rect 181741 530152 181775 530346
rect 181910 530312 181944 530446
rect 181369 530118 181775 530152
rect 181809 530296 181843 530312
rect 181809 530228 181843 530262
rect 181809 530160 181843 530194
rect 181809 530084 181843 530126
rect 181877 530296 181944 530312
rect 181877 530262 181893 530296
rect 181927 530262 181944 530296
rect 181877 530254 181944 530262
rect 181877 530228 181899 530254
rect 181877 530194 181893 530228
rect 181933 530220 181944 530254
rect 181927 530194 181944 530220
rect 181877 530160 181944 530194
rect 181877 530126 181893 530160
rect 181927 530126 181944 530160
rect 181877 530118 181944 530126
rect 181979 530544 182039 530560
rect 181979 530510 181997 530544
rect 182031 530510 182039 530544
rect 181979 530494 182039 530510
rect 182073 530548 182128 530594
rect 182073 530514 182083 530548
rect 182117 530514 182128 530548
rect 182257 530548 182308 530594
rect 182073 530498 182128 530514
rect 182164 530526 182223 530542
rect 181979 530312 182013 530494
rect 182164 530492 182180 530526
rect 182214 530492 182223 530526
rect 182257 530514 182266 530548
rect 182300 530514 182308 530548
rect 182429 530548 182485 530594
rect 182257 530498 182308 530514
rect 182343 530526 182395 530542
rect 182164 530464 182223 530492
rect 182343 530492 182352 530526
rect 182386 530492 182395 530526
rect 182429 530514 182438 530548
rect 182472 530514 182485 530548
rect 182429 530498 182485 530514
rect 182531 530500 182589 530594
rect 182343 530464 182395 530492
rect 182531 530466 182543 530500
rect 182577 530466 182589 530500
rect 182047 530458 182117 530460
rect 182047 530424 182083 530458
rect 182164 530430 182494 530464
rect 182531 530449 182589 530466
rect 182623 530526 182957 530594
rect 182623 530492 182641 530526
rect 182675 530492 182905 530526
rect 182939 530492 182957 530526
rect 182047 530396 182117 530424
rect 182081 530362 182117 530396
rect 182047 530346 182117 530362
rect 182151 530362 182193 530396
rect 182227 530362 182261 530396
rect 182295 530362 182329 530396
rect 182363 530362 182379 530396
rect 182151 530312 182185 530362
rect 182413 530328 182494 530430
rect 182623 530440 182957 530492
rect 183083 530544 183143 530560
rect 183083 530510 183101 530544
rect 183135 530510 183143 530544
rect 183083 530494 183143 530510
rect 183177 530548 183232 530594
rect 183177 530514 183187 530548
rect 183221 530514 183232 530548
rect 183361 530548 183412 530594
rect 183177 530498 183232 530514
rect 183268 530526 183327 530542
rect 182623 530370 182773 530440
rect 182623 530336 182643 530370
rect 182677 530336 182773 530370
rect 182807 530372 182903 530406
rect 182937 530372 182957 530406
rect 181979 530290 182185 530312
rect 181979 530256 181997 530290
rect 182031 530278 182185 530290
rect 182343 530304 182494 530328
rect 182031 530256 182041 530278
rect 181979 530168 182041 530256
rect 182343 530270 182351 530304
rect 182385 530294 182494 530304
rect 182385 530270 182395 530294
rect 182343 530244 182395 530270
rect 182531 530282 182589 530317
rect 182807 530302 182957 530372
rect 181979 530134 181997 530168
rect 182031 530134 182041 530168
rect 181979 530118 182041 530134
rect 182075 530228 182137 530244
rect 182075 530194 182083 530228
rect 182117 530194 182137 530228
rect 182075 530160 182137 530194
rect 182075 530126 182083 530160
rect 182117 530126 182137 530160
rect 182075 530084 182137 530126
rect 182171 530236 182395 530244
rect 182171 530210 182351 530236
rect 182171 530195 182223 530210
rect 182171 530186 182179 530195
rect 182171 530152 182175 530186
rect 182213 530161 182223 530195
rect 182343 530202 182351 530210
rect 182385 530202 182395 530236
rect 182209 530152 182223 530161
rect 182171 530118 182223 530152
rect 182257 530160 182308 530176
rect 182257 530126 182265 530160
rect 182299 530126 182308 530160
rect 182257 530084 182308 530126
rect 182343 530168 182395 530202
rect 182343 530134 182351 530168
rect 182385 530134 182395 530168
rect 182343 530118 182395 530134
rect 182429 530242 182486 530258
rect 182429 530208 182437 530242
rect 182471 530208 182486 530242
rect 182429 530174 182486 530208
rect 182429 530140 182437 530174
rect 182471 530140 182486 530174
rect 182429 530084 182486 530140
rect 182531 530248 182543 530282
rect 182577 530248 182589 530282
rect 182531 530189 182589 530248
rect 182531 530155 182543 530189
rect 182577 530155 182589 530189
rect 182531 530084 182589 530155
rect 182623 530262 182957 530302
rect 182623 530228 182641 530262
rect 182675 530228 182905 530262
rect 182939 530228 182957 530262
rect 182623 530160 182957 530228
rect 182623 530126 182641 530160
rect 182675 530126 182905 530160
rect 182939 530126 182957 530160
rect 182623 530084 182957 530126
rect 183083 530312 183117 530494
rect 183268 530492 183279 530526
rect 183318 530492 183327 530526
rect 183361 530514 183370 530548
rect 183404 530514 183412 530548
rect 183533 530548 183589 530594
rect 183361 530498 183412 530514
rect 183447 530526 183499 530542
rect 183268 530464 183327 530492
rect 183447 530492 183456 530526
rect 183490 530492 183499 530526
rect 183533 530514 183542 530548
rect 183576 530514 183589 530548
rect 183533 530498 183589 530514
rect 183635 530533 184704 530594
rect 183635 530499 183653 530533
rect 183687 530499 184653 530533
rect 184687 530499 184704 530533
rect 183447 530464 183499 530492
rect 183635 530485 184704 530499
rect 184739 530526 185073 530594
rect 184739 530492 184757 530526
rect 184791 530492 185021 530526
rect 185055 530492 185073 530526
rect 183151 530396 183221 530460
rect 183268 530430 183598 530464
rect 183185 530390 183221 530396
rect 183185 530362 183187 530390
rect 183151 530356 183187 530362
rect 183151 530346 183221 530356
rect 183255 530362 183297 530396
rect 183331 530362 183365 530396
rect 183399 530362 183433 530396
rect 183467 530362 183483 530396
rect 183255 530312 183289 530362
rect 183517 530328 183598 530430
rect 183083 530290 183289 530312
rect 183083 530256 183101 530290
rect 183135 530278 183289 530290
rect 183447 530304 183598 530328
rect 183952 530370 184020 530485
rect 184739 530440 185073 530492
rect 185107 530500 185165 530594
rect 185107 530466 185119 530500
rect 185153 530466 185165 530500
rect 185107 530449 185165 530466
rect 185199 530544 185259 530560
rect 185199 530510 185217 530544
rect 185251 530510 185259 530544
rect 185199 530494 185259 530510
rect 185293 530548 185348 530594
rect 185293 530514 185303 530548
rect 185337 530514 185348 530548
rect 185477 530548 185528 530594
rect 185293 530498 185348 530514
rect 185384 530526 185443 530542
rect 183952 530336 183969 530370
rect 184003 530336 184020 530370
rect 183952 530319 184020 530336
rect 184316 530406 184386 530421
rect 184316 530372 184333 530406
rect 184367 530372 184386 530406
rect 183135 530256 183145 530278
rect 183083 530168 183145 530256
rect 183447 530270 183455 530304
rect 183489 530294 183598 530304
rect 183489 530270 183499 530294
rect 183447 530244 183499 530270
rect 183083 530134 183101 530168
rect 183135 530134 183145 530168
rect 183083 530118 183145 530134
rect 183179 530228 183241 530244
rect 183179 530194 183187 530228
rect 183221 530194 183241 530228
rect 183179 530160 183241 530194
rect 183179 530126 183187 530160
rect 183221 530126 183241 530160
rect 183179 530084 183241 530126
rect 183275 530236 183499 530244
rect 183275 530210 183455 530236
rect 183275 530195 183327 530210
rect 183275 530161 183283 530195
rect 183317 530161 183327 530195
rect 183447 530202 183455 530210
rect 183489 530202 183499 530236
rect 183275 530118 183327 530161
rect 183361 530160 183412 530176
rect 183361 530126 183369 530160
rect 183403 530126 183412 530160
rect 183361 530084 183412 530126
rect 183447 530168 183499 530202
rect 183447 530134 183455 530168
rect 183489 530134 183499 530168
rect 183447 530118 183499 530134
rect 183533 530242 183590 530258
rect 183533 530208 183541 530242
rect 183575 530208 183590 530242
rect 183533 530174 183590 530208
rect 183533 530140 183541 530174
rect 183575 530140 183590 530174
rect 184316 530171 184386 530372
rect 184739 530370 184889 530440
rect 184739 530336 184759 530370
rect 184793 530336 184889 530370
rect 184923 530372 185019 530406
rect 185053 530372 185073 530406
rect 184923 530302 185073 530372
rect 184739 530262 185073 530302
rect 184739 530228 184757 530262
rect 184791 530228 185021 530262
rect 185055 530228 185073 530262
rect 183533 530084 183590 530140
rect 183635 530160 184704 530171
rect 183635 530126 183653 530160
rect 183687 530126 184653 530160
rect 184687 530126 184704 530160
rect 183635 530084 184704 530126
rect 184739 530160 185073 530228
rect 184739 530126 184757 530160
rect 184791 530126 185021 530160
rect 185055 530126 185073 530160
rect 184739 530084 185073 530126
rect 185107 530282 185165 530317
rect 185107 530248 185119 530282
rect 185153 530248 185165 530282
rect 185107 530189 185165 530248
rect 185107 530155 185119 530189
rect 185153 530155 185165 530189
rect 185107 530084 185165 530155
rect 185199 530312 185233 530494
rect 185384 530492 185395 530526
rect 185434 530492 185443 530526
rect 185477 530514 185486 530548
rect 185520 530514 185528 530548
rect 185649 530548 185705 530594
rect 185477 530498 185528 530514
rect 185563 530526 185615 530542
rect 185384 530464 185443 530492
rect 185563 530492 185572 530526
rect 185606 530492 185615 530526
rect 185649 530514 185658 530548
rect 185692 530514 185705 530548
rect 185649 530498 185705 530514
rect 185751 530533 186820 530594
rect 187085 530564 187153 530594
rect 185751 530499 185769 530533
rect 185803 530499 186769 530533
rect 186803 530499 186820 530533
rect 185563 530464 185615 530492
rect 185751 530485 186820 530499
rect 186947 530526 187001 530560
rect 187035 530526 187051 530560
rect 186947 530492 187051 530526
rect 185267 530458 185337 530460
rect 185267 530424 185303 530458
rect 185384 530430 185714 530464
rect 185267 530396 185337 530424
rect 185301 530362 185337 530396
rect 185267 530346 185337 530362
rect 185371 530362 185413 530396
rect 185447 530362 185481 530396
rect 185515 530362 185549 530396
rect 185583 530362 185599 530396
rect 185371 530312 185405 530362
rect 185633 530328 185714 530430
rect 185199 530290 185405 530312
rect 185199 530256 185217 530290
rect 185251 530278 185405 530290
rect 185563 530304 185714 530328
rect 186068 530370 186136 530485
rect 186947 530458 187001 530492
rect 187035 530458 187051 530492
rect 187085 530530 187101 530564
rect 187135 530530 187153 530564
rect 187085 530496 187153 530530
rect 187085 530462 187101 530496
rect 187135 530462 187153 530496
rect 187223 530531 187465 530594
rect 187223 530497 187241 530531
rect 187275 530497 187413 530531
rect 187447 530497 187465 530531
rect 186068 530336 186085 530370
rect 186119 530336 186136 530370
rect 186068 530319 186136 530336
rect 186432 530406 186502 530421
rect 186432 530372 186449 530406
rect 186483 530372 186502 530406
rect 185251 530256 185261 530278
rect 185199 530168 185261 530256
rect 185563 530270 185571 530304
rect 185605 530294 185714 530304
rect 185605 530270 185615 530294
rect 185563 530244 185615 530270
rect 185199 530134 185217 530168
rect 185251 530134 185261 530168
rect 185199 530118 185261 530134
rect 185295 530228 185357 530244
rect 185295 530194 185303 530228
rect 185337 530194 185357 530228
rect 185295 530160 185357 530194
rect 185295 530126 185303 530160
rect 185337 530126 185357 530160
rect 185295 530084 185357 530126
rect 185391 530236 185615 530244
rect 185391 530210 185571 530236
rect 185391 530195 185443 530210
rect 185391 530161 185399 530195
rect 185433 530161 185443 530195
rect 185563 530202 185571 530210
rect 185605 530202 185615 530236
rect 185391 530118 185443 530161
rect 185477 530160 185528 530176
rect 185477 530126 185485 530160
rect 185519 530126 185528 530160
rect 185477 530084 185528 530126
rect 185563 530168 185615 530202
rect 185563 530134 185571 530168
rect 185605 530134 185615 530168
rect 185563 530118 185615 530134
rect 185649 530242 185706 530258
rect 185649 530208 185657 530242
rect 185691 530208 185706 530242
rect 185649 530174 185706 530208
rect 185649 530140 185657 530174
rect 185691 530140 185706 530174
rect 186432 530171 186502 530372
rect 186947 530263 187051 530458
rect 187223 530444 187465 530497
rect 187085 530390 187189 530428
rect 187085 530356 187143 530390
rect 187177 530356 187189 530390
rect 187085 530229 187189 530356
rect 186985 530195 187001 530229
rect 187035 530195 187051 530229
rect 185649 530084 185706 530140
rect 185751 530160 186820 530171
rect 185751 530126 185769 530160
rect 185803 530126 186769 530160
rect 186803 530126 186820 530160
rect 185751 530084 186820 530126
rect 186985 530161 187051 530195
rect 186985 530127 187001 530161
rect 187035 530127 187051 530161
rect 186985 530084 187051 530127
rect 187085 530195 187101 530229
rect 187135 530195 187189 530229
rect 187085 530161 187189 530195
rect 187085 530127 187101 530161
rect 187135 530127 187189 530161
rect 187085 530118 187189 530127
rect 187223 530376 187273 530410
rect 187307 530376 187327 530410
rect 187223 530302 187327 530376
rect 187361 530370 187465 530444
rect 187361 530336 187381 530370
rect 187415 530336 187465 530370
rect 187223 530255 187465 530302
rect 187223 530221 187241 530255
rect 187275 530221 187413 530255
rect 187447 530221 187465 530255
rect 187223 530160 187465 530221
rect 187223 530126 187241 530160
rect 187275 530126 187413 530160
rect 187447 530126 187465 530160
rect 187223 530084 187465 530126
rect 172210 530050 172239 530084
rect 172273 530050 172331 530084
rect 172365 530050 172423 530084
rect 172457 530050 172515 530084
rect 172549 530050 172607 530084
rect 172641 530050 172699 530084
rect 172733 530050 172791 530084
rect 172825 530050 172883 530084
rect 172917 530050 172975 530084
rect 173009 530050 173067 530084
rect 173101 530050 173159 530084
rect 173193 530050 173251 530084
rect 173285 530050 173343 530084
rect 173377 530050 173435 530084
rect 173469 530050 173527 530084
rect 173561 530050 173619 530084
rect 173653 530050 173711 530084
rect 173745 530050 173803 530084
rect 173837 530050 173895 530084
rect 173929 530050 173987 530084
rect 174021 530050 174079 530084
rect 174113 530050 174171 530084
rect 174205 530050 174263 530084
rect 174297 530050 174355 530084
rect 174389 530050 174447 530084
rect 174481 530050 174539 530084
rect 174573 530050 174631 530084
rect 174665 530050 174723 530084
rect 174757 530050 174815 530084
rect 174849 530050 174907 530084
rect 174941 530050 174999 530084
rect 175033 530050 175091 530084
rect 175125 530050 175183 530084
rect 175217 530050 175275 530084
rect 175309 530050 175367 530084
rect 175401 530050 175459 530084
rect 175493 530050 175551 530084
rect 175585 530050 175643 530084
rect 175677 530050 175735 530084
rect 175769 530050 175827 530084
rect 175861 530050 175919 530084
rect 175953 530050 176011 530084
rect 176045 530050 176103 530084
rect 176137 530050 176195 530084
rect 176229 530050 176287 530084
rect 176321 530050 176379 530084
rect 176413 530050 176471 530084
rect 176505 530050 176563 530084
rect 176597 530050 176655 530084
rect 176689 530050 176747 530084
rect 176781 530050 176839 530084
rect 176873 530050 176931 530084
rect 176965 530050 177023 530084
rect 177057 530050 177115 530084
rect 177149 530050 177207 530084
rect 177241 530050 177299 530084
rect 177333 530050 177391 530084
rect 177425 530050 177483 530084
rect 177517 530050 177575 530084
rect 177609 530050 177667 530084
rect 177701 530050 177759 530084
rect 177793 530050 177851 530084
rect 177885 530050 177943 530084
rect 177977 530050 178035 530084
rect 178069 530050 178127 530084
rect 178161 530050 178219 530084
rect 178253 530050 178311 530084
rect 178345 530050 178403 530084
rect 178437 530050 178495 530084
rect 178529 530050 178587 530084
rect 178621 530050 178679 530084
rect 178713 530050 178771 530084
rect 178805 530050 178863 530084
rect 178897 530050 178955 530084
rect 178989 530050 179047 530084
rect 179081 530050 179139 530084
rect 179173 530050 179231 530084
rect 179265 530050 179323 530084
rect 179357 530050 179415 530084
rect 179449 530050 179507 530084
rect 179541 530050 179599 530084
rect 179633 530050 179691 530084
rect 179725 530050 179783 530084
rect 179817 530050 179875 530084
rect 179909 530050 179967 530084
rect 180001 530050 180059 530084
rect 180093 530050 180151 530084
rect 180185 530050 180243 530084
rect 180277 530050 180335 530084
rect 180369 530050 180427 530084
rect 180461 530050 180519 530084
rect 180553 530050 180611 530084
rect 180645 530050 180703 530084
rect 180737 530050 180795 530084
rect 180829 530050 180887 530084
rect 180921 530050 180979 530084
rect 181013 530050 181071 530084
rect 181105 530050 181163 530084
rect 181197 530050 181255 530084
rect 181289 530050 181347 530084
rect 181381 530050 181439 530084
rect 181473 530050 181531 530084
rect 181565 530050 181623 530084
rect 181657 530050 181715 530084
rect 181749 530050 181807 530084
rect 181841 530050 181899 530084
rect 181933 530050 181991 530084
rect 182025 530050 182083 530084
rect 182117 530050 182175 530084
rect 182209 530050 182267 530084
rect 182301 530050 182359 530084
rect 182393 530050 182451 530084
rect 182485 530050 182543 530084
rect 182577 530050 182635 530084
rect 182669 530050 182727 530084
rect 182761 530050 182819 530084
rect 182853 530050 182911 530084
rect 182945 530050 183003 530084
rect 183037 530050 183095 530084
rect 183129 530050 183187 530084
rect 183221 530050 183279 530084
rect 183313 530050 183371 530084
rect 183405 530050 183463 530084
rect 183497 530050 183555 530084
rect 183589 530050 183647 530084
rect 183681 530050 183739 530084
rect 183773 530050 183831 530084
rect 183865 530050 183923 530084
rect 183957 530050 184015 530084
rect 184049 530050 184107 530084
rect 184141 530050 184199 530084
rect 184233 530050 184291 530084
rect 184325 530050 184383 530084
rect 184417 530050 184475 530084
rect 184509 530050 184567 530084
rect 184601 530050 184659 530084
rect 184693 530050 184751 530084
rect 184785 530050 184843 530084
rect 184877 530050 184935 530084
rect 184969 530050 185027 530084
rect 185061 530050 185119 530084
rect 185153 530050 185211 530084
rect 185245 530050 185303 530084
rect 185337 530050 185395 530084
rect 185429 530050 185487 530084
rect 185521 530050 185579 530084
rect 185613 530050 185671 530084
rect 185705 530050 185763 530084
rect 185797 530050 185855 530084
rect 185889 530050 185947 530084
rect 185981 530050 186039 530084
rect 186073 530050 186131 530084
rect 186165 530050 186223 530084
rect 186257 530050 186315 530084
rect 186349 530050 186407 530084
rect 186441 530050 186499 530084
rect 186533 530050 186591 530084
rect 186625 530050 186683 530084
rect 186717 530050 186775 530084
rect 186809 530050 186867 530084
rect 186901 530050 186959 530084
rect 186993 530050 187051 530084
rect 187085 530050 187143 530084
rect 187177 530050 187235 530084
rect 187269 530050 187327 530084
rect 187361 530050 187419 530084
rect 187453 530050 187482 530084
rect 172227 530008 172469 530050
rect 172227 529974 172245 530008
rect 172279 529974 172417 530008
rect 172451 529974 172469 530008
rect 172227 529913 172469 529974
rect 172503 530008 173572 530050
rect 172503 529974 172521 530008
rect 172555 529974 173521 530008
rect 173555 529974 173572 530008
rect 172503 529963 173572 529974
rect 173607 530008 174676 530050
rect 173607 529974 173625 530008
rect 173659 529974 174625 530008
rect 174659 529974 174676 530008
rect 173607 529963 174676 529974
rect 174826 529982 174883 530016
rect 172227 529879 172245 529913
rect 172279 529879 172417 529913
rect 172451 529879 172469 529913
rect 172227 529832 172469 529879
rect 172227 529764 172277 529798
rect 172311 529764 172331 529798
rect 172227 529690 172331 529764
rect 172365 529758 172469 529832
rect 172365 529724 172385 529758
rect 172419 529724 172469 529758
rect 172820 529798 172888 529815
rect 172820 529764 172837 529798
rect 172871 529764 172888 529798
rect 172227 529637 172469 529690
rect 172820 529649 172888 529764
rect 173184 529762 173254 529963
rect 173184 529728 173201 529762
rect 173235 529728 173254 529762
rect 173184 529713 173254 529728
rect 173924 529798 173992 529815
rect 173924 529764 173941 529798
rect 173975 529764 173992 529798
rect 173924 529649 173992 529764
rect 174288 529762 174358 529963
rect 174826 529948 174843 529982
rect 174877 529948 174883 529982
rect 174917 530008 174971 530050
rect 174917 529974 174927 530008
rect 174961 529974 174971 530008
rect 174917 529958 174971 529974
rect 175051 529982 175131 530016
rect 174826 529924 174883 529948
rect 175051 529948 175081 529982
rect 175115 529948 175131 529982
rect 174826 529880 175017 529924
rect 174288 529728 174305 529762
rect 174339 529728 174358 529762
rect 174803 529812 174815 529846
rect 174849 529812 174941 529846
rect 174803 529772 174941 529812
rect 174803 529738 174867 529772
rect 174901 529738 174941 529772
rect 174803 529734 174941 529738
rect 174975 529772 175017 529880
rect 174975 529738 174981 529772
rect 175015 529738 175017 529772
rect 174288 529713 174358 529728
rect 174975 529700 175017 529738
rect 174826 529666 175017 529700
rect 175051 529846 175131 529948
rect 175169 529982 175225 530016
rect 175169 529948 175185 529982
rect 175219 529948 175225 529982
rect 175329 530008 175394 530050
rect 175329 529974 175344 530008
rect 175378 529974 175394 530008
rect 175329 529958 175394 529974
rect 175428 529982 175505 530016
rect 175169 529924 175225 529948
rect 175428 529948 175434 529982
rect 175468 529948 175505 529982
rect 175169 529880 175394 529924
rect 175051 529772 175270 529846
rect 175051 529738 175185 529772
rect 175219 529738 175270 529772
rect 175051 529734 175270 529738
rect 175304 529788 175394 529880
rect 175428 529822 175505 529948
rect 175540 530000 175591 530016
rect 175540 529966 175557 530000
rect 175540 529932 175591 529966
rect 175625 529984 175691 530050
rect 175625 529950 175641 529984
rect 175675 529950 175691 529984
rect 175725 530000 175759 530016
rect 175540 529898 175557 529932
rect 175725 529932 175759 529966
rect 175591 529898 175690 529916
rect 175540 529882 175690 529898
rect 175304 529772 175415 529788
rect 175304 529738 175381 529772
rect 172227 529603 172245 529637
rect 172279 529603 172417 529637
rect 172451 529603 172469 529637
rect 172227 529540 172469 529603
rect 172503 529635 173572 529649
rect 172503 529601 172521 529635
rect 172555 529601 173521 529635
rect 173555 529601 173572 529635
rect 172503 529540 173572 529601
rect 173607 529635 174676 529649
rect 173607 529601 173625 529635
rect 173659 529601 174625 529635
rect 174659 529601 174676 529635
rect 173607 529540 174676 529601
rect 174826 529642 174883 529666
rect 174826 529608 174843 529642
rect 174877 529608 174883 529642
rect 175051 529642 175131 529734
rect 175304 529722 175415 529738
rect 175304 529700 175394 529722
rect 174826 529574 174883 529608
rect 174917 529616 174971 529632
rect 174917 529582 174927 529616
rect 174961 529582 174971 529616
rect 174917 529540 174971 529582
rect 175051 529608 175081 529642
rect 175115 529608 175131 529642
rect 175051 529574 175131 529608
rect 175169 529666 175394 529700
rect 175449 529688 175505 529822
rect 175540 529778 175610 529848
rect 175540 529744 175551 529778
rect 175585 529772 175610 529778
rect 175540 529738 175554 529744
rect 175588 529738 175610 529772
rect 175540 529718 175610 529738
rect 175644 529787 175690 529882
rect 175644 529778 175656 529787
rect 175678 529744 175690 529753
rect 175169 529642 175225 529666
rect 175169 529608 175185 529642
rect 175219 529608 175225 529642
rect 175428 529642 175505 529688
rect 175644 529684 175690 529744
rect 175169 529574 175225 529608
rect 175329 529616 175394 529632
rect 175329 529582 175344 529616
rect 175378 529582 175394 529616
rect 175329 529540 175394 529582
rect 175428 529608 175434 529642
rect 175493 529608 175505 529642
rect 175428 529574 175505 529608
rect 175540 529650 175690 529684
rect 175540 529642 175591 529650
rect 175540 529608 175557 529642
rect 175725 529642 175759 529880
rect 175793 529856 175858 530013
rect 175892 530008 175942 530050
rect 175892 529974 175908 530008
rect 175892 529958 175942 529974
rect 175976 530000 176026 530016
rect 175976 529966 175992 530000
rect 175976 529950 176026 529966
rect 176069 530006 176205 530016
rect 176069 529972 176085 530006
rect 176119 529972 176205 530006
rect 176320 529998 176386 530050
rect 176513 530008 176587 530050
rect 176069 529950 176205 529972
rect 175976 529924 176010 529950
rect 175931 529890 176010 529924
rect 176044 529914 176137 529916
rect 175805 529846 175897 529856
rect 175805 529812 175827 529846
rect 175861 529833 175897 529846
rect 175861 529812 175863 529833
rect 175805 529799 175863 529812
rect 175805 529646 175897 529799
rect 175540 529592 175591 529608
rect 175625 529582 175641 529616
rect 175675 529582 175691 529616
rect 175931 529618 175965 529890
rect 176044 529888 176103 529914
rect 176078 529880 176103 529888
rect 176078 529854 176137 529880
rect 176044 529838 176137 529854
rect 175999 529778 176069 529800
rect 175999 529744 176011 529778
rect 176045 529744 176069 529778
rect 175999 529726 176069 529744
rect 175999 529692 176022 529726
rect 176056 529692 176069 529726
rect 175999 529676 176069 529692
rect 176103 529720 176137 529838
rect 176171 529794 176205 529950
rect 176239 529982 176273 529998
rect 176320 529964 176336 529998
rect 176370 529964 176386 529998
rect 176420 529982 176454 529998
rect 176239 529930 176273 529948
rect 176513 529974 176533 530008
rect 176567 529974 176587 530008
rect 176513 529958 176587 529974
rect 176621 530000 176655 530016
rect 176420 529930 176454 529948
rect 176239 529896 176454 529930
rect 176621 529924 176655 529966
rect 176702 530007 176876 530016
rect 176702 529973 176718 530007
rect 176752 529973 176876 530007
rect 176702 529948 176876 529973
rect 176910 530008 176960 530050
rect 176944 529974 176960 530008
rect 177064 530008 177130 530050
rect 176910 529958 176960 529974
rect 176994 529982 177028 529998
rect 176543 529890 176655 529924
rect 176543 529862 176577 529890
rect 176277 529828 176293 529862
rect 176327 529828 176577 529862
rect 176716 529880 176727 529914
rect 176761 529888 176808 529914
rect 176716 529856 176758 529880
rect 176171 529774 176509 529794
rect 176171 529760 176475 529774
rect 176103 529686 176124 529720
rect 176158 529686 176174 529720
rect 176103 529676 176174 529686
rect 176208 529618 176242 529760
rect 176283 529710 176379 529726
rect 176317 529676 176355 529710
rect 176413 529692 176441 529726
rect 176475 529724 176509 529740
rect 176389 529676 176441 529692
rect 176543 529690 176577 529828
rect 175725 529592 175759 529608
rect 175625 529540 175691 529582
rect 175831 529578 175847 529612
rect 175881 529578 175897 529612
rect 175931 529584 175980 529618
rect 176014 529584 176030 529618
rect 176071 529584 176087 529618
rect 176121 529584 176242 529618
rect 176417 529616 176483 529632
rect 175831 529540 175897 529578
rect 176417 529582 176433 529616
rect 176467 529582 176483 529616
rect 176417 529540 176483 529582
rect 176525 529612 176577 529690
rect 176615 529854 176758 529856
rect 176792 529854 176808 529888
rect 176842 529872 176876 529948
rect 177064 529974 177080 530008
rect 177114 529974 177130 530008
rect 177198 530008 177259 530050
rect 177198 529974 177209 530008
rect 177243 529974 177259 530008
rect 176994 529940 177028 529948
rect 177198 529940 177259 529974
rect 176994 529906 177154 529940
rect 176615 529822 176750 529854
rect 176842 529838 177036 529872
rect 177070 529838 177086 529872
rect 176615 529714 176657 529822
rect 176842 529820 176876 529838
rect 176615 529680 176623 529714
rect 176615 529664 176657 529680
rect 176691 529778 176761 529788
rect 176691 529762 176727 529778
rect 176691 529728 176719 529762
rect 176753 529728 176761 529744
rect 176691 529664 176761 529728
rect 176795 529786 176876 529820
rect 176795 529630 176829 529786
rect 176943 529773 177051 529804
rect 177120 529788 177154 529906
rect 177198 529906 177209 529940
rect 177243 529906 177259 529940
rect 177198 529822 177259 529906
rect 177293 529982 177344 529988
rect 177293 529972 177299 529982
rect 177333 529948 177344 529982
rect 177327 529938 177344 529948
rect 177293 529904 177344 529938
rect 177327 529870 177344 529904
rect 177293 529812 177344 529870
rect 177379 529979 177437 530050
rect 177379 529945 177391 529979
rect 177425 529945 177437 529979
rect 177379 529886 177437 529945
rect 177379 529852 177391 529886
rect 177425 529852 177437 529886
rect 177379 529817 177437 529852
rect 177563 529948 177666 529980
rect 177563 529914 177627 529948
rect 177661 529914 177666 529948
rect 177563 529898 177666 529914
rect 177713 529948 177747 530050
rect 177713 529898 177747 529914
rect 177781 529982 178187 530016
rect 177120 529782 177268 529788
rect 176977 529764 177051 529773
rect 176863 529736 176907 529752
rect 176897 529702 176907 529736
rect 176943 529730 176959 529739
rect 176993 529730 177051 529764
rect 176863 529696 176907 529702
rect 177003 529710 177051 529730
rect 176863 529662 176969 529696
rect 176639 529616 176829 529630
rect 176525 529578 176545 529612
rect 176579 529578 176595 529612
rect 176639 529582 176655 529616
rect 176689 529582 176829 529616
rect 176639 529574 176829 529582
rect 176863 529612 176901 529628
rect 176863 529578 176867 529612
rect 176935 529616 176969 529662
rect 177037 529676 177051 529710
rect 177003 529650 177051 529676
rect 177085 529772 177268 529782
rect 177085 529738 177234 529772
rect 177085 529722 177268 529738
rect 177085 529687 177150 529722
rect 177085 529632 177149 529687
rect 177302 529682 177344 529812
rect 177563 529736 177631 529898
rect 177781 529849 177815 529982
rect 177894 529914 177910 529948
rect 177944 529914 177985 529948
rect 178019 529914 178119 529948
rect 177665 529846 177681 529849
rect 177665 529812 177667 529846
rect 177715 529815 177815 529849
rect 177701 529812 177815 529815
rect 177665 529811 177815 529812
rect 177849 529849 178051 529880
rect 177883 529846 178051 529849
rect 177883 529815 177887 529846
rect 177563 529702 177759 529736
rect 177793 529702 177809 529736
rect 177849 529710 177887 529815
rect 177293 529666 177344 529682
rect 177327 529632 177344 529666
rect 176935 529598 177085 529616
rect 177119 529598 177149 529632
rect 176935 529582 177149 529598
rect 177198 529616 177259 529632
rect 177198 529582 177209 529616
rect 177243 529582 177259 529616
rect 176863 529540 176901 529578
rect 177198 529540 177259 529582
rect 177293 529576 177344 529632
rect 177379 529668 177437 529685
rect 177379 529634 177391 529668
rect 177425 529634 177437 529668
rect 177379 529540 177437 529634
rect 177618 529631 177667 529702
rect 177849 529676 177851 529710
rect 177885 529676 177887 529710
rect 177618 529597 177627 529631
rect 177661 529597 177667 529631
rect 177618 529581 177667 529597
rect 177711 529631 177813 529647
rect 177745 529597 177779 529631
rect 177711 529540 177813 529597
rect 177849 529574 177887 529676
rect 177921 529778 177976 529806
rect 177921 529744 177943 529778
rect 177921 529736 177976 529744
rect 177955 529702 177976 529736
rect 177921 529574 177976 529702
rect 178017 529736 178051 529846
rect 178017 529686 178051 529702
rect 178085 529688 178119 529914
rect 178153 529788 178187 529982
rect 178221 530008 178255 530050
rect 178221 529940 178255 529974
rect 178221 529872 178255 529906
rect 178221 529822 178255 529838
rect 178289 530008 178356 530016
rect 178289 529974 178305 530008
rect 178339 529974 178356 530008
rect 178477 530008 178538 530050
rect 178289 529940 178356 529974
rect 178289 529906 178305 529940
rect 178339 529914 178356 529940
rect 178289 529880 178311 529906
rect 178345 529880 178356 529914
rect 178289 529872 178356 529880
rect 178289 529838 178305 529872
rect 178339 529838 178356 529872
rect 178289 529822 178356 529838
rect 178153 529772 178192 529788
rect 178153 529738 178158 529772
rect 178153 529722 178192 529738
rect 178237 529772 178288 529788
rect 178237 529738 178254 529772
rect 178237 529722 178288 529738
rect 178237 529688 178271 529722
rect 178322 529688 178356 529822
rect 178085 529654 178271 529688
rect 178085 529647 178120 529654
rect 178014 529631 178120 529647
rect 178048 529597 178120 529631
rect 178305 529635 178356 529688
rect 178014 529574 178120 529597
rect 178205 529616 178271 529620
rect 178205 529582 178221 529616
rect 178255 529582 178271 529616
rect 178205 529540 178271 529582
rect 178339 529601 178356 529635
rect 178305 529574 178356 529601
rect 178392 529982 178443 529988
rect 178392 529948 178403 529982
rect 178437 529972 178443 529982
rect 178392 529938 178409 529948
rect 178392 529904 178443 529938
rect 178392 529870 178409 529904
rect 178392 529812 178443 529870
rect 178477 529974 178493 530008
rect 178527 529974 178538 530008
rect 178606 530008 178672 530050
rect 178606 529974 178622 530008
rect 178656 529974 178672 530008
rect 178776 530008 178826 530050
rect 178708 529982 178742 529998
rect 178477 529940 178538 529974
rect 178776 529974 178792 530008
rect 178776 529958 178826 529974
rect 178860 530007 179034 530016
rect 178860 529973 178984 530007
rect 179018 529973 179034 530007
rect 178708 529940 178742 529948
rect 178477 529906 178493 529940
rect 178527 529906 178538 529940
rect 178477 529822 178538 529906
rect 178582 529906 178742 529940
rect 178860 529948 179034 529973
rect 179081 530000 179115 530016
rect 178392 529682 178434 529812
rect 178582 529788 178616 529906
rect 178860 529872 178894 529948
rect 179081 529924 179115 529966
rect 179149 530008 179223 530050
rect 179149 529974 179169 530008
rect 179203 529974 179223 530008
rect 179350 529998 179416 530050
rect 179531 530006 179667 530016
rect 179149 529958 179223 529974
rect 179282 529982 179316 529998
rect 179350 529964 179366 529998
rect 179400 529964 179416 529998
rect 179463 529982 179497 529998
rect 179282 529930 179316 529948
rect 179463 529930 179497 529948
rect 178650 529838 178666 529872
rect 178700 529838 178894 529872
rect 178928 529888 178975 529914
rect 178928 529854 178944 529888
rect 179009 529880 179020 529914
rect 179081 529890 179193 529924
rect 179282 529896 179497 529930
rect 179531 529972 179617 530006
rect 179651 529972 179667 530006
rect 179531 529950 179667 529972
rect 179710 530000 179760 530016
rect 179744 529966 179760 530000
rect 179710 529950 179760 529966
rect 179794 530008 179844 530050
rect 179828 529974 179844 530008
rect 179794 529958 179844 529974
rect 178978 529856 179020 529880
rect 179159 529862 179193 529890
rect 178978 529854 179121 529856
rect 178860 529820 178894 529838
rect 178986 529822 179121 529854
rect 178468 529782 178616 529788
rect 178468 529772 178651 529782
rect 178502 529738 178651 529772
rect 178468 529722 178651 529738
rect 178586 529687 178651 529722
rect 178392 529666 178443 529682
rect 178392 529632 178409 529666
rect 178587 529632 178651 529687
rect 178685 529773 178793 529804
rect 178860 529786 178941 529820
rect 178685 529764 178759 529773
rect 178685 529730 178743 529764
rect 178777 529730 178793 529739
rect 178829 529736 178873 529752
rect 178685 529710 178733 529730
rect 178685 529676 178699 529710
rect 178829 529702 178839 529736
rect 178829 529696 178873 529702
rect 178685 529650 178733 529676
rect 178767 529662 178873 529696
rect 178392 529576 178443 529632
rect 178477 529616 178538 529632
rect 178477 529582 178493 529616
rect 178527 529582 178538 529616
rect 178587 529598 178617 529632
rect 178767 529616 178801 529662
rect 178907 529630 178941 529786
rect 178975 529778 179045 529788
rect 179009 529762 179045 529778
rect 178975 529728 178983 529744
rect 179017 529728 179045 529762
rect 178975 529664 179045 529728
rect 179079 529714 179121 529822
rect 179113 529680 179121 529714
rect 179079 529664 179121 529680
rect 179159 529828 179409 529862
rect 179443 529828 179459 529862
rect 179159 529690 179193 529828
rect 179531 529794 179565 529950
rect 179726 529924 179760 529950
rect 179227 529774 179565 529794
rect 179261 529760 179565 529774
rect 179599 529914 179692 529916
rect 179633 529888 179692 529914
rect 179726 529890 179805 529924
rect 179633 529880 179658 529888
rect 179599 529854 179658 529880
rect 179599 529838 179692 529854
rect 179227 529724 179261 529740
rect 179295 529692 179323 529726
rect 179357 529710 179453 529726
rect 178651 529598 178801 529616
rect 178587 529582 178801 529598
rect 178835 529612 178873 529628
rect 178477 529540 178538 529582
rect 178869 529578 178873 529612
rect 178835 529540 178873 529578
rect 178907 529616 179097 529630
rect 178907 529582 179047 529616
rect 179081 529582 179097 529616
rect 179159 529612 179211 529690
rect 179295 529676 179347 529692
rect 179381 529676 179419 529710
rect 178907 529574 179097 529582
rect 179141 529578 179157 529612
rect 179191 529578 179211 529612
rect 179253 529616 179319 529632
rect 179253 529582 179269 529616
rect 179303 529582 179319 529616
rect 179494 529618 179528 529760
rect 179599 529720 179633 529838
rect 179562 529686 179578 529720
rect 179612 529686 179633 529720
rect 179562 529676 179633 529686
rect 179667 529778 179737 529800
rect 179667 529744 179691 529778
rect 179725 529744 179737 529778
rect 179667 529726 179737 529744
rect 179667 529692 179680 529726
rect 179714 529692 179737 529726
rect 179667 529676 179737 529692
rect 179771 529618 179805 529890
rect 179878 529856 179943 530013
rect 179977 530000 180011 530016
rect 179977 529932 180011 529966
rect 180045 529984 180111 530050
rect 180045 529950 180061 529984
rect 180095 529950 180111 529984
rect 180145 530000 180196 530016
rect 180179 529966 180196 530000
rect 180145 529932 180196 529966
rect 179839 529846 179931 529856
rect 179839 529833 179875 529846
rect 179873 529812 179875 529833
rect 179909 529812 179931 529846
rect 179873 529799 179931 529812
rect 179839 529646 179931 529799
rect 179494 529584 179615 529618
rect 179649 529584 179665 529618
rect 179706 529584 179722 529618
rect 179756 529584 179805 529618
rect 179977 529642 180011 529880
rect 180046 529898 180145 529916
rect 180179 529898 180196 529932
rect 180046 529882 180196 529898
rect 180232 530000 180283 530016
rect 180232 529966 180249 530000
rect 180232 529932 180283 529966
rect 180317 529984 180383 530050
rect 180317 529950 180333 529984
rect 180367 529950 180383 529984
rect 180417 530000 180451 530016
rect 180232 529898 180249 529932
rect 180417 529932 180451 529966
rect 180283 529898 180382 529916
rect 180232 529882 180382 529898
rect 180046 529787 180092 529882
rect 180080 529778 180092 529787
rect 180046 529744 180058 529753
rect 180046 529684 180092 529744
rect 180126 529778 180196 529848
rect 180126 529772 180151 529778
rect 180126 529738 180148 529772
rect 180185 529744 180196 529778
rect 180182 529738 180196 529744
rect 180126 529718 180196 529738
rect 180232 529778 180302 529848
rect 180232 529744 180243 529778
rect 180277 529772 180302 529778
rect 180232 529738 180246 529744
rect 180280 529738 180302 529772
rect 180232 529718 180302 529738
rect 180336 529787 180382 529882
rect 180336 529778 180348 529787
rect 180370 529744 180382 529753
rect 180336 529684 180382 529744
rect 180046 529650 180196 529684
rect 179253 529540 179319 529582
rect 179839 529578 179855 529612
rect 179889 529578 179905 529612
rect 180145 529642 180196 529650
rect 179977 529592 180011 529608
rect 179839 529540 179905 529578
rect 180045 529582 180061 529616
rect 180095 529582 180111 529616
rect 180179 529608 180196 529642
rect 180145 529592 180196 529608
rect 180232 529650 180382 529684
rect 180232 529642 180283 529650
rect 180232 529608 180249 529642
rect 180417 529642 180451 529880
rect 180485 529856 180550 530013
rect 180584 530008 180634 530050
rect 180584 529974 180600 530008
rect 180584 529958 180634 529974
rect 180668 530000 180718 530016
rect 180668 529966 180684 530000
rect 180668 529950 180718 529966
rect 180761 530006 180897 530016
rect 180761 529972 180777 530006
rect 180811 529972 180897 530006
rect 181012 529998 181078 530050
rect 181205 530008 181279 530050
rect 180761 529950 180897 529972
rect 180668 529924 180702 529950
rect 180623 529890 180702 529924
rect 180736 529914 180829 529916
rect 180497 529846 180589 529856
rect 180497 529812 180519 529846
rect 180553 529833 180589 529846
rect 180553 529812 180555 529833
rect 180497 529799 180555 529812
rect 180497 529646 180589 529799
rect 180232 529592 180283 529608
rect 180045 529540 180111 529582
rect 180317 529582 180333 529616
rect 180367 529582 180383 529616
rect 180623 529618 180657 529890
rect 180736 529888 180795 529914
rect 180770 529880 180795 529888
rect 180770 529854 180829 529880
rect 180736 529838 180829 529854
rect 180691 529778 180761 529800
rect 180691 529744 180703 529778
rect 180737 529744 180761 529778
rect 180691 529726 180761 529744
rect 180691 529692 180714 529726
rect 180748 529692 180761 529726
rect 180691 529676 180761 529692
rect 180795 529720 180829 529838
rect 180863 529794 180897 529950
rect 180931 529982 180965 529998
rect 181012 529964 181028 529998
rect 181062 529964 181078 529998
rect 181112 529982 181146 529998
rect 180931 529930 180965 529948
rect 181205 529974 181225 530008
rect 181259 529974 181279 530008
rect 181205 529958 181279 529974
rect 181313 530000 181347 530016
rect 181112 529930 181146 529948
rect 180931 529896 181146 529930
rect 181313 529924 181347 529966
rect 181394 530007 181568 530016
rect 181394 529973 181410 530007
rect 181444 529973 181568 530007
rect 181394 529948 181568 529973
rect 181602 530008 181652 530050
rect 181636 529974 181652 530008
rect 181756 530008 181822 530050
rect 181602 529958 181652 529974
rect 181686 529982 181720 529998
rect 181235 529890 181347 529924
rect 181235 529862 181269 529890
rect 180969 529828 180985 529862
rect 181019 529828 181269 529862
rect 181408 529880 181419 529914
rect 181453 529888 181500 529914
rect 181408 529856 181450 529880
rect 180863 529774 181201 529794
rect 180863 529760 181167 529774
rect 180795 529686 180816 529720
rect 180850 529686 180866 529720
rect 180795 529676 180866 529686
rect 180900 529618 180934 529760
rect 180975 529710 181071 529726
rect 181009 529676 181047 529710
rect 181105 529692 181133 529726
rect 181167 529724 181201 529740
rect 181081 529676 181133 529692
rect 181235 529690 181269 529828
rect 180417 529592 180451 529608
rect 180317 529540 180383 529582
rect 180523 529578 180539 529612
rect 180573 529578 180589 529612
rect 180623 529584 180672 529618
rect 180706 529584 180722 529618
rect 180763 529584 180779 529618
rect 180813 529584 180934 529618
rect 181109 529616 181175 529632
rect 180523 529540 180589 529578
rect 181109 529582 181125 529616
rect 181159 529582 181175 529616
rect 181109 529540 181175 529582
rect 181217 529612 181269 529690
rect 181307 529854 181450 529856
rect 181484 529854 181500 529888
rect 181534 529872 181568 529948
rect 181756 529974 181772 530008
rect 181806 529974 181822 530008
rect 181890 530008 181951 530050
rect 181890 529974 181901 530008
rect 181935 529974 181951 530008
rect 182071 530008 182405 530050
rect 181686 529940 181720 529948
rect 181890 529940 181951 529974
rect 181686 529906 181846 529940
rect 181307 529822 181442 529854
rect 181534 529838 181728 529872
rect 181762 529838 181778 529872
rect 181307 529714 181349 529822
rect 181534 529820 181568 529838
rect 181307 529680 181315 529714
rect 181307 529664 181349 529680
rect 181383 529778 181453 529788
rect 181383 529762 181419 529778
rect 181383 529728 181411 529762
rect 181445 529728 181453 529744
rect 181383 529664 181453 529728
rect 181487 529786 181568 529820
rect 181487 529630 181521 529786
rect 181635 529773 181743 529804
rect 181812 529788 181846 529906
rect 181890 529906 181901 529940
rect 181935 529906 181951 529940
rect 181890 529822 181951 529906
rect 181985 529972 182036 529988
rect 182019 529938 182036 529972
rect 181985 529904 182036 529938
rect 182019 529870 182036 529904
rect 181985 529846 182036 529870
rect 181985 529812 181991 529846
rect 182025 529812 182036 529846
rect 182071 529974 182089 530008
rect 182123 529974 182353 530008
rect 182387 529974 182405 530008
rect 182071 529906 182405 529974
rect 182071 529872 182089 529906
rect 182123 529872 182353 529906
rect 182387 529872 182405 529906
rect 182071 529832 182405 529872
rect 181812 529782 181960 529788
rect 181669 529764 181743 529773
rect 181555 529736 181599 529752
rect 181589 529702 181599 529736
rect 181635 529730 181651 529739
rect 181685 529730 181743 529764
rect 181555 529696 181599 529702
rect 181695 529710 181743 529730
rect 181555 529662 181661 529696
rect 181331 529616 181521 529630
rect 181217 529578 181237 529612
rect 181271 529578 181287 529612
rect 181331 529582 181347 529616
rect 181381 529582 181521 529616
rect 181331 529574 181521 529582
rect 181555 529612 181593 529628
rect 181555 529578 181559 529612
rect 181627 529616 181661 529662
rect 181729 529676 181743 529710
rect 181695 529650 181743 529676
rect 181777 529772 181960 529782
rect 181777 529738 181926 529772
rect 181777 529722 181960 529738
rect 181777 529687 181842 529722
rect 181777 529632 181841 529687
rect 181994 529682 182036 529812
rect 181985 529666 182036 529682
rect 182019 529632 182036 529666
rect 181627 529598 181777 529616
rect 181811 529598 181841 529632
rect 181627 529582 181841 529598
rect 181890 529616 181951 529632
rect 181890 529582 181901 529616
rect 181935 529582 181951 529616
rect 181555 529540 181593 529578
rect 181890 529540 181951 529582
rect 181985 529576 182036 529632
rect 182071 529764 182091 529798
rect 182125 529764 182221 529798
rect 182071 529694 182221 529764
rect 182255 529762 182405 529832
rect 182531 529979 182589 530050
rect 182531 529945 182543 529979
rect 182577 529945 182589 529979
rect 182531 529886 182589 529945
rect 182531 529852 182543 529886
rect 182577 529852 182589 529886
rect 182531 529817 182589 529852
rect 182623 529982 182700 530016
rect 182623 529948 182635 529982
rect 182694 529948 182700 529982
rect 182734 530008 182799 530050
rect 182734 529974 182750 530008
rect 182784 529974 182799 530008
rect 182734 529958 182799 529974
rect 182903 529982 182959 530016
rect 182623 529822 182700 529948
rect 182903 529948 182909 529982
rect 182943 529948 182959 529982
rect 182903 529924 182959 529948
rect 182734 529880 182959 529924
rect 182997 529982 183077 530016
rect 182997 529948 183013 529982
rect 183047 529948 183077 529982
rect 183157 530008 183211 530050
rect 183157 529974 183167 530008
rect 183201 529974 183211 530008
rect 183157 529958 183211 529974
rect 183245 529982 183302 530016
rect 182255 529728 182351 529762
rect 182385 529728 182405 529762
rect 182071 529642 182405 529694
rect 182623 529688 182679 529822
rect 182734 529788 182824 529880
rect 182997 529846 183077 529948
rect 183245 529948 183251 529982
rect 183285 529948 183302 529982
rect 183359 530008 184428 530050
rect 183359 529974 183377 530008
rect 183411 529974 184377 530008
rect 184411 529974 184428 530008
rect 183359 529963 184428 529974
rect 184463 530008 185532 530050
rect 184463 529974 184481 530008
rect 184515 529974 185481 530008
rect 185515 529974 185532 530008
rect 184463 529963 185532 529974
rect 185567 530008 186636 530050
rect 185567 529974 185585 530008
rect 185619 529974 186585 530008
rect 186619 529974 186636 530008
rect 185567 529963 186636 529974
rect 186671 530008 187189 530050
rect 186671 529974 186689 530008
rect 186723 529974 187137 530008
rect 187171 529974 187189 530008
rect 183245 529924 183302 529948
rect 182713 529772 182824 529788
rect 182747 529738 182824 529772
rect 182713 529722 182824 529738
rect 182858 529772 183077 529846
rect 182858 529738 182909 529772
rect 182943 529738 183077 529772
rect 182858 529734 183077 529738
rect 182734 529700 182824 529722
rect 182071 529608 182089 529642
rect 182123 529608 182353 529642
rect 182387 529608 182405 529642
rect 182071 529540 182405 529608
rect 182531 529668 182589 529685
rect 182531 529634 182543 529668
rect 182577 529634 182589 529668
rect 182531 529540 182589 529634
rect 182623 529642 182700 529688
rect 182734 529666 182959 529700
rect 182623 529608 182660 529642
rect 182694 529608 182700 529642
rect 182903 529642 182959 529666
rect 182623 529574 182700 529608
rect 182734 529616 182799 529632
rect 182734 529582 182750 529616
rect 182784 529582 182799 529616
rect 182734 529540 182799 529582
rect 182903 529608 182909 529642
rect 182943 529608 182959 529642
rect 182903 529574 182959 529608
rect 182997 529642 183077 529734
rect 183111 529880 183302 529924
rect 183111 529772 183153 529880
rect 183111 529738 183113 529772
rect 183147 529738 183153 529772
rect 183111 529700 183153 529738
rect 183221 529812 183325 529846
rect 183187 529772 183325 529812
rect 183187 529738 183227 529772
rect 183261 529738 183325 529772
rect 183187 529734 183325 529738
rect 183676 529798 183744 529815
rect 183676 529764 183693 529798
rect 183727 529764 183744 529798
rect 183111 529666 183302 529700
rect 182997 529608 183013 529642
rect 183047 529608 183077 529642
rect 183245 529642 183302 529666
rect 183676 529649 183744 529764
rect 184040 529762 184110 529963
rect 184040 529728 184057 529762
rect 184091 529728 184110 529762
rect 184040 529713 184110 529728
rect 184780 529798 184848 529815
rect 184780 529764 184797 529798
rect 184831 529764 184848 529798
rect 184780 529649 184848 529764
rect 185144 529762 185214 529963
rect 185144 529728 185161 529762
rect 185195 529728 185214 529762
rect 185144 529713 185214 529728
rect 185884 529798 185952 529815
rect 185884 529764 185901 529798
rect 185935 529764 185952 529798
rect 185884 529649 185952 529764
rect 186248 529762 186318 529963
rect 186671 529906 187189 529974
rect 186671 529872 186689 529906
rect 186723 529872 187137 529906
rect 187171 529872 187189 529906
rect 186671 529832 187189 529872
rect 186248 529728 186265 529762
rect 186299 529728 186318 529762
rect 186248 529713 186318 529728
rect 186671 529764 186749 529798
rect 186783 529764 186859 529798
rect 186893 529764 186913 529798
rect 186671 529694 186913 529764
rect 186947 529762 187189 529832
rect 186947 529728 186967 529762
rect 187001 529728 187077 529762
rect 187111 529728 187189 529762
rect 187223 530008 187465 530050
rect 187223 529974 187241 530008
rect 187275 529974 187413 530008
rect 187447 529974 187465 530008
rect 187223 529913 187465 529974
rect 187223 529879 187241 529913
rect 187275 529879 187413 529913
rect 187447 529879 187465 529913
rect 187223 529832 187465 529879
rect 187223 529758 187327 529832
rect 187223 529724 187273 529758
rect 187307 529724 187327 529758
rect 187361 529764 187381 529798
rect 187415 529764 187465 529798
rect 182997 529574 183077 529608
rect 183157 529616 183211 529632
rect 183157 529582 183167 529616
rect 183201 529582 183211 529616
rect 183157 529540 183211 529582
rect 183245 529608 183251 529642
rect 183285 529608 183302 529642
rect 183245 529574 183302 529608
rect 183359 529635 184428 529649
rect 183359 529601 183377 529635
rect 183411 529601 184377 529635
rect 184411 529601 184428 529635
rect 183359 529540 184428 529601
rect 184463 529635 185532 529649
rect 184463 529601 184481 529635
rect 184515 529601 185481 529635
rect 185515 529601 185532 529635
rect 184463 529540 185532 529601
rect 185567 529635 186636 529649
rect 185567 529601 185585 529635
rect 185619 529601 186585 529635
rect 186619 529601 186636 529635
rect 185567 529540 186636 529601
rect 186671 529635 187189 529694
rect 187361 529690 187465 529764
rect 186671 529601 186689 529635
rect 186723 529601 187137 529635
rect 187171 529601 187189 529635
rect 186671 529540 187189 529601
rect 187223 529637 187465 529690
rect 187223 529603 187241 529637
rect 187275 529603 187413 529637
rect 187447 529603 187465 529637
rect 187223 529540 187465 529603
rect 172210 529506 172239 529540
rect 172273 529506 172331 529540
rect 172365 529506 172423 529540
rect 172457 529506 172515 529540
rect 172549 529506 172607 529540
rect 172641 529506 172699 529540
rect 172733 529506 172791 529540
rect 172825 529506 172883 529540
rect 172917 529506 172975 529540
rect 173009 529506 173067 529540
rect 173101 529506 173159 529540
rect 173193 529506 173251 529540
rect 173285 529506 173343 529540
rect 173377 529506 173435 529540
rect 173469 529506 173527 529540
rect 173561 529506 173619 529540
rect 173653 529506 173711 529540
rect 173745 529506 173803 529540
rect 173837 529506 173895 529540
rect 173929 529506 173987 529540
rect 174021 529506 174079 529540
rect 174113 529506 174171 529540
rect 174205 529506 174263 529540
rect 174297 529506 174355 529540
rect 174389 529506 174447 529540
rect 174481 529506 174539 529540
rect 174573 529506 174631 529540
rect 174665 529506 174723 529540
rect 174757 529506 174815 529540
rect 174849 529506 174907 529540
rect 174941 529506 174999 529540
rect 175033 529506 175091 529540
rect 175125 529506 175183 529540
rect 175217 529506 175275 529540
rect 175309 529506 175367 529540
rect 175401 529506 175459 529540
rect 175493 529506 175551 529540
rect 175585 529506 175643 529540
rect 175677 529506 175735 529540
rect 175769 529506 175827 529540
rect 175861 529506 175919 529540
rect 175953 529506 176011 529540
rect 176045 529506 176103 529540
rect 176137 529506 176195 529540
rect 176229 529506 176287 529540
rect 176321 529506 176379 529540
rect 176413 529506 176471 529540
rect 176505 529506 176563 529540
rect 176597 529506 176655 529540
rect 176689 529506 176747 529540
rect 176781 529506 176839 529540
rect 176873 529506 176931 529540
rect 176965 529506 177023 529540
rect 177057 529506 177115 529540
rect 177149 529506 177207 529540
rect 177241 529506 177299 529540
rect 177333 529506 177391 529540
rect 177425 529506 177483 529540
rect 177517 529506 177575 529540
rect 177609 529506 177667 529540
rect 177701 529506 177759 529540
rect 177793 529506 177851 529540
rect 177885 529506 177943 529540
rect 177977 529506 178035 529540
rect 178069 529506 178127 529540
rect 178161 529506 178219 529540
rect 178253 529506 178311 529540
rect 178345 529506 178403 529540
rect 178437 529506 178495 529540
rect 178529 529506 178587 529540
rect 178621 529506 178679 529540
rect 178713 529506 178771 529540
rect 178805 529506 178863 529540
rect 178897 529506 178955 529540
rect 178989 529506 179047 529540
rect 179081 529506 179139 529540
rect 179173 529506 179231 529540
rect 179265 529506 179323 529540
rect 179357 529506 179415 529540
rect 179449 529506 179507 529540
rect 179541 529506 179599 529540
rect 179633 529506 179691 529540
rect 179725 529506 179783 529540
rect 179817 529506 179875 529540
rect 179909 529506 179967 529540
rect 180001 529506 180059 529540
rect 180093 529506 180151 529540
rect 180185 529506 180243 529540
rect 180277 529506 180335 529540
rect 180369 529506 180427 529540
rect 180461 529506 180519 529540
rect 180553 529506 180611 529540
rect 180645 529506 180703 529540
rect 180737 529506 180795 529540
rect 180829 529506 180887 529540
rect 180921 529506 180979 529540
rect 181013 529506 181071 529540
rect 181105 529506 181163 529540
rect 181197 529506 181255 529540
rect 181289 529506 181347 529540
rect 181381 529506 181439 529540
rect 181473 529506 181531 529540
rect 181565 529506 181623 529540
rect 181657 529506 181715 529540
rect 181749 529506 181807 529540
rect 181841 529506 181899 529540
rect 181933 529506 181991 529540
rect 182025 529506 182083 529540
rect 182117 529506 182175 529540
rect 182209 529506 182267 529540
rect 182301 529506 182359 529540
rect 182393 529506 182451 529540
rect 182485 529506 182543 529540
rect 182577 529506 182635 529540
rect 182669 529506 182727 529540
rect 182761 529506 182819 529540
rect 182853 529506 182911 529540
rect 182945 529506 183003 529540
rect 183037 529506 183095 529540
rect 183129 529506 183187 529540
rect 183221 529506 183279 529540
rect 183313 529506 183371 529540
rect 183405 529506 183463 529540
rect 183497 529506 183555 529540
rect 183589 529506 183647 529540
rect 183681 529506 183739 529540
rect 183773 529506 183831 529540
rect 183865 529506 183923 529540
rect 183957 529506 184015 529540
rect 184049 529506 184107 529540
rect 184141 529506 184199 529540
rect 184233 529506 184291 529540
rect 184325 529506 184383 529540
rect 184417 529506 184475 529540
rect 184509 529506 184567 529540
rect 184601 529506 184659 529540
rect 184693 529506 184751 529540
rect 184785 529506 184843 529540
rect 184877 529506 184935 529540
rect 184969 529506 185027 529540
rect 185061 529506 185119 529540
rect 185153 529506 185211 529540
rect 185245 529506 185303 529540
rect 185337 529506 185395 529540
rect 185429 529506 185487 529540
rect 185521 529506 185579 529540
rect 185613 529506 185671 529540
rect 185705 529506 185763 529540
rect 185797 529506 185855 529540
rect 185889 529506 185947 529540
rect 185981 529506 186039 529540
rect 186073 529506 186131 529540
rect 186165 529506 186223 529540
rect 186257 529506 186315 529540
rect 186349 529506 186407 529540
rect 186441 529506 186499 529540
rect 186533 529506 186591 529540
rect 186625 529506 186683 529540
rect 186717 529506 186775 529540
rect 186809 529506 186867 529540
rect 186901 529506 186959 529540
rect 186993 529506 187051 529540
rect 187085 529506 187143 529540
rect 187177 529506 187235 529540
rect 187269 529506 187327 529540
rect 187361 529506 187419 529540
rect 187453 529506 187482 529540
rect 172227 529443 172469 529506
rect 172227 529409 172245 529443
rect 172279 529409 172417 529443
rect 172451 529409 172469 529443
rect 172227 529356 172469 529409
rect 172503 529445 173572 529506
rect 172503 529411 172521 529445
rect 172555 529411 173521 529445
rect 173555 529411 173572 529445
rect 172503 529397 173572 529411
rect 173607 529445 174676 529506
rect 173607 529411 173625 529445
rect 173659 529411 174625 529445
rect 174659 529411 174676 529445
rect 173607 529397 174676 529411
rect 174803 529412 174861 529506
rect 172227 529282 172331 529356
rect 172227 529248 172277 529282
rect 172311 529248 172331 529282
rect 172365 529288 172385 529322
rect 172419 529288 172469 529322
rect 172365 529214 172469 529288
rect 172820 529282 172888 529397
rect 172820 529248 172837 529282
rect 172871 529248 172888 529282
rect 172820 529231 172888 529248
rect 173184 529318 173254 529333
rect 173184 529284 173201 529318
rect 173235 529284 173254 529318
rect 172227 529167 172469 529214
rect 172227 529133 172245 529167
rect 172279 529133 172417 529167
rect 172451 529133 172469 529167
rect 172227 529072 172469 529133
rect 173184 529083 173254 529284
rect 173924 529282 173992 529397
rect 174803 529378 174815 529412
rect 174849 529378 174861 529412
rect 174803 529361 174861 529378
rect 175134 529449 175183 529465
rect 175134 529415 175143 529449
rect 175177 529415 175183 529449
rect 175134 529344 175183 529415
rect 175227 529449 175329 529506
rect 175261 529415 175295 529449
rect 175227 529399 175329 529415
rect 175365 529438 175403 529472
rect 175365 529404 175367 529438
rect 175401 529404 175403 529438
rect 173924 529248 173941 529282
rect 173975 529248 173992 529282
rect 173924 529231 173992 529248
rect 174288 529318 174358 529333
rect 174288 529284 174305 529318
rect 174339 529284 174358 529318
rect 174288 529083 174358 529284
rect 175079 529310 175275 529344
rect 175309 529310 175325 529344
rect 174803 529194 174861 529229
rect 174803 529160 174815 529194
rect 174849 529160 174861 529194
rect 174803 529101 174861 529160
rect 172227 529038 172245 529072
rect 172279 529038 172417 529072
rect 172451 529038 172469 529072
rect 172227 528996 172469 529038
rect 172503 529072 173572 529083
rect 172503 529038 172521 529072
rect 172555 529038 173521 529072
rect 173555 529038 173572 529072
rect 172503 528996 173572 529038
rect 173607 529072 174676 529083
rect 173607 529038 173625 529072
rect 173659 529038 174625 529072
rect 174659 529038 174676 529072
rect 173607 528996 174676 529038
rect 174803 529067 174815 529101
rect 174849 529067 174861 529101
rect 174803 528996 174861 529067
rect 175079 529148 175147 529310
rect 175181 529234 175331 529235
rect 175181 529231 175275 529234
rect 175181 529197 175197 529231
rect 175231 529200 175275 529231
rect 175309 529200 175331 529234
rect 175231 529197 175331 529200
rect 175079 529132 175182 529148
rect 175079 529098 175143 529132
rect 175177 529098 175182 529132
rect 175079 529066 175182 529098
rect 175229 529132 175263 529148
rect 175229 528996 175263 529098
rect 175297 529064 175331 529197
rect 175365 529231 175403 529404
rect 175437 529344 175492 529472
rect 175530 529449 175636 529472
rect 175564 529415 175636 529449
rect 175721 529464 175787 529506
rect 175721 529430 175737 529464
rect 175771 529430 175787 529464
rect 175721 529426 175787 529430
rect 175821 529445 175872 529472
rect 175530 529399 175636 529415
rect 175601 529392 175636 529399
rect 175855 529411 175872 529445
rect 175471 529310 175492 529344
rect 175437 529302 175492 529310
rect 175533 529344 175567 529360
rect 175437 529268 175459 529302
rect 175437 529240 175492 529268
rect 175399 529200 175403 529231
rect 175533 529200 175567 529310
rect 175399 529197 175567 529200
rect 175365 529166 175567 529197
rect 175601 529358 175787 529392
rect 175821 529358 175872 529411
rect 175925 529460 175985 529506
rect 175925 529426 175942 529460
rect 175976 529426 175985 529460
rect 175925 529410 175985 529426
rect 176019 529451 176071 529467
rect 176019 529417 176028 529451
rect 176062 529417 176071 529451
rect 176019 529376 176071 529417
rect 176105 529460 176157 529506
rect 176105 529426 176114 529460
rect 176148 529426 176157 529460
rect 176105 529410 176157 529426
rect 176193 529451 176245 529467
rect 176193 529417 176200 529451
rect 176234 529417 176245 529451
rect 176193 529376 176245 529417
rect 176279 529460 176329 529506
rect 176279 529426 176286 529460
rect 176320 529426 176329 529460
rect 176279 529410 176329 529426
rect 176365 529451 176417 529467
rect 176365 529417 176372 529451
rect 176406 529417 176417 529451
rect 176365 529376 176417 529417
rect 176451 529460 176501 529506
rect 176451 529426 176458 529460
rect 176492 529426 176501 529460
rect 176451 529410 176501 529426
rect 176537 529451 176589 529467
rect 176537 529417 176544 529451
rect 176578 529417 176589 529451
rect 176537 529376 176589 529417
rect 176623 529460 176672 529506
rect 176623 529426 176629 529460
rect 176663 529426 176672 529460
rect 176623 529410 176672 529426
rect 176706 529451 176761 529467
rect 176706 529417 176715 529451
rect 176749 529417 176761 529451
rect 176706 529376 176761 529417
rect 176795 529460 176844 529506
rect 176795 529426 176801 529460
rect 176835 529426 176844 529460
rect 176795 529410 176844 529426
rect 176878 529451 176930 529467
rect 176878 529417 176887 529451
rect 176921 529417 176930 529451
rect 176878 529376 176930 529417
rect 176964 529460 177016 529506
rect 176964 529426 176973 529460
rect 177007 529426 177016 529460
rect 176964 529410 177016 529426
rect 177050 529451 177102 529467
rect 177050 529417 177059 529451
rect 177093 529417 177102 529451
rect 177050 529376 177102 529417
rect 177136 529460 177188 529506
rect 177136 529426 177145 529460
rect 177179 529426 177188 529460
rect 177136 529410 177188 529426
rect 177222 529451 177274 529467
rect 177222 529417 177231 529451
rect 177265 529417 177274 529451
rect 177222 529376 177274 529417
rect 177308 529451 177360 529506
rect 177308 529417 177317 529451
rect 177351 529417 177360 529451
rect 177308 529394 177360 529417
rect 177394 529451 177444 529470
rect 177394 529417 177403 529451
rect 177437 529417 177444 529451
rect 175601 529132 175635 529358
rect 175753 529324 175787 529358
rect 175410 529098 175426 529132
rect 175460 529098 175501 529132
rect 175535 529098 175635 529132
rect 175669 529308 175708 529324
rect 175669 529274 175674 529308
rect 175669 529258 175708 529274
rect 175753 529308 175804 529324
rect 175753 529274 175770 529308
rect 175753 529258 175804 529274
rect 175669 529064 175703 529258
rect 175838 529224 175872 529358
rect 175297 529030 175703 529064
rect 175737 529208 175771 529224
rect 175737 529140 175771 529174
rect 175737 529072 175771 529106
rect 175737 528996 175771 529038
rect 175805 529208 175872 529224
rect 175805 529174 175821 529208
rect 175855 529174 175872 529208
rect 175925 529342 177274 529376
rect 175925 529224 176158 529342
rect 177394 529308 177444 529417
rect 177480 529451 177532 529506
rect 177480 529417 177489 529451
rect 177523 529417 177532 529451
rect 177480 529401 177532 529417
rect 177566 529451 177616 529470
rect 177566 529417 177575 529451
rect 177609 529417 177616 529451
rect 177566 529308 177616 529417
rect 177652 529464 177713 529506
rect 177652 529430 177661 529464
rect 177695 529430 177713 529464
rect 177833 529464 177899 529506
rect 177652 529404 177713 529430
rect 177748 529438 177799 529454
rect 177748 529404 177765 529438
rect 177833 529430 177849 529464
rect 177883 529430 177899 529464
rect 178039 529468 178105 529506
rect 177933 529438 177967 529454
rect 177748 529396 177799 529404
rect 178039 529434 178055 529468
rect 178089 529434 178105 529468
rect 178625 529464 178691 529506
rect 176192 529274 176212 529308
rect 176246 529274 176280 529308
rect 176314 529274 176348 529308
rect 176382 529274 176416 529308
rect 176450 529274 176484 529308
rect 176518 529274 176552 529308
rect 176586 529274 176620 529308
rect 176654 529274 176688 529308
rect 176722 529274 176756 529308
rect 176790 529274 176824 529308
rect 176858 529274 176892 529308
rect 176926 529274 176960 529308
rect 176994 529274 177028 529308
rect 177062 529274 177096 529308
rect 177130 529274 177164 529308
rect 177198 529274 177232 529308
rect 177266 529274 177616 529308
rect 176192 529258 177616 529274
rect 177650 529308 177713 529370
rect 177748 529362 177898 529396
rect 177650 529274 177659 529308
rect 177693 529302 177713 529308
rect 177650 529268 177667 529274
rect 177701 529268 177713 529302
rect 177650 529258 177713 529268
rect 177748 529308 177818 529328
rect 177748 529274 177762 529308
rect 177796 529274 177818 529308
rect 175925 529202 177274 529224
rect 175925 529179 176028 529202
rect 175805 529140 175872 529174
rect 176013 529168 176028 529179
rect 176062 529179 176200 529202
rect 176062 529168 176071 529179
rect 175805 529106 175821 529140
rect 175855 529106 175872 529140
rect 175805 529098 175872 529106
rect 175805 529072 175827 529098
rect 175805 529038 175821 529072
rect 175861 529064 175872 529098
rect 175855 529038 175872 529064
rect 175805 529030 175872 529038
rect 175925 529096 175979 529145
rect 175925 529062 175942 529096
rect 175976 529062 175979 529096
rect 175925 528996 175979 529062
rect 176013 529116 176071 529168
rect 176193 529168 176200 529179
rect 176234 529176 176372 529202
rect 176234 529168 176245 529176
rect 176013 529082 176028 529116
rect 176062 529082 176071 529116
rect 176013 529031 176071 529082
rect 176105 529096 176156 529142
rect 176105 529062 176114 529096
rect 176148 529062 176156 529096
rect 176105 528997 176156 529062
rect 176193 529116 176245 529168
rect 176365 529168 176372 529176
rect 176406 529176 176544 529202
rect 176406 529168 176417 529176
rect 176193 529098 176200 529116
rect 176193 529064 176195 529098
rect 176234 529082 176245 529116
rect 176229 529064 176245 529082
rect 176193 529031 176245 529064
rect 176279 529096 176328 529142
rect 176279 529062 176286 529096
rect 176320 529062 176328 529096
rect 176279 528997 176328 529062
rect 176365 529116 176417 529168
rect 176537 529168 176544 529176
rect 176578 529176 176715 529202
rect 176578 529168 176589 529176
rect 176365 529082 176372 529116
rect 176406 529082 176417 529116
rect 176365 529031 176417 529082
rect 176451 529096 176500 529142
rect 176451 529062 176458 529096
rect 176492 529062 176500 529096
rect 176451 528997 176500 529062
rect 176537 529116 176589 529168
rect 176706 529168 176715 529176
rect 176749 529176 176887 529202
rect 176749 529168 176758 529176
rect 176537 529082 176544 529116
rect 176578 529082 176589 529116
rect 176537 529031 176589 529082
rect 176623 529096 176672 529142
rect 176623 529062 176629 529096
rect 176663 529062 176672 529096
rect 176623 528997 176672 529062
rect 176706 529116 176758 529168
rect 176878 529168 176887 529176
rect 176921 529176 177059 529202
rect 176921 529168 176930 529176
rect 176706 529082 176715 529116
rect 176749 529082 176758 529116
rect 176706 529031 176758 529082
rect 176792 529096 176844 529142
rect 176792 529062 176801 529096
rect 176835 529062 176844 529096
rect 176792 528997 176844 529062
rect 176878 529116 176930 529168
rect 177050 529168 177059 529176
rect 177093 529176 177231 529202
rect 177093 529168 177102 529176
rect 176878 529082 176887 529116
rect 176921 529082 176930 529116
rect 176878 529031 176930 529082
rect 176964 529096 177016 529142
rect 176964 529062 176973 529096
rect 177007 529062 177016 529096
rect 176964 528997 177016 529062
rect 177050 529116 177102 529168
rect 177222 529168 177231 529176
rect 177265 529168 177274 529202
rect 177050 529082 177059 529116
rect 177093 529082 177102 529116
rect 177050 529031 177102 529082
rect 177136 529096 177188 529142
rect 177136 529062 177145 529096
rect 177179 529062 177188 529096
rect 177136 528997 177188 529062
rect 177222 529116 177274 529168
rect 177394 529156 177444 529258
rect 177222 529082 177231 529116
rect 177265 529082 177274 529116
rect 177222 529031 177274 529082
rect 177308 529140 177360 529156
rect 177308 529106 177317 529140
rect 177351 529106 177360 529140
rect 177308 529072 177360 529106
rect 177308 529038 177317 529072
rect 177351 529038 177360 529072
rect 177308 528997 177360 529038
rect 177394 529122 177403 529156
rect 177437 529122 177444 529156
rect 177394 529088 177444 529122
rect 177394 529054 177403 529088
rect 177437 529054 177444 529088
rect 177394 529031 177444 529054
rect 177480 529140 177532 529158
rect 177480 529106 177489 529140
rect 177523 529106 177532 529140
rect 177480 529072 177532 529106
rect 177480 529038 177489 529072
rect 177523 529038 177532 529072
rect 176105 528996 177360 528997
rect 177480 528996 177532 529038
rect 177567 529148 177616 529258
rect 177748 529234 177818 529274
rect 177748 529200 177759 529234
rect 177793 529200 177818 529234
rect 177748 529198 177818 529200
rect 177852 529302 177898 529362
rect 177886 529293 177898 529302
rect 177852 529259 177864 529268
rect 177852 529164 177898 529259
rect 177567 529114 177575 529148
rect 177609 529114 177616 529148
rect 177567 529080 177616 529114
rect 177567 529046 177575 529080
rect 177609 529046 177616 529080
rect 177567 529030 177616 529046
rect 177652 529140 177711 529158
rect 177652 529106 177661 529140
rect 177695 529106 177711 529140
rect 177652 529072 177711 529106
rect 177652 529038 177661 529072
rect 177695 529038 177711 529072
rect 177652 528996 177711 529038
rect 177748 529148 177898 529164
rect 177748 529114 177765 529148
rect 177799 529130 177898 529148
rect 177933 529166 177967 529404
rect 178139 529428 178188 529462
rect 178222 529428 178238 529462
rect 178279 529428 178295 529462
rect 178329 529428 178450 529462
rect 178013 529370 178105 529400
rect 178013 529336 178035 529370
rect 178069 529336 178105 529370
rect 178013 529247 178105 529336
rect 178013 529213 178071 529247
rect 178013 529190 178105 529213
rect 177748 529080 177799 529114
rect 177748 529046 177765 529080
rect 177748 529030 177799 529046
rect 177833 529062 177849 529096
rect 177883 529062 177899 529096
rect 177833 528996 177899 529062
rect 177933 529080 177967 529114
rect 177933 529030 177967 529046
rect 178001 529033 178066 529190
rect 178139 529156 178173 529428
rect 178207 529354 178277 529370
rect 178207 529320 178230 529354
rect 178264 529320 178277 529354
rect 178207 529302 178277 529320
rect 178207 529268 178219 529302
rect 178253 529268 178277 529302
rect 178207 529246 178277 529268
rect 178311 529360 178382 529370
rect 178311 529326 178332 529360
rect 178366 529326 178382 529360
rect 178311 529208 178345 529326
rect 178416 529286 178450 529428
rect 178625 529430 178641 529464
rect 178675 529430 178691 529464
rect 178625 529414 178691 529430
rect 178733 529434 178753 529468
rect 178787 529434 178803 529468
rect 178847 529464 179037 529472
rect 178525 529336 178563 529370
rect 178597 529354 178649 529370
rect 178733 529356 178785 529434
rect 178847 529430 178863 529464
rect 178897 529430 179037 529464
rect 178847 529416 179037 529430
rect 179071 529468 179109 529506
rect 179071 529434 179075 529468
rect 179406 529464 179467 529506
rect 179071 529418 179109 529434
rect 179143 529448 179357 529464
rect 179143 529430 179293 529448
rect 178491 529320 178587 529336
rect 178621 529320 178649 529354
rect 178683 529306 178717 529322
rect 178252 529192 178345 529208
rect 178286 529166 178345 529192
rect 178286 529158 178311 529166
rect 178139 529122 178218 529156
rect 178252 529132 178311 529158
rect 178252 529130 178345 529132
rect 178379 529272 178683 529286
rect 178379 529252 178717 529272
rect 178184 529096 178218 529122
rect 178379 529096 178413 529252
rect 178751 529218 178785 529356
rect 178485 529184 178501 529218
rect 178535 529184 178785 529218
rect 178823 529366 178865 529382
rect 178823 529332 178831 529366
rect 178823 529224 178865 529332
rect 178899 529318 178969 529382
rect 178899 529284 178927 529318
rect 178961 529302 178969 529318
rect 178899 529268 178935 529284
rect 178899 529258 178969 529268
rect 179003 529260 179037 529416
rect 179143 529384 179177 529430
rect 179327 529414 179357 529448
rect 179406 529430 179417 529464
rect 179451 529430 179467 529464
rect 179406 529414 179467 529430
rect 179501 529414 179552 529470
rect 179071 529350 179177 529384
rect 179211 529370 179259 529396
rect 179071 529344 179115 529350
rect 179105 529310 179115 529344
rect 179245 529336 179259 529370
rect 179211 529316 179259 529336
rect 179071 529294 179115 529310
rect 179151 529307 179167 529316
rect 179201 529282 179259 529316
rect 179185 529273 179259 529282
rect 179003 529226 179084 529260
rect 179151 529242 179259 529273
rect 179293 529359 179357 529414
rect 179535 529380 179552 529414
rect 179501 529364 179552 529380
rect 179293 529324 179358 529359
rect 179293 529308 179476 529324
rect 179293 529274 179442 529308
rect 179293 529264 179476 529274
rect 179328 529258 179476 529264
rect 178823 529192 178958 529224
rect 179050 529208 179084 529226
rect 178823 529190 178966 529192
rect 178751 529156 178785 529184
rect 178924 529166 178966 529190
rect 178100 529072 178150 529088
rect 178100 529038 178116 529072
rect 178100 528996 178150 529038
rect 178184 529080 178234 529096
rect 178184 529046 178200 529080
rect 178184 529030 178234 529046
rect 178277 529074 178413 529096
rect 178277 529040 178293 529074
rect 178327 529040 178413 529074
rect 178447 529116 178662 529150
rect 178751 529122 178863 529156
rect 178924 529132 178935 529166
rect 179000 529158 179016 529192
rect 178969 529132 179016 529158
rect 179050 529174 179244 529208
rect 179278 529174 179294 529208
rect 178447 529098 178481 529116
rect 178628 529098 178662 529116
rect 178447 529048 178481 529064
rect 178528 529048 178544 529082
rect 178578 529048 178594 529082
rect 178628 529048 178662 529064
rect 178721 529072 178795 529088
rect 178277 529030 178413 529040
rect 178528 528996 178594 529048
rect 178721 529038 178741 529072
rect 178775 529038 178795 529072
rect 178721 528996 178795 529038
rect 178829 529080 178863 529122
rect 179050 529098 179084 529174
rect 179328 529140 179362 529258
rect 179510 529234 179552 529364
rect 179697 529451 179731 529472
rect 179767 529464 179833 529506
rect 179767 529430 179783 529464
rect 179817 529430 179833 529464
rect 179869 529438 179921 529472
rect 179869 529434 179875 529438
rect 179697 529396 179731 529417
rect 179909 529404 179921 529438
rect 179903 529400 179921 529404
rect 179697 529362 179830 529396
rect 179869 529371 179921 529400
rect 179683 529308 179749 529326
rect 179683 529302 179699 529308
rect 179683 529268 179691 529302
rect 179733 529274 179749 529308
rect 179725 529268 179749 529274
rect 179683 529252 179749 529268
rect 179796 529311 179830 529362
rect 179796 529295 179853 529311
rect 179796 529261 179819 529295
rect 178829 529030 178863 529046
rect 178910 529073 179084 529098
rect 179202 529106 179362 529140
rect 179406 529140 179467 529224
rect 179406 529106 179417 529140
rect 179451 529106 179467 529140
rect 179202 529098 179236 529106
rect 178910 529039 178926 529073
rect 178960 529039 179084 529073
rect 178910 529030 179084 529039
rect 179118 529072 179168 529088
rect 179152 529038 179168 529072
rect 179406 529072 179467 529106
rect 179202 529048 179236 529064
rect 179118 528996 179168 529038
rect 179272 529038 179288 529072
rect 179322 529038 179338 529072
rect 179272 528996 179338 529038
rect 179406 529038 179417 529072
rect 179451 529038 179467 529072
rect 179501 529176 179552 529234
rect 179796 529245 179853 529261
rect 179796 529216 179830 529245
rect 179535 529142 179552 529176
rect 179501 529108 179552 529142
rect 179535 529098 179552 529108
rect 179501 529064 179507 529074
rect 179541 529064 179552 529098
rect 179501 529058 179552 529064
rect 179697 529182 179830 529216
rect 179887 529211 179921 529371
rect 179955 529412 180013 529506
rect 179955 529378 179967 529412
rect 180001 529378 180013 529412
rect 179955 529361 180013 529378
rect 180047 529445 180565 529506
rect 180047 529411 180065 529445
rect 180099 529411 180513 529445
rect 180547 529411 180565 529445
rect 180047 529352 180565 529411
rect 180691 529464 180752 529506
rect 180691 529430 180709 529464
rect 180743 529430 180752 529464
rect 180691 529404 180752 529430
rect 180788 529451 180838 529470
rect 180788 529417 180795 529451
rect 180829 529417 180838 529451
rect 180047 529282 180289 529352
rect 180047 529248 180125 529282
rect 180159 529248 180235 529282
rect 180269 529248 180289 529282
rect 180323 529284 180343 529318
rect 180377 529284 180453 529318
rect 180487 529284 180565 529318
rect 179697 529148 179731 529182
rect 179867 529161 179921 529211
rect 179697 529080 179731 529114
rect 179406 528996 179467 529038
rect 179697 529030 179731 529046
rect 179767 529114 179783 529148
rect 179817 529114 179833 529148
rect 179767 529080 179833 529114
rect 179767 529046 179783 529080
rect 179817 529046 179833 529080
rect 179767 528996 179833 529046
rect 179867 529127 179869 529161
rect 179903 529127 179921 529161
rect 179867 529080 179921 529127
rect 179867 529046 179869 529080
rect 179903 529046 179921 529080
rect 179867 529030 179921 529046
rect 179955 529194 180013 529229
rect 180323 529214 180565 529284
rect 180691 529308 180754 529370
rect 180691 529302 180711 529308
rect 180691 529268 180703 529302
rect 180745 529274 180754 529308
rect 180737 529268 180754 529274
rect 180691 529258 180754 529268
rect 180788 529308 180838 529417
rect 180872 529451 180924 529506
rect 180872 529417 180881 529451
rect 180915 529417 180924 529451
rect 180872 529401 180924 529417
rect 180960 529451 181010 529470
rect 180960 529417 180967 529451
rect 181001 529417 181010 529451
rect 180960 529308 181010 529417
rect 181044 529451 181096 529506
rect 181044 529417 181053 529451
rect 181087 529417 181096 529451
rect 181044 529394 181096 529417
rect 181130 529451 181182 529467
rect 181130 529417 181139 529451
rect 181173 529417 181182 529451
rect 181130 529376 181182 529417
rect 181216 529460 181268 529506
rect 181216 529426 181225 529460
rect 181259 529426 181268 529460
rect 181216 529410 181268 529426
rect 181302 529451 181354 529467
rect 181302 529417 181311 529451
rect 181345 529417 181354 529451
rect 181302 529376 181354 529417
rect 181388 529460 181440 529506
rect 181388 529426 181397 529460
rect 181431 529426 181440 529460
rect 181388 529410 181440 529426
rect 181474 529451 181526 529467
rect 181474 529417 181483 529451
rect 181517 529417 181526 529451
rect 181474 529376 181526 529417
rect 181560 529460 181609 529506
rect 181560 529426 181569 529460
rect 181603 529426 181609 529460
rect 181560 529410 181609 529426
rect 181643 529451 181698 529467
rect 181643 529417 181655 529451
rect 181689 529417 181698 529451
rect 181643 529376 181698 529417
rect 181732 529460 181781 529506
rect 181732 529426 181741 529460
rect 181775 529426 181781 529460
rect 181732 529410 181781 529426
rect 181815 529451 181867 529467
rect 181815 529417 181826 529451
rect 181860 529417 181867 529451
rect 181815 529376 181867 529417
rect 181903 529460 181953 529506
rect 181903 529426 181912 529460
rect 181946 529426 181953 529460
rect 181903 529410 181953 529426
rect 181987 529451 182039 529467
rect 181987 529417 181998 529451
rect 182032 529417 182039 529451
rect 181987 529376 182039 529417
rect 182075 529460 182125 529506
rect 182075 529426 182084 529460
rect 182118 529426 182125 529460
rect 182075 529410 182125 529426
rect 182159 529451 182211 529467
rect 182159 529417 182170 529451
rect 182204 529417 182211 529451
rect 182159 529376 182211 529417
rect 182247 529460 182299 529506
rect 182247 529426 182256 529460
rect 182290 529426 182299 529460
rect 182247 529410 182299 529426
rect 182333 529451 182385 529467
rect 182333 529417 182342 529451
rect 182376 529417 182385 529451
rect 182333 529376 182385 529417
rect 182419 529460 182479 529506
rect 182419 529426 182428 529460
rect 182462 529426 182479 529460
rect 182419 529410 182479 529426
rect 182531 529438 182583 529472
rect 182531 529404 182543 529438
rect 182577 529434 182583 529438
rect 182619 529464 182685 529506
rect 182619 529430 182635 529464
rect 182669 529430 182685 529464
rect 182721 529451 182755 529472
rect 182531 529400 182549 529404
rect 181130 529342 182479 529376
rect 180788 529274 181138 529308
rect 181172 529274 181206 529308
rect 181240 529274 181274 529308
rect 181308 529274 181342 529308
rect 181376 529274 181410 529308
rect 181444 529274 181478 529308
rect 181512 529274 181546 529308
rect 181580 529274 181614 529308
rect 181648 529274 181682 529308
rect 181716 529274 181750 529308
rect 181784 529274 181818 529308
rect 181852 529274 181886 529308
rect 181920 529274 181954 529308
rect 181988 529274 182022 529308
rect 182056 529274 182090 529308
rect 182124 529274 182158 529308
rect 182192 529274 182212 529308
rect 180788 529258 182212 529274
rect 179955 529160 179967 529194
rect 180001 529160 180013 529194
rect 179955 529101 180013 529160
rect 179955 529067 179967 529101
rect 180001 529067 180013 529101
rect 179955 528996 180013 529067
rect 180047 529174 180565 529214
rect 180047 529140 180065 529174
rect 180099 529140 180513 529174
rect 180547 529140 180565 529174
rect 180047 529072 180565 529140
rect 180047 529038 180065 529072
rect 180099 529038 180513 529072
rect 180547 529038 180565 529072
rect 180047 528996 180565 529038
rect 180693 529140 180752 529158
rect 180693 529106 180709 529140
rect 180743 529106 180752 529140
rect 180693 529072 180752 529106
rect 180693 529038 180709 529072
rect 180743 529038 180752 529072
rect 180693 528996 180752 529038
rect 180788 529148 180837 529258
rect 180788 529114 180795 529148
rect 180829 529114 180837 529148
rect 180788 529080 180837 529114
rect 180788 529046 180795 529080
rect 180829 529046 180837 529080
rect 180788 529030 180837 529046
rect 180872 529140 180924 529158
rect 180872 529106 180881 529140
rect 180915 529106 180924 529140
rect 180872 529072 180924 529106
rect 180872 529038 180881 529072
rect 180915 529038 180924 529072
rect 180872 528996 180924 529038
rect 180960 529156 181010 529258
rect 182246 529224 182479 529342
rect 181130 529202 182479 529224
rect 181130 529168 181139 529202
rect 181173 529176 181311 529202
rect 181173 529168 181182 529176
rect 180960 529122 180967 529156
rect 181001 529122 181010 529156
rect 180960 529088 181010 529122
rect 180960 529054 180967 529088
rect 181001 529054 181010 529088
rect 180960 529031 181010 529054
rect 181044 529140 181096 529156
rect 181044 529106 181053 529140
rect 181087 529106 181096 529140
rect 181044 529072 181096 529106
rect 181044 529038 181053 529072
rect 181087 529038 181096 529072
rect 181044 528997 181096 529038
rect 181130 529116 181182 529168
rect 181302 529168 181311 529176
rect 181345 529176 181483 529202
rect 181345 529168 181354 529176
rect 181130 529082 181139 529116
rect 181173 529082 181182 529116
rect 181130 529031 181182 529082
rect 181216 529096 181268 529142
rect 181216 529062 181225 529096
rect 181259 529062 181268 529096
rect 181216 528997 181268 529062
rect 181302 529116 181354 529168
rect 181474 529168 181483 529176
rect 181517 529176 181655 529202
rect 181517 529168 181526 529176
rect 181302 529082 181311 529116
rect 181345 529082 181354 529116
rect 181302 529031 181354 529082
rect 181388 529096 181440 529142
rect 181388 529062 181397 529096
rect 181431 529062 181440 529096
rect 181388 528997 181440 529062
rect 181474 529116 181526 529168
rect 181646 529168 181655 529176
rect 181689 529176 181826 529202
rect 181689 529168 181698 529176
rect 181474 529082 181483 529116
rect 181517 529082 181526 529116
rect 181474 529031 181526 529082
rect 181560 529096 181612 529142
rect 181560 529062 181569 529096
rect 181603 529062 181612 529096
rect 181560 528997 181612 529062
rect 181646 529116 181698 529168
rect 181815 529168 181826 529176
rect 181860 529176 181998 529202
rect 181860 529168 181867 529176
rect 181646 529082 181655 529116
rect 181689 529082 181698 529116
rect 181646 529031 181698 529082
rect 181732 529096 181781 529142
rect 181732 529062 181741 529096
rect 181775 529062 181781 529096
rect 181732 528997 181781 529062
rect 181815 529116 181867 529168
rect 181987 529168 181998 529176
rect 182032 529176 182170 529202
rect 182032 529168 182039 529176
rect 181815 529082 181826 529116
rect 181860 529082 181867 529116
rect 181815 529031 181867 529082
rect 181904 529096 181953 529142
rect 181904 529062 181912 529096
rect 181946 529062 181953 529096
rect 181904 528997 181953 529062
rect 181987 529116 182039 529168
rect 182159 529168 182170 529176
rect 182204 529179 182342 529202
rect 182204 529168 182211 529179
rect 181987 529098 181998 529116
rect 181987 529064 181991 529098
rect 182032 529082 182039 529116
rect 182025 529064 182039 529082
rect 181987 529031 182039 529064
rect 182076 529096 182125 529142
rect 182076 529062 182084 529096
rect 182118 529062 182125 529096
rect 182076 528997 182125 529062
rect 182159 529116 182211 529168
rect 182333 529168 182342 529179
rect 182376 529179 182479 529202
rect 182531 529371 182583 529400
rect 182721 529396 182755 529417
rect 182807 529445 183876 529506
rect 182807 529411 182825 529445
rect 182859 529411 183825 529445
rect 183859 529411 183876 529445
rect 182807 529397 183876 529411
rect 183911 529445 184980 529506
rect 183911 529411 183929 529445
rect 183963 529411 184929 529445
rect 184963 529411 184980 529445
rect 183911 529397 184980 529411
rect 185107 529412 185165 529506
rect 182531 529211 182565 529371
rect 182622 529362 182755 529396
rect 182622 529311 182656 529362
rect 182599 529295 182656 529311
rect 182633 529261 182656 529295
rect 182599 529245 182656 529261
rect 182703 529308 182769 529326
rect 182703 529274 182719 529308
rect 182753 529302 182769 529308
rect 182703 529268 182727 529274
rect 182761 529268 182769 529302
rect 182703 529252 182769 529268
rect 183124 529282 183192 529397
rect 182622 529216 182656 529245
rect 183124 529248 183141 529282
rect 183175 529248 183192 529282
rect 183124 529231 183192 529248
rect 183488 529318 183558 529333
rect 183488 529284 183505 529318
rect 183539 529284 183558 529318
rect 182376 529168 182391 529179
rect 182159 529082 182170 529116
rect 182204 529082 182211 529116
rect 182159 529031 182211 529082
rect 182248 529096 182299 529142
rect 182248 529062 182256 529096
rect 182290 529062 182299 529096
rect 182248 528997 182299 529062
rect 182333 529116 182391 529168
rect 182531 529161 182585 529211
rect 182622 529182 182755 529216
rect 182333 529082 182342 529116
rect 182376 529082 182391 529116
rect 182333 529031 182391 529082
rect 182425 529096 182479 529145
rect 182425 529062 182428 529096
rect 182462 529062 182479 529096
rect 181044 528996 182299 528997
rect 182425 528996 182479 529062
rect 182531 529127 182549 529161
rect 182583 529127 182585 529161
rect 182721 529148 182755 529182
rect 182531 529080 182585 529127
rect 182531 529046 182549 529080
rect 182583 529046 182585 529080
rect 182531 529030 182585 529046
rect 182619 529114 182635 529148
rect 182669 529114 182685 529148
rect 182619 529080 182685 529114
rect 182619 529046 182635 529080
rect 182669 529046 182685 529080
rect 182619 528996 182685 529046
rect 182721 529080 182755 529114
rect 183488 529083 183558 529284
rect 184228 529282 184296 529397
rect 185107 529378 185119 529412
rect 185153 529378 185165 529412
rect 185199 529445 186268 529506
rect 185199 529411 185217 529445
rect 185251 529411 186217 529445
rect 186251 529411 186268 529445
rect 185199 529397 186268 529411
rect 186303 529445 187005 529506
rect 186303 529411 186321 529445
rect 186355 529411 186953 529445
rect 186987 529411 187005 529445
rect 185107 529361 185165 529378
rect 184228 529248 184245 529282
rect 184279 529248 184296 529282
rect 184228 529231 184296 529248
rect 184592 529318 184662 529333
rect 184592 529284 184609 529318
rect 184643 529284 184662 529318
rect 184592 529083 184662 529284
rect 185516 529282 185584 529397
rect 186303 529352 187005 529411
rect 187223 529443 187465 529506
rect 187223 529409 187241 529443
rect 187275 529409 187413 529443
rect 187447 529409 187465 529443
rect 187223 529356 187465 529409
rect 185516 529248 185533 529282
rect 185567 529248 185584 529282
rect 185516 529231 185584 529248
rect 185880 529318 185950 529333
rect 185880 529284 185897 529318
rect 185931 529284 185950 529318
rect 185107 529194 185165 529229
rect 185107 529160 185119 529194
rect 185153 529160 185165 529194
rect 185107 529101 185165 529160
rect 182721 529030 182755 529046
rect 182807 529072 183876 529083
rect 182807 529038 182825 529072
rect 182859 529038 183825 529072
rect 183859 529038 183876 529072
rect 182807 528996 183876 529038
rect 183911 529072 184980 529083
rect 183911 529038 183929 529072
rect 183963 529038 184929 529072
rect 184963 529038 184980 529072
rect 183911 528996 184980 529038
rect 185107 529067 185119 529101
rect 185153 529067 185165 529101
rect 185880 529083 185950 529284
rect 186303 529282 186633 529352
rect 186303 529248 186381 529282
rect 186415 529248 186480 529282
rect 186514 529248 186579 529282
rect 186613 529248 186633 529282
rect 186667 529284 186687 529318
rect 186721 529284 186790 529318
rect 186824 529284 186893 529318
rect 186927 529284 187005 529318
rect 186667 529214 187005 529284
rect 186303 529174 187005 529214
rect 186303 529140 186321 529174
rect 186355 529140 186953 529174
rect 186987 529140 187005 529174
rect 185107 528996 185165 529067
rect 185199 529072 186268 529083
rect 185199 529038 185217 529072
rect 185251 529038 186217 529072
rect 186251 529038 186268 529072
rect 185199 528996 186268 529038
rect 186303 529072 187005 529140
rect 186303 529038 186321 529072
rect 186355 529038 186953 529072
rect 186987 529038 187005 529072
rect 186303 528996 187005 529038
rect 187223 529288 187273 529322
rect 187307 529288 187327 529322
rect 187223 529214 187327 529288
rect 187361 529282 187465 529356
rect 187361 529248 187381 529282
rect 187415 529248 187465 529282
rect 187223 529167 187465 529214
rect 187223 529133 187241 529167
rect 187275 529133 187413 529167
rect 187447 529133 187465 529167
rect 187223 529072 187465 529133
rect 187223 529038 187241 529072
rect 187275 529038 187413 529072
rect 187447 529038 187465 529072
rect 187223 528996 187465 529038
rect 172210 528962 172239 528996
rect 172273 528962 172331 528996
rect 172365 528962 172423 528996
rect 172457 528962 172515 528996
rect 172549 528962 172607 528996
rect 172641 528962 172699 528996
rect 172733 528962 172791 528996
rect 172825 528962 172883 528996
rect 172917 528962 172975 528996
rect 173009 528962 173067 528996
rect 173101 528962 173159 528996
rect 173193 528962 173251 528996
rect 173285 528962 173343 528996
rect 173377 528962 173435 528996
rect 173469 528962 173527 528996
rect 173561 528962 173619 528996
rect 173653 528962 173711 528996
rect 173745 528962 173803 528996
rect 173837 528962 173895 528996
rect 173929 528962 173987 528996
rect 174021 528962 174079 528996
rect 174113 528962 174171 528996
rect 174205 528962 174263 528996
rect 174297 528962 174355 528996
rect 174389 528962 174447 528996
rect 174481 528962 174539 528996
rect 174573 528962 174631 528996
rect 174665 528962 174723 528996
rect 174757 528962 174815 528996
rect 174849 528962 174907 528996
rect 174941 528962 174999 528996
rect 175033 528962 175091 528996
rect 175125 528962 175183 528996
rect 175217 528962 175275 528996
rect 175309 528962 175367 528996
rect 175401 528962 175459 528996
rect 175493 528962 175551 528996
rect 175585 528962 175643 528996
rect 175677 528962 175735 528996
rect 175769 528962 175827 528996
rect 175861 528962 175919 528996
rect 175953 528962 176011 528996
rect 176045 528962 176103 528996
rect 176137 528962 176195 528996
rect 176229 528962 176287 528996
rect 176321 528962 176379 528996
rect 176413 528962 176471 528996
rect 176505 528962 176563 528996
rect 176597 528962 176655 528996
rect 176689 528962 176747 528996
rect 176781 528962 176839 528996
rect 176873 528962 176931 528996
rect 176965 528962 177023 528996
rect 177057 528962 177115 528996
rect 177149 528962 177207 528996
rect 177241 528962 177299 528996
rect 177333 528962 177391 528996
rect 177425 528962 177483 528996
rect 177517 528962 177575 528996
rect 177609 528962 177667 528996
rect 177701 528962 177759 528996
rect 177793 528962 177851 528996
rect 177885 528962 177943 528996
rect 177977 528962 178035 528996
rect 178069 528962 178127 528996
rect 178161 528962 178219 528996
rect 178253 528962 178311 528996
rect 178345 528962 178403 528996
rect 178437 528962 178495 528996
rect 178529 528962 178587 528996
rect 178621 528962 178679 528996
rect 178713 528962 178771 528996
rect 178805 528962 178863 528996
rect 178897 528962 178955 528996
rect 178989 528962 179047 528996
rect 179081 528962 179139 528996
rect 179173 528962 179231 528996
rect 179265 528962 179323 528996
rect 179357 528962 179415 528996
rect 179449 528962 179507 528996
rect 179541 528962 179599 528996
rect 179633 528962 179691 528996
rect 179725 528962 179783 528996
rect 179817 528962 179875 528996
rect 179909 528962 179967 528996
rect 180001 528962 180059 528996
rect 180093 528962 180151 528996
rect 180185 528962 180243 528996
rect 180277 528962 180335 528996
rect 180369 528962 180427 528996
rect 180461 528962 180519 528996
rect 180553 528962 180611 528996
rect 180645 528962 180703 528996
rect 180737 528962 180795 528996
rect 180829 528962 180887 528996
rect 180921 528962 180979 528996
rect 181013 528962 181071 528996
rect 181105 528962 181163 528996
rect 181197 528962 181255 528996
rect 181289 528962 181347 528996
rect 181381 528962 181439 528996
rect 181473 528962 181531 528996
rect 181565 528962 181623 528996
rect 181657 528962 181715 528996
rect 181749 528962 181807 528996
rect 181841 528962 181899 528996
rect 181933 528962 181991 528996
rect 182025 528962 182083 528996
rect 182117 528962 182175 528996
rect 182209 528962 182267 528996
rect 182301 528962 182359 528996
rect 182393 528962 182451 528996
rect 182485 528962 182543 528996
rect 182577 528962 182635 528996
rect 182669 528962 182727 528996
rect 182761 528962 182819 528996
rect 182853 528962 182911 528996
rect 182945 528962 183003 528996
rect 183037 528962 183095 528996
rect 183129 528962 183187 528996
rect 183221 528962 183279 528996
rect 183313 528962 183371 528996
rect 183405 528962 183463 528996
rect 183497 528962 183555 528996
rect 183589 528962 183647 528996
rect 183681 528962 183739 528996
rect 183773 528962 183831 528996
rect 183865 528962 183923 528996
rect 183957 528962 184015 528996
rect 184049 528962 184107 528996
rect 184141 528962 184199 528996
rect 184233 528962 184291 528996
rect 184325 528962 184383 528996
rect 184417 528962 184475 528996
rect 184509 528962 184567 528996
rect 184601 528962 184659 528996
rect 184693 528962 184751 528996
rect 184785 528962 184843 528996
rect 184877 528962 184935 528996
rect 184969 528962 185027 528996
rect 185061 528962 185119 528996
rect 185153 528962 185211 528996
rect 185245 528962 185303 528996
rect 185337 528962 185395 528996
rect 185429 528962 185487 528996
rect 185521 528962 185579 528996
rect 185613 528962 185671 528996
rect 185705 528962 185763 528996
rect 185797 528962 185855 528996
rect 185889 528962 185947 528996
rect 185981 528962 186039 528996
rect 186073 528962 186131 528996
rect 186165 528962 186223 528996
rect 186257 528962 186315 528996
rect 186349 528962 186407 528996
rect 186441 528962 186499 528996
rect 186533 528962 186591 528996
rect 186625 528962 186683 528996
rect 186717 528962 186775 528996
rect 186809 528962 186867 528996
rect 186901 528962 186959 528996
rect 186993 528962 187051 528996
rect 187085 528962 187143 528996
rect 187177 528962 187235 528996
rect 187269 528962 187327 528996
rect 187361 528962 187419 528996
rect 187453 528962 187482 528996
rect 172227 528920 172469 528962
rect 172227 528886 172245 528920
rect 172279 528886 172417 528920
rect 172451 528886 172469 528920
rect 172227 528825 172469 528886
rect 172503 528920 173572 528962
rect 172503 528886 172521 528920
rect 172555 528886 173521 528920
rect 173555 528886 173572 528920
rect 172503 528875 173572 528886
rect 173607 528920 174676 528962
rect 173607 528886 173625 528920
rect 173659 528886 174625 528920
rect 174659 528886 174676 528920
rect 173607 528875 174676 528886
rect 174711 528920 175780 528962
rect 174711 528886 174729 528920
rect 174763 528886 175729 528920
rect 175763 528886 175780 528920
rect 174711 528875 175780 528886
rect 175925 528912 175959 528928
rect 172227 528791 172245 528825
rect 172279 528791 172417 528825
rect 172451 528791 172469 528825
rect 172227 528744 172469 528791
rect 172227 528676 172277 528710
rect 172311 528676 172331 528710
rect 172227 528602 172331 528676
rect 172365 528670 172469 528744
rect 172365 528636 172385 528670
rect 172419 528636 172469 528670
rect 172820 528710 172888 528727
rect 172820 528676 172837 528710
rect 172871 528676 172888 528710
rect 172227 528549 172469 528602
rect 172820 528561 172888 528676
rect 173184 528674 173254 528875
rect 173184 528640 173201 528674
rect 173235 528640 173254 528674
rect 173184 528625 173254 528640
rect 173924 528710 173992 528727
rect 173924 528676 173941 528710
rect 173975 528676 173992 528710
rect 173924 528561 173992 528676
rect 174288 528674 174358 528875
rect 174288 528640 174305 528674
rect 174339 528640 174358 528674
rect 174288 528625 174358 528640
rect 175028 528710 175096 528727
rect 175028 528676 175045 528710
rect 175079 528676 175096 528710
rect 175028 528561 175096 528676
rect 175392 528674 175462 528875
rect 175925 528844 175959 528878
rect 175995 528912 176061 528962
rect 175995 528878 176011 528912
rect 176045 528878 176061 528912
rect 175995 528844 176061 528878
rect 175995 528810 176011 528844
rect 176045 528810 176061 528844
rect 176095 528912 176149 528928
rect 176095 528878 176097 528912
rect 176131 528894 176149 528912
rect 176095 528860 176103 528878
rect 176137 528860 176149 528894
rect 176095 528831 176149 528860
rect 175925 528776 175959 528810
rect 176095 528797 176097 528831
rect 176131 528797 176149 528831
rect 175925 528742 176058 528776
rect 176095 528747 176149 528797
rect 176024 528713 176058 528742
rect 175392 528640 175409 528674
rect 175443 528640 175462 528674
rect 175392 528625 175462 528640
rect 175911 528690 175977 528706
rect 175911 528656 175919 528690
rect 175953 528684 175977 528690
rect 175911 528650 175927 528656
rect 175961 528650 175977 528684
rect 175911 528632 175977 528650
rect 176024 528697 176081 528713
rect 176024 528663 176047 528697
rect 176024 528647 176081 528663
rect 176024 528596 176058 528647
rect 175925 528562 176058 528596
rect 176115 528587 176149 528747
rect 176201 528912 176235 528928
rect 176201 528844 176235 528878
rect 176271 528912 176337 528962
rect 176271 528878 176287 528912
rect 176321 528878 176337 528912
rect 176271 528844 176337 528878
rect 176271 528810 176287 528844
rect 176321 528810 176337 528844
rect 176371 528912 176425 528928
rect 176371 528878 176373 528912
rect 176407 528878 176425 528912
rect 176371 528831 176425 528878
rect 176201 528776 176235 528810
rect 176371 528797 176373 528831
rect 176407 528797 176425 528831
rect 176201 528742 176334 528776
rect 176371 528747 176425 528797
rect 176300 528713 176334 528742
rect 176187 528690 176253 528706
rect 176187 528656 176195 528690
rect 176229 528684 176253 528690
rect 176187 528650 176203 528656
rect 176237 528650 176253 528684
rect 176187 528632 176253 528650
rect 176300 528697 176357 528713
rect 176300 528663 176323 528697
rect 176300 528647 176357 528663
rect 176300 528596 176334 528647
rect 172227 528515 172245 528549
rect 172279 528515 172417 528549
rect 172451 528515 172469 528549
rect 172227 528452 172469 528515
rect 172503 528547 173572 528561
rect 172503 528513 172521 528547
rect 172555 528513 173521 528547
rect 173555 528513 173572 528547
rect 172503 528452 173572 528513
rect 173607 528547 174676 528561
rect 173607 528513 173625 528547
rect 173659 528513 174625 528547
rect 174659 528513 174676 528547
rect 173607 528452 174676 528513
rect 174711 528547 175780 528561
rect 174711 528513 174729 528547
rect 174763 528513 175729 528547
rect 175763 528513 175780 528547
rect 174711 528452 175780 528513
rect 175925 528541 175959 528562
rect 176097 528558 176149 528587
rect 175925 528486 175959 528507
rect 175995 528494 176011 528528
rect 176045 528494 176061 528528
rect 175995 528452 176061 528494
rect 176131 528524 176149 528558
rect 176097 528486 176149 528524
rect 176201 528562 176334 528596
rect 176391 528587 176425 528747
rect 176459 528860 176562 528892
rect 176459 528826 176523 528860
rect 176557 528826 176562 528860
rect 176459 528810 176562 528826
rect 176609 528860 176643 528962
rect 176609 528810 176643 528826
rect 176677 528894 177083 528928
rect 176459 528648 176527 528810
rect 176677 528761 176711 528894
rect 176790 528826 176806 528860
rect 176840 528826 176881 528860
rect 176915 528826 177015 528860
rect 176561 528758 176577 528761
rect 176561 528724 176563 528758
rect 176611 528727 176711 528761
rect 176597 528724 176711 528727
rect 176561 528723 176711 528724
rect 176745 528761 176947 528792
rect 176779 528758 176947 528761
rect 176779 528727 176783 528758
rect 176459 528614 176655 528648
rect 176689 528614 176705 528648
rect 176201 528541 176235 528562
rect 176373 528558 176425 528587
rect 176407 528554 176425 528558
rect 176201 528486 176235 528507
rect 176271 528494 176287 528528
rect 176321 528494 176337 528528
rect 176271 528452 176337 528494
rect 176373 528520 176379 528524
rect 176413 528520 176425 528554
rect 176373 528486 176425 528520
rect 176514 528543 176563 528614
rect 176514 528509 176523 528543
rect 176557 528509 176563 528543
rect 176514 528493 176563 528509
rect 176607 528543 176709 528559
rect 176641 528509 176675 528543
rect 176607 528452 176709 528509
rect 176745 528554 176783 528727
rect 176745 528520 176747 528554
rect 176781 528520 176783 528554
rect 176745 528486 176783 528520
rect 176817 528690 176872 528718
rect 176817 528656 176839 528690
rect 176817 528648 176872 528656
rect 176851 528614 176872 528648
rect 176817 528486 176872 528614
rect 176913 528648 176947 528758
rect 176913 528598 176947 528614
rect 176981 528600 177015 528826
rect 177049 528700 177083 528894
rect 177117 528920 177151 528962
rect 177117 528852 177151 528886
rect 177117 528784 177151 528818
rect 177117 528734 177151 528750
rect 177185 528920 177252 528928
rect 177185 528886 177201 528920
rect 177235 528886 177252 528920
rect 177185 528852 177252 528886
rect 177185 528818 177201 528852
rect 177235 528818 177252 528852
rect 177185 528784 177252 528818
rect 177185 528750 177201 528784
rect 177235 528750 177252 528784
rect 177185 528734 177252 528750
rect 177049 528684 177088 528700
rect 177049 528650 177054 528684
rect 177049 528634 177088 528650
rect 177133 528684 177184 528700
rect 177133 528650 177150 528684
rect 177133 528634 177184 528650
rect 177133 528600 177167 528634
rect 177218 528600 177252 528734
rect 177379 528891 177437 528962
rect 177379 528857 177391 528891
rect 177425 528857 177437 528891
rect 177379 528798 177437 528857
rect 177379 528764 177391 528798
rect 177425 528764 177437 528798
rect 177379 528729 177437 528764
rect 177471 528894 177548 528928
rect 177471 528860 177508 528894
rect 177542 528860 177548 528894
rect 177582 528920 177647 528962
rect 177582 528886 177598 528920
rect 177632 528886 177647 528920
rect 177582 528870 177647 528886
rect 177751 528894 177807 528928
rect 177471 528734 177548 528860
rect 177751 528860 177757 528894
rect 177791 528860 177807 528894
rect 177751 528836 177807 528860
rect 177582 528792 177807 528836
rect 177845 528894 177925 528928
rect 177845 528860 177861 528894
rect 177895 528860 177925 528894
rect 178005 528920 178059 528962
rect 178005 528886 178015 528920
rect 178049 528886 178059 528920
rect 178005 528870 178059 528886
rect 178093 528894 178150 528928
rect 176981 528566 177167 528600
rect 176981 528559 177016 528566
rect 176910 528543 177016 528559
rect 176944 528509 177016 528543
rect 177201 528554 177252 528600
rect 177471 528690 177527 528734
rect 177582 528700 177672 528792
rect 177845 528758 177925 528860
rect 178093 528860 178099 528894
rect 178133 528860 178150 528894
rect 178093 528836 178150 528860
rect 177471 528656 177483 528690
rect 177517 528656 177527 528690
rect 177471 528600 177527 528656
rect 177561 528684 177672 528700
rect 177595 528650 177672 528684
rect 177561 528634 177672 528650
rect 177706 528684 177925 528758
rect 177706 528650 177757 528684
rect 177791 528650 177925 528684
rect 177706 528646 177925 528650
rect 177582 528612 177672 528634
rect 177201 528547 177207 528554
rect 176910 528486 177016 528509
rect 177101 528528 177167 528532
rect 177101 528494 177117 528528
rect 177151 528494 177167 528528
rect 177101 528452 177167 528494
rect 177241 528520 177252 528554
rect 177235 528513 177252 528520
rect 177201 528486 177252 528513
rect 177379 528580 177437 528597
rect 177379 528546 177391 528580
rect 177425 528546 177437 528580
rect 177379 528452 177437 528546
rect 177471 528554 177548 528600
rect 177582 528578 177807 528612
rect 177471 528520 177508 528554
rect 177542 528520 177548 528554
rect 177751 528554 177807 528578
rect 177471 528486 177548 528520
rect 177582 528528 177647 528544
rect 177582 528494 177598 528528
rect 177632 528494 177647 528528
rect 177582 528452 177647 528494
rect 177751 528520 177757 528554
rect 177791 528520 177807 528554
rect 177751 528486 177807 528520
rect 177845 528554 177925 528646
rect 177959 528792 178150 528836
rect 178393 528920 178452 528962
rect 178393 528886 178409 528920
rect 178443 528886 178452 528920
rect 178393 528852 178452 528886
rect 178393 528818 178409 528852
rect 178443 528818 178452 528852
rect 178393 528800 178452 528818
rect 178488 528912 178537 528928
rect 178488 528878 178495 528912
rect 178529 528878 178537 528912
rect 178488 528844 178537 528878
rect 178488 528810 178495 528844
rect 178529 528810 178537 528844
rect 177959 528684 178001 528792
rect 177959 528650 177961 528684
rect 177995 528650 178001 528684
rect 177959 528612 178001 528650
rect 178035 528724 178127 528758
rect 178161 528724 178173 528758
rect 178035 528684 178173 528724
rect 178488 528700 178537 528810
rect 178572 528920 178624 528962
rect 178744 528961 179999 528962
rect 178572 528886 178581 528920
rect 178615 528886 178624 528920
rect 178572 528852 178624 528886
rect 178572 528818 178581 528852
rect 178615 528818 178624 528852
rect 178572 528800 178624 528818
rect 178660 528904 178710 528927
rect 178660 528870 178667 528904
rect 178701 528870 178710 528904
rect 178660 528836 178710 528870
rect 178660 528802 178667 528836
rect 178701 528802 178710 528836
rect 178744 528920 178796 528961
rect 178744 528886 178753 528920
rect 178787 528886 178796 528920
rect 178744 528852 178796 528886
rect 178744 528818 178753 528852
rect 178787 528818 178796 528852
rect 178744 528802 178796 528818
rect 178830 528876 178882 528927
rect 178830 528842 178839 528876
rect 178873 528842 178882 528876
rect 178660 528700 178710 528802
rect 178830 528790 178882 528842
rect 178916 528896 178968 528961
rect 178916 528862 178925 528896
rect 178959 528862 178968 528896
rect 178916 528816 178968 528862
rect 179002 528876 179054 528927
rect 179002 528842 179011 528876
rect 179045 528842 179054 528876
rect 178830 528756 178839 528790
rect 178873 528782 178882 528790
rect 179002 528790 179054 528842
rect 179088 528896 179140 528961
rect 179088 528862 179097 528896
rect 179131 528862 179140 528896
rect 179088 528816 179140 528862
rect 179174 528876 179226 528927
rect 179174 528842 179183 528876
rect 179217 528842 179226 528876
rect 179002 528782 179011 528790
rect 178873 528756 179011 528782
rect 179045 528782 179054 528790
rect 179174 528790 179226 528842
rect 179260 528896 179312 528961
rect 179260 528862 179269 528896
rect 179303 528862 179312 528896
rect 179260 528816 179312 528862
rect 179346 528876 179398 528927
rect 179346 528842 179355 528876
rect 179389 528842 179398 528876
rect 179174 528782 179183 528790
rect 179045 528756 179183 528782
rect 179217 528782 179226 528790
rect 179346 528790 179398 528842
rect 179432 528896 179481 528961
rect 179432 528862 179441 528896
rect 179475 528862 179481 528896
rect 179432 528816 179481 528862
rect 179515 528876 179567 528927
rect 179515 528842 179526 528876
rect 179560 528842 179567 528876
rect 179346 528782 179355 528790
rect 179217 528756 179355 528782
rect 179389 528782 179398 528790
rect 179515 528790 179567 528842
rect 179604 528896 179653 528961
rect 179604 528862 179612 528896
rect 179646 528862 179653 528896
rect 179604 528816 179653 528862
rect 179687 528894 179739 528927
rect 179687 528860 179691 528894
rect 179725 528876 179739 528894
rect 179687 528842 179698 528860
rect 179732 528842 179739 528876
rect 179515 528782 179526 528790
rect 179389 528756 179526 528782
rect 179560 528782 179567 528790
rect 179687 528790 179739 528842
rect 179776 528896 179825 528961
rect 179776 528862 179784 528896
rect 179818 528862 179825 528896
rect 179776 528816 179825 528862
rect 179859 528876 179911 528927
rect 179859 528842 179870 528876
rect 179904 528842 179911 528876
rect 179687 528782 179698 528790
rect 179560 528756 179698 528782
rect 179732 528782 179739 528790
rect 179859 528790 179911 528842
rect 179948 528896 179999 528961
rect 179948 528862 179956 528896
rect 179990 528862 179999 528896
rect 179948 528816 179999 528862
rect 180033 528876 180091 528927
rect 180033 528842 180042 528876
rect 180076 528842 180091 528876
rect 179859 528782 179870 528790
rect 179732 528756 179870 528782
rect 179904 528779 179911 528790
rect 180033 528790 180091 528842
rect 180125 528896 180179 528962
rect 180125 528862 180128 528896
rect 180162 528862 180179 528896
rect 180125 528813 180179 528862
rect 180249 528912 180283 528928
rect 180249 528844 180283 528878
rect 180033 528779 180042 528790
rect 179904 528756 180042 528779
rect 180076 528779 180091 528790
rect 180319 528912 180385 528962
rect 180319 528878 180335 528912
rect 180369 528878 180385 528912
rect 180319 528844 180385 528878
rect 180319 528810 180335 528844
rect 180369 528810 180385 528844
rect 180419 528912 180473 528928
rect 180419 528878 180421 528912
rect 180455 528878 180473 528912
rect 180419 528831 180473 528878
rect 180076 528756 180179 528779
rect 178830 528734 180179 528756
rect 180249 528776 180283 528810
rect 180419 528797 180421 528831
rect 180455 528826 180473 528831
rect 180419 528792 180427 528797
rect 180461 528792 180473 528826
rect 180508 528912 180559 528928
rect 180508 528878 180525 528912
rect 180508 528844 180559 528878
rect 180593 528896 180659 528962
rect 180593 528862 180609 528896
rect 180643 528862 180659 528896
rect 180693 528912 180727 528928
rect 180508 528810 180525 528844
rect 180693 528844 180727 528878
rect 180559 528810 180658 528828
rect 180508 528794 180658 528810
rect 180249 528742 180382 528776
rect 180419 528747 180473 528792
rect 178035 528650 178075 528684
rect 178109 528650 178173 528684
rect 178035 528646 178173 528650
rect 178391 528684 178454 528700
rect 178391 528650 178411 528684
rect 178445 528650 178454 528684
rect 178391 528622 178454 528650
rect 177959 528578 178150 528612
rect 178391 528588 178403 528622
rect 178437 528588 178454 528622
rect 178488 528684 179912 528700
rect 178488 528650 178838 528684
rect 178872 528650 178906 528684
rect 178940 528650 178974 528684
rect 179008 528650 179042 528684
rect 179076 528650 179110 528684
rect 179144 528650 179178 528684
rect 179212 528650 179246 528684
rect 179280 528650 179314 528684
rect 179348 528650 179382 528684
rect 179416 528650 179450 528684
rect 179484 528650 179518 528684
rect 179552 528650 179586 528684
rect 179620 528650 179654 528684
rect 179688 528650 179722 528684
rect 179756 528650 179790 528684
rect 179824 528650 179858 528684
rect 179892 528650 179912 528684
rect 177845 528520 177861 528554
rect 177895 528520 177925 528554
rect 178093 528554 178150 528578
rect 177845 528486 177925 528520
rect 178005 528528 178059 528544
rect 178005 528494 178015 528528
rect 178049 528494 178059 528528
rect 178005 528452 178059 528494
rect 178093 528520 178099 528554
rect 178133 528520 178150 528554
rect 178093 528486 178150 528520
rect 178391 528528 178452 528554
rect 178391 528494 178409 528528
rect 178443 528494 178452 528528
rect 178391 528452 178452 528494
rect 178488 528541 178538 528650
rect 178488 528507 178495 528541
rect 178529 528507 178538 528541
rect 178488 528488 178538 528507
rect 178572 528541 178624 528557
rect 178572 528507 178581 528541
rect 178615 528507 178624 528541
rect 178572 528452 178624 528507
rect 178660 528541 178710 528650
rect 179946 528616 180179 528734
rect 180348 528713 180382 528742
rect 180235 528690 180301 528706
rect 180235 528656 180243 528690
rect 180277 528684 180301 528690
rect 180235 528650 180251 528656
rect 180285 528650 180301 528684
rect 180235 528632 180301 528650
rect 180348 528697 180405 528713
rect 180348 528663 180371 528697
rect 180348 528647 180405 528663
rect 178830 528582 180179 528616
rect 180348 528596 180382 528647
rect 178660 528507 178667 528541
rect 178701 528507 178710 528541
rect 178660 528488 178710 528507
rect 178744 528541 178796 528564
rect 178744 528507 178753 528541
rect 178787 528507 178796 528541
rect 178744 528452 178796 528507
rect 178830 528541 178882 528582
rect 178830 528507 178839 528541
rect 178873 528507 178882 528541
rect 178830 528491 178882 528507
rect 178916 528532 178968 528548
rect 178916 528498 178925 528532
rect 178959 528498 178968 528532
rect 178916 528452 178968 528498
rect 179002 528541 179054 528582
rect 179002 528507 179011 528541
rect 179045 528507 179054 528541
rect 179002 528491 179054 528507
rect 179088 528532 179140 528548
rect 179088 528498 179097 528532
rect 179131 528498 179140 528532
rect 179088 528452 179140 528498
rect 179174 528541 179226 528582
rect 179174 528507 179183 528541
rect 179217 528507 179226 528541
rect 179174 528491 179226 528507
rect 179260 528532 179309 528548
rect 179260 528498 179269 528532
rect 179303 528498 179309 528532
rect 179260 528452 179309 528498
rect 179343 528541 179398 528582
rect 179343 528507 179355 528541
rect 179389 528507 179398 528541
rect 179343 528491 179398 528507
rect 179432 528532 179481 528548
rect 179432 528498 179441 528532
rect 179475 528498 179481 528532
rect 179432 528452 179481 528498
rect 179515 528541 179567 528582
rect 179515 528507 179526 528541
rect 179560 528507 179567 528541
rect 179515 528491 179567 528507
rect 179603 528532 179653 528548
rect 179603 528498 179612 528532
rect 179646 528498 179653 528532
rect 179603 528452 179653 528498
rect 179687 528541 179739 528582
rect 179687 528507 179698 528541
rect 179732 528507 179739 528541
rect 179687 528491 179739 528507
rect 179775 528532 179825 528548
rect 179775 528498 179784 528532
rect 179818 528498 179825 528532
rect 179775 528452 179825 528498
rect 179859 528541 179911 528582
rect 179859 528507 179870 528541
rect 179904 528507 179911 528541
rect 179859 528491 179911 528507
rect 179947 528532 179999 528548
rect 179947 528498 179956 528532
rect 179990 528498 179999 528532
rect 179947 528452 179999 528498
rect 180033 528541 180085 528582
rect 180249 528562 180382 528596
rect 180439 528587 180473 528747
rect 180508 528758 180578 528760
rect 180508 528724 180519 528758
rect 180553 528724 180578 528758
rect 180508 528684 180578 528724
rect 180508 528650 180522 528684
rect 180556 528650 180578 528684
rect 180508 528630 180578 528650
rect 180612 528699 180658 528794
rect 180612 528690 180624 528699
rect 180646 528656 180658 528665
rect 180612 528596 180658 528656
rect 180033 528507 180042 528541
rect 180076 528507 180085 528541
rect 180033 528491 180085 528507
rect 180119 528532 180179 528548
rect 180119 528498 180128 528532
rect 180162 528498 180179 528532
rect 180119 528452 180179 528498
rect 180249 528541 180283 528562
rect 180421 528558 180473 528587
rect 180249 528486 180283 528507
rect 180319 528494 180335 528528
rect 180369 528494 180385 528528
rect 180319 528452 180385 528494
rect 180455 528524 180473 528558
rect 180421 528486 180473 528524
rect 180508 528562 180658 528596
rect 180508 528554 180559 528562
rect 180508 528520 180525 528554
rect 180693 528554 180727 528792
rect 180761 528768 180826 528925
rect 180860 528920 180910 528962
rect 180860 528886 180876 528920
rect 180860 528870 180910 528886
rect 180944 528912 180994 528928
rect 180944 528878 180960 528912
rect 180944 528862 180994 528878
rect 181037 528918 181173 528928
rect 181037 528884 181053 528918
rect 181087 528884 181173 528918
rect 181288 528910 181354 528962
rect 181481 528920 181555 528962
rect 181037 528862 181173 528884
rect 180944 528836 180978 528862
rect 180899 528802 180978 528836
rect 181012 528826 181105 528828
rect 180773 528758 180865 528768
rect 180773 528724 180795 528758
rect 180829 528745 180865 528758
rect 180829 528724 180831 528745
rect 180773 528711 180831 528724
rect 180773 528558 180865 528711
rect 180508 528504 180559 528520
rect 180593 528494 180609 528528
rect 180643 528494 180659 528528
rect 180899 528530 180933 528802
rect 181012 528800 181071 528826
rect 181046 528792 181071 528800
rect 181046 528766 181105 528792
rect 181012 528750 181105 528766
rect 180967 528690 181037 528712
rect 180967 528656 180979 528690
rect 181013 528656 181037 528690
rect 180967 528638 181037 528656
rect 180967 528604 180990 528638
rect 181024 528604 181037 528638
rect 180967 528588 181037 528604
rect 181071 528632 181105 528750
rect 181139 528706 181173 528862
rect 181207 528894 181241 528910
rect 181288 528876 181304 528910
rect 181338 528876 181354 528910
rect 181388 528894 181422 528910
rect 181207 528842 181241 528860
rect 181481 528886 181501 528920
rect 181535 528886 181555 528920
rect 181481 528870 181555 528886
rect 181589 528912 181623 528928
rect 181388 528842 181422 528860
rect 181207 528808 181422 528842
rect 181589 528836 181623 528878
rect 181670 528919 181844 528928
rect 181670 528885 181686 528919
rect 181720 528885 181844 528919
rect 181670 528860 181844 528885
rect 181878 528920 181928 528962
rect 181912 528886 181928 528920
rect 182032 528920 182098 528962
rect 181878 528870 181928 528886
rect 181962 528894 181996 528910
rect 181511 528802 181623 528836
rect 181511 528774 181545 528802
rect 181245 528740 181261 528774
rect 181295 528740 181545 528774
rect 181684 528792 181695 528826
rect 181729 528800 181776 528826
rect 181684 528768 181726 528792
rect 181139 528686 181477 528706
rect 181139 528672 181443 528686
rect 181071 528598 181092 528632
rect 181126 528598 181142 528632
rect 181071 528588 181142 528598
rect 181176 528530 181210 528672
rect 181251 528622 181347 528638
rect 181285 528588 181323 528622
rect 181381 528604 181409 528638
rect 181443 528636 181477 528652
rect 181357 528588 181409 528604
rect 181511 528602 181545 528740
rect 180693 528504 180727 528520
rect 180593 528452 180659 528494
rect 180799 528490 180815 528524
rect 180849 528490 180865 528524
rect 180899 528496 180948 528530
rect 180982 528496 180998 528530
rect 181039 528496 181055 528530
rect 181089 528496 181210 528530
rect 181385 528528 181451 528544
rect 180799 528452 180865 528490
rect 181385 528494 181401 528528
rect 181435 528494 181451 528528
rect 181385 528452 181451 528494
rect 181493 528524 181545 528602
rect 181583 528766 181726 528768
rect 181760 528766 181776 528800
rect 181810 528784 181844 528860
rect 182032 528886 182048 528920
rect 182082 528886 182098 528920
rect 182166 528920 182227 528962
rect 182166 528886 182177 528920
rect 182211 528886 182227 528920
rect 181962 528852 181996 528860
rect 182166 528852 182227 528886
rect 181962 528818 182122 528852
rect 181583 528734 181718 528766
rect 181810 528750 182004 528784
rect 182038 528750 182054 528784
rect 181583 528626 181625 528734
rect 181810 528732 181844 528750
rect 181583 528592 181591 528626
rect 181583 528576 181625 528592
rect 181659 528690 181729 528700
rect 181659 528674 181695 528690
rect 181659 528640 181687 528674
rect 181721 528640 181729 528656
rect 181659 528576 181729 528640
rect 181763 528698 181844 528732
rect 181763 528542 181797 528698
rect 181911 528685 182019 528716
rect 182088 528700 182122 528818
rect 182166 528818 182177 528852
rect 182211 528818 182227 528852
rect 182166 528734 182227 528818
rect 182261 528894 182312 528900
rect 182261 528884 182267 528894
rect 182301 528860 182312 528894
rect 182295 528850 182312 528860
rect 182261 528816 182312 528850
rect 182295 528782 182312 528816
rect 182261 528724 182312 528782
rect 182531 528891 182589 528962
rect 182531 528857 182543 528891
rect 182577 528857 182589 528891
rect 182623 528920 183692 528962
rect 182623 528886 182641 528920
rect 182675 528886 183641 528920
rect 183675 528886 183692 528920
rect 182623 528875 183692 528886
rect 183727 528920 184796 528962
rect 183727 528886 183745 528920
rect 183779 528886 184745 528920
rect 184779 528886 184796 528920
rect 183727 528875 184796 528886
rect 184831 528920 185900 528962
rect 184831 528886 184849 528920
rect 184883 528886 185849 528920
rect 185883 528886 185900 528920
rect 184831 528875 185900 528886
rect 185935 528920 187004 528962
rect 185935 528886 185953 528920
rect 185987 528886 186953 528920
rect 186987 528886 187004 528920
rect 185935 528875 187004 528886
rect 187223 528920 187465 528962
rect 187223 528886 187241 528920
rect 187275 528886 187413 528920
rect 187447 528886 187465 528920
rect 182531 528798 182589 528857
rect 182531 528764 182543 528798
rect 182577 528764 182589 528798
rect 182531 528729 182589 528764
rect 182088 528694 182236 528700
rect 181945 528676 182019 528685
rect 181831 528648 181875 528664
rect 181865 528614 181875 528648
rect 181911 528642 181927 528651
rect 181961 528642 182019 528676
rect 181831 528608 181875 528614
rect 181971 528622 182019 528642
rect 181831 528574 181937 528608
rect 181607 528528 181797 528542
rect 181493 528490 181513 528524
rect 181547 528490 181563 528524
rect 181607 528494 181623 528528
rect 181657 528494 181797 528528
rect 181607 528486 181797 528494
rect 181831 528524 181869 528540
rect 181831 528490 181835 528524
rect 181903 528528 181937 528574
rect 182005 528588 182019 528622
rect 181971 528562 182019 528588
rect 182053 528684 182236 528694
rect 182053 528650 182202 528684
rect 182053 528634 182236 528650
rect 182053 528599 182118 528634
rect 182053 528544 182117 528599
rect 182270 528594 182312 528724
rect 182940 528710 183008 528727
rect 182940 528676 182957 528710
rect 182991 528676 183008 528710
rect 182261 528578 182312 528594
rect 182295 528544 182312 528578
rect 181903 528510 182053 528528
rect 182087 528510 182117 528544
rect 181903 528494 182117 528510
rect 182166 528528 182227 528544
rect 182166 528494 182177 528528
rect 182211 528494 182227 528528
rect 181831 528452 181869 528490
rect 182166 528452 182227 528494
rect 182261 528488 182312 528544
rect 182531 528580 182589 528597
rect 182531 528546 182543 528580
rect 182577 528546 182589 528580
rect 182940 528561 183008 528676
rect 183304 528674 183374 528875
rect 183304 528640 183321 528674
rect 183355 528640 183374 528674
rect 183304 528625 183374 528640
rect 184044 528710 184112 528727
rect 184044 528676 184061 528710
rect 184095 528676 184112 528710
rect 184044 528561 184112 528676
rect 184408 528674 184478 528875
rect 184408 528640 184425 528674
rect 184459 528640 184478 528674
rect 184408 528625 184478 528640
rect 185148 528710 185216 528727
rect 185148 528676 185165 528710
rect 185199 528676 185216 528710
rect 185148 528561 185216 528676
rect 185512 528674 185582 528875
rect 185512 528640 185529 528674
rect 185563 528640 185582 528674
rect 185512 528625 185582 528640
rect 186252 528710 186320 528727
rect 186252 528676 186269 528710
rect 186303 528676 186320 528710
rect 186252 528561 186320 528676
rect 186616 528674 186686 528875
rect 186616 528640 186633 528674
rect 186667 528640 186686 528674
rect 186616 528625 186686 528640
rect 187223 528825 187465 528886
rect 187223 528791 187241 528825
rect 187275 528791 187413 528825
rect 187447 528791 187465 528825
rect 187223 528744 187465 528791
rect 187223 528670 187327 528744
rect 187223 528636 187273 528670
rect 187307 528636 187327 528670
rect 187361 528676 187381 528710
rect 187415 528676 187465 528710
rect 187361 528602 187465 528676
rect 182531 528452 182589 528546
rect 182623 528547 183692 528561
rect 182623 528513 182641 528547
rect 182675 528513 183641 528547
rect 183675 528513 183692 528547
rect 182623 528452 183692 528513
rect 183727 528547 184796 528561
rect 183727 528513 183745 528547
rect 183779 528513 184745 528547
rect 184779 528513 184796 528547
rect 183727 528452 184796 528513
rect 184831 528547 185900 528561
rect 184831 528513 184849 528547
rect 184883 528513 185849 528547
rect 185883 528513 185900 528547
rect 184831 528452 185900 528513
rect 185935 528547 187004 528561
rect 185935 528513 185953 528547
rect 185987 528513 186953 528547
rect 186987 528513 187004 528547
rect 185935 528452 187004 528513
rect 187223 528549 187465 528602
rect 187223 528515 187241 528549
rect 187275 528515 187413 528549
rect 187447 528515 187465 528549
rect 187223 528452 187465 528515
rect 172210 528418 172239 528452
rect 172273 528418 172331 528452
rect 172365 528418 172423 528452
rect 172457 528418 172515 528452
rect 172549 528418 172607 528452
rect 172641 528418 172699 528452
rect 172733 528418 172791 528452
rect 172825 528418 172883 528452
rect 172917 528418 172975 528452
rect 173009 528418 173067 528452
rect 173101 528418 173159 528452
rect 173193 528418 173251 528452
rect 173285 528418 173343 528452
rect 173377 528418 173435 528452
rect 173469 528418 173527 528452
rect 173561 528418 173619 528452
rect 173653 528418 173711 528452
rect 173745 528418 173803 528452
rect 173837 528418 173895 528452
rect 173929 528418 173987 528452
rect 174021 528418 174079 528452
rect 174113 528418 174171 528452
rect 174205 528418 174263 528452
rect 174297 528418 174355 528452
rect 174389 528418 174447 528452
rect 174481 528418 174539 528452
rect 174573 528418 174631 528452
rect 174665 528418 174723 528452
rect 174757 528418 174815 528452
rect 174849 528418 174907 528452
rect 174941 528418 174999 528452
rect 175033 528418 175091 528452
rect 175125 528418 175183 528452
rect 175217 528418 175275 528452
rect 175309 528418 175367 528452
rect 175401 528418 175459 528452
rect 175493 528418 175551 528452
rect 175585 528418 175643 528452
rect 175677 528418 175735 528452
rect 175769 528418 175827 528452
rect 175861 528418 175919 528452
rect 175953 528418 176011 528452
rect 176045 528418 176103 528452
rect 176137 528418 176195 528452
rect 176229 528418 176287 528452
rect 176321 528418 176379 528452
rect 176413 528418 176471 528452
rect 176505 528418 176563 528452
rect 176597 528418 176655 528452
rect 176689 528418 176747 528452
rect 176781 528418 176839 528452
rect 176873 528418 176931 528452
rect 176965 528418 177023 528452
rect 177057 528418 177115 528452
rect 177149 528418 177207 528452
rect 177241 528418 177299 528452
rect 177333 528418 177391 528452
rect 177425 528418 177483 528452
rect 177517 528418 177575 528452
rect 177609 528418 177667 528452
rect 177701 528418 177759 528452
rect 177793 528418 177851 528452
rect 177885 528418 177943 528452
rect 177977 528418 178035 528452
rect 178069 528418 178127 528452
rect 178161 528418 178219 528452
rect 178253 528418 178311 528452
rect 178345 528418 178403 528452
rect 178437 528418 178495 528452
rect 178529 528418 178587 528452
rect 178621 528418 178679 528452
rect 178713 528418 178771 528452
rect 178805 528418 178863 528452
rect 178897 528418 178955 528452
rect 178989 528418 179047 528452
rect 179081 528418 179139 528452
rect 179173 528418 179231 528452
rect 179265 528418 179323 528452
rect 179357 528418 179415 528452
rect 179449 528418 179507 528452
rect 179541 528418 179599 528452
rect 179633 528418 179691 528452
rect 179725 528418 179783 528452
rect 179817 528418 179875 528452
rect 179909 528418 179967 528452
rect 180001 528418 180059 528452
rect 180093 528418 180151 528452
rect 180185 528418 180243 528452
rect 180277 528418 180335 528452
rect 180369 528418 180427 528452
rect 180461 528418 180519 528452
rect 180553 528418 180611 528452
rect 180645 528418 180703 528452
rect 180737 528418 180795 528452
rect 180829 528418 180887 528452
rect 180921 528418 180979 528452
rect 181013 528418 181071 528452
rect 181105 528418 181163 528452
rect 181197 528418 181255 528452
rect 181289 528418 181347 528452
rect 181381 528418 181439 528452
rect 181473 528418 181531 528452
rect 181565 528418 181623 528452
rect 181657 528418 181715 528452
rect 181749 528418 181807 528452
rect 181841 528418 181899 528452
rect 181933 528418 181991 528452
rect 182025 528418 182083 528452
rect 182117 528418 182175 528452
rect 182209 528418 182267 528452
rect 182301 528418 182359 528452
rect 182393 528418 182451 528452
rect 182485 528418 182543 528452
rect 182577 528418 182635 528452
rect 182669 528418 182727 528452
rect 182761 528418 182819 528452
rect 182853 528418 182911 528452
rect 182945 528418 183003 528452
rect 183037 528418 183095 528452
rect 183129 528418 183187 528452
rect 183221 528418 183279 528452
rect 183313 528418 183371 528452
rect 183405 528418 183463 528452
rect 183497 528418 183555 528452
rect 183589 528418 183647 528452
rect 183681 528418 183739 528452
rect 183773 528418 183831 528452
rect 183865 528418 183923 528452
rect 183957 528418 184015 528452
rect 184049 528418 184107 528452
rect 184141 528418 184199 528452
rect 184233 528418 184291 528452
rect 184325 528418 184383 528452
rect 184417 528418 184475 528452
rect 184509 528418 184567 528452
rect 184601 528418 184659 528452
rect 184693 528418 184751 528452
rect 184785 528418 184843 528452
rect 184877 528418 184935 528452
rect 184969 528418 185027 528452
rect 185061 528418 185119 528452
rect 185153 528418 185211 528452
rect 185245 528418 185303 528452
rect 185337 528418 185395 528452
rect 185429 528418 185487 528452
rect 185521 528418 185579 528452
rect 185613 528418 185671 528452
rect 185705 528418 185763 528452
rect 185797 528418 185855 528452
rect 185889 528418 185947 528452
rect 185981 528418 186039 528452
rect 186073 528418 186131 528452
rect 186165 528418 186223 528452
rect 186257 528418 186315 528452
rect 186349 528418 186407 528452
rect 186441 528418 186499 528452
rect 186533 528418 186591 528452
rect 186625 528418 186683 528452
rect 186717 528418 186775 528452
rect 186809 528418 186867 528452
rect 186901 528418 186959 528452
rect 186993 528418 187051 528452
rect 187085 528418 187143 528452
rect 187177 528418 187235 528452
rect 187269 528418 187327 528452
rect 187361 528418 187419 528452
rect 187453 528418 187482 528452
rect 172227 528355 172469 528418
rect 172227 528321 172245 528355
rect 172279 528321 172417 528355
rect 172451 528321 172469 528355
rect 172227 528268 172469 528321
rect 172503 528357 173572 528418
rect 172503 528323 172521 528357
rect 172555 528323 173521 528357
rect 173555 528323 173572 528357
rect 172503 528309 173572 528323
rect 173607 528357 174676 528418
rect 173607 528323 173625 528357
rect 173659 528323 174625 528357
rect 174659 528323 174676 528357
rect 173607 528309 174676 528323
rect 174803 528324 174861 528418
rect 172227 528194 172331 528268
rect 172227 528160 172277 528194
rect 172311 528160 172331 528194
rect 172365 528200 172385 528234
rect 172419 528200 172469 528234
rect 172365 528126 172469 528200
rect 172820 528194 172888 528309
rect 172820 528160 172837 528194
rect 172871 528160 172888 528194
rect 172820 528143 172888 528160
rect 173184 528230 173254 528245
rect 173184 528196 173201 528230
rect 173235 528196 173254 528230
rect 172227 528079 172469 528126
rect 172227 528045 172245 528079
rect 172279 528045 172417 528079
rect 172451 528045 172469 528079
rect 172227 527984 172469 528045
rect 173184 527995 173254 528196
rect 173924 528194 173992 528309
rect 174803 528290 174815 528324
rect 174849 528290 174861 528324
rect 174895 528357 175964 528418
rect 176177 528376 176243 528418
rect 174895 528323 174913 528357
rect 174947 528323 175913 528357
rect 175947 528323 175964 528357
rect 174895 528309 175964 528323
rect 176092 528350 176143 528366
rect 176092 528316 176109 528350
rect 176177 528342 176193 528376
rect 176227 528342 176243 528376
rect 176383 528380 176449 528418
rect 176277 528350 176311 528366
rect 174803 528273 174861 528290
rect 173924 528160 173941 528194
rect 173975 528160 173992 528194
rect 173924 528143 173992 528160
rect 174288 528230 174358 528245
rect 174288 528196 174305 528230
rect 174339 528196 174358 528230
rect 174288 527995 174358 528196
rect 175212 528194 175280 528309
rect 176092 528308 176143 528316
rect 176383 528346 176399 528380
rect 176433 528346 176449 528380
rect 176969 528376 177035 528418
rect 176092 528274 176242 528308
rect 175212 528160 175229 528194
rect 175263 528160 175280 528194
rect 175212 528143 175280 528160
rect 175576 528230 175646 528245
rect 175576 528196 175593 528230
rect 175627 528196 175646 528230
rect 174803 528106 174861 528141
rect 174803 528072 174815 528106
rect 174849 528072 174861 528106
rect 174803 528013 174861 528072
rect 172227 527950 172245 527984
rect 172279 527950 172417 527984
rect 172451 527950 172469 527984
rect 172227 527908 172469 527950
rect 172503 527984 173572 527995
rect 172503 527950 172521 527984
rect 172555 527950 173521 527984
rect 173555 527950 173572 527984
rect 172503 527908 173572 527950
rect 173607 527984 174676 527995
rect 173607 527950 173625 527984
rect 173659 527950 174625 527984
rect 174659 527950 174676 527984
rect 173607 527908 174676 527950
rect 174803 527979 174815 528013
rect 174849 527979 174861 528013
rect 175576 527995 175646 528196
rect 176092 528220 176162 528240
rect 176092 528214 176106 528220
rect 176092 528180 176103 528214
rect 176140 528186 176162 528220
rect 176137 528180 176162 528186
rect 176092 528110 176162 528180
rect 176196 528214 176242 528274
rect 176230 528205 176242 528214
rect 176196 528171 176208 528180
rect 176196 528076 176242 528171
rect 176092 528060 176242 528076
rect 176092 528026 176109 528060
rect 176143 528042 176242 528060
rect 176277 528078 176311 528316
rect 176483 528340 176532 528374
rect 176566 528340 176582 528374
rect 176623 528340 176639 528374
rect 176673 528340 176794 528374
rect 176357 528282 176449 528312
rect 176357 528248 176379 528282
rect 176413 528248 176449 528282
rect 176357 528159 176449 528248
rect 176357 528125 176415 528159
rect 176357 528102 176449 528125
rect 174803 527908 174861 527979
rect 174895 527984 175964 527995
rect 174895 527950 174913 527984
rect 174947 527950 175913 527984
rect 175947 527950 175964 527984
rect 174895 527908 175964 527950
rect 176092 527992 176143 528026
rect 176092 527958 176109 527992
rect 176092 527942 176143 527958
rect 176177 527974 176193 528008
rect 176227 527974 176243 528008
rect 176177 527908 176243 527974
rect 176277 527992 176311 528026
rect 176277 527942 176311 527958
rect 176345 527945 176410 528102
rect 176483 528068 176517 528340
rect 176551 528266 176621 528282
rect 176551 528232 176574 528266
rect 176608 528232 176621 528266
rect 176551 528214 176621 528232
rect 176551 528180 176563 528214
rect 176597 528180 176621 528214
rect 176551 528158 176621 528180
rect 176655 528272 176726 528282
rect 176655 528238 176676 528272
rect 176710 528238 176726 528272
rect 176655 528120 176689 528238
rect 176760 528198 176794 528340
rect 176969 528342 176985 528376
rect 177019 528342 177035 528376
rect 176969 528326 177035 528342
rect 177077 528346 177097 528380
rect 177131 528346 177147 528380
rect 177191 528376 177381 528384
rect 176869 528248 176907 528282
rect 176941 528266 176993 528282
rect 177077 528268 177129 528346
rect 177191 528342 177207 528376
rect 177241 528342 177381 528376
rect 177191 528328 177381 528342
rect 177415 528380 177453 528418
rect 177415 528346 177419 528380
rect 177750 528376 177811 528418
rect 177415 528330 177453 528346
rect 177487 528360 177701 528376
rect 177487 528342 177637 528360
rect 176835 528232 176931 528248
rect 176965 528232 176993 528266
rect 177027 528218 177061 528234
rect 176596 528104 176689 528120
rect 176630 528078 176689 528104
rect 176630 528070 176655 528078
rect 176483 528034 176562 528068
rect 176596 528044 176655 528070
rect 176596 528042 176689 528044
rect 176723 528184 177027 528198
rect 176723 528164 177061 528184
rect 176528 528008 176562 528034
rect 176723 528008 176757 528164
rect 177095 528130 177129 528268
rect 176829 528096 176845 528130
rect 176879 528096 177129 528130
rect 177167 528278 177209 528294
rect 177167 528244 177175 528278
rect 177167 528136 177209 528244
rect 177243 528230 177313 528294
rect 177243 528196 177271 528230
rect 177305 528214 177313 528230
rect 177243 528180 177279 528196
rect 177243 528170 177313 528180
rect 177347 528172 177381 528328
rect 177487 528296 177521 528342
rect 177671 528326 177701 528360
rect 177750 528342 177761 528376
rect 177795 528342 177811 528376
rect 177750 528326 177811 528342
rect 177845 528350 177896 528382
rect 177845 528326 177851 528350
rect 177415 528262 177521 528296
rect 177555 528282 177603 528308
rect 177415 528256 177459 528262
rect 177449 528222 177459 528256
rect 177589 528248 177603 528282
rect 177555 528228 177603 528248
rect 177415 528206 177459 528222
rect 177495 528219 177511 528228
rect 177545 528194 177603 528228
rect 177529 528185 177603 528194
rect 177347 528138 177428 528172
rect 177495 528154 177603 528185
rect 177637 528271 177701 528326
rect 177885 528316 177896 528350
rect 177879 528292 177896 528316
rect 177845 528276 177896 528292
rect 177637 528236 177702 528271
rect 177637 528220 177820 528236
rect 177637 528186 177786 528220
rect 177637 528176 177820 528186
rect 177672 528170 177820 528176
rect 177167 528104 177302 528136
rect 177394 528120 177428 528138
rect 177167 528102 177310 528104
rect 177095 528068 177129 528096
rect 177268 528078 177310 528102
rect 176444 527984 176494 528000
rect 176444 527950 176460 527984
rect 176444 527908 176494 527950
rect 176528 527992 176578 528008
rect 176528 527958 176544 527992
rect 176528 527942 176578 527958
rect 176621 527986 176757 528008
rect 176621 527952 176637 527986
rect 176671 527952 176757 527986
rect 176791 528028 177006 528062
rect 177095 528034 177207 528068
rect 177268 528044 177279 528078
rect 177344 528070 177360 528104
rect 177313 528044 177360 528070
rect 177394 528086 177588 528120
rect 177622 528086 177638 528120
rect 176791 528010 176825 528028
rect 176972 528010 177006 528028
rect 176791 527960 176825 527976
rect 176872 527960 176888 527994
rect 176922 527960 176938 527994
rect 176972 527960 177006 527976
rect 177065 527984 177139 528000
rect 176621 527942 176757 527952
rect 176872 527908 176938 527960
rect 177065 527950 177085 527984
rect 177119 527950 177139 527984
rect 177065 527908 177139 527950
rect 177173 527992 177207 528034
rect 177394 528010 177428 528086
rect 177672 528052 177706 528170
rect 177854 528146 177896 528276
rect 177173 527942 177207 527958
rect 177254 527985 177428 528010
rect 177546 528018 177706 528052
rect 177750 528052 177811 528136
rect 177750 528018 177761 528052
rect 177795 528018 177811 528052
rect 177546 528010 177580 528018
rect 177254 527951 177270 527985
rect 177304 527951 177428 527985
rect 177254 527942 177428 527951
rect 177462 527984 177512 528000
rect 177496 527950 177512 527984
rect 177750 527984 177811 528018
rect 177546 527960 177580 527976
rect 177462 527908 177512 527950
rect 177616 527950 177632 527984
rect 177666 527950 177682 527984
rect 177616 527908 177682 527950
rect 177750 527950 177761 527984
rect 177795 527950 177811 527984
rect 177845 528088 177896 528146
rect 177879 528054 177896 528088
rect 177845 528020 177896 528054
rect 177879 527986 177896 528020
rect 177845 527970 177896 527986
rect 177931 528346 177983 528384
rect 177931 528312 177949 528346
rect 178019 528376 178085 528418
rect 178019 528342 178035 528376
rect 178069 528342 178085 528376
rect 178121 528363 178155 528384
rect 177931 528283 177983 528312
rect 178121 528308 178155 528329
rect 177931 528123 177965 528283
rect 178022 528274 178155 528308
rect 178207 528357 178909 528418
rect 178207 528323 178225 528357
rect 178259 528323 178857 528357
rect 178891 528323 178909 528357
rect 178022 528223 178056 528274
rect 178207 528264 178909 528323
rect 178944 528357 178995 528384
rect 178944 528350 178961 528357
rect 178944 528316 178955 528350
rect 179029 528376 179095 528418
rect 179029 528342 179045 528376
rect 179079 528342 179095 528376
rect 179029 528338 179095 528342
rect 179180 528361 179286 528384
rect 178989 528316 178995 528323
rect 178944 528270 178995 528316
rect 179180 528327 179252 528361
rect 179180 528311 179286 528327
rect 179180 528304 179215 528311
rect 179029 528270 179215 528304
rect 177999 528207 178056 528223
rect 178033 528173 178056 528207
rect 177999 528157 178056 528173
rect 178103 528220 178169 528238
rect 178103 528186 178119 528220
rect 178153 528214 178169 528220
rect 178103 528180 178127 528186
rect 178161 528180 178169 528214
rect 178103 528164 178169 528180
rect 178207 528194 178537 528264
rect 178207 528160 178285 528194
rect 178319 528160 178384 528194
rect 178418 528160 178483 528194
rect 178517 528160 178537 528194
rect 178571 528196 178591 528230
rect 178625 528196 178694 528230
rect 178728 528196 178797 528230
rect 178831 528196 178909 528230
rect 178022 528128 178056 528157
rect 177931 528078 177985 528123
rect 178022 528094 178155 528128
rect 178571 528126 178909 528196
rect 177931 528044 177943 528078
rect 177977 528073 177985 528078
rect 177931 528039 177949 528044
rect 177983 528039 177985 528073
rect 178121 528060 178155 528094
rect 177931 527992 177985 528039
rect 177750 527908 177811 527950
rect 177931 527958 177949 527992
rect 177983 527958 177985 527992
rect 177931 527942 177985 527958
rect 178019 528026 178035 528060
rect 178069 528026 178085 528060
rect 178019 527992 178085 528026
rect 178019 527958 178035 527992
rect 178069 527958 178085 527992
rect 178019 527908 178085 527958
rect 178121 527992 178155 528026
rect 178121 527942 178155 527958
rect 178207 528086 178909 528126
rect 178207 528052 178225 528086
rect 178259 528052 178857 528086
rect 178891 528052 178909 528086
rect 178207 527984 178909 528052
rect 178207 527950 178225 527984
rect 178259 527950 178857 527984
rect 178891 527950 178909 527984
rect 178207 527908 178909 527950
rect 178944 528136 178978 528270
rect 179029 528236 179063 528270
rect 179012 528220 179063 528236
rect 179046 528186 179063 528220
rect 179012 528170 179063 528186
rect 179108 528220 179147 528236
rect 179142 528186 179147 528220
rect 179108 528170 179147 528186
rect 178944 528120 179011 528136
rect 178944 528086 178961 528120
rect 178995 528086 179011 528120
rect 178944 528052 179011 528086
rect 178944 528018 178961 528052
rect 178995 528018 179011 528052
rect 178944 527984 179011 528018
rect 178944 527950 178961 527984
rect 178995 527950 179011 527984
rect 178944 527942 179011 527950
rect 179045 528120 179079 528136
rect 179045 528052 179079 528086
rect 179045 527984 179079 528018
rect 179045 527908 179079 527950
rect 179113 527976 179147 528170
rect 179181 528044 179215 528270
rect 179249 528256 179283 528272
rect 179249 528112 179283 528222
rect 179324 528256 179379 528384
rect 179324 528222 179345 528256
rect 179324 528214 179379 528222
rect 179357 528180 179379 528214
rect 179324 528152 179379 528180
rect 179413 528350 179451 528384
rect 179413 528316 179415 528350
rect 179449 528316 179451 528350
rect 179413 528143 179451 528316
rect 179487 528361 179589 528418
rect 179521 528327 179555 528361
rect 179487 528311 179589 528327
rect 179633 528361 179682 528377
rect 179633 528327 179639 528361
rect 179673 528327 179682 528361
rect 179633 528256 179682 528327
rect 179955 528324 180013 528418
rect 179955 528290 179967 528324
rect 180001 528290 180013 528324
rect 179955 528273 180013 528290
rect 180047 528357 180749 528418
rect 180047 528323 180065 528357
rect 180099 528323 180697 528357
rect 180731 528323 180749 528357
rect 180047 528264 180749 528323
rect 180968 528357 181019 528384
rect 180968 528350 180985 528357
rect 180968 528316 180979 528350
rect 181053 528376 181119 528418
rect 181053 528342 181069 528376
rect 181103 528342 181119 528376
rect 181053 528338 181119 528342
rect 181204 528361 181310 528384
rect 181013 528316 181019 528323
rect 180968 528270 181019 528316
rect 181204 528327 181276 528361
rect 181204 528311 181310 528327
rect 181204 528304 181239 528311
rect 181053 528270 181239 528304
rect 179491 528222 179507 528256
rect 179541 528222 179737 528256
rect 179413 528112 179417 528143
rect 179249 528109 179417 528112
rect 179249 528078 179451 528109
rect 179485 528146 179635 528147
rect 179485 528112 179507 528146
rect 179541 528143 179635 528146
rect 179541 528112 179585 528143
rect 179485 528109 179585 528112
rect 179619 528109 179635 528143
rect 179181 528010 179281 528044
rect 179315 528010 179356 528044
rect 179390 528010 179406 528044
rect 179485 527976 179519 528109
rect 179669 528060 179737 528222
rect 180047 528194 180377 528264
rect 180047 528160 180125 528194
rect 180159 528160 180224 528194
rect 180258 528160 180323 528194
rect 180357 528160 180377 528194
rect 180411 528196 180431 528230
rect 180465 528196 180534 528230
rect 180568 528196 180637 528230
rect 180671 528196 180749 528230
rect 179113 527942 179519 527976
rect 179553 528044 179587 528060
rect 179553 527908 179587 528010
rect 179634 528044 179737 528060
rect 179634 528010 179639 528044
rect 179673 528010 179737 528044
rect 179634 527978 179737 528010
rect 179955 528106 180013 528141
rect 180411 528126 180749 528196
rect 179955 528072 179967 528106
rect 180001 528072 180013 528106
rect 179955 528013 180013 528072
rect 179955 527979 179967 528013
rect 180001 527979 180013 528013
rect 179955 527908 180013 527979
rect 180047 528086 180749 528126
rect 180047 528052 180065 528086
rect 180099 528052 180697 528086
rect 180731 528052 180749 528086
rect 180047 527984 180749 528052
rect 180047 527950 180065 527984
rect 180099 527950 180697 527984
rect 180731 527950 180749 527984
rect 180047 527908 180749 527950
rect 180968 528136 181002 528270
rect 181053 528236 181087 528270
rect 181036 528220 181087 528236
rect 181070 528186 181087 528220
rect 181036 528170 181087 528186
rect 181132 528220 181171 528236
rect 181166 528186 181171 528220
rect 181132 528170 181171 528186
rect 180968 528120 181035 528136
rect 180968 528086 180985 528120
rect 181019 528086 181035 528120
rect 180968 528052 181035 528086
rect 180968 528018 180985 528052
rect 181019 528018 181035 528052
rect 180968 527984 181035 528018
rect 180968 527950 180985 527984
rect 181019 527950 181035 527984
rect 180968 527942 181035 527950
rect 181069 528120 181103 528136
rect 181069 528052 181103 528086
rect 181069 527984 181103 528018
rect 181069 527908 181103 527950
rect 181137 527976 181171 528170
rect 181205 528044 181239 528270
rect 181273 528256 181307 528272
rect 181273 528112 181307 528222
rect 181348 528256 181403 528384
rect 181348 528222 181369 528256
rect 181348 528214 181403 528222
rect 181381 528180 181403 528214
rect 181348 528152 181403 528180
rect 181437 528350 181475 528384
rect 181437 528316 181439 528350
rect 181473 528316 181475 528350
rect 181437 528143 181475 528316
rect 181511 528361 181613 528418
rect 181545 528327 181579 528361
rect 181511 528311 181613 528327
rect 181657 528361 181706 528377
rect 181657 528327 181663 528361
rect 181697 528327 181706 528361
rect 181657 528256 181706 528327
rect 181795 528357 182864 528418
rect 181795 528323 181813 528357
rect 181847 528323 182813 528357
rect 182847 528323 182864 528357
rect 181795 528309 182864 528323
rect 182899 528357 183968 528418
rect 182899 528323 182917 528357
rect 182951 528323 183917 528357
rect 183951 528323 183968 528357
rect 182899 528309 183968 528323
rect 184003 528357 185072 528418
rect 184003 528323 184021 528357
rect 184055 528323 185021 528357
rect 185055 528323 185072 528357
rect 184003 528309 185072 528323
rect 185107 528324 185165 528418
rect 181515 528222 181531 528256
rect 181565 528222 181761 528256
rect 181437 528112 181441 528143
rect 181273 528109 181441 528112
rect 181273 528078 181475 528109
rect 181509 528146 181659 528147
rect 181509 528112 181531 528146
rect 181565 528143 181659 528146
rect 181565 528112 181609 528143
rect 181509 528109 181609 528112
rect 181643 528109 181659 528143
rect 181205 528010 181305 528044
rect 181339 528010 181380 528044
rect 181414 528010 181430 528044
rect 181509 527976 181543 528109
rect 181693 528060 181761 528222
rect 182112 528194 182180 528309
rect 182112 528160 182129 528194
rect 182163 528160 182180 528194
rect 182112 528143 182180 528160
rect 182476 528230 182546 528245
rect 182476 528196 182493 528230
rect 182527 528196 182546 528230
rect 181137 527942 181543 527976
rect 181577 528044 181611 528060
rect 181577 527908 181611 528010
rect 181658 528044 181761 528060
rect 181658 528010 181663 528044
rect 181697 528010 181761 528044
rect 181658 527978 181761 528010
rect 182476 527995 182546 528196
rect 183216 528194 183284 528309
rect 183216 528160 183233 528194
rect 183267 528160 183284 528194
rect 183216 528143 183284 528160
rect 183580 528230 183650 528245
rect 183580 528196 183597 528230
rect 183631 528196 183650 528230
rect 183580 527995 183650 528196
rect 184320 528194 184388 528309
rect 185107 528290 185119 528324
rect 185153 528290 185165 528324
rect 185199 528357 186268 528418
rect 185199 528323 185217 528357
rect 185251 528323 186217 528357
rect 186251 528323 186268 528357
rect 185199 528309 186268 528323
rect 186303 528357 187005 528418
rect 186303 528323 186321 528357
rect 186355 528323 186953 528357
rect 186987 528323 187005 528357
rect 185107 528273 185165 528290
rect 184320 528160 184337 528194
rect 184371 528160 184388 528194
rect 184320 528143 184388 528160
rect 184684 528230 184754 528245
rect 184684 528196 184701 528230
rect 184735 528196 184754 528230
rect 184684 527995 184754 528196
rect 185516 528194 185584 528309
rect 186303 528264 187005 528323
rect 187223 528355 187465 528418
rect 187223 528321 187241 528355
rect 187275 528321 187413 528355
rect 187447 528321 187465 528355
rect 187223 528268 187465 528321
rect 185516 528160 185533 528194
rect 185567 528160 185584 528194
rect 185516 528143 185584 528160
rect 185880 528230 185950 528245
rect 185880 528196 185897 528230
rect 185931 528196 185950 528230
rect 185107 528106 185165 528141
rect 185107 528072 185119 528106
rect 185153 528072 185165 528106
rect 185107 528013 185165 528072
rect 181795 527984 182864 527995
rect 181795 527950 181813 527984
rect 181847 527950 182813 527984
rect 182847 527950 182864 527984
rect 181795 527908 182864 527950
rect 182899 527984 183968 527995
rect 182899 527950 182917 527984
rect 182951 527950 183917 527984
rect 183951 527950 183968 527984
rect 182899 527908 183968 527950
rect 184003 527984 185072 527995
rect 184003 527950 184021 527984
rect 184055 527950 185021 527984
rect 185055 527950 185072 527984
rect 184003 527908 185072 527950
rect 185107 527979 185119 528013
rect 185153 527979 185165 528013
rect 185880 527995 185950 528196
rect 186303 528194 186633 528264
rect 186303 528160 186381 528194
rect 186415 528160 186480 528194
rect 186514 528160 186579 528194
rect 186613 528160 186633 528194
rect 186667 528196 186687 528230
rect 186721 528196 186790 528230
rect 186824 528196 186893 528230
rect 186927 528196 187005 528230
rect 186667 528126 187005 528196
rect 186303 528086 187005 528126
rect 186303 528052 186321 528086
rect 186355 528052 186953 528086
rect 186987 528052 187005 528086
rect 185107 527908 185165 527979
rect 185199 527984 186268 527995
rect 185199 527950 185217 527984
rect 185251 527950 186217 527984
rect 186251 527950 186268 527984
rect 185199 527908 186268 527950
rect 186303 527984 187005 528052
rect 186303 527950 186321 527984
rect 186355 527950 186953 527984
rect 186987 527950 187005 527984
rect 186303 527908 187005 527950
rect 187223 528200 187273 528234
rect 187307 528200 187327 528234
rect 187223 528126 187327 528200
rect 187361 528194 187465 528268
rect 187361 528160 187381 528194
rect 187415 528160 187465 528194
rect 187223 528079 187465 528126
rect 187223 528045 187241 528079
rect 187275 528045 187413 528079
rect 187447 528045 187465 528079
rect 187223 527984 187465 528045
rect 187223 527950 187241 527984
rect 187275 527950 187413 527984
rect 187447 527950 187465 527984
rect 187223 527908 187465 527950
rect 172210 527874 172239 527908
rect 172273 527874 172331 527908
rect 172365 527874 172423 527908
rect 172457 527874 172515 527908
rect 172549 527874 172607 527908
rect 172641 527874 172699 527908
rect 172733 527874 172791 527908
rect 172825 527874 172883 527908
rect 172917 527874 172975 527908
rect 173009 527874 173067 527908
rect 173101 527874 173159 527908
rect 173193 527874 173251 527908
rect 173285 527874 173343 527908
rect 173377 527874 173435 527908
rect 173469 527874 173527 527908
rect 173561 527874 173619 527908
rect 173653 527874 173711 527908
rect 173745 527874 173803 527908
rect 173837 527874 173895 527908
rect 173929 527874 173987 527908
rect 174021 527874 174079 527908
rect 174113 527874 174171 527908
rect 174205 527874 174263 527908
rect 174297 527874 174355 527908
rect 174389 527874 174447 527908
rect 174481 527874 174539 527908
rect 174573 527874 174631 527908
rect 174665 527874 174723 527908
rect 174757 527874 174815 527908
rect 174849 527874 174907 527908
rect 174941 527874 174999 527908
rect 175033 527874 175091 527908
rect 175125 527874 175183 527908
rect 175217 527874 175275 527908
rect 175309 527874 175367 527908
rect 175401 527874 175459 527908
rect 175493 527874 175551 527908
rect 175585 527874 175643 527908
rect 175677 527874 175735 527908
rect 175769 527874 175827 527908
rect 175861 527874 175919 527908
rect 175953 527874 176011 527908
rect 176045 527874 176103 527908
rect 176137 527874 176195 527908
rect 176229 527874 176287 527908
rect 176321 527874 176379 527908
rect 176413 527874 176471 527908
rect 176505 527874 176563 527908
rect 176597 527874 176655 527908
rect 176689 527874 176747 527908
rect 176781 527874 176839 527908
rect 176873 527874 176931 527908
rect 176965 527874 177023 527908
rect 177057 527874 177115 527908
rect 177149 527874 177207 527908
rect 177241 527874 177299 527908
rect 177333 527874 177391 527908
rect 177425 527874 177483 527908
rect 177517 527874 177575 527908
rect 177609 527874 177667 527908
rect 177701 527874 177759 527908
rect 177793 527874 177851 527908
rect 177885 527874 177943 527908
rect 177977 527874 178035 527908
rect 178069 527874 178127 527908
rect 178161 527874 178219 527908
rect 178253 527874 178311 527908
rect 178345 527874 178403 527908
rect 178437 527874 178495 527908
rect 178529 527874 178587 527908
rect 178621 527874 178679 527908
rect 178713 527874 178771 527908
rect 178805 527874 178863 527908
rect 178897 527874 178955 527908
rect 178989 527874 179047 527908
rect 179081 527874 179139 527908
rect 179173 527874 179231 527908
rect 179265 527874 179323 527908
rect 179357 527874 179415 527908
rect 179449 527874 179507 527908
rect 179541 527874 179599 527908
rect 179633 527874 179691 527908
rect 179725 527874 179783 527908
rect 179817 527874 179875 527908
rect 179909 527874 179967 527908
rect 180001 527874 180059 527908
rect 180093 527874 180151 527908
rect 180185 527874 180243 527908
rect 180277 527874 180335 527908
rect 180369 527874 180427 527908
rect 180461 527874 180519 527908
rect 180553 527874 180611 527908
rect 180645 527874 180703 527908
rect 180737 527874 180795 527908
rect 180829 527874 180887 527908
rect 180921 527874 180979 527908
rect 181013 527874 181071 527908
rect 181105 527874 181163 527908
rect 181197 527874 181255 527908
rect 181289 527874 181347 527908
rect 181381 527874 181439 527908
rect 181473 527874 181531 527908
rect 181565 527874 181623 527908
rect 181657 527874 181715 527908
rect 181749 527874 181807 527908
rect 181841 527874 181899 527908
rect 181933 527874 181991 527908
rect 182025 527874 182083 527908
rect 182117 527874 182175 527908
rect 182209 527874 182267 527908
rect 182301 527874 182359 527908
rect 182393 527874 182451 527908
rect 182485 527874 182543 527908
rect 182577 527874 182635 527908
rect 182669 527874 182727 527908
rect 182761 527874 182819 527908
rect 182853 527874 182911 527908
rect 182945 527874 183003 527908
rect 183037 527874 183095 527908
rect 183129 527874 183187 527908
rect 183221 527874 183279 527908
rect 183313 527874 183371 527908
rect 183405 527874 183463 527908
rect 183497 527874 183555 527908
rect 183589 527874 183647 527908
rect 183681 527874 183739 527908
rect 183773 527874 183831 527908
rect 183865 527874 183923 527908
rect 183957 527874 184015 527908
rect 184049 527874 184107 527908
rect 184141 527874 184199 527908
rect 184233 527874 184291 527908
rect 184325 527874 184383 527908
rect 184417 527874 184475 527908
rect 184509 527874 184567 527908
rect 184601 527874 184659 527908
rect 184693 527874 184751 527908
rect 184785 527874 184843 527908
rect 184877 527874 184935 527908
rect 184969 527874 185027 527908
rect 185061 527874 185119 527908
rect 185153 527874 185211 527908
rect 185245 527874 185303 527908
rect 185337 527874 185395 527908
rect 185429 527874 185487 527908
rect 185521 527874 185579 527908
rect 185613 527874 185671 527908
rect 185705 527874 185763 527908
rect 185797 527874 185855 527908
rect 185889 527874 185947 527908
rect 185981 527874 186039 527908
rect 186073 527874 186131 527908
rect 186165 527874 186223 527908
rect 186257 527874 186315 527908
rect 186349 527874 186407 527908
rect 186441 527874 186499 527908
rect 186533 527874 186591 527908
rect 186625 527874 186683 527908
rect 186717 527874 186775 527908
rect 186809 527874 186867 527908
rect 186901 527874 186959 527908
rect 186993 527874 187051 527908
rect 187085 527874 187143 527908
rect 187177 527874 187235 527908
rect 187269 527874 187327 527908
rect 187361 527874 187419 527908
rect 187453 527874 187482 527908
rect 172227 527832 172469 527874
rect 172227 527798 172245 527832
rect 172279 527798 172417 527832
rect 172451 527798 172469 527832
rect 172227 527737 172469 527798
rect 172503 527832 173572 527874
rect 172503 527798 172521 527832
rect 172555 527798 173521 527832
rect 173555 527798 173572 527832
rect 172503 527787 173572 527798
rect 173607 527832 174676 527874
rect 173607 527798 173625 527832
rect 173659 527798 174625 527832
rect 174659 527798 174676 527832
rect 173607 527787 174676 527798
rect 174711 527832 175780 527874
rect 174711 527798 174729 527832
rect 174763 527798 175729 527832
rect 175763 527798 175780 527832
rect 174711 527787 175780 527798
rect 175815 527832 176333 527874
rect 175815 527798 175833 527832
rect 175867 527798 176281 527832
rect 176315 527798 176333 527832
rect 172227 527703 172245 527737
rect 172279 527703 172417 527737
rect 172451 527703 172469 527737
rect 172227 527656 172469 527703
rect 172227 527588 172277 527622
rect 172311 527588 172331 527622
rect 172227 527514 172331 527588
rect 172365 527582 172469 527656
rect 172365 527548 172385 527582
rect 172419 527548 172469 527582
rect 172820 527622 172888 527639
rect 172820 527588 172837 527622
rect 172871 527588 172888 527622
rect 172227 527461 172469 527514
rect 172820 527473 172888 527588
rect 173184 527586 173254 527787
rect 173184 527552 173201 527586
rect 173235 527552 173254 527586
rect 173184 527537 173254 527552
rect 173924 527622 173992 527639
rect 173924 527588 173941 527622
rect 173975 527588 173992 527622
rect 173924 527473 173992 527588
rect 174288 527586 174358 527787
rect 174288 527552 174305 527586
rect 174339 527552 174358 527586
rect 174288 527537 174358 527552
rect 175028 527622 175096 527639
rect 175028 527588 175045 527622
rect 175079 527588 175096 527622
rect 175028 527473 175096 527588
rect 175392 527586 175462 527787
rect 175815 527730 176333 527798
rect 175815 527696 175833 527730
rect 175867 527696 176281 527730
rect 176315 527696 176333 527730
rect 175815 527656 176333 527696
rect 175392 527552 175409 527586
rect 175443 527552 175462 527586
rect 175392 527537 175462 527552
rect 175815 527588 175893 527622
rect 175927 527588 176003 527622
rect 176037 527588 176057 527622
rect 175815 527518 176057 527588
rect 176091 527586 176333 527656
rect 176091 527552 176111 527586
rect 176145 527552 176221 527586
rect 176255 527552 176333 527586
rect 176367 527806 176444 527840
rect 176367 527772 176379 527806
rect 176438 527772 176444 527806
rect 176478 527832 176543 527874
rect 176478 527798 176494 527832
rect 176528 527798 176543 527832
rect 176478 527782 176543 527798
rect 176647 527806 176703 527840
rect 176367 527646 176444 527772
rect 176647 527772 176653 527806
rect 176687 527772 176703 527806
rect 176647 527748 176703 527772
rect 176478 527704 176703 527748
rect 176741 527806 176821 527840
rect 176741 527772 176757 527806
rect 176791 527772 176821 527806
rect 176901 527832 176955 527874
rect 176901 527798 176911 527832
rect 176945 527798 176955 527832
rect 176901 527782 176955 527798
rect 176989 527806 177046 527840
rect 172227 527427 172245 527461
rect 172279 527427 172417 527461
rect 172451 527427 172469 527461
rect 172227 527364 172469 527427
rect 172503 527459 173572 527473
rect 172503 527425 172521 527459
rect 172555 527425 173521 527459
rect 173555 527425 173572 527459
rect 172503 527364 173572 527425
rect 173607 527459 174676 527473
rect 173607 527425 173625 527459
rect 173659 527425 174625 527459
rect 174659 527425 174676 527459
rect 173607 527364 174676 527425
rect 174711 527459 175780 527473
rect 174711 527425 174729 527459
rect 174763 527425 175729 527459
rect 175763 527425 175780 527459
rect 174711 527364 175780 527425
rect 175815 527459 176333 527518
rect 175815 527425 175833 527459
rect 175867 527425 176281 527459
rect 176315 527425 176333 527459
rect 175815 527364 176333 527425
rect 176367 527512 176423 527646
rect 176478 527612 176568 527704
rect 176741 527670 176821 527772
rect 176989 527772 176995 527806
rect 177029 527772 177046 527806
rect 176989 527748 177046 527772
rect 176457 527596 176568 527612
rect 176491 527562 176568 527596
rect 176457 527546 176568 527562
rect 176602 527596 176821 527670
rect 176602 527562 176653 527596
rect 176687 527562 176821 527596
rect 176602 527558 176821 527562
rect 176478 527524 176568 527546
rect 176367 527466 176444 527512
rect 176478 527490 176703 527524
rect 176367 527432 176404 527466
rect 176438 527432 176444 527466
rect 176647 527466 176703 527490
rect 176367 527398 176444 527432
rect 176478 527440 176543 527456
rect 176478 527406 176494 527440
rect 176528 527406 176543 527440
rect 176478 527364 176543 527406
rect 176647 527432 176653 527466
rect 176687 527432 176703 527466
rect 176647 527398 176703 527432
rect 176741 527466 176821 527558
rect 176855 527704 177046 527748
rect 177103 527832 177345 527874
rect 177103 527798 177121 527832
rect 177155 527798 177293 527832
rect 177327 527798 177345 527832
rect 177103 527737 177345 527798
rect 176855 527596 176897 527704
rect 177103 527703 177121 527737
rect 177155 527703 177293 527737
rect 177327 527703 177345 527737
rect 176855 527562 176857 527596
rect 176891 527562 176897 527596
rect 176855 527524 176897 527562
rect 176931 527636 177023 527670
rect 177057 527636 177069 527670
rect 177103 527656 177345 527703
rect 176931 527596 177069 527636
rect 176931 527562 176971 527596
rect 177005 527562 177069 527596
rect 176931 527558 177069 527562
rect 177103 527588 177153 527622
rect 177187 527588 177207 527622
rect 176855 527490 177046 527524
rect 176741 527432 176757 527466
rect 176791 527432 176821 527466
rect 176989 527466 177046 527490
rect 176741 527398 176821 527432
rect 176901 527440 176955 527456
rect 176901 527406 176911 527440
rect 176945 527406 176955 527440
rect 176901 527364 176955 527406
rect 176989 527432 176995 527466
rect 177029 527432 177046 527466
rect 176989 527398 177046 527432
rect 177103 527514 177207 527588
rect 177241 527582 177345 527656
rect 177379 527803 177437 527874
rect 177379 527769 177391 527803
rect 177425 527769 177437 527803
rect 177471 527832 178540 527874
rect 177471 527798 177489 527832
rect 177523 527798 178489 527832
rect 178523 527798 178540 527832
rect 177471 527787 178540 527798
rect 178575 527832 178909 527874
rect 178575 527798 178593 527832
rect 178627 527798 178857 527832
rect 178891 527798 178909 527832
rect 177379 527710 177437 527769
rect 177379 527676 177391 527710
rect 177425 527676 177437 527710
rect 177379 527641 177437 527676
rect 177241 527548 177261 527582
rect 177295 527548 177345 527582
rect 177788 527622 177856 527639
rect 177788 527588 177805 527622
rect 177839 527588 177856 527622
rect 177103 527461 177345 527514
rect 177103 527427 177121 527461
rect 177155 527427 177293 527461
rect 177327 527427 177345 527461
rect 177103 527364 177345 527427
rect 177379 527492 177437 527509
rect 177379 527458 177391 527492
rect 177425 527458 177437 527492
rect 177788 527473 177856 527588
rect 178152 527586 178222 527787
rect 178575 527730 178909 527798
rect 178575 527696 178593 527730
rect 178627 527696 178857 527730
rect 178891 527696 178909 527730
rect 178575 527656 178909 527696
rect 178152 527552 178169 527586
rect 178203 527552 178222 527586
rect 178152 527537 178222 527552
rect 178575 527588 178595 527622
rect 178629 527588 178725 527622
rect 178575 527518 178725 527588
rect 178759 527586 178909 527656
rect 178759 527552 178855 527586
rect 178889 527552 178909 527586
rect 178943 527806 179020 527840
rect 178943 527772 178955 527806
rect 179014 527772 179020 527806
rect 179054 527832 179119 527874
rect 179054 527798 179070 527832
rect 179104 527798 179119 527832
rect 179054 527782 179119 527798
rect 179223 527806 179279 527840
rect 178943 527646 179020 527772
rect 179223 527772 179229 527806
rect 179263 527772 179279 527806
rect 179223 527748 179279 527772
rect 179054 527704 179279 527748
rect 179317 527806 179397 527840
rect 179317 527772 179333 527806
rect 179367 527772 179397 527806
rect 179477 527832 179531 527874
rect 179477 527798 179487 527832
rect 179521 527798 179531 527832
rect 179477 527782 179531 527798
rect 179565 527806 179622 527840
rect 177379 527364 177437 527458
rect 177471 527459 178540 527473
rect 177471 527425 177489 527459
rect 177523 527425 178489 527459
rect 178523 527425 178540 527459
rect 177471 527364 178540 527425
rect 178575 527466 178909 527518
rect 178575 527432 178593 527466
rect 178627 527432 178857 527466
rect 178891 527432 178909 527466
rect 178575 527364 178909 527432
rect 178943 527512 178999 527646
rect 179054 527612 179144 527704
rect 179317 527670 179397 527772
rect 179565 527772 179571 527806
rect 179605 527772 179622 527806
rect 179679 527832 180748 527874
rect 179679 527798 179697 527832
rect 179731 527798 180697 527832
rect 180731 527798 180748 527832
rect 179679 527787 180748 527798
rect 180783 527832 181852 527874
rect 180783 527798 180801 527832
rect 180835 527798 181801 527832
rect 181835 527798 181852 527832
rect 180783 527787 181852 527798
rect 181887 527832 182405 527874
rect 181887 527798 181905 527832
rect 181939 527798 182353 527832
rect 182387 527798 182405 527832
rect 179565 527748 179622 527772
rect 179033 527596 179144 527612
rect 179067 527562 179144 527596
rect 179033 527546 179144 527562
rect 179178 527596 179397 527670
rect 179178 527562 179229 527596
rect 179263 527562 179397 527596
rect 179178 527558 179397 527562
rect 179054 527524 179144 527546
rect 178943 527466 179020 527512
rect 179054 527490 179279 527524
rect 178943 527432 178980 527466
rect 179014 527432 179020 527466
rect 179223 527466 179279 527490
rect 178943 527398 179020 527432
rect 179054 527440 179119 527456
rect 179054 527406 179070 527440
rect 179104 527406 179119 527440
rect 179054 527364 179119 527406
rect 179223 527432 179229 527466
rect 179263 527432 179279 527466
rect 179223 527398 179279 527432
rect 179317 527466 179397 527558
rect 179431 527704 179622 527748
rect 179431 527596 179473 527704
rect 179431 527562 179433 527596
rect 179467 527562 179473 527596
rect 179431 527524 179473 527562
rect 179541 527636 179645 527670
rect 179507 527596 179645 527636
rect 179507 527562 179547 527596
rect 179581 527562 179645 527596
rect 179507 527558 179645 527562
rect 179996 527622 180064 527639
rect 179996 527588 180013 527622
rect 180047 527588 180064 527622
rect 179431 527490 179622 527524
rect 179317 527432 179333 527466
rect 179367 527432 179397 527466
rect 179565 527466 179622 527490
rect 179996 527473 180064 527588
rect 180360 527586 180430 527787
rect 180360 527552 180377 527586
rect 180411 527552 180430 527586
rect 180360 527537 180430 527552
rect 181100 527622 181168 527639
rect 181100 527588 181117 527622
rect 181151 527588 181168 527622
rect 181100 527473 181168 527588
rect 181464 527586 181534 527787
rect 181887 527730 182405 527798
rect 181887 527696 181905 527730
rect 181939 527696 182353 527730
rect 182387 527696 182405 527730
rect 181887 527656 182405 527696
rect 181464 527552 181481 527586
rect 181515 527552 181534 527586
rect 181464 527537 181534 527552
rect 181887 527588 181965 527622
rect 181999 527588 182075 527622
rect 182109 527588 182129 527622
rect 181887 527518 182129 527588
rect 182163 527586 182405 527656
rect 182531 527803 182589 527874
rect 182531 527769 182543 527803
rect 182577 527769 182589 527803
rect 182623 527832 183692 527874
rect 182623 527798 182641 527832
rect 182675 527798 183641 527832
rect 183675 527798 183692 527832
rect 182623 527787 183692 527798
rect 183727 527832 184796 527874
rect 183727 527798 183745 527832
rect 183779 527798 184745 527832
rect 184779 527798 184796 527832
rect 183727 527787 184796 527798
rect 184831 527832 185900 527874
rect 184831 527798 184849 527832
rect 184883 527798 185849 527832
rect 185883 527798 185900 527832
rect 184831 527787 185900 527798
rect 185935 527832 187004 527874
rect 185935 527798 185953 527832
rect 185987 527798 186953 527832
rect 186987 527798 187004 527832
rect 185935 527787 187004 527798
rect 187223 527832 187465 527874
rect 187223 527798 187241 527832
rect 187275 527798 187413 527832
rect 187447 527798 187465 527832
rect 182531 527710 182589 527769
rect 182531 527676 182543 527710
rect 182577 527676 182589 527710
rect 182531 527641 182589 527676
rect 182163 527552 182183 527586
rect 182217 527552 182293 527586
rect 182327 527552 182405 527586
rect 182940 527622 183008 527639
rect 182940 527588 182957 527622
rect 182991 527588 183008 527622
rect 179317 527398 179397 527432
rect 179477 527440 179531 527456
rect 179477 527406 179487 527440
rect 179521 527406 179531 527440
rect 179477 527364 179531 527406
rect 179565 527432 179571 527466
rect 179605 527432 179622 527466
rect 179565 527398 179622 527432
rect 179679 527459 180748 527473
rect 179679 527425 179697 527459
rect 179731 527425 180697 527459
rect 180731 527425 180748 527459
rect 179679 527364 180748 527425
rect 180783 527459 181852 527473
rect 180783 527425 180801 527459
rect 180835 527425 181801 527459
rect 181835 527425 181852 527459
rect 180783 527364 181852 527425
rect 181887 527459 182405 527518
rect 181887 527425 181905 527459
rect 181939 527425 182353 527459
rect 182387 527425 182405 527459
rect 181887 527364 182405 527425
rect 182531 527492 182589 527509
rect 182531 527458 182543 527492
rect 182577 527458 182589 527492
rect 182940 527473 183008 527588
rect 183304 527586 183374 527787
rect 183304 527552 183321 527586
rect 183355 527552 183374 527586
rect 183304 527537 183374 527552
rect 184044 527622 184112 527639
rect 184044 527588 184061 527622
rect 184095 527588 184112 527622
rect 184044 527473 184112 527588
rect 184408 527586 184478 527787
rect 184408 527552 184425 527586
rect 184459 527552 184478 527586
rect 184408 527537 184478 527552
rect 185148 527622 185216 527639
rect 185148 527588 185165 527622
rect 185199 527588 185216 527622
rect 185148 527473 185216 527588
rect 185512 527586 185582 527787
rect 185512 527552 185529 527586
rect 185563 527552 185582 527586
rect 185512 527537 185582 527552
rect 186252 527622 186320 527639
rect 186252 527588 186269 527622
rect 186303 527588 186320 527622
rect 186252 527473 186320 527588
rect 186616 527586 186686 527787
rect 186616 527552 186633 527586
rect 186667 527552 186686 527586
rect 186616 527537 186686 527552
rect 187223 527737 187465 527798
rect 187223 527703 187241 527737
rect 187275 527703 187413 527737
rect 187447 527703 187465 527737
rect 187223 527656 187465 527703
rect 187223 527582 187327 527656
rect 187223 527548 187273 527582
rect 187307 527548 187327 527582
rect 187361 527588 187381 527622
rect 187415 527588 187465 527622
rect 187361 527514 187465 527588
rect 182531 527364 182589 527458
rect 182623 527459 183692 527473
rect 182623 527425 182641 527459
rect 182675 527425 183641 527459
rect 183675 527425 183692 527459
rect 182623 527364 183692 527425
rect 183727 527459 184796 527473
rect 183727 527425 183745 527459
rect 183779 527425 184745 527459
rect 184779 527425 184796 527459
rect 183727 527364 184796 527425
rect 184831 527459 185900 527473
rect 184831 527425 184849 527459
rect 184883 527425 185849 527459
rect 185883 527425 185900 527459
rect 184831 527364 185900 527425
rect 185935 527459 187004 527473
rect 185935 527425 185953 527459
rect 185987 527425 186953 527459
rect 186987 527425 187004 527459
rect 185935 527364 187004 527425
rect 187223 527461 187465 527514
rect 187223 527427 187241 527461
rect 187275 527427 187413 527461
rect 187447 527427 187465 527461
rect 187223 527364 187465 527427
rect 172210 527330 172239 527364
rect 172273 527330 172331 527364
rect 172365 527330 172423 527364
rect 172457 527330 172515 527364
rect 172549 527330 172607 527364
rect 172641 527330 172699 527364
rect 172733 527330 172791 527364
rect 172825 527330 172883 527364
rect 172917 527330 172975 527364
rect 173009 527330 173067 527364
rect 173101 527330 173159 527364
rect 173193 527330 173251 527364
rect 173285 527330 173343 527364
rect 173377 527330 173435 527364
rect 173469 527330 173527 527364
rect 173561 527330 173619 527364
rect 173653 527330 173711 527364
rect 173745 527330 173803 527364
rect 173837 527330 173895 527364
rect 173929 527330 173987 527364
rect 174021 527330 174079 527364
rect 174113 527330 174171 527364
rect 174205 527330 174263 527364
rect 174297 527330 174355 527364
rect 174389 527330 174447 527364
rect 174481 527330 174539 527364
rect 174573 527330 174631 527364
rect 174665 527330 174723 527364
rect 174757 527330 174815 527364
rect 174849 527330 174907 527364
rect 174941 527330 174999 527364
rect 175033 527330 175091 527364
rect 175125 527330 175183 527364
rect 175217 527330 175275 527364
rect 175309 527330 175367 527364
rect 175401 527330 175459 527364
rect 175493 527330 175551 527364
rect 175585 527330 175643 527364
rect 175677 527330 175735 527364
rect 175769 527330 175827 527364
rect 175861 527330 175919 527364
rect 175953 527330 176011 527364
rect 176045 527330 176103 527364
rect 176137 527330 176195 527364
rect 176229 527330 176287 527364
rect 176321 527330 176379 527364
rect 176413 527330 176471 527364
rect 176505 527330 176563 527364
rect 176597 527330 176655 527364
rect 176689 527330 176747 527364
rect 176781 527330 176839 527364
rect 176873 527330 176931 527364
rect 176965 527330 177023 527364
rect 177057 527330 177115 527364
rect 177149 527330 177207 527364
rect 177241 527330 177299 527364
rect 177333 527330 177391 527364
rect 177425 527330 177483 527364
rect 177517 527330 177575 527364
rect 177609 527330 177667 527364
rect 177701 527330 177759 527364
rect 177793 527330 177851 527364
rect 177885 527330 177943 527364
rect 177977 527330 178035 527364
rect 178069 527330 178127 527364
rect 178161 527330 178219 527364
rect 178253 527330 178311 527364
rect 178345 527330 178403 527364
rect 178437 527330 178495 527364
rect 178529 527330 178587 527364
rect 178621 527330 178679 527364
rect 178713 527330 178771 527364
rect 178805 527330 178863 527364
rect 178897 527330 178955 527364
rect 178989 527330 179047 527364
rect 179081 527330 179139 527364
rect 179173 527330 179231 527364
rect 179265 527330 179323 527364
rect 179357 527330 179415 527364
rect 179449 527330 179507 527364
rect 179541 527330 179599 527364
rect 179633 527330 179691 527364
rect 179725 527330 179783 527364
rect 179817 527330 179875 527364
rect 179909 527330 179967 527364
rect 180001 527330 180059 527364
rect 180093 527330 180151 527364
rect 180185 527330 180243 527364
rect 180277 527330 180335 527364
rect 180369 527330 180427 527364
rect 180461 527330 180519 527364
rect 180553 527330 180611 527364
rect 180645 527330 180703 527364
rect 180737 527330 180795 527364
rect 180829 527330 180887 527364
rect 180921 527330 180979 527364
rect 181013 527330 181071 527364
rect 181105 527330 181163 527364
rect 181197 527330 181255 527364
rect 181289 527330 181347 527364
rect 181381 527330 181439 527364
rect 181473 527330 181531 527364
rect 181565 527330 181623 527364
rect 181657 527330 181715 527364
rect 181749 527330 181807 527364
rect 181841 527330 181899 527364
rect 181933 527330 181991 527364
rect 182025 527330 182083 527364
rect 182117 527330 182175 527364
rect 182209 527330 182267 527364
rect 182301 527330 182359 527364
rect 182393 527330 182451 527364
rect 182485 527330 182543 527364
rect 182577 527330 182635 527364
rect 182669 527330 182727 527364
rect 182761 527330 182819 527364
rect 182853 527330 182911 527364
rect 182945 527330 183003 527364
rect 183037 527330 183095 527364
rect 183129 527330 183187 527364
rect 183221 527330 183279 527364
rect 183313 527330 183371 527364
rect 183405 527330 183463 527364
rect 183497 527330 183555 527364
rect 183589 527330 183647 527364
rect 183681 527330 183739 527364
rect 183773 527330 183831 527364
rect 183865 527330 183923 527364
rect 183957 527330 184015 527364
rect 184049 527330 184107 527364
rect 184141 527330 184199 527364
rect 184233 527330 184291 527364
rect 184325 527330 184383 527364
rect 184417 527330 184475 527364
rect 184509 527330 184567 527364
rect 184601 527330 184659 527364
rect 184693 527330 184751 527364
rect 184785 527330 184843 527364
rect 184877 527330 184935 527364
rect 184969 527330 185027 527364
rect 185061 527330 185119 527364
rect 185153 527330 185211 527364
rect 185245 527330 185303 527364
rect 185337 527330 185395 527364
rect 185429 527330 185487 527364
rect 185521 527330 185579 527364
rect 185613 527330 185671 527364
rect 185705 527330 185763 527364
rect 185797 527330 185855 527364
rect 185889 527330 185947 527364
rect 185981 527330 186039 527364
rect 186073 527330 186131 527364
rect 186165 527330 186223 527364
rect 186257 527330 186315 527364
rect 186349 527330 186407 527364
rect 186441 527330 186499 527364
rect 186533 527330 186591 527364
rect 186625 527330 186683 527364
rect 186717 527330 186775 527364
rect 186809 527330 186867 527364
rect 186901 527330 186959 527364
rect 186993 527330 187051 527364
rect 187085 527330 187143 527364
rect 187177 527330 187235 527364
rect 187269 527330 187327 527364
rect 187361 527330 187419 527364
rect 187453 527330 187482 527364
rect 172227 527267 172469 527330
rect 172227 527233 172245 527267
rect 172279 527233 172417 527267
rect 172451 527233 172469 527267
rect 172227 527180 172469 527233
rect 172503 527269 173572 527330
rect 172503 527235 172521 527269
rect 172555 527235 173521 527269
rect 173555 527235 173572 527269
rect 172503 527221 173572 527235
rect 173607 527269 174676 527330
rect 173607 527235 173625 527269
rect 173659 527235 174625 527269
rect 174659 527235 174676 527269
rect 173607 527221 174676 527235
rect 174803 527236 174861 527330
rect 172227 527106 172331 527180
rect 172227 527072 172277 527106
rect 172311 527072 172331 527106
rect 172365 527112 172385 527146
rect 172419 527112 172469 527146
rect 172365 527038 172469 527112
rect 172820 527106 172888 527221
rect 172820 527072 172837 527106
rect 172871 527072 172888 527106
rect 172820 527055 172888 527072
rect 173184 527142 173254 527157
rect 173184 527108 173201 527142
rect 173235 527108 173254 527142
rect 172227 526991 172469 527038
rect 172227 526957 172245 526991
rect 172279 526957 172417 526991
rect 172451 526957 172469 526991
rect 172227 526896 172469 526957
rect 173184 526907 173254 527108
rect 173924 527106 173992 527221
rect 174803 527202 174815 527236
rect 174849 527202 174861 527236
rect 174895 527269 175964 527330
rect 174895 527235 174913 527269
rect 174947 527235 175913 527269
rect 175947 527235 175964 527269
rect 174895 527221 175964 527235
rect 175999 527269 177068 527330
rect 175999 527235 176017 527269
rect 176051 527235 177017 527269
rect 177051 527235 177068 527269
rect 175999 527221 177068 527235
rect 177103 527269 178172 527330
rect 177103 527235 177121 527269
rect 177155 527235 178121 527269
rect 178155 527235 178172 527269
rect 177103 527221 178172 527235
rect 178207 527269 179276 527330
rect 178207 527235 178225 527269
rect 178259 527235 179225 527269
rect 179259 527235 179276 527269
rect 178207 527221 179276 527235
rect 179311 527269 179829 527330
rect 179311 527235 179329 527269
rect 179363 527235 179777 527269
rect 179811 527235 179829 527269
rect 174803 527185 174861 527202
rect 173924 527072 173941 527106
rect 173975 527072 173992 527106
rect 173924 527055 173992 527072
rect 174288 527142 174358 527157
rect 174288 527108 174305 527142
rect 174339 527108 174358 527142
rect 174288 526907 174358 527108
rect 175212 527106 175280 527221
rect 175212 527072 175229 527106
rect 175263 527072 175280 527106
rect 175212 527055 175280 527072
rect 175576 527142 175646 527157
rect 175576 527108 175593 527142
rect 175627 527108 175646 527142
rect 174803 527018 174861 527053
rect 174803 526984 174815 527018
rect 174849 526984 174861 527018
rect 174803 526925 174861 526984
rect 172227 526862 172245 526896
rect 172279 526862 172417 526896
rect 172451 526862 172469 526896
rect 172227 526820 172469 526862
rect 172503 526896 173572 526907
rect 172503 526862 172521 526896
rect 172555 526862 173521 526896
rect 173555 526862 173572 526896
rect 172503 526820 173572 526862
rect 173607 526896 174676 526907
rect 173607 526862 173625 526896
rect 173659 526862 174625 526896
rect 174659 526862 174676 526896
rect 173607 526820 174676 526862
rect 174803 526891 174815 526925
rect 174849 526891 174861 526925
rect 175576 526907 175646 527108
rect 176316 527106 176384 527221
rect 176316 527072 176333 527106
rect 176367 527072 176384 527106
rect 176316 527055 176384 527072
rect 176680 527142 176750 527157
rect 176680 527108 176697 527142
rect 176731 527108 176750 527142
rect 176680 526907 176750 527108
rect 177420 527106 177488 527221
rect 177420 527072 177437 527106
rect 177471 527072 177488 527106
rect 177420 527055 177488 527072
rect 177784 527142 177854 527157
rect 177784 527108 177801 527142
rect 177835 527108 177854 527142
rect 177784 526907 177854 527108
rect 178524 527106 178592 527221
rect 179311 527176 179829 527235
rect 179955 527236 180013 527330
rect 179955 527202 179967 527236
rect 180001 527202 180013 527236
rect 180047 527269 181116 527330
rect 180047 527235 180065 527269
rect 180099 527235 181065 527269
rect 181099 527235 181116 527269
rect 180047 527221 181116 527235
rect 181151 527269 182220 527330
rect 181151 527235 181169 527269
rect 181203 527235 182169 527269
rect 182203 527235 182220 527269
rect 181151 527221 182220 527235
rect 182255 527269 183324 527330
rect 182255 527235 182273 527269
rect 182307 527235 183273 527269
rect 183307 527235 183324 527269
rect 182255 527221 183324 527235
rect 183359 527269 184428 527330
rect 183359 527235 183377 527269
rect 183411 527235 184377 527269
rect 184411 527235 184428 527269
rect 183359 527221 184428 527235
rect 184463 527269 184981 527330
rect 184463 527235 184481 527269
rect 184515 527235 184929 527269
rect 184963 527235 184981 527269
rect 179955 527185 180013 527202
rect 178524 527072 178541 527106
rect 178575 527072 178592 527106
rect 178524 527055 178592 527072
rect 178888 527142 178958 527157
rect 178888 527108 178905 527142
rect 178939 527108 178958 527142
rect 178888 526907 178958 527108
rect 179311 527106 179553 527176
rect 179311 527072 179389 527106
rect 179423 527072 179499 527106
rect 179533 527072 179553 527106
rect 179587 527108 179607 527142
rect 179641 527108 179717 527142
rect 179751 527108 179829 527142
rect 179587 527038 179829 527108
rect 180364 527106 180432 527221
rect 180364 527072 180381 527106
rect 180415 527072 180432 527106
rect 180364 527055 180432 527072
rect 180728 527142 180798 527157
rect 180728 527108 180745 527142
rect 180779 527108 180798 527142
rect 179311 526998 179829 527038
rect 179311 526964 179329 526998
rect 179363 526964 179777 526998
rect 179811 526964 179829 526998
rect 174803 526820 174861 526891
rect 174895 526896 175964 526907
rect 174895 526862 174913 526896
rect 174947 526862 175913 526896
rect 175947 526862 175964 526896
rect 174895 526820 175964 526862
rect 175999 526896 177068 526907
rect 175999 526862 176017 526896
rect 176051 526862 177017 526896
rect 177051 526862 177068 526896
rect 175999 526820 177068 526862
rect 177103 526896 178172 526907
rect 177103 526862 177121 526896
rect 177155 526862 178121 526896
rect 178155 526862 178172 526896
rect 177103 526820 178172 526862
rect 178207 526896 179276 526907
rect 178207 526862 178225 526896
rect 178259 526862 179225 526896
rect 179259 526862 179276 526896
rect 178207 526820 179276 526862
rect 179311 526896 179829 526964
rect 179311 526862 179329 526896
rect 179363 526862 179777 526896
rect 179811 526862 179829 526896
rect 179311 526820 179829 526862
rect 179955 527018 180013 527053
rect 179955 526984 179967 527018
rect 180001 526984 180013 527018
rect 179955 526925 180013 526984
rect 179955 526891 179967 526925
rect 180001 526891 180013 526925
rect 180728 526907 180798 527108
rect 181468 527106 181536 527221
rect 181468 527072 181485 527106
rect 181519 527072 181536 527106
rect 181468 527055 181536 527072
rect 181832 527142 181902 527157
rect 181832 527108 181849 527142
rect 181883 527108 181902 527142
rect 181832 526907 181902 527108
rect 182572 527106 182640 527221
rect 182572 527072 182589 527106
rect 182623 527072 182640 527106
rect 182572 527055 182640 527072
rect 182936 527142 183006 527157
rect 182936 527108 182953 527142
rect 182987 527108 183006 527142
rect 182936 526907 183006 527108
rect 183676 527106 183744 527221
rect 184463 527176 184981 527235
rect 185107 527236 185165 527330
rect 185107 527202 185119 527236
rect 185153 527202 185165 527236
rect 185199 527269 186268 527330
rect 185199 527235 185217 527269
rect 185251 527235 186217 527269
rect 186251 527235 186268 527269
rect 185199 527221 186268 527235
rect 186303 527269 187005 527330
rect 186303 527235 186321 527269
rect 186355 527235 186953 527269
rect 186987 527235 187005 527269
rect 185107 527185 185165 527202
rect 183676 527072 183693 527106
rect 183727 527072 183744 527106
rect 183676 527055 183744 527072
rect 184040 527142 184110 527157
rect 184040 527108 184057 527142
rect 184091 527108 184110 527142
rect 184040 526907 184110 527108
rect 184463 527106 184705 527176
rect 184463 527072 184541 527106
rect 184575 527072 184651 527106
rect 184685 527072 184705 527106
rect 184739 527108 184759 527142
rect 184793 527108 184869 527142
rect 184903 527108 184981 527142
rect 184739 527038 184981 527108
rect 185516 527106 185584 527221
rect 186303 527176 187005 527235
rect 187223 527267 187465 527330
rect 187223 527233 187241 527267
rect 187275 527233 187413 527267
rect 187447 527233 187465 527267
rect 187223 527180 187465 527233
rect 185516 527072 185533 527106
rect 185567 527072 185584 527106
rect 185516 527055 185584 527072
rect 185880 527142 185950 527157
rect 185880 527108 185897 527142
rect 185931 527108 185950 527142
rect 184463 526998 184981 527038
rect 184463 526964 184481 526998
rect 184515 526964 184929 526998
rect 184963 526964 184981 526998
rect 179955 526820 180013 526891
rect 180047 526896 181116 526907
rect 180047 526862 180065 526896
rect 180099 526862 181065 526896
rect 181099 526862 181116 526896
rect 180047 526820 181116 526862
rect 181151 526896 182220 526907
rect 181151 526862 181169 526896
rect 181203 526862 182169 526896
rect 182203 526862 182220 526896
rect 181151 526820 182220 526862
rect 182255 526896 183324 526907
rect 182255 526862 182273 526896
rect 182307 526862 183273 526896
rect 183307 526862 183324 526896
rect 182255 526820 183324 526862
rect 183359 526896 184428 526907
rect 183359 526862 183377 526896
rect 183411 526862 184377 526896
rect 184411 526862 184428 526896
rect 183359 526820 184428 526862
rect 184463 526896 184981 526964
rect 184463 526862 184481 526896
rect 184515 526862 184929 526896
rect 184963 526862 184981 526896
rect 184463 526820 184981 526862
rect 185107 527018 185165 527053
rect 185107 526984 185119 527018
rect 185153 526984 185165 527018
rect 185107 526925 185165 526984
rect 185107 526891 185119 526925
rect 185153 526891 185165 526925
rect 185880 526907 185950 527108
rect 186303 527106 186633 527176
rect 186303 527072 186381 527106
rect 186415 527072 186480 527106
rect 186514 527072 186579 527106
rect 186613 527072 186633 527106
rect 186667 527108 186687 527142
rect 186721 527108 186790 527142
rect 186824 527108 186893 527142
rect 186927 527108 187005 527142
rect 186667 527038 187005 527108
rect 186303 526998 187005 527038
rect 186303 526964 186321 526998
rect 186355 526964 186953 526998
rect 186987 526964 187005 526998
rect 185107 526820 185165 526891
rect 185199 526896 186268 526907
rect 185199 526862 185217 526896
rect 185251 526862 186217 526896
rect 186251 526862 186268 526896
rect 185199 526820 186268 526862
rect 186303 526896 187005 526964
rect 186303 526862 186321 526896
rect 186355 526862 186953 526896
rect 186987 526862 187005 526896
rect 186303 526820 187005 526862
rect 187223 527112 187273 527146
rect 187307 527112 187327 527146
rect 187223 527038 187327 527112
rect 187361 527106 187465 527180
rect 187361 527072 187381 527106
rect 187415 527072 187465 527106
rect 187223 526991 187465 527038
rect 187223 526957 187241 526991
rect 187275 526957 187413 526991
rect 187447 526957 187465 526991
rect 187223 526896 187465 526957
rect 187223 526862 187241 526896
rect 187275 526862 187413 526896
rect 187447 526862 187465 526896
rect 187223 526820 187465 526862
rect 172210 526786 172239 526820
rect 172273 526786 172331 526820
rect 172365 526786 172423 526820
rect 172457 526786 172515 526820
rect 172549 526786 172607 526820
rect 172641 526786 172699 526820
rect 172733 526786 172791 526820
rect 172825 526786 172883 526820
rect 172917 526786 172975 526820
rect 173009 526786 173067 526820
rect 173101 526786 173159 526820
rect 173193 526786 173251 526820
rect 173285 526786 173343 526820
rect 173377 526786 173435 526820
rect 173469 526786 173527 526820
rect 173561 526786 173619 526820
rect 173653 526786 173711 526820
rect 173745 526786 173803 526820
rect 173837 526786 173895 526820
rect 173929 526786 173987 526820
rect 174021 526786 174079 526820
rect 174113 526786 174171 526820
rect 174205 526786 174263 526820
rect 174297 526786 174355 526820
rect 174389 526786 174447 526820
rect 174481 526786 174539 526820
rect 174573 526786 174631 526820
rect 174665 526786 174723 526820
rect 174757 526786 174815 526820
rect 174849 526786 174907 526820
rect 174941 526786 174999 526820
rect 175033 526786 175091 526820
rect 175125 526786 175183 526820
rect 175217 526786 175275 526820
rect 175309 526786 175367 526820
rect 175401 526786 175459 526820
rect 175493 526786 175551 526820
rect 175585 526786 175643 526820
rect 175677 526786 175735 526820
rect 175769 526786 175827 526820
rect 175861 526786 175919 526820
rect 175953 526786 176011 526820
rect 176045 526786 176103 526820
rect 176137 526786 176195 526820
rect 176229 526786 176287 526820
rect 176321 526786 176379 526820
rect 176413 526786 176471 526820
rect 176505 526786 176563 526820
rect 176597 526786 176655 526820
rect 176689 526786 176747 526820
rect 176781 526786 176839 526820
rect 176873 526786 176931 526820
rect 176965 526786 177023 526820
rect 177057 526786 177115 526820
rect 177149 526786 177207 526820
rect 177241 526786 177299 526820
rect 177333 526786 177391 526820
rect 177425 526786 177483 526820
rect 177517 526786 177575 526820
rect 177609 526786 177667 526820
rect 177701 526786 177759 526820
rect 177793 526786 177851 526820
rect 177885 526786 177943 526820
rect 177977 526786 178035 526820
rect 178069 526786 178127 526820
rect 178161 526786 178219 526820
rect 178253 526786 178311 526820
rect 178345 526786 178403 526820
rect 178437 526786 178495 526820
rect 178529 526786 178587 526820
rect 178621 526786 178679 526820
rect 178713 526786 178771 526820
rect 178805 526786 178863 526820
rect 178897 526786 178955 526820
rect 178989 526786 179047 526820
rect 179081 526786 179139 526820
rect 179173 526786 179231 526820
rect 179265 526786 179323 526820
rect 179357 526786 179415 526820
rect 179449 526786 179507 526820
rect 179541 526786 179599 526820
rect 179633 526786 179691 526820
rect 179725 526786 179783 526820
rect 179817 526786 179875 526820
rect 179909 526786 179967 526820
rect 180001 526786 180059 526820
rect 180093 526786 180151 526820
rect 180185 526786 180243 526820
rect 180277 526786 180335 526820
rect 180369 526786 180427 526820
rect 180461 526786 180519 526820
rect 180553 526786 180611 526820
rect 180645 526786 180703 526820
rect 180737 526786 180795 526820
rect 180829 526786 180887 526820
rect 180921 526786 180979 526820
rect 181013 526786 181071 526820
rect 181105 526786 181163 526820
rect 181197 526786 181255 526820
rect 181289 526786 181347 526820
rect 181381 526786 181439 526820
rect 181473 526786 181531 526820
rect 181565 526786 181623 526820
rect 181657 526786 181715 526820
rect 181749 526786 181807 526820
rect 181841 526786 181899 526820
rect 181933 526786 181991 526820
rect 182025 526786 182083 526820
rect 182117 526786 182175 526820
rect 182209 526786 182267 526820
rect 182301 526786 182359 526820
rect 182393 526786 182451 526820
rect 182485 526786 182543 526820
rect 182577 526786 182635 526820
rect 182669 526786 182727 526820
rect 182761 526786 182819 526820
rect 182853 526786 182911 526820
rect 182945 526786 183003 526820
rect 183037 526786 183095 526820
rect 183129 526786 183187 526820
rect 183221 526786 183279 526820
rect 183313 526786 183371 526820
rect 183405 526786 183463 526820
rect 183497 526786 183555 526820
rect 183589 526786 183647 526820
rect 183681 526786 183739 526820
rect 183773 526786 183831 526820
rect 183865 526786 183923 526820
rect 183957 526786 184015 526820
rect 184049 526786 184107 526820
rect 184141 526786 184199 526820
rect 184233 526786 184291 526820
rect 184325 526786 184383 526820
rect 184417 526786 184475 526820
rect 184509 526786 184567 526820
rect 184601 526786 184659 526820
rect 184693 526786 184751 526820
rect 184785 526786 184843 526820
rect 184877 526786 184935 526820
rect 184969 526786 185027 526820
rect 185061 526786 185119 526820
rect 185153 526786 185211 526820
rect 185245 526786 185303 526820
rect 185337 526786 185395 526820
rect 185429 526786 185487 526820
rect 185521 526786 185579 526820
rect 185613 526786 185671 526820
rect 185705 526786 185763 526820
rect 185797 526786 185855 526820
rect 185889 526786 185947 526820
rect 185981 526786 186039 526820
rect 186073 526786 186131 526820
rect 186165 526786 186223 526820
rect 186257 526786 186315 526820
rect 186349 526786 186407 526820
rect 186441 526786 186499 526820
rect 186533 526786 186591 526820
rect 186625 526786 186683 526820
rect 186717 526786 186775 526820
rect 186809 526786 186867 526820
rect 186901 526786 186959 526820
rect 186993 526786 187051 526820
rect 187085 526786 187143 526820
rect 187177 526786 187235 526820
rect 187269 526786 187327 526820
rect 187361 526786 187419 526820
rect 187453 526786 187482 526820
rect 172227 526744 172469 526786
rect 172227 526710 172245 526744
rect 172279 526710 172417 526744
rect 172451 526710 172469 526744
rect 172227 526649 172469 526710
rect 172503 526744 173572 526786
rect 172503 526710 172521 526744
rect 172555 526710 173521 526744
rect 173555 526710 173572 526744
rect 172503 526699 173572 526710
rect 173607 526744 174676 526786
rect 173607 526710 173625 526744
rect 173659 526710 174625 526744
rect 174659 526710 174676 526744
rect 173607 526699 174676 526710
rect 174711 526744 175780 526786
rect 174711 526710 174729 526744
rect 174763 526710 175729 526744
rect 175763 526710 175780 526744
rect 174711 526699 175780 526710
rect 175815 526744 176884 526786
rect 175815 526710 175833 526744
rect 175867 526710 176833 526744
rect 176867 526710 176884 526744
rect 175815 526699 176884 526710
rect 176919 526744 177253 526786
rect 176919 526710 176937 526744
rect 176971 526710 177201 526744
rect 177235 526710 177253 526744
rect 172227 526615 172245 526649
rect 172279 526615 172417 526649
rect 172451 526615 172469 526649
rect 172227 526568 172469 526615
rect 172227 526500 172277 526534
rect 172311 526500 172331 526534
rect 172227 526426 172331 526500
rect 172365 526494 172469 526568
rect 172365 526460 172385 526494
rect 172419 526460 172469 526494
rect 172820 526534 172888 526551
rect 172820 526500 172837 526534
rect 172871 526500 172888 526534
rect 172227 526373 172469 526426
rect 172820 526385 172888 526500
rect 173184 526498 173254 526699
rect 173184 526464 173201 526498
rect 173235 526464 173254 526498
rect 173184 526449 173254 526464
rect 173924 526534 173992 526551
rect 173924 526500 173941 526534
rect 173975 526500 173992 526534
rect 173924 526385 173992 526500
rect 174288 526498 174358 526699
rect 174288 526464 174305 526498
rect 174339 526464 174358 526498
rect 174288 526449 174358 526464
rect 175028 526534 175096 526551
rect 175028 526500 175045 526534
rect 175079 526500 175096 526534
rect 175028 526385 175096 526500
rect 175392 526498 175462 526699
rect 175392 526464 175409 526498
rect 175443 526464 175462 526498
rect 175392 526449 175462 526464
rect 176132 526534 176200 526551
rect 176132 526500 176149 526534
rect 176183 526500 176200 526534
rect 176132 526385 176200 526500
rect 176496 526498 176566 526699
rect 176919 526642 177253 526710
rect 176919 526608 176937 526642
rect 176971 526608 177201 526642
rect 177235 526608 177253 526642
rect 176919 526568 177253 526608
rect 176496 526464 176513 526498
rect 176547 526464 176566 526498
rect 176496 526449 176566 526464
rect 176919 526500 176939 526534
rect 176973 526500 177069 526534
rect 176919 526430 177069 526500
rect 177103 526498 177253 526568
rect 177379 526715 177437 526786
rect 177379 526681 177391 526715
rect 177425 526681 177437 526715
rect 177471 526744 178540 526786
rect 177471 526710 177489 526744
rect 177523 526710 178489 526744
rect 178523 526710 178540 526744
rect 177471 526699 178540 526710
rect 178575 526744 179644 526786
rect 178575 526710 178593 526744
rect 178627 526710 179593 526744
rect 179627 526710 179644 526744
rect 178575 526699 179644 526710
rect 179679 526744 180748 526786
rect 179679 526710 179697 526744
rect 179731 526710 180697 526744
rect 180731 526710 180748 526744
rect 179679 526699 180748 526710
rect 180783 526744 181852 526786
rect 180783 526710 180801 526744
rect 180835 526710 181801 526744
rect 181835 526710 181852 526744
rect 180783 526699 181852 526710
rect 181887 526744 182405 526786
rect 181887 526710 181905 526744
rect 181939 526710 182353 526744
rect 182387 526710 182405 526744
rect 177379 526622 177437 526681
rect 177379 526588 177391 526622
rect 177425 526588 177437 526622
rect 177379 526553 177437 526588
rect 177103 526464 177199 526498
rect 177233 526464 177253 526498
rect 177788 526534 177856 526551
rect 177788 526500 177805 526534
rect 177839 526500 177856 526534
rect 172227 526339 172245 526373
rect 172279 526339 172417 526373
rect 172451 526339 172469 526373
rect 172227 526276 172469 526339
rect 172503 526371 173572 526385
rect 172503 526337 172521 526371
rect 172555 526337 173521 526371
rect 173555 526337 173572 526371
rect 172503 526276 173572 526337
rect 173607 526371 174676 526385
rect 173607 526337 173625 526371
rect 173659 526337 174625 526371
rect 174659 526337 174676 526371
rect 173607 526276 174676 526337
rect 174711 526371 175780 526385
rect 174711 526337 174729 526371
rect 174763 526337 175729 526371
rect 175763 526337 175780 526371
rect 174711 526276 175780 526337
rect 175815 526371 176884 526385
rect 175815 526337 175833 526371
rect 175867 526337 176833 526371
rect 176867 526337 176884 526371
rect 175815 526276 176884 526337
rect 176919 526378 177253 526430
rect 176919 526344 176937 526378
rect 176971 526344 177201 526378
rect 177235 526344 177253 526378
rect 176919 526276 177253 526344
rect 177379 526404 177437 526421
rect 177379 526370 177391 526404
rect 177425 526370 177437 526404
rect 177788 526385 177856 526500
rect 178152 526498 178222 526699
rect 178152 526464 178169 526498
rect 178203 526464 178222 526498
rect 178152 526449 178222 526464
rect 178892 526534 178960 526551
rect 178892 526500 178909 526534
rect 178943 526500 178960 526534
rect 178892 526385 178960 526500
rect 179256 526498 179326 526699
rect 179256 526464 179273 526498
rect 179307 526464 179326 526498
rect 179256 526449 179326 526464
rect 179996 526534 180064 526551
rect 179996 526500 180013 526534
rect 180047 526500 180064 526534
rect 179996 526385 180064 526500
rect 180360 526498 180430 526699
rect 180360 526464 180377 526498
rect 180411 526464 180430 526498
rect 180360 526449 180430 526464
rect 181100 526534 181168 526551
rect 181100 526500 181117 526534
rect 181151 526500 181168 526534
rect 181100 526385 181168 526500
rect 181464 526498 181534 526699
rect 181887 526642 182405 526710
rect 181887 526608 181905 526642
rect 181939 526608 182353 526642
rect 182387 526608 182405 526642
rect 181887 526568 182405 526608
rect 181464 526464 181481 526498
rect 181515 526464 181534 526498
rect 181464 526449 181534 526464
rect 181887 526500 181965 526534
rect 181999 526500 182075 526534
rect 182109 526500 182129 526534
rect 181887 526430 182129 526500
rect 182163 526498 182405 526568
rect 182531 526715 182589 526786
rect 182531 526681 182543 526715
rect 182577 526681 182589 526715
rect 182623 526744 183692 526786
rect 182623 526710 182641 526744
rect 182675 526710 183641 526744
rect 183675 526710 183692 526744
rect 182623 526699 183692 526710
rect 183727 526744 184796 526786
rect 183727 526710 183745 526744
rect 183779 526710 184745 526744
rect 184779 526710 184796 526744
rect 183727 526699 184796 526710
rect 184831 526744 185900 526786
rect 184831 526710 184849 526744
rect 184883 526710 185849 526744
rect 185883 526710 185900 526744
rect 184831 526699 185900 526710
rect 185935 526744 187004 526786
rect 185935 526710 185953 526744
rect 185987 526710 186953 526744
rect 186987 526710 187004 526744
rect 185935 526699 187004 526710
rect 187223 526744 187465 526786
rect 187223 526710 187241 526744
rect 187275 526710 187413 526744
rect 187447 526710 187465 526744
rect 182531 526622 182589 526681
rect 182531 526588 182543 526622
rect 182577 526588 182589 526622
rect 182531 526553 182589 526588
rect 182163 526464 182183 526498
rect 182217 526464 182293 526498
rect 182327 526464 182405 526498
rect 182940 526534 183008 526551
rect 182940 526500 182957 526534
rect 182991 526500 183008 526534
rect 177379 526276 177437 526370
rect 177471 526371 178540 526385
rect 177471 526337 177489 526371
rect 177523 526337 178489 526371
rect 178523 526337 178540 526371
rect 177471 526276 178540 526337
rect 178575 526371 179644 526385
rect 178575 526337 178593 526371
rect 178627 526337 179593 526371
rect 179627 526337 179644 526371
rect 178575 526276 179644 526337
rect 179679 526371 180748 526385
rect 179679 526337 179697 526371
rect 179731 526337 180697 526371
rect 180731 526337 180748 526371
rect 179679 526276 180748 526337
rect 180783 526371 181852 526385
rect 180783 526337 180801 526371
rect 180835 526337 181801 526371
rect 181835 526337 181852 526371
rect 180783 526276 181852 526337
rect 181887 526371 182405 526430
rect 181887 526337 181905 526371
rect 181939 526337 182353 526371
rect 182387 526337 182405 526371
rect 181887 526276 182405 526337
rect 182531 526404 182589 526421
rect 182531 526370 182543 526404
rect 182577 526370 182589 526404
rect 182940 526385 183008 526500
rect 183304 526498 183374 526699
rect 183304 526464 183321 526498
rect 183355 526464 183374 526498
rect 183304 526449 183374 526464
rect 184044 526534 184112 526551
rect 184044 526500 184061 526534
rect 184095 526500 184112 526534
rect 184044 526385 184112 526500
rect 184408 526498 184478 526699
rect 184408 526464 184425 526498
rect 184459 526464 184478 526498
rect 184408 526449 184478 526464
rect 185148 526534 185216 526551
rect 185148 526500 185165 526534
rect 185199 526500 185216 526534
rect 185148 526385 185216 526500
rect 185512 526498 185582 526699
rect 185512 526464 185529 526498
rect 185563 526464 185582 526498
rect 185512 526449 185582 526464
rect 186252 526534 186320 526551
rect 186252 526500 186269 526534
rect 186303 526500 186320 526534
rect 186252 526385 186320 526500
rect 186616 526498 186686 526699
rect 186616 526464 186633 526498
rect 186667 526464 186686 526498
rect 186616 526449 186686 526464
rect 187223 526649 187465 526710
rect 187223 526615 187241 526649
rect 187275 526615 187413 526649
rect 187447 526615 187465 526649
rect 187223 526568 187465 526615
rect 187223 526494 187327 526568
rect 187223 526460 187273 526494
rect 187307 526460 187327 526494
rect 187361 526500 187381 526534
rect 187415 526500 187465 526534
rect 187361 526426 187465 526500
rect 182531 526276 182589 526370
rect 182623 526371 183692 526385
rect 182623 526337 182641 526371
rect 182675 526337 183641 526371
rect 183675 526337 183692 526371
rect 182623 526276 183692 526337
rect 183727 526371 184796 526385
rect 183727 526337 183745 526371
rect 183779 526337 184745 526371
rect 184779 526337 184796 526371
rect 183727 526276 184796 526337
rect 184831 526371 185900 526385
rect 184831 526337 184849 526371
rect 184883 526337 185849 526371
rect 185883 526337 185900 526371
rect 184831 526276 185900 526337
rect 185935 526371 187004 526385
rect 185935 526337 185953 526371
rect 185987 526337 186953 526371
rect 186987 526337 187004 526371
rect 185935 526276 187004 526337
rect 187223 526373 187465 526426
rect 187223 526339 187241 526373
rect 187275 526339 187413 526373
rect 187447 526339 187465 526373
rect 187223 526276 187465 526339
rect 172210 526242 172239 526276
rect 172273 526242 172331 526276
rect 172365 526242 172423 526276
rect 172457 526242 172515 526276
rect 172549 526242 172607 526276
rect 172641 526242 172699 526276
rect 172733 526242 172791 526276
rect 172825 526242 172883 526276
rect 172917 526242 172975 526276
rect 173009 526242 173067 526276
rect 173101 526242 173159 526276
rect 173193 526242 173251 526276
rect 173285 526242 173343 526276
rect 173377 526242 173435 526276
rect 173469 526242 173527 526276
rect 173561 526242 173619 526276
rect 173653 526242 173711 526276
rect 173745 526242 173803 526276
rect 173837 526242 173895 526276
rect 173929 526242 173987 526276
rect 174021 526242 174079 526276
rect 174113 526242 174171 526276
rect 174205 526242 174263 526276
rect 174297 526242 174355 526276
rect 174389 526242 174447 526276
rect 174481 526242 174539 526276
rect 174573 526242 174631 526276
rect 174665 526242 174723 526276
rect 174757 526242 174815 526276
rect 174849 526242 174907 526276
rect 174941 526242 174999 526276
rect 175033 526242 175091 526276
rect 175125 526242 175183 526276
rect 175217 526242 175275 526276
rect 175309 526242 175367 526276
rect 175401 526242 175459 526276
rect 175493 526242 175551 526276
rect 175585 526242 175643 526276
rect 175677 526242 175735 526276
rect 175769 526242 175827 526276
rect 175861 526242 175919 526276
rect 175953 526242 176011 526276
rect 176045 526242 176103 526276
rect 176137 526242 176195 526276
rect 176229 526242 176287 526276
rect 176321 526242 176379 526276
rect 176413 526242 176471 526276
rect 176505 526242 176563 526276
rect 176597 526242 176655 526276
rect 176689 526242 176747 526276
rect 176781 526242 176839 526276
rect 176873 526242 176931 526276
rect 176965 526242 177023 526276
rect 177057 526242 177115 526276
rect 177149 526242 177207 526276
rect 177241 526242 177299 526276
rect 177333 526242 177391 526276
rect 177425 526242 177483 526276
rect 177517 526242 177575 526276
rect 177609 526242 177667 526276
rect 177701 526242 177759 526276
rect 177793 526242 177851 526276
rect 177885 526242 177943 526276
rect 177977 526242 178035 526276
rect 178069 526242 178127 526276
rect 178161 526242 178219 526276
rect 178253 526242 178311 526276
rect 178345 526242 178403 526276
rect 178437 526242 178495 526276
rect 178529 526242 178587 526276
rect 178621 526242 178679 526276
rect 178713 526242 178771 526276
rect 178805 526242 178863 526276
rect 178897 526242 178955 526276
rect 178989 526242 179047 526276
rect 179081 526242 179139 526276
rect 179173 526242 179231 526276
rect 179265 526242 179323 526276
rect 179357 526242 179415 526276
rect 179449 526242 179507 526276
rect 179541 526242 179599 526276
rect 179633 526242 179691 526276
rect 179725 526242 179783 526276
rect 179817 526242 179875 526276
rect 179909 526242 179967 526276
rect 180001 526242 180059 526276
rect 180093 526242 180151 526276
rect 180185 526242 180243 526276
rect 180277 526242 180335 526276
rect 180369 526242 180427 526276
rect 180461 526242 180519 526276
rect 180553 526242 180611 526276
rect 180645 526242 180703 526276
rect 180737 526242 180795 526276
rect 180829 526242 180887 526276
rect 180921 526242 180979 526276
rect 181013 526242 181071 526276
rect 181105 526242 181163 526276
rect 181197 526242 181255 526276
rect 181289 526242 181347 526276
rect 181381 526242 181439 526276
rect 181473 526242 181531 526276
rect 181565 526242 181623 526276
rect 181657 526242 181715 526276
rect 181749 526242 181807 526276
rect 181841 526242 181899 526276
rect 181933 526242 181991 526276
rect 182025 526242 182083 526276
rect 182117 526242 182175 526276
rect 182209 526242 182267 526276
rect 182301 526242 182359 526276
rect 182393 526242 182451 526276
rect 182485 526242 182543 526276
rect 182577 526242 182635 526276
rect 182669 526242 182727 526276
rect 182761 526242 182819 526276
rect 182853 526242 182911 526276
rect 182945 526242 183003 526276
rect 183037 526242 183095 526276
rect 183129 526242 183187 526276
rect 183221 526242 183279 526276
rect 183313 526242 183371 526276
rect 183405 526242 183463 526276
rect 183497 526242 183555 526276
rect 183589 526242 183647 526276
rect 183681 526242 183739 526276
rect 183773 526242 183831 526276
rect 183865 526242 183923 526276
rect 183957 526242 184015 526276
rect 184049 526242 184107 526276
rect 184141 526242 184199 526276
rect 184233 526242 184291 526276
rect 184325 526242 184383 526276
rect 184417 526242 184475 526276
rect 184509 526242 184567 526276
rect 184601 526242 184659 526276
rect 184693 526242 184751 526276
rect 184785 526242 184843 526276
rect 184877 526242 184935 526276
rect 184969 526242 185027 526276
rect 185061 526242 185119 526276
rect 185153 526242 185211 526276
rect 185245 526242 185303 526276
rect 185337 526242 185395 526276
rect 185429 526242 185487 526276
rect 185521 526242 185579 526276
rect 185613 526242 185671 526276
rect 185705 526242 185763 526276
rect 185797 526242 185855 526276
rect 185889 526242 185947 526276
rect 185981 526242 186039 526276
rect 186073 526242 186131 526276
rect 186165 526242 186223 526276
rect 186257 526242 186315 526276
rect 186349 526242 186407 526276
rect 186441 526242 186499 526276
rect 186533 526242 186591 526276
rect 186625 526242 186683 526276
rect 186717 526242 186775 526276
rect 186809 526242 186867 526276
rect 186901 526242 186959 526276
rect 186993 526242 187051 526276
rect 187085 526242 187143 526276
rect 187177 526242 187235 526276
rect 187269 526242 187327 526276
rect 187361 526242 187419 526276
rect 187453 526242 187482 526276
rect 172227 526179 172469 526242
rect 172227 526145 172245 526179
rect 172279 526145 172417 526179
rect 172451 526145 172469 526179
rect 172227 526092 172469 526145
rect 172503 526181 173572 526242
rect 172503 526147 172521 526181
rect 172555 526147 173521 526181
rect 173555 526147 173572 526181
rect 172503 526133 173572 526147
rect 173607 526181 174676 526242
rect 173607 526147 173625 526181
rect 173659 526147 174625 526181
rect 174659 526147 174676 526181
rect 173607 526133 174676 526147
rect 174803 526148 174861 526242
rect 172227 526018 172331 526092
rect 172227 525984 172277 526018
rect 172311 525984 172331 526018
rect 172365 526024 172385 526058
rect 172419 526024 172469 526058
rect 172365 525950 172469 526024
rect 172820 526018 172888 526133
rect 172820 525984 172837 526018
rect 172871 525984 172888 526018
rect 172820 525967 172888 525984
rect 173184 526054 173254 526069
rect 173184 526020 173201 526054
rect 173235 526020 173254 526054
rect 172227 525903 172469 525950
rect 172227 525869 172245 525903
rect 172279 525869 172417 525903
rect 172451 525869 172469 525903
rect 172227 525808 172469 525869
rect 173184 525819 173254 526020
rect 173924 526018 173992 526133
rect 174803 526114 174815 526148
rect 174849 526114 174861 526148
rect 174895 526181 175964 526242
rect 174895 526147 174913 526181
rect 174947 526147 175913 526181
rect 175947 526147 175964 526181
rect 174895 526133 175964 526147
rect 175999 526181 177068 526242
rect 175999 526147 176017 526181
rect 176051 526147 177017 526181
rect 177051 526147 177068 526181
rect 175999 526133 177068 526147
rect 177103 526181 178172 526242
rect 177103 526147 177121 526181
rect 177155 526147 178121 526181
rect 178155 526147 178172 526181
rect 177103 526133 178172 526147
rect 178207 526181 179276 526242
rect 178207 526147 178225 526181
rect 178259 526147 179225 526181
rect 179259 526147 179276 526181
rect 178207 526133 179276 526147
rect 179311 526181 179829 526242
rect 179311 526147 179329 526181
rect 179363 526147 179777 526181
rect 179811 526147 179829 526181
rect 174803 526097 174861 526114
rect 173924 525984 173941 526018
rect 173975 525984 173992 526018
rect 173924 525967 173992 525984
rect 174288 526054 174358 526069
rect 174288 526020 174305 526054
rect 174339 526020 174358 526054
rect 174288 525819 174358 526020
rect 175212 526018 175280 526133
rect 175212 525984 175229 526018
rect 175263 525984 175280 526018
rect 175212 525967 175280 525984
rect 175576 526054 175646 526069
rect 175576 526020 175593 526054
rect 175627 526020 175646 526054
rect 174803 525930 174861 525965
rect 174803 525896 174815 525930
rect 174849 525896 174861 525930
rect 174803 525837 174861 525896
rect 172227 525774 172245 525808
rect 172279 525774 172417 525808
rect 172451 525774 172469 525808
rect 172227 525732 172469 525774
rect 172503 525808 173572 525819
rect 172503 525774 172521 525808
rect 172555 525774 173521 525808
rect 173555 525774 173572 525808
rect 172503 525732 173572 525774
rect 173607 525808 174676 525819
rect 173607 525774 173625 525808
rect 173659 525774 174625 525808
rect 174659 525774 174676 525808
rect 173607 525732 174676 525774
rect 174803 525803 174815 525837
rect 174849 525803 174861 525837
rect 175576 525819 175646 526020
rect 176316 526018 176384 526133
rect 176316 525984 176333 526018
rect 176367 525984 176384 526018
rect 176316 525967 176384 525984
rect 176680 526054 176750 526069
rect 176680 526020 176697 526054
rect 176731 526020 176750 526054
rect 176680 525819 176750 526020
rect 177420 526018 177488 526133
rect 177420 525984 177437 526018
rect 177471 525984 177488 526018
rect 177420 525967 177488 525984
rect 177784 526054 177854 526069
rect 177784 526020 177801 526054
rect 177835 526020 177854 526054
rect 177784 525819 177854 526020
rect 178524 526018 178592 526133
rect 179311 526088 179829 526147
rect 179955 526148 180013 526242
rect 179955 526114 179967 526148
rect 180001 526114 180013 526148
rect 180047 526181 181116 526242
rect 180047 526147 180065 526181
rect 180099 526147 181065 526181
rect 181099 526147 181116 526181
rect 180047 526133 181116 526147
rect 181151 526181 182220 526242
rect 181151 526147 181169 526181
rect 181203 526147 182169 526181
rect 182203 526147 182220 526181
rect 181151 526133 182220 526147
rect 182255 526181 183324 526242
rect 182255 526147 182273 526181
rect 182307 526147 183273 526181
rect 183307 526147 183324 526181
rect 182255 526133 183324 526147
rect 183359 526181 184428 526242
rect 183359 526147 183377 526181
rect 183411 526147 184377 526181
rect 184411 526147 184428 526181
rect 183359 526133 184428 526147
rect 184463 526181 184981 526242
rect 184463 526147 184481 526181
rect 184515 526147 184929 526181
rect 184963 526147 184981 526181
rect 179955 526097 180013 526114
rect 178524 525984 178541 526018
rect 178575 525984 178592 526018
rect 178524 525967 178592 525984
rect 178888 526054 178958 526069
rect 178888 526020 178905 526054
rect 178939 526020 178958 526054
rect 178888 525819 178958 526020
rect 179311 526018 179553 526088
rect 179311 525984 179389 526018
rect 179423 525984 179499 526018
rect 179533 525984 179553 526018
rect 179587 526020 179607 526054
rect 179641 526020 179717 526054
rect 179751 526020 179829 526054
rect 179587 525950 179829 526020
rect 180364 526018 180432 526133
rect 180364 525984 180381 526018
rect 180415 525984 180432 526018
rect 180364 525967 180432 525984
rect 180728 526054 180798 526069
rect 180728 526020 180745 526054
rect 180779 526020 180798 526054
rect 179311 525910 179829 525950
rect 179311 525876 179329 525910
rect 179363 525876 179777 525910
rect 179811 525876 179829 525910
rect 174803 525732 174861 525803
rect 174895 525808 175964 525819
rect 174895 525774 174913 525808
rect 174947 525774 175913 525808
rect 175947 525774 175964 525808
rect 174895 525732 175964 525774
rect 175999 525808 177068 525819
rect 175999 525774 176017 525808
rect 176051 525774 177017 525808
rect 177051 525774 177068 525808
rect 175999 525732 177068 525774
rect 177103 525808 178172 525819
rect 177103 525774 177121 525808
rect 177155 525774 178121 525808
rect 178155 525774 178172 525808
rect 177103 525732 178172 525774
rect 178207 525808 179276 525819
rect 178207 525774 178225 525808
rect 178259 525774 179225 525808
rect 179259 525774 179276 525808
rect 178207 525732 179276 525774
rect 179311 525808 179829 525876
rect 179311 525774 179329 525808
rect 179363 525774 179777 525808
rect 179811 525774 179829 525808
rect 179311 525732 179829 525774
rect 179955 525930 180013 525965
rect 179955 525896 179967 525930
rect 180001 525896 180013 525930
rect 179955 525837 180013 525896
rect 179955 525803 179967 525837
rect 180001 525803 180013 525837
rect 180728 525819 180798 526020
rect 181468 526018 181536 526133
rect 181468 525984 181485 526018
rect 181519 525984 181536 526018
rect 181468 525967 181536 525984
rect 181832 526054 181902 526069
rect 181832 526020 181849 526054
rect 181883 526020 181902 526054
rect 181832 525819 181902 526020
rect 182572 526018 182640 526133
rect 182572 525984 182589 526018
rect 182623 525984 182640 526018
rect 182572 525967 182640 525984
rect 182936 526054 183006 526069
rect 182936 526020 182953 526054
rect 182987 526020 183006 526054
rect 182936 525819 183006 526020
rect 183676 526018 183744 526133
rect 184463 526088 184981 526147
rect 185107 526148 185165 526242
rect 185107 526114 185119 526148
rect 185153 526114 185165 526148
rect 185199 526181 186268 526242
rect 185199 526147 185217 526181
rect 185251 526147 186217 526181
rect 186251 526147 186268 526181
rect 185199 526133 186268 526147
rect 186303 526181 187005 526242
rect 186303 526147 186321 526181
rect 186355 526147 186953 526181
rect 186987 526147 187005 526181
rect 185107 526097 185165 526114
rect 183676 525984 183693 526018
rect 183727 525984 183744 526018
rect 183676 525967 183744 525984
rect 184040 526054 184110 526069
rect 184040 526020 184057 526054
rect 184091 526020 184110 526054
rect 184040 525819 184110 526020
rect 184463 526018 184705 526088
rect 184463 525984 184541 526018
rect 184575 525984 184651 526018
rect 184685 525984 184705 526018
rect 184739 526020 184759 526054
rect 184793 526020 184869 526054
rect 184903 526020 184981 526054
rect 184739 525950 184981 526020
rect 185516 526018 185584 526133
rect 186303 526088 187005 526147
rect 187223 526179 187465 526242
rect 187223 526145 187241 526179
rect 187275 526145 187413 526179
rect 187447 526145 187465 526179
rect 187223 526092 187465 526145
rect 185516 525984 185533 526018
rect 185567 525984 185584 526018
rect 185516 525967 185584 525984
rect 185880 526054 185950 526069
rect 185880 526020 185897 526054
rect 185931 526020 185950 526054
rect 184463 525910 184981 525950
rect 184463 525876 184481 525910
rect 184515 525876 184929 525910
rect 184963 525876 184981 525910
rect 179955 525732 180013 525803
rect 180047 525808 181116 525819
rect 180047 525774 180065 525808
rect 180099 525774 181065 525808
rect 181099 525774 181116 525808
rect 180047 525732 181116 525774
rect 181151 525808 182220 525819
rect 181151 525774 181169 525808
rect 181203 525774 182169 525808
rect 182203 525774 182220 525808
rect 181151 525732 182220 525774
rect 182255 525808 183324 525819
rect 182255 525774 182273 525808
rect 182307 525774 183273 525808
rect 183307 525774 183324 525808
rect 182255 525732 183324 525774
rect 183359 525808 184428 525819
rect 183359 525774 183377 525808
rect 183411 525774 184377 525808
rect 184411 525774 184428 525808
rect 183359 525732 184428 525774
rect 184463 525808 184981 525876
rect 184463 525774 184481 525808
rect 184515 525774 184929 525808
rect 184963 525774 184981 525808
rect 184463 525732 184981 525774
rect 185107 525930 185165 525965
rect 185107 525896 185119 525930
rect 185153 525896 185165 525930
rect 185107 525837 185165 525896
rect 185107 525803 185119 525837
rect 185153 525803 185165 525837
rect 185880 525819 185950 526020
rect 186303 526018 186633 526088
rect 186303 525984 186381 526018
rect 186415 525984 186480 526018
rect 186514 525984 186579 526018
rect 186613 525984 186633 526018
rect 186667 526020 186687 526054
rect 186721 526020 186790 526054
rect 186824 526020 186893 526054
rect 186927 526020 187005 526054
rect 186667 525950 187005 526020
rect 186303 525910 187005 525950
rect 186303 525876 186321 525910
rect 186355 525876 186953 525910
rect 186987 525876 187005 525910
rect 185107 525732 185165 525803
rect 185199 525808 186268 525819
rect 185199 525774 185217 525808
rect 185251 525774 186217 525808
rect 186251 525774 186268 525808
rect 185199 525732 186268 525774
rect 186303 525808 187005 525876
rect 186303 525774 186321 525808
rect 186355 525774 186953 525808
rect 186987 525774 187005 525808
rect 186303 525732 187005 525774
rect 187223 526024 187273 526058
rect 187307 526024 187327 526058
rect 187223 525950 187327 526024
rect 187361 526018 187465 526092
rect 187361 525984 187381 526018
rect 187415 525984 187465 526018
rect 187223 525903 187465 525950
rect 187223 525869 187241 525903
rect 187275 525869 187413 525903
rect 187447 525869 187465 525903
rect 187223 525808 187465 525869
rect 187223 525774 187241 525808
rect 187275 525774 187413 525808
rect 187447 525774 187465 525808
rect 187223 525732 187465 525774
rect 172210 525698 172239 525732
rect 172273 525698 172331 525732
rect 172365 525698 172423 525732
rect 172457 525698 172515 525732
rect 172549 525698 172607 525732
rect 172641 525698 172699 525732
rect 172733 525698 172791 525732
rect 172825 525698 172883 525732
rect 172917 525698 172975 525732
rect 173009 525698 173067 525732
rect 173101 525698 173159 525732
rect 173193 525698 173251 525732
rect 173285 525698 173343 525732
rect 173377 525698 173435 525732
rect 173469 525698 173527 525732
rect 173561 525698 173619 525732
rect 173653 525698 173711 525732
rect 173745 525698 173803 525732
rect 173837 525698 173895 525732
rect 173929 525698 173987 525732
rect 174021 525698 174079 525732
rect 174113 525698 174171 525732
rect 174205 525698 174263 525732
rect 174297 525698 174355 525732
rect 174389 525698 174447 525732
rect 174481 525698 174539 525732
rect 174573 525698 174631 525732
rect 174665 525698 174723 525732
rect 174757 525698 174815 525732
rect 174849 525698 174907 525732
rect 174941 525698 174999 525732
rect 175033 525698 175091 525732
rect 175125 525698 175183 525732
rect 175217 525698 175275 525732
rect 175309 525698 175367 525732
rect 175401 525698 175459 525732
rect 175493 525698 175551 525732
rect 175585 525698 175643 525732
rect 175677 525698 175735 525732
rect 175769 525698 175827 525732
rect 175861 525698 175919 525732
rect 175953 525698 176011 525732
rect 176045 525698 176103 525732
rect 176137 525698 176195 525732
rect 176229 525698 176287 525732
rect 176321 525698 176379 525732
rect 176413 525698 176471 525732
rect 176505 525698 176563 525732
rect 176597 525698 176655 525732
rect 176689 525698 176747 525732
rect 176781 525698 176839 525732
rect 176873 525698 176931 525732
rect 176965 525698 177023 525732
rect 177057 525698 177115 525732
rect 177149 525698 177207 525732
rect 177241 525698 177299 525732
rect 177333 525698 177391 525732
rect 177425 525698 177483 525732
rect 177517 525698 177575 525732
rect 177609 525698 177667 525732
rect 177701 525698 177759 525732
rect 177793 525698 177851 525732
rect 177885 525698 177943 525732
rect 177977 525698 178035 525732
rect 178069 525698 178127 525732
rect 178161 525698 178219 525732
rect 178253 525698 178311 525732
rect 178345 525698 178403 525732
rect 178437 525698 178495 525732
rect 178529 525698 178587 525732
rect 178621 525698 178679 525732
rect 178713 525698 178771 525732
rect 178805 525698 178863 525732
rect 178897 525698 178955 525732
rect 178989 525698 179047 525732
rect 179081 525698 179139 525732
rect 179173 525698 179231 525732
rect 179265 525698 179323 525732
rect 179357 525698 179415 525732
rect 179449 525698 179507 525732
rect 179541 525698 179599 525732
rect 179633 525698 179691 525732
rect 179725 525698 179783 525732
rect 179817 525698 179875 525732
rect 179909 525698 179967 525732
rect 180001 525698 180059 525732
rect 180093 525698 180151 525732
rect 180185 525698 180243 525732
rect 180277 525698 180335 525732
rect 180369 525698 180427 525732
rect 180461 525698 180519 525732
rect 180553 525698 180611 525732
rect 180645 525698 180703 525732
rect 180737 525698 180795 525732
rect 180829 525698 180887 525732
rect 180921 525698 180979 525732
rect 181013 525698 181071 525732
rect 181105 525698 181163 525732
rect 181197 525698 181255 525732
rect 181289 525698 181347 525732
rect 181381 525698 181439 525732
rect 181473 525698 181531 525732
rect 181565 525698 181623 525732
rect 181657 525698 181715 525732
rect 181749 525698 181807 525732
rect 181841 525698 181899 525732
rect 181933 525698 181991 525732
rect 182025 525698 182083 525732
rect 182117 525698 182175 525732
rect 182209 525698 182267 525732
rect 182301 525698 182359 525732
rect 182393 525698 182451 525732
rect 182485 525698 182543 525732
rect 182577 525698 182635 525732
rect 182669 525698 182727 525732
rect 182761 525698 182819 525732
rect 182853 525698 182911 525732
rect 182945 525698 183003 525732
rect 183037 525698 183095 525732
rect 183129 525698 183187 525732
rect 183221 525698 183279 525732
rect 183313 525698 183371 525732
rect 183405 525698 183463 525732
rect 183497 525698 183555 525732
rect 183589 525698 183647 525732
rect 183681 525698 183739 525732
rect 183773 525698 183831 525732
rect 183865 525698 183923 525732
rect 183957 525698 184015 525732
rect 184049 525698 184107 525732
rect 184141 525698 184199 525732
rect 184233 525698 184291 525732
rect 184325 525698 184383 525732
rect 184417 525698 184475 525732
rect 184509 525698 184567 525732
rect 184601 525698 184659 525732
rect 184693 525698 184751 525732
rect 184785 525698 184843 525732
rect 184877 525698 184935 525732
rect 184969 525698 185027 525732
rect 185061 525698 185119 525732
rect 185153 525698 185211 525732
rect 185245 525698 185303 525732
rect 185337 525698 185395 525732
rect 185429 525698 185487 525732
rect 185521 525698 185579 525732
rect 185613 525698 185671 525732
rect 185705 525698 185763 525732
rect 185797 525698 185855 525732
rect 185889 525698 185947 525732
rect 185981 525698 186039 525732
rect 186073 525698 186131 525732
rect 186165 525698 186223 525732
rect 186257 525698 186315 525732
rect 186349 525698 186407 525732
rect 186441 525698 186499 525732
rect 186533 525698 186591 525732
rect 186625 525698 186683 525732
rect 186717 525698 186775 525732
rect 186809 525698 186867 525732
rect 186901 525698 186959 525732
rect 186993 525698 187051 525732
rect 187085 525698 187143 525732
rect 187177 525698 187235 525732
rect 187269 525698 187327 525732
rect 187361 525698 187419 525732
rect 187453 525698 187482 525732
rect 172227 525656 172469 525698
rect 172227 525622 172245 525656
rect 172279 525622 172417 525656
rect 172451 525622 172469 525656
rect 172227 525561 172469 525622
rect 172503 525656 173572 525698
rect 172503 525622 172521 525656
rect 172555 525622 173521 525656
rect 173555 525622 173572 525656
rect 172503 525611 173572 525622
rect 173607 525656 174676 525698
rect 173607 525622 173625 525656
rect 173659 525622 174625 525656
rect 174659 525622 174676 525656
rect 173607 525611 174676 525622
rect 174711 525656 175780 525698
rect 174711 525622 174729 525656
rect 174763 525622 175729 525656
rect 175763 525622 175780 525656
rect 174711 525611 175780 525622
rect 175815 525656 176884 525698
rect 175815 525622 175833 525656
rect 175867 525622 176833 525656
rect 176867 525622 176884 525656
rect 175815 525611 176884 525622
rect 176919 525656 177253 525698
rect 176919 525622 176937 525656
rect 176971 525622 177201 525656
rect 177235 525622 177253 525656
rect 172227 525527 172245 525561
rect 172279 525527 172417 525561
rect 172451 525527 172469 525561
rect 172227 525480 172469 525527
rect 172227 525412 172277 525446
rect 172311 525412 172331 525446
rect 172227 525338 172331 525412
rect 172365 525406 172469 525480
rect 172365 525372 172385 525406
rect 172419 525372 172469 525406
rect 172820 525446 172888 525463
rect 172820 525412 172837 525446
rect 172871 525412 172888 525446
rect 172227 525285 172469 525338
rect 172820 525297 172888 525412
rect 173184 525410 173254 525611
rect 173184 525376 173201 525410
rect 173235 525376 173254 525410
rect 173184 525361 173254 525376
rect 173924 525446 173992 525463
rect 173924 525412 173941 525446
rect 173975 525412 173992 525446
rect 173924 525297 173992 525412
rect 174288 525410 174358 525611
rect 174288 525376 174305 525410
rect 174339 525376 174358 525410
rect 174288 525361 174358 525376
rect 175028 525446 175096 525463
rect 175028 525412 175045 525446
rect 175079 525412 175096 525446
rect 175028 525297 175096 525412
rect 175392 525410 175462 525611
rect 175392 525376 175409 525410
rect 175443 525376 175462 525410
rect 175392 525361 175462 525376
rect 176132 525446 176200 525463
rect 176132 525412 176149 525446
rect 176183 525412 176200 525446
rect 176132 525297 176200 525412
rect 176496 525410 176566 525611
rect 176919 525554 177253 525622
rect 176919 525520 176937 525554
rect 176971 525520 177201 525554
rect 177235 525520 177253 525554
rect 176919 525480 177253 525520
rect 176496 525376 176513 525410
rect 176547 525376 176566 525410
rect 176496 525361 176566 525376
rect 176919 525412 176939 525446
rect 176973 525412 177069 525446
rect 176919 525342 177069 525412
rect 177103 525410 177253 525480
rect 177379 525627 177437 525698
rect 177379 525593 177391 525627
rect 177425 525593 177437 525627
rect 177471 525656 178540 525698
rect 177471 525622 177489 525656
rect 177523 525622 178489 525656
rect 178523 525622 178540 525656
rect 177471 525611 178540 525622
rect 178575 525656 179644 525698
rect 178575 525622 178593 525656
rect 178627 525622 179593 525656
rect 179627 525622 179644 525656
rect 178575 525611 179644 525622
rect 179679 525656 180748 525698
rect 179679 525622 179697 525656
rect 179731 525622 180697 525656
rect 180731 525622 180748 525656
rect 179679 525611 180748 525622
rect 180783 525656 181852 525698
rect 180783 525622 180801 525656
rect 180835 525622 181801 525656
rect 181835 525622 181852 525656
rect 180783 525611 181852 525622
rect 181887 525656 182405 525698
rect 181887 525622 181905 525656
rect 181939 525622 182353 525656
rect 182387 525622 182405 525656
rect 177379 525534 177437 525593
rect 177379 525500 177391 525534
rect 177425 525500 177437 525534
rect 177379 525465 177437 525500
rect 177103 525376 177199 525410
rect 177233 525376 177253 525410
rect 177788 525446 177856 525463
rect 177788 525412 177805 525446
rect 177839 525412 177856 525446
rect 172227 525251 172245 525285
rect 172279 525251 172417 525285
rect 172451 525251 172469 525285
rect 172227 525188 172469 525251
rect 172503 525283 173572 525297
rect 172503 525249 172521 525283
rect 172555 525249 173521 525283
rect 173555 525249 173572 525283
rect 172503 525188 173572 525249
rect 173607 525283 174676 525297
rect 173607 525249 173625 525283
rect 173659 525249 174625 525283
rect 174659 525249 174676 525283
rect 173607 525188 174676 525249
rect 174711 525283 175780 525297
rect 174711 525249 174729 525283
rect 174763 525249 175729 525283
rect 175763 525249 175780 525283
rect 174711 525188 175780 525249
rect 175815 525283 176884 525297
rect 175815 525249 175833 525283
rect 175867 525249 176833 525283
rect 176867 525249 176884 525283
rect 175815 525188 176884 525249
rect 176919 525290 177253 525342
rect 176919 525256 176937 525290
rect 176971 525256 177201 525290
rect 177235 525256 177253 525290
rect 176919 525188 177253 525256
rect 177379 525316 177437 525333
rect 177379 525282 177391 525316
rect 177425 525282 177437 525316
rect 177788 525297 177856 525412
rect 178152 525410 178222 525611
rect 178152 525376 178169 525410
rect 178203 525376 178222 525410
rect 178152 525361 178222 525376
rect 178892 525446 178960 525463
rect 178892 525412 178909 525446
rect 178943 525412 178960 525446
rect 178892 525297 178960 525412
rect 179256 525410 179326 525611
rect 179256 525376 179273 525410
rect 179307 525376 179326 525410
rect 179256 525361 179326 525376
rect 179996 525446 180064 525463
rect 179996 525412 180013 525446
rect 180047 525412 180064 525446
rect 179996 525297 180064 525412
rect 180360 525410 180430 525611
rect 180360 525376 180377 525410
rect 180411 525376 180430 525410
rect 180360 525361 180430 525376
rect 181100 525446 181168 525463
rect 181100 525412 181117 525446
rect 181151 525412 181168 525446
rect 181100 525297 181168 525412
rect 181464 525410 181534 525611
rect 181887 525554 182405 525622
rect 181887 525520 181905 525554
rect 181939 525520 182353 525554
rect 182387 525520 182405 525554
rect 181887 525480 182405 525520
rect 181464 525376 181481 525410
rect 181515 525376 181534 525410
rect 181464 525361 181534 525376
rect 181887 525412 181965 525446
rect 181999 525412 182075 525446
rect 182109 525412 182129 525446
rect 181887 525342 182129 525412
rect 182163 525410 182405 525480
rect 182531 525627 182589 525698
rect 182531 525593 182543 525627
rect 182577 525593 182589 525627
rect 182623 525656 183692 525698
rect 182623 525622 182641 525656
rect 182675 525622 183641 525656
rect 183675 525622 183692 525656
rect 182623 525611 183692 525622
rect 183727 525656 184796 525698
rect 183727 525622 183745 525656
rect 183779 525622 184745 525656
rect 184779 525622 184796 525656
rect 183727 525611 184796 525622
rect 184831 525656 185900 525698
rect 184831 525622 184849 525656
rect 184883 525622 185849 525656
rect 185883 525622 185900 525656
rect 184831 525611 185900 525622
rect 185935 525656 187004 525698
rect 185935 525622 185953 525656
rect 185987 525622 186953 525656
rect 186987 525622 187004 525656
rect 185935 525611 187004 525622
rect 187223 525656 187465 525698
rect 187223 525622 187241 525656
rect 187275 525622 187413 525656
rect 187447 525622 187465 525656
rect 182531 525534 182589 525593
rect 182531 525500 182543 525534
rect 182577 525500 182589 525534
rect 182531 525465 182589 525500
rect 182163 525376 182183 525410
rect 182217 525376 182293 525410
rect 182327 525376 182405 525410
rect 182940 525446 183008 525463
rect 182940 525412 182957 525446
rect 182991 525412 183008 525446
rect 177379 525188 177437 525282
rect 177471 525283 178540 525297
rect 177471 525249 177489 525283
rect 177523 525249 178489 525283
rect 178523 525249 178540 525283
rect 177471 525188 178540 525249
rect 178575 525283 179644 525297
rect 178575 525249 178593 525283
rect 178627 525249 179593 525283
rect 179627 525249 179644 525283
rect 178575 525188 179644 525249
rect 179679 525283 180748 525297
rect 179679 525249 179697 525283
rect 179731 525249 180697 525283
rect 180731 525249 180748 525283
rect 179679 525188 180748 525249
rect 180783 525283 181852 525297
rect 180783 525249 180801 525283
rect 180835 525249 181801 525283
rect 181835 525249 181852 525283
rect 180783 525188 181852 525249
rect 181887 525283 182405 525342
rect 181887 525249 181905 525283
rect 181939 525249 182353 525283
rect 182387 525249 182405 525283
rect 181887 525188 182405 525249
rect 182531 525316 182589 525333
rect 182531 525282 182543 525316
rect 182577 525282 182589 525316
rect 182940 525297 183008 525412
rect 183304 525410 183374 525611
rect 183304 525376 183321 525410
rect 183355 525376 183374 525410
rect 183304 525361 183374 525376
rect 184044 525446 184112 525463
rect 184044 525412 184061 525446
rect 184095 525412 184112 525446
rect 184044 525297 184112 525412
rect 184408 525410 184478 525611
rect 184408 525376 184425 525410
rect 184459 525376 184478 525410
rect 184408 525361 184478 525376
rect 185148 525446 185216 525463
rect 185148 525412 185165 525446
rect 185199 525412 185216 525446
rect 185148 525297 185216 525412
rect 185512 525410 185582 525611
rect 185512 525376 185529 525410
rect 185563 525376 185582 525410
rect 185512 525361 185582 525376
rect 186252 525446 186320 525463
rect 186252 525412 186269 525446
rect 186303 525412 186320 525446
rect 186252 525297 186320 525412
rect 186616 525410 186686 525611
rect 186616 525376 186633 525410
rect 186667 525376 186686 525410
rect 186616 525361 186686 525376
rect 187223 525561 187465 525622
rect 187223 525527 187241 525561
rect 187275 525527 187413 525561
rect 187447 525527 187465 525561
rect 187223 525480 187465 525527
rect 187223 525406 187327 525480
rect 187223 525372 187273 525406
rect 187307 525372 187327 525406
rect 187361 525412 187381 525446
rect 187415 525412 187465 525446
rect 187361 525338 187465 525412
rect 182531 525188 182589 525282
rect 182623 525283 183692 525297
rect 182623 525249 182641 525283
rect 182675 525249 183641 525283
rect 183675 525249 183692 525283
rect 182623 525188 183692 525249
rect 183727 525283 184796 525297
rect 183727 525249 183745 525283
rect 183779 525249 184745 525283
rect 184779 525249 184796 525283
rect 183727 525188 184796 525249
rect 184831 525283 185900 525297
rect 184831 525249 184849 525283
rect 184883 525249 185849 525283
rect 185883 525249 185900 525283
rect 184831 525188 185900 525249
rect 185935 525283 187004 525297
rect 185935 525249 185953 525283
rect 185987 525249 186953 525283
rect 186987 525249 187004 525283
rect 185935 525188 187004 525249
rect 187223 525285 187465 525338
rect 187223 525251 187241 525285
rect 187275 525251 187413 525285
rect 187447 525251 187465 525285
rect 187223 525188 187465 525251
rect 172210 525154 172239 525188
rect 172273 525154 172331 525188
rect 172365 525154 172423 525188
rect 172457 525154 172515 525188
rect 172549 525154 172607 525188
rect 172641 525154 172699 525188
rect 172733 525154 172791 525188
rect 172825 525154 172883 525188
rect 172917 525154 172975 525188
rect 173009 525154 173067 525188
rect 173101 525154 173159 525188
rect 173193 525154 173251 525188
rect 173285 525154 173343 525188
rect 173377 525154 173435 525188
rect 173469 525154 173527 525188
rect 173561 525154 173619 525188
rect 173653 525154 173711 525188
rect 173745 525154 173803 525188
rect 173837 525154 173895 525188
rect 173929 525154 173987 525188
rect 174021 525154 174079 525188
rect 174113 525154 174171 525188
rect 174205 525154 174263 525188
rect 174297 525154 174355 525188
rect 174389 525154 174447 525188
rect 174481 525154 174539 525188
rect 174573 525154 174631 525188
rect 174665 525154 174723 525188
rect 174757 525154 174815 525188
rect 174849 525154 174907 525188
rect 174941 525154 174999 525188
rect 175033 525154 175091 525188
rect 175125 525154 175183 525188
rect 175217 525154 175275 525188
rect 175309 525154 175367 525188
rect 175401 525154 175459 525188
rect 175493 525154 175551 525188
rect 175585 525154 175643 525188
rect 175677 525154 175735 525188
rect 175769 525154 175827 525188
rect 175861 525154 175919 525188
rect 175953 525154 176011 525188
rect 176045 525154 176103 525188
rect 176137 525154 176195 525188
rect 176229 525154 176287 525188
rect 176321 525154 176379 525188
rect 176413 525154 176471 525188
rect 176505 525154 176563 525188
rect 176597 525154 176655 525188
rect 176689 525154 176747 525188
rect 176781 525154 176839 525188
rect 176873 525154 176931 525188
rect 176965 525154 177023 525188
rect 177057 525154 177115 525188
rect 177149 525154 177207 525188
rect 177241 525154 177299 525188
rect 177333 525154 177391 525188
rect 177425 525154 177483 525188
rect 177517 525154 177575 525188
rect 177609 525154 177667 525188
rect 177701 525154 177759 525188
rect 177793 525154 177851 525188
rect 177885 525154 177943 525188
rect 177977 525154 178035 525188
rect 178069 525154 178127 525188
rect 178161 525154 178219 525188
rect 178253 525154 178311 525188
rect 178345 525154 178403 525188
rect 178437 525154 178495 525188
rect 178529 525154 178587 525188
rect 178621 525154 178679 525188
rect 178713 525154 178771 525188
rect 178805 525154 178863 525188
rect 178897 525154 178955 525188
rect 178989 525154 179047 525188
rect 179081 525154 179139 525188
rect 179173 525154 179231 525188
rect 179265 525154 179323 525188
rect 179357 525154 179415 525188
rect 179449 525154 179507 525188
rect 179541 525154 179599 525188
rect 179633 525154 179691 525188
rect 179725 525154 179783 525188
rect 179817 525154 179875 525188
rect 179909 525154 179967 525188
rect 180001 525154 180059 525188
rect 180093 525154 180151 525188
rect 180185 525154 180243 525188
rect 180277 525154 180335 525188
rect 180369 525154 180427 525188
rect 180461 525154 180519 525188
rect 180553 525154 180611 525188
rect 180645 525154 180703 525188
rect 180737 525154 180795 525188
rect 180829 525154 180887 525188
rect 180921 525154 180979 525188
rect 181013 525154 181071 525188
rect 181105 525154 181163 525188
rect 181197 525154 181255 525188
rect 181289 525154 181347 525188
rect 181381 525154 181439 525188
rect 181473 525154 181531 525188
rect 181565 525154 181623 525188
rect 181657 525154 181715 525188
rect 181749 525154 181807 525188
rect 181841 525154 181899 525188
rect 181933 525154 181991 525188
rect 182025 525154 182083 525188
rect 182117 525154 182175 525188
rect 182209 525154 182267 525188
rect 182301 525154 182359 525188
rect 182393 525154 182451 525188
rect 182485 525154 182543 525188
rect 182577 525154 182635 525188
rect 182669 525154 182727 525188
rect 182761 525154 182819 525188
rect 182853 525154 182911 525188
rect 182945 525154 183003 525188
rect 183037 525154 183095 525188
rect 183129 525154 183187 525188
rect 183221 525154 183279 525188
rect 183313 525154 183371 525188
rect 183405 525154 183463 525188
rect 183497 525154 183555 525188
rect 183589 525154 183647 525188
rect 183681 525154 183739 525188
rect 183773 525154 183831 525188
rect 183865 525154 183923 525188
rect 183957 525154 184015 525188
rect 184049 525154 184107 525188
rect 184141 525154 184199 525188
rect 184233 525154 184291 525188
rect 184325 525154 184383 525188
rect 184417 525154 184475 525188
rect 184509 525154 184567 525188
rect 184601 525154 184659 525188
rect 184693 525154 184751 525188
rect 184785 525154 184843 525188
rect 184877 525154 184935 525188
rect 184969 525154 185027 525188
rect 185061 525154 185119 525188
rect 185153 525154 185211 525188
rect 185245 525154 185303 525188
rect 185337 525154 185395 525188
rect 185429 525154 185487 525188
rect 185521 525154 185579 525188
rect 185613 525154 185671 525188
rect 185705 525154 185763 525188
rect 185797 525154 185855 525188
rect 185889 525154 185947 525188
rect 185981 525154 186039 525188
rect 186073 525154 186131 525188
rect 186165 525154 186223 525188
rect 186257 525154 186315 525188
rect 186349 525154 186407 525188
rect 186441 525154 186499 525188
rect 186533 525154 186591 525188
rect 186625 525154 186683 525188
rect 186717 525154 186775 525188
rect 186809 525154 186867 525188
rect 186901 525154 186959 525188
rect 186993 525154 187051 525188
rect 187085 525154 187143 525188
rect 187177 525154 187235 525188
rect 187269 525154 187327 525188
rect 187361 525154 187419 525188
rect 187453 525154 187482 525188
rect 172227 525091 172469 525154
rect 172227 525057 172245 525091
rect 172279 525057 172417 525091
rect 172451 525057 172469 525091
rect 172227 525004 172469 525057
rect 172503 525093 173572 525154
rect 172503 525059 172521 525093
rect 172555 525059 173521 525093
rect 173555 525059 173572 525093
rect 172503 525045 173572 525059
rect 173607 525093 174676 525154
rect 173607 525059 173625 525093
rect 173659 525059 174625 525093
rect 174659 525059 174676 525093
rect 173607 525045 174676 525059
rect 174803 525060 174861 525154
rect 172227 524930 172331 525004
rect 172227 524896 172277 524930
rect 172311 524896 172331 524930
rect 172365 524936 172385 524970
rect 172419 524936 172469 524970
rect 172365 524862 172469 524936
rect 172820 524930 172888 525045
rect 172820 524896 172837 524930
rect 172871 524896 172888 524930
rect 172820 524879 172888 524896
rect 173184 524966 173254 524981
rect 173184 524932 173201 524966
rect 173235 524932 173254 524966
rect 172227 524815 172469 524862
rect 172227 524781 172245 524815
rect 172279 524781 172417 524815
rect 172451 524781 172469 524815
rect 172227 524720 172469 524781
rect 173184 524731 173254 524932
rect 173924 524930 173992 525045
rect 174803 525026 174815 525060
rect 174849 525026 174861 525060
rect 174895 525093 175964 525154
rect 174895 525059 174913 525093
rect 174947 525059 175913 525093
rect 175947 525059 175964 525093
rect 174895 525045 175964 525059
rect 175999 525093 177068 525154
rect 175999 525059 176017 525093
rect 176051 525059 177017 525093
rect 177051 525059 177068 525093
rect 175999 525045 177068 525059
rect 177103 525093 178172 525154
rect 177103 525059 177121 525093
rect 177155 525059 178121 525093
rect 178155 525059 178172 525093
rect 177103 525045 178172 525059
rect 178207 525093 179276 525154
rect 178207 525059 178225 525093
rect 178259 525059 179225 525093
rect 179259 525059 179276 525093
rect 178207 525045 179276 525059
rect 179311 525093 179829 525154
rect 179311 525059 179329 525093
rect 179363 525059 179777 525093
rect 179811 525059 179829 525093
rect 174803 525009 174861 525026
rect 173924 524896 173941 524930
rect 173975 524896 173992 524930
rect 173924 524879 173992 524896
rect 174288 524966 174358 524981
rect 174288 524932 174305 524966
rect 174339 524932 174358 524966
rect 174288 524731 174358 524932
rect 175212 524930 175280 525045
rect 175212 524896 175229 524930
rect 175263 524896 175280 524930
rect 175212 524879 175280 524896
rect 175576 524966 175646 524981
rect 175576 524932 175593 524966
rect 175627 524932 175646 524966
rect 174803 524842 174861 524877
rect 174803 524808 174815 524842
rect 174849 524808 174861 524842
rect 174803 524749 174861 524808
rect 172227 524686 172245 524720
rect 172279 524686 172417 524720
rect 172451 524686 172469 524720
rect 172227 524644 172469 524686
rect 172503 524720 173572 524731
rect 172503 524686 172521 524720
rect 172555 524686 173521 524720
rect 173555 524686 173572 524720
rect 172503 524644 173572 524686
rect 173607 524720 174676 524731
rect 173607 524686 173625 524720
rect 173659 524686 174625 524720
rect 174659 524686 174676 524720
rect 173607 524644 174676 524686
rect 174803 524715 174815 524749
rect 174849 524715 174861 524749
rect 175576 524731 175646 524932
rect 176316 524930 176384 525045
rect 176316 524896 176333 524930
rect 176367 524896 176384 524930
rect 176316 524879 176384 524896
rect 176680 524966 176750 524981
rect 176680 524932 176697 524966
rect 176731 524932 176750 524966
rect 176680 524731 176750 524932
rect 177420 524930 177488 525045
rect 177420 524896 177437 524930
rect 177471 524896 177488 524930
rect 177420 524879 177488 524896
rect 177784 524966 177854 524981
rect 177784 524932 177801 524966
rect 177835 524932 177854 524966
rect 177784 524731 177854 524932
rect 178524 524930 178592 525045
rect 179311 525000 179829 525059
rect 179955 525060 180013 525154
rect 179955 525026 179967 525060
rect 180001 525026 180013 525060
rect 180047 525093 181116 525154
rect 180047 525059 180065 525093
rect 180099 525059 181065 525093
rect 181099 525059 181116 525093
rect 180047 525045 181116 525059
rect 181151 525093 182220 525154
rect 181151 525059 181169 525093
rect 181203 525059 182169 525093
rect 182203 525059 182220 525093
rect 181151 525045 182220 525059
rect 182255 525093 183324 525154
rect 182255 525059 182273 525093
rect 182307 525059 183273 525093
rect 183307 525059 183324 525093
rect 182255 525045 183324 525059
rect 183359 525093 184428 525154
rect 183359 525059 183377 525093
rect 183411 525059 184377 525093
rect 184411 525059 184428 525093
rect 183359 525045 184428 525059
rect 184463 525093 184981 525154
rect 184463 525059 184481 525093
rect 184515 525059 184929 525093
rect 184963 525059 184981 525093
rect 179955 525009 180013 525026
rect 178524 524896 178541 524930
rect 178575 524896 178592 524930
rect 178524 524879 178592 524896
rect 178888 524966 178958 524981
rect 178888 524932 178905 524966
rect 178939 524932 178958 524966
rect 178888 524731 178958 524932
rect 179311 524930 179553 525000
rect 179311 524896 179389 524930
rect 179423 524896 179499 524930
rect 179533 524896 179553 524930
rect 179587 524932 179607 524966
rect 179641 524932 179717 524966
rect 179751 524932 179829 524966
rect 179587 524862 179829 524932
rect 180364 524930 180432 525045
rect 180364 524896 180381 524930
rect 180415 524896 180432 524930
rect 180364 524879 180432 524896
rect 180728 524966 180798 524981
rect 180728 524932 180745 524966
rect 180779 524932 180798 524966
rect 179311 524822 179829 524862
rect 179311 524788 179329 524822
rect 179363 524788 179777 524822
rect 179811 524788 179829 524822
rect 174803 524644 174861 524715
rect 174895 524720 175964 524731
rect 174895 524686 174913 524720
rect 174947 524686 175913 524720
rect 175947 524686 175964 524720
rect 174895 524644 175964 524686
rect 175999 524720 177068 524731
rect 175999 524686 176017 524720
rect 176051 524686 177017 524720
rect 177051 524686 177068 524720
rect 175999 524644 177068 524686
rect 177103 524720 178172 524731
rect 177103 524686 177121 524720
rect 177155 524686 178121 524720
rect 178155 524686 178172 524720
rect 177103 524644 178172 524686
rect 178207 524720 179276 524731
rect 178207 524686 178225 524720
rect 178259 524686 179225 524720
rect 179259 524686 179276 524720
rect 178207 524644 179276 524686
rect 179311 524720 179829 524788
rect 179311 524686 179329 524720
rect 179363 524686 179777 524720
rect 179811 524686 179829 524720
rect 179311 524644 179829 524686
rect 179955 524842 180013 524877
rect 179955 524808 179967 524842
rect 180001 524808 180013 524842
rect 179955 524749 180013 524808
rect 179955 524715 179967 524749
rect 180001 524715 180013 524749
rect 180728 524731 180798 524932
rect 181468 524930 181536 525045
rect 181468 524896 181485 524930
rect 181519 524896 181536 524930
rect 181468 524879 181536 524896
rect 181832 524966 181902 524981
rect 181832 524932 181849 524966
rect 181883 524932 181902 524966
rect 181832 524731 181902 524932
rect 182572 524930 182640 525045
rect 182572 524896 182589 524930
rect 182623 524896 182640 524930
rect 182572 524879 182640 524896
rect 182936 524966 183006 524981
rect 182936 524932 182953 524966
rect 182987 524932 183006 524966
rect 182936 524731 183006 524932
rect 183676 524930 183744 525045
rect 184463 525000 184981 525059
rect 185107 525060 185165 525154
rect 185107 525026 185119 525060
rect 185153 525026 185165 525060
rect 185199 525093 186268 525154
rect 185199 525059 185217 525093
rect 185251 525059 186217 525093
rect 186251 525059 186268 525093
rect 185199 525045 186268 525059
rect 186303 525093 187005 525154
rect 186303 525059 186321 525093
rect 186355 525059 186953 525093
rect 186987 525059 187005 525093
rect 185107 525009 185165 525026
rect 183676 524896 183693 524930
rect 183727 524896 183744 524930
rect 183676 524879 183744 524896
rect 184040 524966 184110 524981
rect 184040 524932 184057 524966
rect 184091 524932 184110 524966
rect 184040 524731 184110 524932
rect 184463 524930 184705 525000
rect 184463 524896 184541 524930
rect 184575 524896 184651 524930
rect 184685 524896 184705 524930
rect 184739 524932 184759 524966
rect 184793 524932 184869 524966
rect 184903 524932 184981 524966
rect 184739 524862 184981 524932
rect 185516 524930 185584 525045
rect 186303 525000 187005 525059
rect 187223 525091 187465 525154
rect 187223 525057 187241 525091
rect 187275 525057 187413 525091
rect 187447 525057 187465 525091
rect 187223 525004 187465 525057
rect 185516 524896 185533 524930
rect 185567 524896 185584 524930
rect 185516 524879 185584 524896
rect 185880 524966 185950 524981
rect 185880 524932 185897 524966
rect 185931 524932 185950 524966
rect 184463 524822 184981 524862
rect 184463 524788 184481 524822
rect 184515 524788 184929 524822
rect 184963 524788 184981 524822
rect 179955 524644 180013 524715
rect 180047 524720 181116 524731
rect 180047 524686 180065 524720
rect 180099 524686 181065 524720
rect 181099 524686 181116 524720
rect 180047 524644 181116 524686
rect 181151 524720 182220 524731
rect 181151 524686 181169 524720
rect 181203 524686 182169 524720
rect 182203 524686 182220 524720
rect 181151 524644 182220 524686
rect 182255 524720 183324 524731
rect 182255 524686 182273 524720
rect 182307 524686 183273 524720
rect 183307 524686 183324 524720
rect 182255 524644 183324 524686
rect 183359 524720 184428 524731
rect 183359 524686 183377 524720
rect 183411 524686 184377 524720
rect 184411 524686 184428 524720
rect 183359 524644 184428 524686
rect 184463 524720 184981 524788
rect 184463 524686 184481 524720
rect 184515 524686 184929 524720
rect 184963 524686 184981 524720
rect 184463 524644 184981 524686
rect 185107 524842 185165 524877
rect 185107 524808 185119 524842
rect 185153 524808 185165 524842
rect 185107 524749 185165 524808
rect 185107 524715 185119 524749
rect 185153 524715 185165 524749
rect 185880 524731 185950 524932
rect 186303 524930 186633 525000
rect 186303 524896 186381 524930
rect 186415 524896 186480 524930
rect 186514 524896 186579 524930
rect 186613 524896 186633 524930
rect 186667 524932 186687 524966
rect 186721 524932 186790 524966
rect 186824 524932 186893 524966
rect 186927 524932 187005 524966
rect 186667 524862 187005 524932
rect 186303 524822 187005 524862
rect 186303 524788 186321 524822
rect 186355 524788 186953 524822
rect 186987 524788 187005 524822
rect 185107 524644 185165 524715
rect 185199 524720 186268 524731
rect 185199 524686 185217 524720
rect 185251 524686 186217 524720
rect 186251 524686 186268 524720
rect 185199 524644 186268 524686
rect 186303 524720 187005 524788
rect 186303 524686 186321 524720
rect 186355 524686 186953 524720
rect 186987 524686 187005 524720
rect 186303 524644 187005 524686
rect 187223 524936 187273 524970
rect 187307 524936 187327 524970
rect 187223 524862 187327 524936
rect 187361 524930 187465 525004
rect 187361 524896 187381 524930
rect 187415 524896 187465 524930
rect 187223 524815 187465 524862
rect 187223 524781 187241 524815
rect 187275 524781 187413 524815
rect 187447 524781 187465 524815
rect 187223 524720 187465 524781
rect 187223 524686 187241 524720
rect 187275 524686 187413 524720
rect 187447 524686 187465 524720
rect 187223 524644 187465 524686
rect 172210 524610 172239 524644
rect 172273 524610 172331 524644
rect 172365 524610 172423 524644
rect 172457 524610 172515 524644
rect 172549 524610 172607 524644
rect 172641 524610 172699 524644
rect 172733 524610 172791 524644
rect 172825 524610 172883 524644
rect 172917 524610 172975 524644
rect 173009 524610 173067 524644
rect 173101 524610 173159 524644
rect 173193 524610 173251 524644
rect 173285 524610 173343 524644
rect 173377 524610 173435 524644
rect 173469 524610 173527 524644
rect 173561 524610 173619 524644
rect 173653 524610 173711 524644
rect 173745 524610 173803 524644
rect 173837 524610 173895 524644
rect 173929 524610 173987 524644
rect 174021 524610 174079 524644
rect 174113 524610 174171 524644
rect 174205 524610 174263 524644
rect 174297 524610 174355 524644
rect 174389 524610 174447 524644
rect 174481 524610 174539 524644
rect 174573 524610 174631 524644
rect 174665 524610 174723 524644
rect 174757 524610 174815 524644
rect 174849 524610 174907 524644
rect 174941 524610 174999 524644
rect 175033 524610 175091 524644
rect 175125 524610 175183 524644
rect 175217 524610 175275 524644
rect 175309 524610 175367 524644
rect 175401 524610 175459 524644
rect 175493 524610 175551 524644
rect 175585 524610 175643 524644
rect 175677 524610 175735 524644
rect 175769 524610 175827 524644
rect 175861 524610 175919 524644
rect 175953 524610 176011 524644
rect 176045 524610 176103 524644
rect 176137 524610 176195 524644
rect 176229 524610 176287 524644
rect 176321 524610 176379 524644
rect 176413 524610 176471 524644
rect 176505 524610 176563 524644
rect 176597 524610 176655 524644
rect 176689 524610 176747 524644
rect 176781 524610 176839 524644
rect 176873 524610 176931 524644
rect 176965 524610 177023 524644
rect 177057 524610 177115 524644
rect 177149 524610 177207 524644
rect 177241 524610 177299 524644
rect 177333 524610 177391 524644
rect 177425 524610 177483 524644
rect 177517 524610 177575 524644
rect 177609 524610 177667 524644
rect 177701 524610 177759 524644
rect 177793 524610 177851 524644
rect 177885 524610 177943 524644
rect 177977 524610 178035 524644
rect 178069 524610 178127 524644
rect 178161 524610 178219 524644
rect 178253 524610 178311 524644
rect 178345 524610 178403 524644
rect 178437 524610 178495 524644
rect 178529 524610 178587 524644
rect 178621 524610 178679 524644
rect 178713 524610 178771 524644
rect 178805 524610 178863 524644
rect 178897 524610 178955 524644
rect 178989 524610 179047 524644
rect 179081 524610 179139 524644
rect 179173 524610 179231 524644
rect 179265 524610 179323 524644
rect 179357 524610 179415 524644
rect 179449 524610 179507 524644
rect 179541 524610 179599 524644
rect 179633 524610 179691 524644
rect 179725 524610 179783 524644
rect 179817 524610 179875 524644
rect 179909 524610 179967 524644
rect 180001 524610 180059 524644
rect 180093 524610 180151 524644
rect 180185 524610 180243 524644
rect 180277 524610 180335 524644
rect 180369 524610 180427 524644
rect 180461 524610 180519 524644
rect 180553 524610 180611 524644
rect 180645 524610 180703 524644
rect 180737 524610 180795 524644
rect 180829 524610 180887 524644
rect 180921 524610 180979 524644
rect 181013 524610 181071 524644
rect 181105 524610 181163 524644
rect 181197 524610 181255 524644
rect 181289 524610 181347 524644
rect 181381 524610 181439 524644
rect 181473 524610 181531 524644
rect 181565 524610 181623 524644
rect 181657 524610 181715 524644
rect 181749 524610 181807 524644
rect 181841 524610 181899 524644
rect 181933 524610 181991 524644
rect 182025 524610 182083 524644
rect 182117 524610 182175 524644
rect 182209 524610 182267 524644
rect 182301 524610 182359 524644
rect 182393 524610 182451 524644
rect 182485 524610 182543 524644
rect 182577 524610 182635 524644
rect 182669 524610 182727 524644
rect 182761 524610 182819 524644
rect 182853 524610 182911 524644
rect 182945 524610 183003 524644
rect 183037 524610 183095 524644
rect 183129 524610 183187 524644
rect 183221 524610 183279 524644
rect 183313 524610 183371 524644
rect 183405 524610 183463 524644
rect 183497 524610 183555 524644
rect 183589 524610 183647 524644
rect 183681 524610 183739 524644
rect 183773 524610 183831 524644
rect 183865 524610 183923 524644
rect 183957 524610 184015 524644
rect 184049 524610 184107 524644
rect 184141 524610 184199 524644
rect 184233 524610 184291 524644
rect 184325 524610 184383 524644
rect 184417 524610 184475 524644
rect 184509 524610 184567 524644
rect 184601 524610 184659 524644
rect 184693 524610 184751 524644
rect 184785 524610 184843 524644
rect 184877 524610 184935 524644
rect 184969 524610 185027 524644
rect 185061 524610 185119 524644
rect 185153 524610 185211 524644
rect 185245 524610 185303 524644
rect 185337 524610 185395 524644
rect 185429 524610 185487 524644
rect 185521 524610 185579 524644
rect 185613 524610 185671 524644
rect 185705 524610 185763 524644
rect 185797 524610 185855 524644
rect 185889 524610 185947 524644
rect 185981 524610 186039 524644
rect 186073 524610 186131 524644
rect 186165 524610 186223 524644
rect 186257 524610 186315 524644
rect 186349 524610 186407 524644
rect 186441 524610 186499 524644
rect 186533 524610 186591 524644
rect 186625 524610 186683 524644
rect 186717 524610 186775 524644
rect 186809 524610 186867 524644
rect 186901 524610 186959 524644
rect 186993 524610 187051 524644
rect 187085 524610 187143 524644
rect 187177 524610 187235 524644
rect 187269 524610 187327 524644
rect 187361 524610 187419 524644
rect 187453 524610 187482 524644
rect 172227 524568 172469 524610
rect 172227 524534 172245 524568
rect 172279 524534 172417 524568
rect 172451 524534 172469 524568
rect 172227 524473 172469 524534
rect 172503 524568 173572 524610
rect 172503 524534 172521 524568
rect 172555 524534 173521 524568
rect 173555 524534 173572 524568
rect 172503 524523 173572 524534
rect 173607 524568 174676 524610
rect 173607 524534 173625 524568
rect 173659 524534 174625 524568
rect 174659 524534 174676 524568
rect 173607 524523 174676 524534
rect 174711 524568 175780 524610
rect 174711 524534 174729 524568
rect 174763 524534 175729 524568
rect 175763 524534 175780 524568
rect 174711 524523 175780 524534
rect 175815 524568 176884 524610
rect 175815 524534 175833 524568
rect 175867 524534 176833 524568
rect 176867 524534 176884 524568
rect 175815 524523 176884 524534
rect 176919 524568 177253 524610
rect 176919 524534 176937 524568
rect 176971 524534 177201 524568
rect 177235 524534 177253 524568
rect 172227 524439 172245 524473
rect 172279 524439 172417 524473
rect 172451 524439 172469 524473
rect 172227 524392 172469 524439
rect 172227 524324 172277 524358
rect 172311 524324 172331 524358
rect 172227 524250 172331 524324
rect 172365 524318 172469 524392
rect 172365 524284 172385 524318
rect 172419 524284 172469 524318
rect 172820 524358 172888 524375
rect 172820 524324 172837 524358
rect 172871 524324 172888 524358
rect 172227 524197 172469 524250
rect 172820 524209 172888 524324
rect 173184 524322 173254 524523
rect 173184 524288 173201 524322
rect 173235 524288 173254 524322
rect 173184 524273 173254 524288
rect 173924 524358 173992 524375
rect 173924 524324 173941 524358
rect 173975 524324 173992 524358
rect 173924 524209 173992 524324
rect 174288 524322 174358 524523
rect 174288 524288 174305 524322
rect 174339 524288 174358 524322
rect 174288 524273 174358 524288
rect 175028 524358 175096 524375
rect 175028 524324 175045 524358
rect 175079 524324 175096 524358
rect 175028 524209 175096 524324
rect 175392 524322 175462 524523
rect 175392 524288 175409 524322
rect 175443 524288 175462 524322
rect 175392 524273 175462 524288
rect 176132 524358 176200 524375
rect 176132 524324 176149 524358
rect 176183 524324 176200 524358
rect 176132 524209 176200 524324
rect 176496 524322 176566 524523
rect 176919 524466 177253 524534
rect 176919 524432 176937 524466
rect 176971 524432 177201 524466
rect 177235 524432 177253 524466
rect 176919 524392 177253 524432
rect 176496 524288 176513 524322
rect 176547 524288 176566 524322
rect 176496 524273 176566 524288
rect 176919 524324 176939 524358
rect 176973 524324 177069 524358
rect 176919 524254 177069 524324
rect 177103 524322 177253 524392
rect 177379 524539 177437 524610
rect 177379 524505 177391 524539
rect 177425 524505 177437 524539
rect 177471 524568 178540 524610
rect 177471 524534 177489 524568
rect 177523 524534 178489 524568
rect 178523 524534 178540 524568
rect 177471 524523 178540 524534
rect 178575 524568 179644 524610
rect 178575 524534 178593 524568
rect 178627 524534 179593 524568
rect 179627 524534 179644 524568
rect 178575 524523 179644 524534
rect 179679 524568 180748 524610
rect 179679 524534 179697 524568
rect 179731 524534 180697 524568
rect 180731 524534 180748 524568
rect 179679 524523 180748 524534
rect 180783 524568 181852 524610
rect 180783 524534 180801 524568
rect 180835 524534 181801 524568
rect 181835 524534 181852 524568
rect 180783 524523 181852 524534
rect 181887 524568 182405 524610
rect 181887 524534 181905 524568
rect 181939 524534 182353 524568
rect 182387 524534 182405 524568
rect 177379 524446 177437 524505
rect 177379 524412 177391 524446
rect 177425 524412 177437 524446
rect 177379 524377 177437 524412
rect 177103 524288 177199 524322
rect 177233 524288 177253 524322
rect 177788 524358 177856 524375
rect 177788 524324 177805 524358
rect 177839 524324 177856 524358
rect 172227 524163 172245 524197
rect 172279 524163 172417 524197
rect 172451 524163 172469 524197
rect 172227 524100 172469 524163
rect 172503 524195 173572 524209
rect 172503 524161 172521 524195
rect 172555 524161 173521 524195
rect 173555 524161 173572 524195
rect 172503 524100 173572 524161
rect 173607 524195 174676 524209
rect 173607 524161 173625 524195
rect 173659 524161 174625 524195
rect 174659 524161 174676 524195
rect 173607 524100 174676 524161
rect 174711 524195 175780 524209
rect 174711 524161 174729 524195
rect 174763 524161 175729 524195
rect 175763 524161 175780 524195
rect 174711 524100 175780 524161
rect 175815 524195 176884 524209
rect 175815 524161 175833 524195
rect 175867 524161 176833 524195
rect 176867 524161 176884 524195
rect 175815 524100 176884 524161
rect 176919 524202 177253 524254
rect 176919 524168 176937 524202
rect 176971 524168 177201 524202
rect 177235 524168 177253 524202
rect 176919 524100 177253 524168
rect 177379 524228 177437 524245
rect 177379 524194 177391 524228
rect 177425 524194 177437 524228
rect 177788 524209 177856 524324
rect 178152 524322 178222 524523
rect 178152 524288 178169 524322
rect 178203 524288 178222 524322
rect 178152 524273 178222 524288
rect 178892 524358 178960 524375
rect 178892 524324 178909 524358
rect 178943 524324 178960 524358
rect 178892 524209 178960 524324
rect 179256 524322 179326 524523
rect 179256 524288 179273 524322
rect 179307 524288 179326 524322
rect 179256 524273 179326 524288
rect 179996 524358 180064 524375
rect 179996 524324 180013 524358
rect 180047 524324 180064 524358
rect 179996 524209 180064 524324
rect 180360 524322 180430 524523
rect 180360 524288 180377 524322
rect 180411 524288 180430 524322
rect 180360 524273 180430 524288
rect 181100 524358 181168 524375
rect 181100 524324 181117 524358
rect 181151 524324 181168 524358
rect 181100 524209 181168 524324
rect 181464 524322 181534 524523
rect 181887 524466 182405 524534
rect 181887 524432 181905 524466
rect 181939 524432 182353 524466
rect 182387 524432 182405 524466
rect 181887 524392 182405 524432
rect 181464 524288 181481 524322
rect 181515 524288 181534 524322
rect 181464 524273 181534 524288
rect 181887 524324 181965 524358
rect 181999 524324 182075 524358
rect 182109 524324 182129 524358
rect 181887 524254 182129 524324
rect 182163 524322 182405 524392
rect 182531 524539 182589 524610
rect 182531 524505 182543 524539
rect 182577 524505 182589 524539
rect 182623 524568 183692 524610
rect 182623 524534 182641 524568
rect 182675 524534 183641 524568
rect 183675 524534 183692 524568
rect 182623 524523 183692 524534
rect 183727 524568 184796 524610
rect 183727 524534 183745 524568
rect 183779 524534 184745 524568
rect 184779 524534 184796 524568
rect 183727 524523 184796 524534
rect 184831 524568 185900 524610
rect 184831 524534 184849 524568
rect 184883 524534 185849 524568
rect 185883 524534 185900 524568
rect 184831 524523 185900 524534
rect 185935 524568 187004 524610
rect 185935 524534 185953 524568
rect 185987 524534 186953 524568
rect 186987 524534 187004 524568
rect 185935 524523 187004 524534
rect 187223 524568 187465 524610
rect 187223 524534 187241 524568
rect 187275 524534 187413 524568
rect 187447 524534 187465 524568
rect 182531 524446 182589 524505
rect 182531 524412 182543 524446
rect 182577 524412 182589 524446
rect 182531 524377 182589 524412
rect 182163 524288 182183 524322
rect 182217 524288 182293 524322
rect 182327 524288 182405 524322
rect 182940 524358 183008 524375
rect 182940 524324 182957 524358
rect 182991 524324 183008 524358
rect 177379 524100 177437 524194
rect 177471 524195 178540 524209
rect 177471 524161 177489 524195
rect 177523 524161 178489 524195
rect 178523 524161 178540 524195
rect 177471 524100 178540 524161
rect 178575 524195 179644 524209
rect 178575 524161 178593 524195
rect 178627 524161 179593 524195
rect 179627 524161 179644 524195
rect 178575 524100 179644 524161
rect 179679 524195 180748 524209
rect 179679 524161 179697 524195
rect 179731 524161 180697 524195
rect 180731 524161 180748 524195
rect 179679 524100 180748 524161
rect 180783 524195 181852 524209
rect 180783 524161 180801 524195
rect 180835 524161 181801 524195
rect 181835 524161 181852 524195
rect 180783 524100 181852 524161
rect 181887 524195 182405 524254
rect 181887 524161 181905 524195
rect 181939 524161 182353 524195
rect 182387 524161 182405 524195
rect 181887 524100 182405 524161
rect 182531 524228 182589 524245
rect 182531 524194 182543 524228
rect 182577 524194 182589 524228
rect 182940 524209 183008 524324
rect 183304 524322 183374 524523
rect 183304 524288 183321 524322
rect 183355 524288 183374 524322
rect 183304 524273 183374 524288
rect 184044 524358 184112 524375
rect 184044 524324 184061 524358
rect 184095 524324 184112 524358
rect 184044 524209 184112 524324
rect 184408 524322 184478 524523
rect 184408 524288 184425 524322
rect 184459 524288 184478 524322
rect 184408 524273 184478 524288
rect 185148 524358 185216 524375
rect 185148 524324 185165 524358
rect 185199 524324 185216 524358
rect 185148 524209 185216 524324
rect 185512 524322 185582 524523
rect 185512 524288 185529 524322
rect 185563 524288 185582 524322
rect 185512 524273 185582 524288
rect 186252 524358 186320 524375
rect 186252 524324 186269 524358
rect 186303 524324 186320 524358
rect 186252 524209 186320 524324
rect 186616 524322 186686 524523
rect 186616 524288 186633 524322
rect 186667 524288 186686 524322
rect 186616 524273 186686 524288
rect 187223 524473 187465 524534
rect 187223 524439 187241 524473
rect 187275 524439 187413 524473
rect 187447 524439 187465 524473
rect 187223 524392 187465 524439
rect 187223 524318 187327 524392
rect 187223 524284 187273 524318
rect 187307 524284 187327 524318
rect 187361 524324 187381 524358
rect 187415 524324 187465 524358
rect 187361 524250 187465 524324
rect 182531 524100 182589 524194
rect 182623 524195 183692 524209
rect 182623 524161 182641 524195
rect 182675 524161 183641 524195
rect 183675 524161 183692 524195
rect 182623 524100 183692 524161
rect 183727 524195 184796 524209
rect 183727 524161 183745 524195
rect 183779 524161 184745 524195
rect 184779 524161 184796 524195
rect 183727 524100 184796 524161
rect 184831 524195 185900 524209
rect 184831 524161 184849 524195
rect 184883 524161 185849 524195
rect 185883 524161 185900 524195
rect 184831 524100 185900 524161
rect 185935 524195 187004 524209
rect 185935 524161 185953 524195
rect 185987 524161 186953 524195
rect 186987 524161 187004 524195
rect 185935 524100 187004 524161
rect 187223 524197 187465 524250
rect 187223 524163 187241 524197
rect 187275 524163 187413 524197
rect 187447 524163 187465 524197
rect 187223 524100 187465 524163
rect 172210 524066 172239 524100
rect 172273 524066 172331 524100
rect 172365 524066 172423 524100
rect 172457 524066 172515 524100
rect 172549 524066 172607 524100
rect 172641 524066 172699 524100
rect 172733 524066 172791 524100
rect 172825 524066 172883 524100
rect 172917 524066 172975 524100
rect 173009 524066 173067 524100
rect 173101 524066 173159 524100
rect 173193 524066 173251 524100
rect 173285 524066 173343 524100
rect 173377 524066 173435 524100
rect 173469 524066 173527 524100
rect 173561 524066 173619 524100
rect 173653 524066 173711 524100
rect 173745 524066 173803 524100
rect 173837 524066 173895 524100
rect 173929 524066 173987 524100
rect 174021 524066 174079 524100
rect 174113 524066 174171 524100
rect 174205 524066 174263 524100
rect 174297 524066 174355 524100
rect 174389 524066 174447 524100
rect 174481 524066 174539 524100
rect 174573 524066 174631 524100
rect 174665 524066 174723 524100
rect 174757 524066 174815 524100
rect 174849 524066 174907 524100
rect 174941 524066 174999 524100
rect 175033 524066 175091 524100
rect 175125 524066 175183 524100
rect 175217 524066 175275 524100
rect 175309 524066 175367 524100
rect 175401 524066 175459 524100
rect 175493 524066 175551 524100
rect 175585 524066 175643 524100
rect 175677 524066 175735 524100
rect 175769 524066 175827 524100
rect 175861 524066 175919 524100
rect 175953 524066 176011 524100
rect 176045 524066 176103 524100
rect 176137 524066 176195 524100
rect 176229 524066 176287 524100
rect 176321 524066 176379 524100
rect 176413 524066 176471 524100
rect 176505 524066 176563 524100
rect 176597 524066 176655 524100
rect 176689 524066 176747 524100
rect 176781 524066 176839 524100
rect 176873 524066 176931 524100
rect 176965 524066 177023 524100
rect 177057 524066 177115 524100
rect 177149 524066 177207 524100
rect 177241 524066 177299 524100
rect 177333 524066 177391 524100
rect 177425 524066 177483 524100
rect 177517 524066 177575 524100
rect 177609 524066 177667 524100
rect 177701 524066 177759 524100
rect 177793 524066 177851 524100
rect 177885 524066 177943 524100
rect 177977 524066 178035 524100
rect 178069 524066 178127 524100
rect 178161 524066 178219 524100
rect 178253 524066 178311 524100
rect 178345 524066 178403 524100
rect 178437 524066 178495 524100
rect 178529 524066 178587 524100
rect 178621 524066 178679 524100
rect 178713 524066 178771 524100
rect 178805 524066 178863 524100
rect 178897 524066 178955 524100
rect 178989 524066 179047 524100
rect 179081 524066 179139 524100
rect 179173 524066 179231 524100
rect 179265 524066 179323 524100
rect 179357 524066 179415 524100
rect 179449 524066 179507 524100
rect 179541 524066 179599 524100
rect 179633 524066 179691 524100
rect 179725 524066 179783 524100
rect 179817 524066 179875 524100
rect 179909 524066 179967 524100
rect 180001 524066 180059 524100
rect 180093 524066 180151 524100
rect 180185 524066 180243 524100
rect 180277 524066 180335 524100
rect 180369 524066 180427 524100
rect 180461 524066 180519 524100
rect 180553 524066 180611 524100
rect 180645 524066 180703 524100
rect 180737 524066 180795 524100
rect 180829 524066 180887 524100
rect 180921 524066 180979 524100
rect 181013 524066 181071 524100
rect 181105 524066 181163 524100
rect 181197 524066 181255 524100
rect 181289 524066 181347 524100
rect 181381 524066 181439 524100
rect 181473 524066 181531 524100
rect 181565 524066 181623 524100
rect 181657 524066 181715 524100
rect 181749 524066 181807 524100
rect 181841 524066 181899 524100
rect 181933 524066 181991 524100
rect 182025 524066 182083 524100
rect 182117 524066 182175 524100
rect 182209 524066 182267 524100
rect 182301 524066 182359 524100
rect 182393 524066 182451 524100
rect 182485 524066 182543 524100
rect 182577 524066 182635 524100
rect 182669 524066 182727 524100
rect 182761 524066 182819 524100
rect 182853 524066 182911 524100
rect 182945 524066 183003 524100
rect 183037 524066 183095 524100
rect 183129 524066 183187 524100
rect 183221 524066 183279 524100
rect 183313 524066 183371 524100
rect 183405 524066 183463 524100
rect 183497 524066 183555 524100
rect 183589 524066 183647 524100
rect 183681 524066 183739 524100
rect 183773 524066 183831 524100
rect 183865 524066 183923 524100
rect 183957 524066 184015 524100
rect 184049 524066 184107 524100
rect 184141 524066 184199 524100
rect 184233 524066 184291 524100
rect 184325 524066 184383 524100
rect 184417 524066 184475 524100
rect 184509 524066 184567 524100
rect 184601 524066 184659 524100
rect 184693 524066 184751 524100
rect 184785 524066 184843 524100
rect 184877 524066 184935 524100
rect 184969 524066 185027 524100
rect 185061 524066 185119 524100
rect 185153 524066 185211 524100
rect 185245 524066 185303 524100
rect 185337 524066 185395 524100
rect 185429 524066 185487 524100
rect 185521 524066 185579 524100
rect 185613 524066 185671 524100
rect 185705 524066 185763 524100
rect 185797 524066 185855 524100
rect 185889 524066 185947 524100
rect 185981 524066 186039 524100
rect 186073 524066 186131 524100
rect 186165 524066 186223 524100
rect 186257 524066 186315 524100
rect 186349 524066 186407 524100
rect 186441 524066 186499 524100
rect 186533 524066 186591 524100
rect 186625 524066 186683 524100
rect 186717 524066 186775 524100
rect 186809 524066 186867 524100
rect 186901 524066 186959 524100
rect 186993 524066 187051 524100
rect 187085 524066 187143 524100
rect 187177 524066 187235 524100
rect 187269 524066 187327 524100
rect 187361 524066 187419 524100
rect 187453 524066 187482 524100
rect 172227 524003 172469 524066
rect 172227 523969 172245 524003
rect 172279 523969 172417 524003
rect 172451 523969 172469 524003
rect 172227 523916 172469 523969
rect 172503 524005 173572 524066
rect 172503 523971 172521 524005
rect 172555 523971 173521 524005
rect 173555 523971 173572 524005
rect 172503 523957 173572 523971
rect 173607 524005 174676 524066
rect 173607 523971 173625 524005
rect 173659 523971 174625 524005
rect 174659 523971 174676 524005
rect 173607 523957 174676 523971
rect 174803 523972 174861 524066
rect 172227 523842 172331 523916
rect 172227 523808 172277 523842
rect 172311 523808 172331 523842
rect 172365 523848 172385 523882
rect 172419 523848 172469 523882
rect 172365 523774 172469 523848
rect 172820 523842 172888 523957
rect 172820 523808 172837 523842
rect 172871 523808 172888 523842
rect 172820 523791 172888 523808
rect 173184 523878 173254 523893
rect 173184 523844 173201 523878
rect 173235 523844 173254 523878
rect 172227 523727 172469 523774
rect 172227 523693 172245 523727
rect 172279 523693 172417 523727
rect 172451 523693 172469 523727
rect 172227 523632 172469 523693
rect 173184 523643 173254 523844
rect 173924 523842 173992 523957
rect 174803 523938 174815 523972
rect 174849 523938 174861 523972
rect 174895 524005 175964 524066
rect 174895 523971 174913 524005
rect 174947 523971 175913 524005
rect 175947 523971 175964 524005
rect 174895 523957 175964 523971
rect 175999 524005 177068 524066
rect 175999 523971 176017 524005
rect 176051 523971 177017 524005
rect 177051 523971 177068 524005
rect 175999 523957 177068 523971
rect 177103 524005 178172 524066
rect 177103 523971 177121 524005
rect 177155 523971 178121 524005
rect 178155 523971 178172 524005
rect 177103 523957 178172 523971
rect 178207 524005 179276 524066
rect 178207 523971 178225 524005
rect 178259 523971 179225 524005
rect 179259 523971 179276 524005
rect 178207 523957 179276 523971
rect 179311 524005 179829 524066
rect 179311 523971 179329 524005
rect 179363 523971 179777 524005
rect 179811 523971 179829 524005
rect 174803 523921 174861 523938
rect 173924 523808 173941 523842
rect 173975 523808 173992 523842
rect 173924 523791 173992 523808
rect 174288 523878 174358 523893
rect 174288 523844 174305 523878
rect 174339 523844 174358 523878
rect 174288 523643 174358 523844
rect 175212 523842 175280 523957
rect 175212 523808 175229 523842
rect 175263 523808 175280 523842
rect 175212 523791 175280 523808
rect 175576 523878 175646 523893
rect 175576 523844 175593 523878
rect 175627 523844 175646 523878
rect 174803 523754 174861 523789
rect 174803 523720 174815 523754
rect 174849 523720 174861 523754
rect 174803 523661 174861 523720
rect 172227 523598 172245 523632
rect 172279 523598 172417 523632
rect 172451 523598 172469 523632
rect 172227 523556 172469 523598
rect 172503 523632 173572 523643
rect 172503 523598 172521 523632
rect 172555 523598 173521 523632
rect 173555 523598 173572 523632
rect 172503 523556 173572 523598
rect 173607 523632 174676 523643
rect 173607 523598 173625 523632
rect 173659 523598 174625 523632
rect 174659 523598 174676 523632
rect 173607 523556 174676 523598
rect 174803 523627 174815 523661
rect 174849 523627 174861 523661
rect 175576 523643 175646 523844
rect 176316 523842 176384 523957
rect 176316 523808 176333 523842
rect 176367 523808 176384 523842
rect 176316 523791 176384 523808
rect 176680 523878 176750 523893
rect 176680 523844 176697 523878
rect 176731 523844 176750 523878
rect 176680 523643 176750 523844
rect 177420 523842 177488 523957
rect 177420 523808 177437 523842
rect 177471 523808 177488 523842
rect 177420 523791 177488 523808
rect 177784 523878 177854 523893
rect 177784 523844 177801 523878
rect 177835 523844 177854 523878
rect 177784 523643 177854 523844
rect 178524 523842 178592 523957
rect 179311 523912 179829 523971
rect 179955 523972 180013 524066
rect 179955 523938 179967 523972
rect 180001 523938 180013 523972
rect 180047 524005 181116 524066
rect 180047 523971 180065 524005
rect 180099 523971 181065 524005
rect 181099 523971 181116 524005
rect 180047 523957 181116 523971
rect 181151 524005 182220 524066
rect 181151 523971 181169 524005
rect 181203 523971 182169 524005
rect 182203 523971 182220 524005
rect 181151 523957 182220 523971
rect 182255 524005 183324 524066
rect 182255 523971 182273 524005
rect 182307 523971 183273 524005
rect 183307 523971 183324 524005
rect 182255 523957 183324 523971
rect 183359 524005 184428 524066
rect 183359 523971 183377 524005
rect 183411 523971 184377 524005
rect 184411 523971 184428 524005
rect 183359 523957 184428 523971
rect 184463 524005 184981 524066
rect 184463 523971 184481 524005
rect 184515 523971 184929 524005
rect 184963 523971 184981 524005
rect 179955 523921 180013 523938
rect 178524 523808 178541 523842
rect 178575 523808 178592 523842
rect 178524 523791 178592 523808
rect 178888 523878 178958 523893
rect 178888 523844 178905 523878
rect 178939 523844 178958 523878
rect 178888 523643 178958 523844
rect 179311 523842 179553 523912
rect 179311 523808 179389 523842
rect 179423 523808 179499 523842
rect 179533 523808 179553 523842
rect 179587 523844 179607 523878
rect 179641 523844 179717 523878
rect 179751 523844 179829 523878
rect 179587 523774 179829 523844
rect 180364 523842 180432 523957
rect 180364 523808 180381 523842
rect 180415 523808 180432 523842
rect 180364 523791 180432 523808
rect 180728 523878 180798 523893
rect 180728 523844 180745 523878
rect 180779 523844 180798 523878
rect 179311 523734 179829 523774
rect 179311 523700 179329 523734
rect 179363 523700 179777 523734
rect 179811 523700 179829 523734
rect 174803 523556 174861 523627
rect 174895 523632 175964 523643
rect 174895 523598 174913 523632
rect 174947 523598 175913 523632
rect 175947 523598 175964 523632
rect 174895 523556 175964 523598
rect 175999 523632 177068 523643
rect 175999 523598 176017 523632
rect 176051 523598 177017 523632
rect 177051 523598 177068 523632
rect 175999 523556 177068 523598
rect 177103 523632 178172 523643
rect 177103 523598 177121 523632
rect 177155 523598 178121 523632
rect 178155 523598 178172 523632
rect 177103 523556 178172 523598
rect 178207 523632 179276 523643
rect 178207 523598 178225 523632
rect 178259 523598 179225 523632
rect 179259 523598 179276 523632
rect 178207 523556 179276 523598
rect 179311 523632 179829 523700
rect 179311 523598 179329 523632
rect 179363 523598 179777 523632
rect 179811 523598 179829 523632
rect 179311 523556 179829 523598
rect 179955 523754 180013 523789
rect 179955 523720 179967 523754
rect 180001 523720 180013 523754
rect 179955 523661 180013 523720
rect 179955 523627 179967 523661
rect 180001 523627 180013 523661
rect 180728 523643 180798 523844
rect 181468 523842 181536 523957
rect 181468 523808 181485 523842
rect 181519 523808 181536 523842
rect 181468 523791 181536 523808
rect 181832 523878 181902 523893
rect 181832 523844 181849 523878
rect 181883 523844 181902 523878
rect 181832 523643 181902 523844
rect 182572 523842 182640 523957
rect 182572 523808 182589 523842
rect 182623 523808 182640 523842
rect 182572 523791 182640 523808
rect 182936 523878 183006 523893
rect 182936 523844 182953 523878
rect 182987 523844 183006 523878
rect 182936 523643 183006 523844
rect 183676 523842 183744 523957
rect 184463 523912 184981 523971
rect 185107 523972 185165 524066
rect 185107 523938 185119 523972
rect 185153 523938 185165 523972
rect 185199 524005 186268 524066
rect 185199 523971 185217 524005
rect 185251 523971 186217 524005
rect 186251 523971 186268 524005
rect 185199 523957 186268 523971
rect 186303 524005 187005 524066
rect 186303 523971 186321 524005
rect 186355 523971 186953 524005
rect 186987 523971 187005 524005
rect 185107 523921 185165 523938
rect 183676 523808 183693 523842
rect 183727 523808 183744 523842
rect 183676 523791 183744 523808
rect 184040 523878 184110 523893
rect 184040 523844 184057 523878
rect 184091 523844 184110 523878
rect 184040 523643 184110 523844
rect 184463 523842 184705 523912
rect 184463 523808 184541 523842
rect 184575 523808 184651 523842
rect 184685 523808 184705 523842
rect 184739 523844 184759 523878
rect 184793 523844 184869 523878
rect 184903 523844 184981 523878
rect 184739 523774 184981 523844
rect 185516 523842 185584 523957
rect 186303 523912 187005 523971
rect 187223 524003 187465 524066
rect 187223 523969 187241 524003
rect 187275 523969 187413 524003
rect 187447 523969 187465 524003
rect 187223 523916 187465 523969
rect 185516 523808 185533 523842
rect 185567 523808 185584 523842
rect 185516 523791 185584 523808
rect 185880 523878 185950 523893
rect 185880 523844 185897 523878
rect 185931 523844 185950 523878
rect 184463 523734 184981 523774
rect 184463 523700 184481 523734
rect 184515 523700 184929 523734
rect 184963 523700 184981 523734
rect 179955 523556 180013 523627
rect 180047 523632 181116 523643
rect 180047 523598 180065 523632
rect 180099 523598 181065 523632
rect 181099 523598 181116 523632
rect 180047 523556 181116 523598
rect 181151 523632 182220 523643
rect 181151 523598 181169 523632
rect 181203 523598 182169 523632
rect 182203 523598 182220 523632
rect 181151 523556 182220 523598
rect 182255 523632 183324 523643
rect 182255 523598 182273 523632
rect 182307 523598 183273 523632
rect 183307 523598 183324 523632
rect 182255 523556 183324 523598
rect 183359 523632 184428 523643
rect 183359 523598 183377 523632
rect 183411 523598 184377 523632
rect 184411 523598 184428 523632
rect 183359 523556 184428 523598
rect 184463 523632 184981 523700
rect 184463 523598 184481 523632
rect 184515 523598 184929 523632
rect 184963 523598 184981 523632
rect 184463 523556 184981 523598
rect 185107 523754 185165 523789
rect 185107 523720 185119 523754
rect 185153 523720 185165 523754
rect 185107 523661 185165 523720
rect 185107 523627 185119 523661
rect 185153 523627 185165 523661
rect 185880 523643 185950 523844
rect 186303 523842 186633 523912
rect 186303 523808 186381 523842
rect 186415 523808 186480 523842
rect 186514 523808 186579 523842
rect 186613 523808 186633 523842
rect 186667 523844 186687 523878
rect 186721 523844 186790 523878
rect 186824 523844 186893 523878
rect 186927 523844 187005 523878
rect 186667 523774 187005 523844
rect 186303 523734 187005 523774
rect 186303 523700 186321 523734
rect 186355 523700 186953 523734
rect 186987 523700 187005 523734
rect 185107 523556 185165 523627
rect 185199 523632 186268 523643
rect 185199 523598 185217 523632
rect 185251 523598 186217 523632
rect 186251 523598 186268 523632
rect 185199 523556 186268 523598
rect 186303 523632 187005 523700
rect 186303 523598 186321 523632
rect 186355 523598 186953 523632
rect 186987 523598 187005 523632
rect 186303 523556 187005 523598
rect 187223 523848 187273 523882
rect 187307 523848 187327 523882
rect 187223 523774 187327 523848
rect 187361 523842 187465 523916
rect 187361 523808 187381 523842
rect 187415 523808 187465 523842
rect 187223 523727 187465 523774
rect 187223 523693 187241 523727
rect 187275 523693 187413 523727
rect 187447 523693 187465 523727
rect 187223 523632 187465 523693
rect 187223 523598 187241 523632
rect 187275 523598 187413 523632
rect 187447 523598 187465 523632
rect 187223 523556 187465 523598
rect 172210 523522 172239 523556
rect 172273 523522 172331 523556
rect 172365 523522 172423 523556
rect 172457 523522 172515 523556
rect 172549 523522 172607 523556
rect 172641 523522 172699 523556
rect 172733 523522 172791 523556
rect 172825 523522 172883 523556
rect 172917 523522 172975 523556
rect 173009 523522 173067 523556
rect 173101 523522 173159 523556
rect 173193 523522 173251 523556
rect 173285 523522 173343 523556
rect 173377 523522 173435 523556
rect 173469 523522 173527 523556
rect 173561 523522 173619 523556
rect 173653 523522 173711 523556
rect 173745 523522 173803 523556
rect 173837 523522 173895 523556
rect 173929 523522 173987 523556
rect 174021 523522 174079 523556
rect 174113 523522 174171 523556
rect 174205 523522 174263 523556
rect 174297 523522 174355 523556
rect 174389 523522 174447 523556
rect 174481 523522 174539 523556
rect 174573 523522 174631 523556
rect 174665 523522 174723 523556
rect 174757 523522 174815 523556
rect 174849 523522 174907 523556
rect 174941 523522 174999 523556
rect 175033 523522 175091 523556
rect 175125 523522 175183 523556
rect 175217 523522 175275 523556
rect 175309 523522 175367 523556
rect 175401 523522 175459 523556
rect 175493 523522 175551 523556
rect 175585 523522 175643 523556
rect 175677 523522 175735 523556
rect 175769 523522 175827 523556
rect 175861 523522 175919 523556
rect 175953 523522 176011 523556
rect 176045 523522 176103 523556
rect 176137 523522 176195 523556
rect 176229 523522 176287 523556
rect 176321 523522 176379 523556
rect 176413 523522 176471 523556
rect 176505 523522 176563 523556
rect 176597 523522 176655 523556
rect 176689 523522 176747 523556
rect 176781 523522 176839 523556
rect 176873 523522 176931 523556
rect 176965 523522 177023 523556
rect 177057 523522 177115 523556
rect 177149 523522 177207 523556
rect 177241 523522 177299 523556
rect 177333 523522 177391 523556
rect 177425 523522 177483 523556
rect 177517 523522 177575 523556
rect 177609 523522 177667 523556
rect 177701 523522 177759 523556
rect 177793 523522 177851 523556
rect 177885 523522 177943 523556
rect 177977 523522 178035 523556
rect 178069 523522 178127 523556
rect 178161 523522 178219 523556
rect 178253 523522 178311 523556
rect 178345 523522 178403 523556
rect 178437 523522 178495 523556
rect 178529 523522 178587 523556
rect 178621 523522 178679 523556
rect 178713 523522 178771 523556
rect 178805 523522 178863 523556
rect 178897 523522 178955 523556
rect 178989 523522 179047 523556
rect 179081 523522 179139 523556
rect 179173 523522 179231 523556
rect 179265 523522 179323 523556
rect 179357 523522 179415 523556
rect 179449 523522 179507 523556
rect 179541 523522 179599 523556
rect 179633 523522 179691 523556
rect 179725 523522 179783 523556
rect 179817 523522 179875 523556
rect 179909 523522 179967 523556
rect 180001 523522 180059 523556
rect 180093 523522 180151 523556
rect 180185 523522 180243 523556
rect 180277 523522 180335 523556
rect 180369 523522 180427 523556
rect 180461 523522 180519 523556
rect 180553 523522 180611 523556
rect 180645 523522 180703 523556
rect 180737 523522 180795 523556
rect 180829 523522 180887 523556
rect 180921 523522 180979 523556
rect 181013 523522 181071 523556
rect 181105 523522 181163 523556
rect 181197 523522 181255 523556
rect 181289 523522 181347 523556
rect 181381 523522 181439 523556
rect 181473 523522 181531 523556
rect 181565 523522 181623 523556
rect 181657 523522 181715 523556
rect 181749 523522 181807 523556
rect 181841 523522 181899 523556
rect 181933 523522 181991 523556
rect 182025 523522 182083 523556
rect 182117 523522 182175 523556
rect 182209 523522 182267 523556
rect 182301 523522 182359 523556
rect 182393 523522 182451 523556
rect 182485 523522 182543 523556
rect 182577 523522 182635 523556
rect 182669 523522 182727 523556
rect 182761 523522 182819 523556
rect 182853 523522 182911 523556
rect 182945 523522 183003 523556
rect 183037 523522 183095 523556
rect 183129 523522 183187 523556
rect 183221 523522 183279 523556
rect 183313 523522 183371 523556
rect 183405 523522 183463 523556
rect 183497 523522 183555 523556
rect 183589 523522 183647 523556
rect 183681 523522 183739 523556
rect 183773 523522 183831 523556
rect 183865 523522 183923 523556
rect 183957 523522 184015 523556
rect 184049 523522 184107 523556
rect 184141 523522 184199 523556
rect 184233 523522 184291 523556
rect 184325 523522 184383 523556
rect 184417 523522 184475 523556
rect 184509 523522 184567 523556
rect 184601 523522 184659 523556
rect 184693 523522 184751 523556
rect 184785 523522 184843 523556
rect 184877 523522 184935 523556
rect 184969 523522 185027 523556
rect 185061 523522 185119 523556
rect 185153 523522 185211 523556
rect 185245 523522 185303 523556
rect 185337 523522 185395 523556
rect 185429 523522 185487 523556
rect 185521 523522 185579 523556
rect 185613 523522 185671 523556
rect 185705 523522 185763 523556
rect 185797 523522 185855 523556
rect 185889 523522 185947 523556
rect 185981 523522 186039 523556
rect 186073 523522 186131 523556
rect 186165 523522 186223 523556
rect 186257 523522 186315 523556
rect 186349 523522 186407 523556
rect 186441 523522 186499 523556
rect 186533 523522 186591 523556
rect 186625 523522 186683 523556
rect 186717 523522 186775 523556
rect 186809 523522 186867 523556
rect 186901 523522 186959 523556
rect 186993 523522 187051 523556
rect 187085 523522 187143 523556
rect 187177 523522 187235 523556
rect 187269 523522 187327 523556
rect 187361 523522 187419 523556
rect 187453 523522 187482 523556
rect 172227 523480 172469 523522
rect 172227 523446 172245 523480
rect 172279 523446 172417 523480
rect 172451 523446 172469 523480
rect 172227 523385 172469 523446
rect 172503 523480 173572 523522
rect 172503 523446 172521 523480
rect 172555 523446 173521 523480
rect 173555 523446 173572 523480
rect 172503 523435 173572 523446
rect 173607 523480 174676 523522
rect 173607 523446 173625 523480
rect 173659 523446 174625 523480
rect 174659 523446 174676 523480
rect 173607 523435 174676 523446
rect 174711 523480 175780 523522
rect 174711 523446 174729 523480
rect 174763 523446 175729 523480
rect 175763 523446 175780 523480
rect 174711 523435 175780 523446
rect 175815 523480 176884 523522
rect 175815 523446 175833 523480
rect 175867 523446 176833 523480
rect 176867 523446 176884 523480
rect 175815 523435 176884 523446
rect 176919 523480 177253 523522
rect 176919 523446 176937 523480
rect 176971 523446 177201 523480
rect 177235 523446 177253 523480
rect 172227 523351 172245 523385
rect 172279 523351 172417 523385
rect 172451 523351 172469 523385
rect 172227 523304 172469 523351
rect 172227 523236 172277 523270
rect 172311 523236 172331 523270
rect 172227 523162 172331 523236
rect 172365 523230 172469 523304
rect 172365 523196 172385 523230
rect 172419 523196 172469 523230
rect 172820 523270 172888 523287
rect 172820 523236 172837 523270
rect 172871 523236 172888 523270
rect 172227 523109 172469 523162
rect 172820 523121 172888 523236
rect 173184 523234 173254 523435
rect 173184 523200 173201 523234
rect 173235 523200 173254 523234
rect 173184 523185 173254 523200
rect 173924 523270 173992 523287
rect 173924 523236 173941 523270
rect 173975 523236 173992 523270
rect 173924 523121 173992 523236
rect 174288 523234 174358 523435
rect 174288 523200 174305 523234
rect 174339 523200 174358 523234
rect 174288 523185 174358 523200
rect 175028 523270 175096 523287
rect 175028 523236 175045 523270
rect 175079 523236 175096 523270
rect 175028 523121 175096 523236
rect 175392 523234 175462 523435
rect 175392 523200 175409 523234
rect 175443 523200 175462 523234
rect 175392 523185 175462 523200
rect 176132 523270 176200 523287
rect 176132 523236 176149 523270
rect 176183 523236 176200 523270
rect 176132 523121 176200 523236
rect 176496 523234 176566 523435
rect 176919 523378 177253 523446
rect 176919 523344 176937 523378
rect 176971 523344 177201 523378
rect 177235 523344 177253 523378
rect 176919 523304 177253 523344
rect 176496 523200 176513 523234
rect 176547 523200 176566 523234
rect 176496 523185 176566 523200
rect 176919 523236 176939 523270
rect 176973 523236 177069 523270
rect 176919 523166 177069 523236
rect 177103 523234 177253 523304
rect 177379 523451 177437 523522
rect 177379 523417 177391 523451
rect 177425 523417 177437 523451
rect 177471 523480 178540 523522
rect 177471 523446 177489 523480
rect 177523 523446 178489 523480
rect 178523 523446 178540 523480
rect 177471 523435 178540 523446
rect 178575 523480 179644 523522
rect 178575 523446 178593 523480
rect 178627 523446 179593 523480
rect 179627 523446 179644 523480
rect 178575 523435 179644 523446
rect 179679 523480 180748 523522
rect 179679 523446 179697 523480
rect 179731 523446 180697 523480
rect 180731 523446 180748 523480
rect 179679 523435 180748 523446
rect 180783 523480 181852 523522
rect 180783 523446 180801 523480
rect 180835 523446 181801 523480
rect 181835 523446 181852 523480
rect 180783 523435 181852 523446
rect 181887 523480 182405 523522
rect 181887 523446 181905 523480
rect 181939 523446 182353 523480
rect 182387 523446 182405 523480
rect 177379 523358 177437 523417
rect 177379 523324 177391 523358
rect 177425 523324 177437 523358
rect 177379 523289 177437 523324
rect 177103 523200 177199 523234
rect 177233 523200 177253 523234
rect 177788 523270 177856 523287
rect 177788 523236 177805 523270
rect 177839 523236 177856 523270
rect 172227 523075 172245 523109
rect 172279 523075 172417 523109
rect 172451 523075 172469 523109
rect 172227 523012 172469 523075
rect 172503 523107 173572 523121
rect 172503 523073 172521 523107
rect 172555 523073 173521 523107
rect 173555 523073 173572 523107
rect 172503 523012 173572 523073
rect 173607 523107 174676 523121
rect 173607 523073 173625 523107
rect 173659 523073 174625 523107
rect 174659 523073 174676 523107
rect 173607 523012 174676 523073
rect 174711 523107 175780 523121
rect 174711 523073 174729 523107
rect 174763 523073 175729 523107
rect 175763 523073 175780 523107
rect 174711 523012 175780 523073
rect 175815 523107 176884 523121
rect 175815 523073 175833 523107
rect 175867 523073 176833 523107
rect 176867 523073 176884 523107
rect 175815 523012 176884 523073
rect 176919 523114 177253 523166
rect 176919 523080 176937 523114
rect 176971 523080 177201 523114
rect 177235 523080 177253 523114
rect 176919 523012 177253 523080
rect 177379 523140 177437 523157
rect 177379 523106 177391 523140
rect 177425 523106 177437 523140
rect 177788 523121 177856 523236
rect 178152 523234 178222 523435
rect 178152 523200 178169 523234
rect 178203 523200 178222 523234
rect 178152 523185 178222 523200
rect 178892 523270 178960 523287
rect 178892 523236 178909 523270
rect 178943 523236 178960 523270
rect 178892 523121 178960 523236
rect 179256 523234 179326 523435
rect 179256 523200 179273 523234
rect 179307 523200 179326 523234
rect 179256 523185 179326 523200
rect 179996 523270 180064 523287
rect 179996 523236 180013 523270
rect 180047 523236 180064 523270
rect 179996 523121 180064 523236
rect 180360 523234 180430 523435
rect 180360 523200 180377 523234
rect 180411 523200 180430 523234
rect 180360 523185 180430 523200
rect 181100 523270 181168 523287
rect 181100 523236 181117 523270
rect 181151 523236 181168 523270
rect 181100 523121 181168 523236
rect 181464 523234 181534 523435
rect 181887 523378 182405 523446
rect 181887 523344 181905 523378
rect 181939 523344 182353 523378
rect 182387 523344 182405 523378
rect 181887 523304 182405 523344
rect 181464 523200 181481 523234
rect 181515 523200 181534 523234
rect 181464 523185 181534 523200
rect 181887 523236 181965 523270
rect 181999 523236 182075 523270
rect 182109 523236 182129 523270
rect 181887 523166 182129 523236
rect 182163 523234 182405 523304
rect 182531 523451 182589 523522
rect 182531 523417 182543 523451
rect 182577 523417 182589 523451
rect 182623 523480 183692 523522
rect 182623 523446 182641 523480
rect 182675 523446 183641 523480
rect 183675 523446 183692 523480
rect 182623 523435 183692 523446
rect 183727 523480 184796 523522
rect 183727 523446 183745 523480
rect 183779 523446 184745 523480
rect 184779 523446 184796 523480
rect 183727 523435 184796 523446
rect 184831 523480 185900 523522
rect 184831 523446 184849 523480
rect 184883 523446 185849 523480
rect 185883 523446 185900 523480
rect 184831 523435 185900 523446
rect 185935 523480 187004 523522
rect 185935 523446 185953 523480
rect 185987 523446 186953 523480
rect 186987 523446 187004 523480
rect 185935 523435 187004 523446
rect 187223 523480 187465 523522
rect 187223 523446 187241 523480
rect 187275 523446 187413 523480
rect 187447 523446 187465 523480
rect 182531 523358 182589 523417
rect 182531 523324 182543 523358
rect 182577 523324 182589 523358
rect 182531 523289 182589 523324
rect 182163 523200 182183 523234
rect 182217 523200 182293 523234
rect 182327 523200 182405 523234
rect 182940 523270 183008 523287
rect 182940 523236 182957 523270
rect 182991 523236 183008 523270
rect 177379 523012 177437 523106
rect 177471 523107 178540 523121
rect 177471 523073 177489 523107
rect 177523 523073 178489 523107
rect 178523 523073 178540 523107
rect 177471 523012 178540 523073
rect 178575 523107 179644 523121
rect 178575 523073 178593 523107
rect 178627 523073 179593 523107
rect 179627 523073 179644 523107
rect 178575 523012 179644 523073
rect 179679 523107 180748 523121
rect 179679 523073 179697 523107
rect 179731 523073 180697 523107
rect 180731 523073 180748 523107
rect 179679 523012 180748 523073
rect 180783 523107 181852 523121
rect 180783 523073 180801 523107
rect 180835 523073 181801 523107
rect 181835 523073 181852 523107
rect 180783 523012 181852 523073
rect 181887 523107 182405 523166
rect 181887 523073 181905 523107
rect 181939 523073 182353 523107
rect 182387 523073 182405 523107
rect 181887 523012 182405 523073
rect 182531 523140 182589 523157
rect 182531 523106 182543 523140
rect 182577 523106 182589 523140
rect 182940 523121 183008 523236
rect 183304 523234 183374 523435
rect 183304 523200 183321 523234
rect 183355 523200 183374 523234
rect 183304 523185 183374 523200
rect 184044 523270 184112 523287
rect 184044 523236 184061 523270
rect 184095 523236 184112 523270
rect 184044 523121 184112 523236
rect 184408 523234 184478 523435
rect 184408 523200 184425 523234
rect 184459 523200 184478 523234
rect 184408 523185 184478 523200
rect 185148 523270 185216 523287
rect 185148 523236 185165 523270
rect 185199 523236 185216 523270
rect 185148 523121 185216 523236
rect 185512 523234 185582 523435
rect 185512 523200 185529 523234
rect 185563 523200 185582 523234
rect 185512 523185 185582 523200
rect 186252 523270 186320 523287
rect 186252 523236 186269 523270
rect 186303 523236 186320 523270
rect 186252 523121 186320 523236
rect 186616 523234 186686 523435
rect 186616 523200 186633 523234
rect 186667 523200 186686 523234
rect 186616 523185 186686 523200
rect 187223 523385 187465 523446
rect 187223 523351 187241 523385
rect 187275 523351 187413 523385
rect 187447 523351 187465 523385
rect 187223 523304 187465 523351
rect 187223 523230 187327 523304
rect 187223 523196 187273 523230
rect 187307 523196 187327 523230
rect 187361 523236 187381 523270
rect 187415 523236 187465 523270
rect 187361 523162 187465 523236
rect 182531 523012 182589 523106
rect 182623 523107 183692 523121
rect 182623 523073 182641 523107
rect 182675 523073 183641 523107
rect 183675 523073 183692 523107
rect 182623 523012 183692 523073
rect 183727 523107 184796 523121
rect 183727 523073 183745 523107
rect 183779 523073 184745 523107
rect 184779 523073 184796 523107
rect 183727 523012 184796 523073
rect 184831 523107 185900 523121
rect 184831 523073 184849 523107
rect 184883 523073 185849 523107
rect 185883 523073 185900 523107
rect 184831 523012 185900 523073
rect 185935 523107 187004 523121
rect 185935 523073 185953 523107
rect 185987 523073 186953 523107
rect 186987 523073 187004 523107
rect 185935 523012 187004 523073
rect 187223 523109 187465 523162
rect 187223 523075 187241 523109
rect 187275 523075 187413 523109
rect 187447 523075 187465 523109
rect 187223 523012 187465 523075
rect 172210 522978 172239 523012
rect 172273 522978 172331 523012
rect 172365 522978 172423 523012
rect 172457 522978 172515 523012
rect 172549 522978 172607 523012
rect 172641 522978 172699 523012
rect 172733 522978 172791 523012
rect 172825 522978 172883 523012
rect 172917 522978 172975 523012
rect 173009 522978 173067 523012
rect 173101 522978 173159 523012
rect 173193 522978 173251 523012
rect 173285 522978 173343 523012
rect 173377 522978 173435 523012
rect 173469 522978 173527 523012
rect 173561 522978 173619 523012
rect 173653 522978 173711 523012
rect 173745 522978 173803 523012
rect 173837 522978 173895 523012
rect 173929 522978 173987 523012
rect 174021 522978 174079 523012
rect 174113 522978 174171 523012
rect 174205 522978 174263 523012
rect 174297 522978 174355 523012
rect 174389 522978 174447 523012
rect 174481 522978 174539 523012
rect 174573 522978 174631 523012
rect 174665 522978 174723 523012
rect 174757 522978 174815 523012
rect 174849 522978 174907 523012
rect 174941 522978 174999 523012
rect 175033 522978 175091 523012
rect 175125 522978 175183 523012
rect 175217 522978 175275 523012
rect 175309 522978 175367 523012
rect 175401 522978 175459 523012
rect 175493 522978 175551 523012
rect 175585 522978 175643 523012
rect 175677 522978 175735 523012
rect 175769 522978 175827 523012
rect 175861 522978 175919 523012
rect 175953 522978 176011 523012
rect 176045 522978 176103 523012
rect 176137 522978 176195 523012
rect 176229 522978 176287 523012
rect 176321 522978 176379 523012
rect 176413 522978 176471 523012
rect 176505 522978 176563 523012
rect 176597 522978 176655 523012
rect 176689 522978 176747 523012
rect 176781 522978 176839 523012
rect 176873 522978 176931 523012
rect 176965 522978 177023 523012
rect 177057 522978 177115 523012
rect 177149 522978 177207 523012
rect 177241 522978 177299 523012
rect 177333 522978 177391 523012
rect 177425 522978 177483 523012
rect 177517 522978 177575 523012
rect 177609 522978 177667 523012
rect 177701 522978 177759 523012
rect 177793 522978 177851 523012
rect 177885 522978 177943 523012
rect 177977 522978 178035 523012
rect 178069 522978 178127 523012
rect 178161 522978 178219 523012
rect 178253 522978 178311 523012
rect 178345 522978 178403 523012
rect 178437 522978 178495 523012
rect 178529 522978 178587 523012
rect 178621 522978 178679 523012
rect 178713 522978 178771 523012
rect 178805 522978 178863 523012
rect 178897 522978 178955 523012
rect 178989 522978 179047 523012
rect 179081 522978 179139 523012
rect 179173 522978 179231 523012
rect 179265 522978 179323 523012
rect 179357 522978 179415 523012
rect 179449 522978 179507 523012
rect 179541 522978 179599 523012
rect 179633 522978 179691 523012
rect 179725 522978 179783 523012
rect 179817 522978 179875 523012
rect 179909 522978 179967 523012
rect 180001 522978 180059 523012
rect 180093 522978 180151 523012
rect 180185 522978 180243 523012
rect 180277 522978 180335 523012
rect 180369 522978 180427 523012
rect 180461 522978 180519 523012
rect 180553 522978 180611 523012
rect 180645 522978 180703 523012
rect 180737 522978 180795 523012
rect 180829 522978 180887 523012
rect 180921 522978 180979 523012
rect 181013 522978 181071 523012
rect 181105 522978 181163 523012
rect 181197 522978 181255 523012
rect 181289 522978 181347 523012
rect 181381 522978 181439 523012
rect 181473 522978 181531 523012
rect 181565 522978 181623 523012
rect 181657 522978 181715 523012
rect 181749 522978 181807 523012
rect 181841 522978 181899 523012
rect 181933 522978 181991 523012
rect 182025 522978 182083 523012
rect 182117 522978 182175 523012
rect 182209 522978 182267 523012
rect 182301 522978 182359 523012
rect 182393 522978 182451 523012
rect 182485 522978 182543 523012
rect 182577 522978 182635 523012
rect 182669 522978 182727 523012
rect 182761 522978 182819 523012
rect 182853 522978 182911 523012
rect 182945 522978 183003 523012
rect 183037 522978 183095 523012
rect 183129 522978 183187 523012
rect 183221 522978 183279 523012
rect 183313 522978 183371 523012
rect 183405 522978 183463 523012
rect 183497 522978 183555 523012
rect 183589 522978 183647 523012
rect 183681 522978 183739 523012
rect 183773 522978 183831 523012
rect 183865 522978 183923 523012
rect 183957 522978 184015 523012
rect 184049 522978 184107 523012
rect 184141 522978 184199 523012
rect 184233 522978 184291 523012
rect 184325 522978 184383 523012
rect 184417 522978 184475 523012
rect 184509 522978 184567 523012
rect 184601 522978 184659 523012
rect 184693 522978 184751 523012
rect 184785 522978 184843 523012
rect 184877 522978 184935 523012
rect 184969 522978 185027 523012
rect 185061 522978 185119 523012
rect 185153 522978 185211 523012
rect 185245 522978 185303 523012
rect 185337 522978 185395 523012
rect 185429 522978 185487 523012
rect 185521 522978 185579 523012
rect 185613 522978 185671 523012
rect 185705 522978 185763 523012
rect 185797 522978 185855 523012
rect 185889 522978 185947 523012
rect 185981 522978 186039 523012
rect 186073 522978 186131 523012
rect 186165 522978 186223 523012
rect 186257 522978 186315 523012
rect 186349 522978 186407 523012
rect 186441 522978 186499 523012
rect 186533 522978 186591 523012
rect 186625 522978 186683 523012
rect 186717 522978 186775 523012
rect 186809 522978 186867 523012
rect 186901 522978 186959 523012
rect 186993 522978 187051 523012
rect 187085 522978 187143 523012
rect 187177 522978 187235 523012
rect 187269 522978 187327 523012
rect 187361 522978 187419 523012
rect 187453 522978 187482 523012
rect 172227 522915 172469 522978
rect 172227 522881 172245 522915
rect 172279 522881 172417 522915
rect 172451 522881 172469 522915
rect 172227 522828 172469 522881
rect 172503 522917 173572 522978
rect 172503 522883 172521 522917
rect 172555 522883 173521 522917
rect 173555 522883 173572 522917
rect 172503 522869 173572 522883
rect 173607 522917 174676 522978
rect 173607 522883 173625 522917
rect 173659 522883 174625 522917
rect 174659 522883 174676 522917
rect 173607 522869 174676 522883
rect 174803 522884 174861 522978
rect 172227 522754 172331 522828
rect 172227 522720 172277 522754
rect 172311 522720 172331 522754
rect 172365 522760 172385 522794
rect 172419 522760 172469 522794
rect 172365 522686 172469 522760
rect 172820 522754 172888 522869
rect 172820 522720 172837 522754
rect 172871 522720 172888 522754
rect 172820 522703 172888 522720
rect 173184 522790 173254 522805
rect 173184 522756 173201 522790
rect 173235 522756 173254 522790
rect 172227 522639 172469 522686
rect 172227 522605 172245 522639
rect 172279 522605 172417 522639
rect 172451 522605 172469 522639
rect 172227 522544 172469 522605
rect 173184 522555 173254 522756
rect 173924 522754 173992 522869
rect 174803 522850 174815 522884
rect 174849 522850 174861 522884
rect 174895 522917 175964 522978
rect 174895 522883 174913 522917
rect 174947 522883 175913 522917
rect 175947 522883 175964 522917
rect 174895 522869 175964 522883
rect 175999 522917 177068 522978
rect 175999 522883 176017 522917
rect 176051 522883 177017 522917
rect 177051 522883 177068 522917
rect 175999 522869 177068 522883
rect 177103 522917 178172 522978
rect 177103 522883 177121 522917
rect 177155 522883 178121 522917
rect 178155 522883 178172 522917
rect 177103 522869 178172 522883
rect 178207 522917 179276 522978
rect 178207 522883 178225 522917
rect 178259 522883 179225 522917
rect 179259 522883 179276 522917
rect 178207 522869 179276 522883
rect 179311 522917 179829 522978
rect 179311 522883 179329 522917
rect 179363 522883 179777 522917
rect 179811 522883 179829 522917
rect 174803 522833 174861 522850
rect 173924 522720 173941 522754
rect 173975 522720 173992 522754
rect 173924 522703 173992 522720
rect 174288 522790 174358 522805
rect 174288 522756 174305 522790
rect 174339 522756 174358 522790
rect 174288 522555 174358 522756
rect 175212 522754 175280 522869
rect 175212 522720 175229 522754
rect 175263 522720 175280 522754
rect 175212 522703 175280 522720
rect 175576 522790 175646 522805
rect 175576 522756 175593 522790
rect 175627 522756 175646 522790
rect 174803 522666 174861 522701
rect 174803 522632 174815 522666
rect 174849 522632 174861 522666
rect 174803 522573 174861 522632
rect 172227 522510 172245 522544
rect 172279 522510 172417 522544
rect 172451 522510 172469 522544
rect 172227 522468 172469 522510
rect 172503 522544 173572 522555
rect 172503 522510 172521 522544
rect 172555 522510 173521 522544
rect 173555 522510 173572 522544
rect 172503 522468 173572 522510
rect 173607 522544 174676 522555
rect 173607 522510 173625 522544
rect 173659 522510 174625 522544
rect 174659 522510 174676 522544
rect 173607 522468 174676 522510
rect 174803 522539 174815 522573
rect 174849 522539 174861 522573
rect 175576 522555 175646 522756
rect 176316 522754 176384 522869
rect 176316 522720 176333 522754
rect 176367 522720 176384 522754
rect 176316 522703 176384 522720
rect 176680 522790 176750 522805
rect 176680 522756 176697 522790
rect 176731 522756 176750 522790
rect 176680 522555 176750 522756
rect 177420 522754 177488 522869
rect 177420 522720 177437 522754
rect 177471 522720 177488 522754
rect 177420 522703 177488 522720
rect 177784 522790 177854 522805
rect 177784 522756 177801 522790
rect 177835 522756 177854 522790
rect 177784 522555 177854 522756
rect 178524 522754 178592 522869
rect 179311 522824 179829 522883
rect 179955 522884 180013 522978
rect 179955 522850 179967 522884
rect 180001 522850 180013 522884
rect 180047 522917 181116 522978
rect 180047 522883 180065 522917
rect 180099 522883 181065 522917
rect 181099 522883 181116 522917
rect 180047 522869 181116 522883
rect 181151 522917 182220 522978
rect 181151 522883 181169 522917
rect 181203 522883 182169 522917
rect 182203 522883 182220 522917
rect 181151 522869 182220 522883
rect 182255 522917 183324 522978
rect 182255 522883 182273 522917
rect 182307 522883 183273 522917
rect 183307 522883 183324 522917
rect 182255 522869 183324 522883
rect 183359 522917 184428 522978
rect 183359 522883 183377 522917
rect 183411 522883 184377 522917
rect 184411 522883 184428 522917
rect 183359 522869 184428 522883
rect 184463 522917 184981 522978
rect 184463 522883 184481 522917
rect 184515 522883 184929 522917
rect 184963 522883 184981 522917
rect 179955 522833 180013 522850
rect 178524 522720 178541 522754
rect 178575 522720 178592 522754
rect 178524 522703 178592 522720
rect 178888 522790 178958 522805
rect 178888 522756 178905 522790
rect 178939 522756 178958 522790
rect 178888 522555 178958 522756
rect 179311 522754 179553 522824
rect 179311 522720 179389 522754
rect 179423 522720 179499 522754
rect 179533 522720 179553 522754
rect 179587 522756 179607 522790
rect 179641 522756 179717 522790
rect 179751 522756 179829 522790
rect 179587 522686 179829 522756
rect 180364 522754 180432 522869
rect 180364 522720 180381 522754
rect 180415 522720 180432 522754
rect 180364 522703 180432 522720
rect 180728 522790 180798 522805
rect 180728 522756 180745 522790
rect 180779 522756 180798 522790
rect 179311 522646 179829 522686
rect 179311 522612 179329 522646
rect 179363 522612 179777 522646
rect 179811 522612 179829 522646
rect 174803 522468 174861 522539
rect 174895 522544 175964 522555
rect 174895 522510 174913 522544
rect 174947 522510 175913 522544
rect 175947 522510 175964 522544
rect 174895 522468 175964 522510
rect 175999 522544 177068 522555
rect 175999 522510 176017 522544
rect 176051 522510 177017 522544
rect 177051 522510 177068 522544
rect 175999 522468 177068 522510
rect 177103 522544 178172 522555
rect 177103 522510 177121 522544
rect 177155 522510 178121 522544
rect 178155 522510 178172 522544
rect 177103 522468 178172 522510
rect 178207 522544 179276 522555
rect 178207 522510 178225 522544
rect 178259 522510 179225 522544
rect 179259 522510 179276 522544
rect 178207 522468 179276 522510
rect 179311 522544 179829 522612
rect 179311 522510 179329 522544
rect 179363 522510 179777 522544
rect 179811 522510 179829 522544
rect 179311 522468 179829 522510
rect 179955 522666 180013 522701
rect 179955 522632 179967 522666
rect 180001 522632 180013 522666
rect 179955 522573 180013 522632
rect 179955 522539 179967 522573
rect 180001 522539 180013 522573
rect 180728 522555 180798 522756
rect 181468 522754 181536 522869
rect 181468 522720 181485 522754
rect 181519 522720 181536 522754
rect 181468 522703 181536 522720
rect 181832 522790 181902 522805
rect 181832 522756 181849 522790
rect 181883 522756 181902 522790
rect 181832 522555 181902 522756
rect 182572 522754 182640 522869
rect 182572 522720 182589 522754
rect 182623 522720 182640 522754
rect 182572 522703 182640 522720
rect 182936 522790 183006 522805
rect 182936 522756 182953 522790
rect 182987 522756 183006 522790
rect 182936 522555 183006 522756
rect 183676 522754 183744 522869
rect 184463 522824 184981 522883
rect 185107 522884 185165 522978
rect 185107 522850 185119 522884
rect 185153 522850 185165 522884
rect 185199 522917 186268 522978
rect 185199 522883 185217 522917
rect 185251 522883 186217 522917
rect 186251 522883 186268 522917
rect 185199 522869 186268 522883
rect 186303 522917 187005 522978
rect 186303 522883 186321 522917
rect 186355 522883 186953 522917
rect 186987 522883 187005 522917
rect 185107 522833 185165 522850
rect 183676 522720 183693 522754
rect 183727 522720 183744 522754
rect 183676 522703 183744 522720
rect 184040 522790 184110 522805
rect 184040 522756 184057 522790
rect 184091 522756 184110 522790
rect 184040 522555 184110 522756
rect 184463 522754 184705 522824
rect 184463 522720 184541 522754
rect 184575 522720 184651 522754
rect 184685 522720 184705 522754
rect 184739 522756 184759 522790
rect 184793 522756 184869 522790
rect 184903 522756 184981 522790
rect 184739 522686 184981 522756
rect 185516 522754 185584 522869
rect 186303 522824 187005 522883
rect 187223 522915 187465 522978
rect 187223 522881 187241 522915
rect 187275 522881 187413 522915
rect 187447 522881 187465 522915
rect 187223 522828 187465 522881
rect 185516 522720 185533 522754
rect 185567 522720 185584 522754
rect 185516 522703 185584 522720
rect 185880 522790 185950 522805
rect 185880 522756 185897 522790
rect 185931 522756 185950 522790
rect 184463 522646 184981 522686
rect 184463 522612 184481 522646
rect 184515 522612 184929 522646
rect 184963 522612 184981 522646
rect 179955 522468 180013 522539
rect 180047 522544 181116 522555
rect 180047 522510 180065 522544
rect 180099 522510 181065 522544
rect 181099 522510 181116 522544
rect 180047 522468 181116 522510
rect 181151 522544 182220 522555
rect 181151 522510 181169 522544
rect 181203 522510 182169 522544
rect 182203 522510 182220 522544
rect 181151 522468 182220 522510
rect 182255 522544 183324 522555
rect 182255 522510 182273 522544
rect 182307 522510 183273 522544
rect 183307 522510 183324 522544
rect 182255 522468 183324 522510
rect 183359 522544 184428 522555
rect 183359 522510 183377 522544
rect 183411 522510 184377 522544
rect 184411 522510 184428 522544
rect 183359 522468 184428 522510
rect 184463 522544 184981 522612
rect 184463 522510 184481 522544
rect 184515 522510 184929 522544
rect 184963 522510 184981 522544
rect 184463 522468 184981 522510
rect 185107 522666 185165 522701
rect 185107 522632 185119 522666
rect 185153 522632 185165 522666
rect 185107 522573 185165 522632
rect 185107 522539 185119 522573
rect 185153 522539 185165 522573
rect 185880 522555 185950 522756
rect 186303 522754 186633 522824
rect 186303 522720 186381 522754
rect 186415 522720 186480 522754
rect 186514 522720 186579 522754
rect 186613 522720 186633 522754
rect 186667 522756 186687 522790
rect 186721 522756 186790 522790
rect 186824 522756 186893 522790
rect 186927 522756 187005 522790
rect 186667 522686 187005 522756
rect 186303 522646 187005 522686
rect 186303 522612 186321 522646
rect 186355 522612 186953 522646
rect 186987 522612 187005 522646
rect 185107 522468 185165 522539
rect 185199 522544 186268 522555
rect 185199 522510 185217 522544
rect 185251 522510 186217 522544
rect 186251 522510 186268 522544
rect 185199 522468 186268 522510
rect 186303 522544 187005 522612
rect 186303 522510 186321 522544
rect 186355 522510 186953 522544
rect 186987 522510 187005 522544
rect 186303 522468 187005 522510
rect 187223 522760 187273 522794
rect 187307 522760 187327 522794
rect 187223 522686 187327 522760
rect 187361 522754 187465 522828
rect 187361 522720 187381 522754
rect 187415 522720 187465 522754
rect 187223 522639 187465 522686
rect 187223 522605 187241 522639
rect 187275 522605 187413 522639
rect 187447 522605 187465 522639
rect 187223 522544 187465 522605
rect 187223 522510 187241 522544
rect 187275 522510 187413 522544
rect 187447 522510 187465 522544
rect 187223 522468 187465 522510
rect 172210 522434 172239 522468
rect 172273 522434 172331 522468
rect 172365 522434 172423 522468
rect 172457 522434 172515 522468
rect 172549 522434 172607 522468
rect 172641 522434 172699 522468
rect 172733 522434 172791 522468
rect 172825 522434 172883 522468
rect 172917 522434 172975 522468
rect 173009 522434 173067 522468
rect 173101 522434 173159 522468
rect 173193 522434 173251 522468
rect 173285 522434 173343 522468
rect 173377 522434 173435 522468
rect 173469 522434 173527 522468
rect 173561 522434 173619 522468
rect 173653 522434 173711 522468
rect 173745 522434 173803 522468
rect 173837 522434 173895 522468
rect 173929 522434 173987 522468
rect 174021 522434 174079 522468
rect 174113 522434 174171 522468
rect 174205 522434 174263 522468
rect 174297 522434 174355 522468
rect 174389 522434 174447 522468
rect 174481 522434 174539 522468
rect 174573 522434 174631 522468
rect 174665 522434 174723 522468
rect 174757 522434 174815 522468
rect 174849 522434 174907 522468
rect 174941 522434 174999 522468
rect 175033 522434 175091 522468
rect 175125 522434 175183 522468
rect 175217 522434 175275 522468
rect 175309 522434 175367 522468
rect 175401 522434 175459 522468
rect 175493 522434 175551 522468
rect 175585 522434 175643 522468
rect 175677 522434 175735 522468
rect 175769 522434 175827 522468
rect 175861 522434 175919 522468
rect 175953 522434 176011 522468
rect 176045 522434 176103 522468
rect 176137 522434 176195 522468
rect 176229 522434 176287 522468
rect 176321 522434 176379 522468
rect 176413 522434 176471 522468
rect 176505 522434 176563 522468
rect 176597 522434 176655 522468
rect 176689 522434 176747 522468
rect 176781 522434 176839 522468
rect 176873 522434 176931 522468
rect 176965 522434 177023 522468
rect 177057 522434 177115 522468
rect 177149 522434 177207 522468
rect 177241 522434 177299 522468
rect 177333 522434 177391 522468
rect 177425 522434 177483 522468
rect 177517 522434 177575 522468
rect 177609 522434 177667 522468
rect 177701 522434 177759 522468
rect 177793 522434 177851 522468
rect 177885 522434 177943 522468
rect 177977 522434 178035 522468
rect 178069 522434 178127 522468
rect 178161 522434 178219 522468
rect 178253 522434 178311 522468
rect 178345 522434 178403 522468
rect 178437 522434 178495 522468
rect 178529 522434 178587 522468
rect 178621 522434 178679 522468
rect 178713 522434 178771 522468
rect 178805 522434 178863 522468
rect 178897 522434 178955 522468
rect 178989 522434 179047 522468
rect 179081 522434 179139 522468
rect 179173 522434 179231 522468
rect 179265 522434 179323 522468
rect 179357 522434 179415 522468
rect 179449 522434 179507 522468
rect 179541 522434 179599 522468
rect 179633 522434 179691 522468
rect 179725 522434 179783 522468
rect 179817 522434 179875 522468
rect 179909 522434 179967 522468
rect 180001 522434 180059 522468
rect 180093 522434 180151 522468
rect 180185 522434 180243 522468
rect 180277 522434 180335 522468
rect 180369 522434 180427 522468
rect 180461 522434 180519 522468
rect 180553 522434 180611 522468
rect 180645 522434 180703 522468
rect 180737 522434 180795 522468
rect 180829 522434 180887 522468
rect 180921 522434 180979 522468
rect 181013 522434 181071 522468
rect 181105 522434 181163 522468
rect 181197 522434 181255 522468
rect 181289 522434 181347 522468
rect 181381 522434 181439 522468
rect 181473 522434 181531 522468
rect 181565 522434 181623 522468
rect 181657 522434 181715 522468
rect 181749 522434 181807 522468
rect 181841 522434 181899 522468
rect 181933 522434 181991 522468
rect 182025 522434 182083 522468
rect 182117 522434 182175 522468
rect 182209 522434 182267 522468
rect 182301 522434 182359 522468
rect 182393 522434 182451 522468
rect 182485 522434 182543 522468
rect 182577 522434 182635 522468
rect 182669 522434 182727 522468
rect 182761 522434 182819 522468
rect 182853 522434 182911 522468
rect 182945 522434 183003 522468
rect 183037 522434 183095 522468
rect 183129 522434 183187 522468
rect 183221 522434 183279 522468
rect 183313 522434 183371 522468
rect 183405 522434 183463 522468
rect 183497 522434 183555 522468
rect 183589 522434 183647 522468
rect 183681 522434 183739 522468
rect 183773 522434 183831 522468
rect 183865 522434 183923 522468
rect 183957 522434 184015 522468
rect 184049 522434 184107 522468
rect 184141 522434 184199 522468
rect 184233 522434 184291 522468
rect 184325 522434 184383 522468
rect 184417 522434 184475 522468
rect 184509 522434 184567 522468
rect 184601 522434 184659 522468
rect 184693 522434 184751 522468
rect 184785 522434 184843 522468
rect 184877 522434 184935 522468
rect 184969 522434 185027 522468
rect 185061 522434 185119 522468
rect 185153 522434 185211 522468
rect 185245 522434 185303 522468
rect 185337 522434 185395 522468
rect 185429 522434 185487 522468
rect 185521 522434 185579 522468
rect 185613 522434 185671 522468
rect 185705 522434 185763 522468
rect 185797 522434 185855 522468
rect 185889 522434 185947 522468
rect 185981 522434 186039 522468
rect 186073 522434 186131 522468
rect 186165 522434 186223 522468
rect 186257 522434 186315 522468
rect 186349 522434 186407 522468
rect 186441 522434 186499 522468
rect 186533 522434 186591 522468
rect 186625 522434 186683 522468
rect 186717 522434 186775 522468
rect 186809 522434 186867 522468
rect 186901 522434 186959 522468
rect 186993 522434 187051 522468
rect 187085 522434 187143 522468
rect 187177 522434 187235 522468
rect 187269 522434 187327 522468
rect 187361 522434 187419 522468
rect 187453 522434 187482 522468
rect 172227 522392 172469 522434
rect 172227 522358 172245 522392
rect 172279 522358 172417 522392
rect 172451 522358 172469 522392
rect 172227 522297 172469 522358
rect 172503 522392 173572 522434
rect 172503 522358 172521 522392
rect 172555 522358 173521 522392
rect 173555 522358 173572 522392
rect 172503 522347 173572 522358
rect 173607 522392 174676 522434
rect 173607 522358 173625 522392
rect 173659 522358 174625 522392
rect 174659 522358 174676 522392
rect 173607 522347 174676 522358
rect 174711 522392 175780 522434
rect 174711 522358 174729 522392
rect 174763 522358 175729 522392
rect 175763 522358 175780 522392
rect 174711 522347 175780 522358
rect 175815 522392 176884 522434
rect 175815 522358 175833 522392
rect 175867 522358 176833 522392
rect 176867 522358 176884 522392
rect 175815 522347 176884 522358
rect 176919 522392 177253 522434
rect 176919 522358 176937 522392
rect 176971 522358 177201 522392
rect 177235 522358 177253 522392
rect 172227 522263 172245 522297
rect 172279 522263 172417 522297
rect 172451 522263 172469 522297
rect 172227 522216 172469 522263
rect 172227 522148 172277 522182
rect 172311 522148 172331 522182
rect 172227 522074 172331 522148
rect 172365 522142 172469 522216
rect 172365 522108 172385 522142
rect 172419 522108 172469 522142
rect 172820 522182 172888 522199
rect 172820 522148 172837 522182
rect 172871 522148 172888 522182
rect 172227 522021 172469 522074
rect 172820 522033 172888 522148
rect 173184 522146 173254 522347
rect 173184 522112 173201 522146
rect 173235 522112 173254 522146
rect 173184 522097 173254 522112
rect 173924 522182 173992 522199
rect 173924 522148 173941 522182
rect 173975 522148 173992 522182
rect 173924 522033 173992 522148
rect 174288 522146 174358 522347
rect 174288 522112 174305 522146
rect 174339 522112 174358 522146
rect 174288 522097 174358 522112
rect 175028 522182 175096 522199
rect 175028 522148 175045 522182
rect 175079 522148 175096 522182
rect 175028 522033 175096 522148
rect 175392 522146 175462 522347
rect 175392 522112 175409 522146
rect 175443 522112 175462 522146
rect 175392 522097 175462 522112
rect 176132 522182 176200 522199
rect 176132 522148 176149 522182
rect 176183 522148 176200 522182
rect 176132 522033 176200 522148
rect 176496 522146 176566 522347
rect 176919 522290 177253 522358
rect 176919 522256 176937 522290
rect 176971 522256 177201 522290
rect 177235 522256 177253 522290
rect 176919 522216 177253 522256
rect 176496 522112 176513 522146
rect 176547 522112 176566 522146
rect 176496 522097 176566 522112
rect 176919 522148 176939 522182
rect 176973 522148 177069 522182
rect 176919 522078 177069 522148
rect 177103 522146 177253 522216
rect 177379 522363 177437 522434
rect 177379 522329 177391 522363
rect 177425 522329 177437 522363
rect 177471 522392 178540 522434
rect 177471 522358 177489 522392
rect 177523 522358 178489 522392
rect 178523 522358 178540 522392
rect 177471 522347 178540 522358
rect 178575 522392 179644 522434
rect 178575 522358 178593 522392
rect 178627 522358 179593 522392
rect 179627 522358 179644 522392
rect 178575 522347 179644 522358
rect 179679 522392 180748 522434
rect 179679 522358 179697 522392
rect 179731 522358 180697 522392
rect 180731 522358 180748 522392
rect 179679 522347 180748 522358
rect 180783 522392 181852 522434
rect 180783 522358 180801 522392
rect 180835 522358 181801 522392
rect 181835 522358 181852 522392
rect 180783 522347 181852 522358
rect 181887 522392 182405 522434
rect 181887 522358 181905 522392
rect 181939 522358 182353 522392
rect 182387 522358 182405 522392
rect 177379 522270 177437 522329
rect 177379 522236 177391 522270
rect 177425 522236 177437 522270
rect 177379 522201 177437 522236
rect 177103 522112 177199 522146
rect 177233 522112 177253 522146
rect 177788 522182 177856 522199
rect 177788 522148 177805 522182
rect 177839 522148 177856 522182
rect 172227 521987 172245 522021
rect 172279 521987 172417 522021
rect 172451 521987 172469 522021
rect 172227 521924 172469 521987
rect 172503 522019 173572 522033
rect 172503 521985 172521 522019
rect 172555 521985 173521 522019
rect 173555 521985 173572 522019
rect 172503 521924 173572 521985
rect 173607 522019 174676 522033
rect 173607 521985 173625 522019
rect 173659 521985 174625 522019
rect 174659 521985 174676 522019
rect 173607 521924 174676 521985
rect 174711 522019 175780 522033
rect 174711 521985 174729 522019
rect 174763 521985 175729 522019
rect 175763 521985 175780 522019
rect 174711 521924 175780 521985
rect 175815 522019 176884 522033
rect 175815 521985 175833 522019
rect 175867 521985 176833 522019
rect 176867 521985 176884 522019
rect 175815 521924 176884 521985
rect 176919 522026 177253 522078
rect 176919 521992 176937 522026
rect 176971 521992 177201 522026
rect 177235 521992 177253 522026
rect 176919 521924 177253 521992
rect 177379 522052 177437 522069
rect 177379 522018 177391 522052
rect 177425 522018 177437 522052
rect 177788 522033 177856 522148
rect 178152 522146 178222 522347
rect 178152 522112 178169 522146
rect 178203 522112 178222 522146
rect 178152 522097 178222 522112
rect 178892 522182 178960 522199
rect 178892 522148 178909 522182
rect 178943 522148 178960 522182
rect 178892 522033 178960 522148
rect 179256 522146 179326 522347
rect 179256 522112 179273 522146
rect 179307 522112 179326 522146
rect 179256 522097 179326 522112
rect 179996 522182 180064 522199
rect 179996 522148 180013 522182
rect 180047 522148 180064 522182
rect 179996 522033 180064 522148
rect 180360 522146 180430 522347
rect 180360 522112 180377 522146
rect 180411 522112 180430 522146
rect 180360 522097 180430 522112
rect 181100 522182 181168 522199
rect 181100 522148 181117 522182
rect 181151 522148 181168 522182
rect 181100 522033 181168 522148
rect 181464 522146 181534 522347
rect 181887 522290 182405 522358
rect 181887 522256 181905 522290
rect 181939 522256 182353 522290
rect 182387 522256 182405 522290
rect 181887 522216 182405 522256
rect 181464 522112 181481 522146
rect 181515 522112 181534 522146
rect 181464 522097 181534 522112
rect 181887 522148 181965 522182
rect 181999 522148 182075 522182
rect 182109 522148 182129 522182
rect 181887 522078 182129 522148
rect 182163 522146 182405 522216
rect 182531 522363 182589 522434
rect 182531 522329 182543 522363
rect 182577 522329 182589 522363
rect 182623 522392 183692 522434
rect 182623 522358 182641 522392
rect 182675 522358 183641 522392
rect 183675 522358 183692 522392
rect 182623 522347 183692 522358
rect 183727 522392 184796 522434
rect 183727 522358 183745 522392
rect 183779 522358 184745 522392
rect 184779 522358 184796 522392
rect 183727 522347 184796 522358
rect 184831 522392 185900 522434
rect 184831 522358 184849 522392
rect 184883 522358 185849 522392
rect 185883 522358 185900 522392
rect 184831 522347 185900 522358
rect 185935 522392 187004 522434
rect 185935 522358 185953 522392
rect 185987 522358 186953 522392
rect 186987 522358 187004 522392
rect 185935 522347 187004 522358
rect 187223 522392 187465 522434
rect 187223 522358 187241 522392
rect 187275 522358 187413 522392
rect 187447 522358 187465 522392
rect 182531 522270 182589 522329
rect 182531 522236 182543 522270
rect 182577 522236 182589 522270
rect 182531 522201 182589 522236
rect 182163 522112 182183 522146
rect 182217 522112 182293 522146
rect 182327 522112 182405 522146
rect 182940 522182 183008 522199
rect 182940 522148 182957 522182
rect 182991 522148 183008 522182
rect 177379 521924 177437 522018
rect 177471 522019 178540 522033
rect 177471 521985 177489 522019
rect 177523 521985 178489 522019
rect 178523 521985 178540 522019
rect 177471 521924 178540 521985
rect 178575 522019 179644 522033
rect 178575 521985 178593 522019
rect 178627 521985 179593 522019
rect 179627 521985 179644 522019
rect 178575 521924 179644 521985
rect 179679 522019 180748 522033
rect 179679 521985 179697 522019
rect 179731 521985 180697 522019
rect 180731 521985 180748 522019
rect 179679 521924 180748 521985
rect 180783 522019 181852 522033
rect 180783 521985 180801 522019
rect 180835 521985 181801 522019
rect 181835 521985 181852 522019
rect 180783 521924 181852 521985
rect 181887 522019 182405 522078
rect 181887 521985 181905 522019
rect 181939 521985 182353 522019
rect 182387 521985 182405 522019
rect 181887 521924 182405 521985
rect 182531 522052 182589 522069
rect 182531 522018 182543 522052
rect 182577 522018 182589 522052
rect 182940 522033 183008 522148
rect 183304 522146 183374 522347
rect 183304 522112 183321 522146
rect 183355 522112 183374 522146
rect 183304 522097 183374 522112
rect 184044 522182 184112 522199
rect 184044 522148 184061 522182
rect 184095 522148 184112 522182
rect 184044 522033 184112 522148
rect 184408 522146 184478 522347
rect 184408 522112 184425 522146
rect 184459 522112 184478 522146
rect 184408 522097 184478 522112
rect 185148 522182 185216 522199
rect 185148 522148 185165 522182
rect 185199 522148 185216 522182
rect 185148 522033 185216 522148
rect 185512 522146 185582 522347
rect 185512 522112 185529 522146
rect 185563 522112 185582 522146
rect 185512 522097 185582 522112
rect 186252 522182 186320 522199
rect 186252 522148 186269 522182
rect 186303 522148 186320 522182
rect 186252 522033 186320 522148
rect 186616 522146 186686 522347
rect 186616 522112 186633 522146
rect 186667 522112 186686 522146
rect 186616 522097 186686 522112
rect 187223 522297 187465 522358
rect 187223 522263 187241 522297
rect 187275 522263 187413 522297
rect 187447 522263 187465 522297
rect 187223 522216 187465 522263
rect 187223 522142 187327 522216
rect 187223 522108 187273 522142
rect 187307 522108 187327 522142
rect 187361 522148 187381 522182
rect 187415 522148 187465 522182
rect 187361 522074 187465 522148
rect 182531 521924 182589 522018
rect 182623 522019 183692 522033
rect 182623 521985 182641 522019
rect 182675 521985 183641 522019
rect 183675 521985 183692 522019
rect 182623 521924 183692 521985
rect 183727 522019 184796 522033
rect 183727 521985 183745 522019
rect 183779 521985 184745 522019
rect 184779 521985 184796 522019
rect 183727 521924 184796 521985
rect 184831 522019 185900 522033
rect 184831 521985 184849 522019
rect 184883 521985 185849 522019
rect 185883 521985 185900 522019
rect 184831 521924 185900 521985
rect 185935 522019 187004 522033
rect 185935 521985 185953 522019
rect 185987 521985 186953 522019
rect 186987 521985 187004 522019
rect 185935 521924 187004 521985
rect 187223 522021 187465 522074
rect 187223 521987 187241 522021
rect 187275 521987 187413 522021
rect 187447 521987 187465 522021
rect 187223 521924 187465 521987
rect 172210 521890 172239 521924
rect 172273 521890 172331 521924
rect 172365 521890 172423 521924
rect 172457 521890 172515 521924
rect 172549 521890 172607 521924
rect 172641 521890 172699 521924
rect 172733 521890 172791 521924
rect 172825 521890 172883 521924
rect 172917 521890 172975 521924
rect 173009 521890 173067 521924
rect 173101 521890 173159 521924
rect 173193 521890 173251 521924
rect 173285 521890 173343 521924
rect 173377 521890 173435 521924
rect 173469 521890 173527 521924
rect 173561 521890 173619 521924
rect 173653 521890 173711 521924
rect 173745 521890 173803 521924
rect 173837 521890 173895 521924
rect 173929 521890 173987 521924
rect 174021 521890 174079 521924
rect 174113 521890 174171 521924
rect 174205 521890 174263 521924
rect 174297 521890 174355 521924
rect 174389 521890 174447 521924
rect 174481 521890 174539 521924
rect 174573 521890 174631 521924
rect 174665 521890 174723 521924
rect 174757 521890 174815 521924
rect 174849 521890 174907 521924
rect 174941 521890 174999 521924
rect 175033 521890 175091 521924
rect 175125 521890 175183 521924
rect 175217 521890 175275 521924
rect 175309 521890 175367 521924
rect 175401 521890 175459 521924
rect 175493 521890 175551 521924
rect 175585 521890 175643 521924
rect 175677 521890 175735 521924
rect 175769 521890 175827 521924
rect 175861 521890 175919 521924
rect 175953 521890 176011 521924
rect 176045 521890 176103 521924
rect 176137 521890 176195 521924
rect 176229 521890 176287 521924
rect 176321 521890 176379 521924
rect 176413 521890 176471 521924
rect 176505 521890 176563 521924
rect 176597 521890 176655 521924
rect 176689 521890 176747 521924
rect 176781 521890 176839 521924
rect 176873 521890 176931 521924
rect 176965 521890 177023 521924
rect 177057 521890 177115 521924
rect 177149 521890 177207 521924
rect 177241 521890 177299 521924
rect 177333 521890 177391 521924
rect 177425 521890 177483 521924
rect 177517 521890 177575 521924
rect 177609 521890 177667 521924
rect 177701 521890 177759 521924
rect 177793 521890 177851 521924
rect 177885 521890 177943 521924
rect 177977 521890 178035 521924
rect 178069 521890 178127 521924
rect 178161 521890 178219 521924
rect 178253 521890 178311 521924
rect 178345 521890 178403 521924
rect 178437 521890 178495 521924
rect 178529 521890 178587 521924
rect 178621 521890 178679 521924
rect 178713 521890 178771 521924
rect 178805 521890 178863 521924
rect 178897 521890 178955 521924
rect 178989 521890 179047 521924
rect 179081 521890 179139 521924
rect 179173 521890 179231 521924
rect 179265 521890 179323 521924
rect 179357 521890 179415 521924
rect 179449 521890 179507 521924
rect 179541 521890 179599 521924
rect 179633 521890 179691 521924
rect 179725 521890 179783 521924
rect 179817 521890 179875 521924
rect 179909 521890 179967 521924
rect 180001 521890 180059 521924
rect 180093 521890 180151 521924
rect 180185 521890 180243 521924
rect 180277 521890 180335 521924
rect 180369 521890 180427 521924
rect 180461 521890 180519 521924
rect 180553 521890 180611 521924
rect 180645 521890 180703 521924
rect 180737 521890 180795 521924
rect 180829 521890 180887 521924
rect 180921 521890 180979 521924
rect 181013 521890 181071 521924
rect 181105 521890 181163 521924
rect 181197 521890 181255 521924
rect 181289 521890 181347 521924
rect 181381 521890 181439 521924
rect 181473 521890 181531 521924
rect 181565 521890 181623 521924
rect 181657 521890 181715 521924
rect 181749 521890 181807 521924
rect 181841 521890 181899 521924
rect 181933 521890 181991 521924
rect 182025 521890 182083 521924
rect 182117 521890 182175 521924
rect 182209 521890 182267 521924
rect 182301 521890 182359 521924
rect 182393 521890 182451 521924
rect 182485 521890 182543 521924
rect 182577 521890 182635 521924
rect 182669 521890 182727 521924
rect 182761 521890 182819 521924
rect 182853 521890 182911 521924
rect 182945 521890 183003 521924
rect 183037 521890 183095 521924
rect 183129 521890 183187 521924
rect 183221 521890 183279 521924
rect 183313 521890 183371 521924
rect 183405 521890 183463 521924
rect 183497 521890 183555 521924
rect 183589 521890 183647 521924
rect 183681 521890 183739 521924
rect 183773 521890 183831 521924
rect 183865 521890 183923 521924
rect 183957 521890 184015 521924
rect 184049 521890 184107 521924
rect 184141 521890 184199 521924
rect 184233 521890 184291 521924
rect 184325 521890 184383 521924
rect 184417 521890 184475 521924
rect 184509 521890 184567 521924
rect 184601 521890 184659 521924
rect 184693 521890 184751 521924
rect 184785 521890 184843 521924
rect 184877 521890 184935 521924
rect 184969 521890 185027 521924
rect 185061 521890 185119 521924
rect 185153 521890 185211 521924
rect 185245 521890 185303 521924
rect 185337 521890 185395 521924
rect 185429 521890 185487 521924
rect 185521 521890 185579 521924
rect 185613 521890 185671 521924
rect 185705 521890 185763 521924
rect 185797 521890 185855 521924
rect 185889 521890 185947 521924
rect 185981 521890 186039 521924
rect 186073 521890 186131 521924
rect 186165 521890 186223 521924
rect 186257 521890 186315 521924
rect 186349 521890 186407 521924
rect 186441 521890 186499 521924
rect 186533 521890 186591 521924
rect 186625 521890 186683 521924
rect 186717 521890 186775 521924
rect 186809 521890 186867 521924
rect 186901 521890 186959 521924
rect 186993 521890 187051 521924
rect 187085 521890 187143 521924
rect 187177 521890 187235 521924
rect 187269 521890 187327 521924
rect 187361 521890 187419 521924
rect 187453 521890 187482 521924
rect 172227 521827 172469 521890
rect 172227 521793 172245 521827
rect 172279 521793 172417 521827
rect 172451 521793 172469 521827
rect 172227 521740 172469 521793
rect 172503 521829 173572 521890
rect 172503 521795 172521 521829
rect 172555 521795 173521 521829
rect 173555 521795 173572 521829
rect 172503 521781 173572 521795
rect 173607 521829 174676 521890
rect 173607 521795 173625 521829
rect 173659 521795 174625 521829
rect 174659 521795 174676 521829
rect 173607 521781 174676 521795
rect 174803 521796 174861 521890
rect 172227 521666 172331 521740
rect 172227 521632 172277 521666
rect 172311 521632 172331 521666
rect 172365 521672 172385 521706
rect 172419 521672 172469 521706
rect 172365 521598 172469 521672
rect 172820 521666 172888 521781
rect 172820 521632 172837 521666
rect 172871 521632 172888 521666
rect 172820 521615 172888 521632
rect 173184 521702 173254 521717
rect 173184 521668 173201 521702
rect 173235 521668 173254 521702
rect 172227 521551 172469 521598
rect 172227 521517 172245 521551
rect 172279 521517 172417 521551
rect 172451 521517 172469 521551
rect 172227 521456 172469 521517
rect 173184 521467 173254 521668
rect 173924 521666 173992 521781
rect 174803 521762 174815 521796
rect 174849 521762 174861 521796
rect 174895 521829 175964 521890
rect 174895 521795 174913 521829
rect 174947 521795 175913 521829
rect 175947 521795 175964 521829
rect 174895 521781 175964 521795
rect 175999 521829 177068 521890
rect 175999 521795 176017 521829
rect 176051 521795 177017 521829
rect 177051 521795 177068 521829
rect 175999 521781 177068 521795
rect 177103 521829 178172 521890
rect 177103 521795 177121 521829
rect 177155 521795 178121 521829
rect 178155 521795 178172 521829
rect 177103 521781 178172 521795
rect 178207 521829 179276 521890
rect 178207 521795 178225 521829
rect 178259 521795 179225 521829
rect 179259 521795 179276 521829
rect 178207 521781 179276 521795
rect 179311 521829 179829 521890
rect 179311 521795 179329 521829
rect 179363 521795 179777 521829
rect 179811 521795 179829 521829
rect 174803 521745 174861 521762
rect 173924 521632 173941 521666
rect 173975 521632 173992 521666
rect 173924 521615 173992 521632
rect 174288 521702 174358 521717
rect 174288 521668 174305 521702
rect 174339 521668 174358 521702
rect 174288 521467 174358 521668
rect 175212 521666 175280 521781
rect 175212 521632 175229 521666
rect 175263 521632 175280 521666
rect 175212 521615 175280 521632
rect 175576 521702 175646 521717
rect 175576 521668 175593 521702
rect 175627 521668 175646 521702
rect 174803 521578 174861 521613
rect 174803 521544 174815 521578
rect 174849 521544 174861 521578
rect 174803 521485 174861 521544
rect 172227 521422 172245 521456
rect 172279 521422 172417 521456
rect 172451 521422 172469 521456
rect 172227 521380 172469 521422
rect 172503 521456 173572 521467
rect 172503 521422 172521 521456
rect 172555 521422 173521 521456
rect 173555 521422 173572 521456
rect 172503 521380 173572 521422
rect 173607 521456 174676 521467
rect 173607 521422 173625 521456
rect 173659 521422 174625 521456
rect 174659 521422 174676 521456
rect 173607 521380 174676 521422
rect 174803 521451 174815 521485
rect 174849 521451 174861 521485
rect 175576 521467 175646 521668
rect 176316 521666 176384 521781
rect 176316 521632 176333 521666
rect 176367 521632 176384 521666
rect 176316 521615 176384 521632
rect 176680 521702 176750 521717
rect 176680 521668 176697 521702
rect 176731 521668 176750 521702
rect 176680 521467 176750 521668
rect 177420 521666 177488 521781
rect 177420 521632 177437 521666
rect 177471 521632 177488 521666
rect 177420 521615 177488 521632
rect 177784 521702 177854 521717
rect 177784 521668 177801 521702
rect 177835 521668 177854 521702
rect 177784 521467 177854 521668
rect 178524 521666 178592 521781
rect 179311 521736 179829 521795
rect 179955 521796 180013 521890
rect 179955 521762 179967 521796
rect 180001 521762 180013 521796
rect 180047 521829 181116 521890
rect 180047 521795 180065 521829
rect 180099 521795 181065 521829
rect 181099 521795 181116 521829
rect 180047 521781 181116 521795
rect 181151 521829 182220 521890
rect 181151 521795 181169 521829
rect 181203 521795 182169 521829
rect 182203 521795 182220 521829
rect 181151 521781 182220 521795
rect 182255 521829 183324 521890
rect 182255 521795 182273 521829
rect 182307 521795 183273 521829
rect 183307 521795 183324 521829
rect 182255 521781 183324 521795
rect 183359 521829 184428 521890
rect 183359 521795 183377 521829
rect 183411 521795 184377 521829
rect 184411 521795 184428 521829
rect 183359 521781 184428 521795
rect 184463 521829 184981 521890
rect 184463 521795 184481 521829
rect 184515 521795 184929 521829
rect 184963 521795 184981 521829
rect 179955 521745 180013 521762
rect 178524 521632 178541 521666
rect 178575 521632 178592 521666
rect 178524 521615 178592 521632
rect 178888 521702 178958 521717
rect 178888 521668 178905 521702
rect 178939 521668 178958 521702
rect 178888 521467 178958 521668
rect 179311 521666 179553 521736
rect 179311 521632 179389 521666
rect 179423 521632 179499 521666
rect 179533 521632 179553 521666
rect 179587 521668 179607 521702
rect 179641 521668 179717 521702
rect 179751 521668 179829 521702
rect 179587 521598 179829 521668
rect 180364 521666 180432 521781
rect 180364 521632 180381 521666
rect 180415 521632 180432 521666
rect 180364 521615 180432 521632
rect 180728 521702 180798 521717
rect 180728 521668 180745 521702
rect 180779 521668 180798 521702
rect 179311 521558 179829 521598
rect 179311 521524 179329 521558
rect 179363 521524 179777 521558
rect 179811 521524 179829 521558
rect 174803 521380 174861 521451
rect 174895 521456 175964 521467
rect 174895 521422 174913 521456
rect 174947 521422 175913 521456
rect 175947 521422 175964 521456
rect 174895 521380 175964 521422
rect 175999 521456 177068 521467
rect 175999 521422 176017 521456
rect 176051 521422 177017 521456
rect 177051 521422 177068 521456
rect 175999 521380 177068 521422
rect 177103 521456 178172 521467
rect 177103 521422 177121 521456
rect 177155 521422 178121 521456
rect 178155 521422 178172 521456
rect 177103 521380 178172 521422
rect 178207 521456 179276 521467
rect 178207 521422 178225 521456
rect 178259 521422 179225 521456
rect 179259 521422 179276 521456
rect 178207 521380 179276 521422
rect 179311 521456 179829 521524
rect 179311 521422 179329 521456
rect 179363 521422 179777 521456
rect 179811 521422 179829 521456
rect 179311 521380 179829 521422
rect 179955 521578 180013 521613
rect 179955 521544 179967 521578
rect 180001 521544 180013 521578
rect 179955 521485 180013 521544
rect 179955 521451 179967 521485
rect 180001 521451 180013 521485
rect 180728 521467 180798 521668
rect 181468 521666 181536 521781
rect 181468 521632 181485 521666
rect 181519 521632 181536 521666
rect 181468 521615 181536 521632
rect 181832 521702 181902 521717
rect 181832 521668 181849 521702
rect 181883 521668 181902 521702
rect 181832 521467 181902 521668
rect 182572 521666 182640 521781
rect 182572 521632 182589 521666
rect 182623 521632 182640 521666
rect 182572 521615 182640 521632
rect 182936 521702 183006 521717
rect 182936 521668 182953 521702
rect 182987 521668 183006 521702
rect 182936 521467 183006 521668
rect 183676 521666 183744 521781
rect 184463 521736 184981 521795
rect 185107 521796 185165 521890
rect 185107 521762 185119 521796
rect 185153 521762 185165 521796
rect 185199 521829 186268 521890
rect 185199 521795 185217 521829
rect 185251 521795 186217 521829
rect 186251 521795 186268 521829
rect 185199 521781 186268 521795
rect 186303 521829 187005 521890
rect 186303 521795 186321 521829
rect 186355 521795 186953 521829
rect 186987 521795 187005 521829
rect 185107 521745 185165 521762
rect 183676 521632 183693 521666
rect 183727 521632 183744 521666
rect 183676 521615 183744 521632
rect 184040 521702 184110 521717
rect 184040 521668 184057 521702
rect 184091 521668 184110 521702
rect 184040 521467 184110 521668
rect 184463 521666 184705 521736
rect 184463 521632 184541 521666
rect 184575 521632 184651 521666
rect 184685 521632 184705 521666
rect 184739 521668 184759 521702
rect 184793 521668 184869 521702
rect 184903 521668 184981 521702
rect 184739 521598 184981 521668
rect 185516 521666 185584 521781
rect 186303 521736 187005 521795
rect 187223 521827 187465 521890
rect 187223 521793 187241 521827
rect 187275 521793 187413 521827
rect 187447 521793 187465 521827
rect 187223 521740 187465 521793
rect 185516 521632 185533 521666
rect 185567 521632 185584 521666
rect 185516 521615 185584 521632
rect 185880 521702 185950 521717
rect 185880 521668 185897 521702
rect 185931 521668 185950 521702
rect 184463 521558 184981 521598
rect 184463 521524 184481 521558
rect 184515 521524 184929 521558
rect 184963 521524 184981 521558
rect 179955 521380 180013 521451
rect 180047 521456 181116 521467
rect 180047 521422 180065 521456
rect 180099 521422 181065 521456
rect 181099 521422 181116 521456
rect 180047 521380 181116 521422
rect 181151 521456 182220 521467
rect 181151 521422 181169 521456
rect 181203 521422 182169 521456
rect 182203 521422 182220 521456
rect 181151 521380 182220 521422
rect 182255 521456 183324 521467
rect 182255 521422 182273 521456
rect 182307 521422 183273 521456
rect 183307 521422 183324 521456
rect 182255 521380 183324 521422
rect 183359 521456 184428 521467
rect 183359 521422 183377 521456
rect 183411 521422 184377 521456
rect 184411 521422 184428 521456
rect 183359 521380 184428 521422
rect 184463 521456 184981 521524
rect 184463 521422 184481 521456
rect 184515 521422 184929 521456
rect 184963 521422 184981 521456
rect 184463 521380 184981 521422
rect 185107 521578 185165 521613
rect 185107 521544 185119 521578
rect 185153 521544 185165 521578
rect 185107 521485 185165 521544
rect 185107 521451 185119 521485
rect 185153 521451 185165 521485
rect 185880 521467 185950 521668
rect 186303 521666 186633 521736
rect 186303 521632 186381 521666
rect 186415 521632 186480 521666
rect 186514 521632 186579 521666
rect 186613 521632 186633 521666
rect 186667 521668 186687 521702
rect 186721 521668 186790 521702
rect 186824 521668 186893 521702
rect 186927 521668 187005 521702
rect 186667 521598 187005 521668
rect 186303 521558 187005 521598
rect 186303 521524 186321 521558
rect 186355 521524 186953 521558
rect 186987 521524 187005 521558
rect 185107 521380 185165 521451
rect 185199 521456 186268 521467
rect 185199 521422 185217 521456
rect 185251 521422 186217 521456
rect 186251 521422 186268 521456
rect 185199 521380 186268 521422
rect 186303 521456 187005 521524
rect 186303 521422 186321 521456
rect 186355 521422 186953 521456
rect 186987 521422 187005 521456
rect 186303 521380 187005 521422
rect 187223 521672 187273 521706
rect 187307 521672 187327 521706
rect 187223 521598 187327 521672
rect 187361 521666 187465 521740
rect 187361 521632 187381 521666
rect 187415 521632 187465 521666
rect 187223 521551 187465 521598
rect 187223 521517 187241 521551
rect 187275 521517 187413 521551
rect 187447 521517 187465 521551
rect 187223 521456 187465 521517
rect 187223 521422 187241 521456
rect 187275 521422 187413 521456
rect 187447 521422 187465 521456
rect 187223 521380 187465 521422
rect 172210 521346 172239 521380
rect 172273 521346 172331 521380
rect 172365 521346 172423 521380
rect 172457 521346 172515 521380
rect 172549 521346 172607 521380
rect 172641 521346 172699 521380
rect 172733 521346 172791 521380
rect 172825 521346 172883 521380
rect 172917 521346 172975 521380
rect 173009 521346 173067 521380
rect 173101 521346 173159 521380
rect 173193 521346 173251 521380
rect 173285 521346 173343 521380
rect 173377 521346 173435 521380
rect 173469 521346 173527 521380
rect 173561 521346 173619 521380
rect 173653 521346 173711 521380
rect 173745 521346 173803 521380
rect 173837 521346 173895 521380
rect 173929 521346 173987 521380
rect 174021 521346 174079 521380
rect 174113 521346 174171 521380
rect 174205 521346 174263 521380
rect 174297 521346 174355 521380
rect 174389 521346 174447 521380
rect 174481 521346 174539 521380
rect 174573 521346 174631 521380
rect 174665 521346 174723 521380
rect 174757 521346 174815 521380
rect 174849 521346 174907 521380
rect 174941 521346 174999 521380
rect 175033 521346 175091 521380
rect 175125 521346 175183 521380
rect 175217 521346 175275 521380
rect 175309 521346 175367 521380
rect 175401 521346 175459 521380
rect 175493 521346 175551 521380
rect 175585 521346 175643 521380
rect 175677 521346 175735 521380
rect 175769 521346 175827 521380
rect 175861 521346 175919 521380
rect 175953 521346 176011 521380
rect 176045 521346 176103 521380
rect 176137 521346 176195 521380
rect 176229 521346 176287 521380
rect 176321 521346 176379 521380
rect 176413 521346 176471 521380
rect 176505 521346 176563 521380
rect 176597 521346 176655 521380
rect 176689 521346 176747 521380
rect 176781 521346 176839 521380
rect 176873 521346 176931 521380
rect 176965 521346 177023 521380
rect 177057 521346 177115 521380
rect 177149 521346 177207 521380
rect 177241 521346 177299 521380
rect 177333 521346 177391 521380
rect 177425 521346 177483 521380
rect 177517 521346 177575 521380
rect 177609 521346 177667 521380
rect 177701 521346 177759 521380
rect 177793 521346 177851 521380
rect 177885 521346 177943 521380
rect 177977 521346 178035 521380
rect 178069 521346 178127 521380
rect 178161 521346 178219 521380
rect 178253 521346 178311 521380
rect 178345 521346 178403 521380
rect 178437 521346 178495 521380
rect 178529 521346 178587 521380
rect 178621 521346 178679 521380
rect 178713 521346 178771 521380
rect 178805 521346 178863 521380
rect 178897 521346 178955 521380
rect 178989 521346 179047 521380
rect 179081 521346 179139 521380
rect 179173 521346 179231 521380
rect 179265 521346 179323 521380
rect 179357 521346 179415 521380
rect 179449 521346 179507 521380
rect 179541 521346 179599 521380
rect 179633 521346 179691 521380
rect 179725 521346 179783 521380
rect 179817 521346 179875 521380
rect 179909 521346 179967 521380
rect 180001 521346 180059 521380
rect 180093 521346 180151 521380
rect 180185 521346 180243 521380
rect 180277 521346 180335 521380
rect 180369 521346 180427 521380
rect 180461 521346 180519 521380
rect 180553 521346 180611 521380
rect 180645 521346 180703 521380
rect 180737 521346 180795 521380
rect 180829 521346 180887 521380
rect 180921 521346 180979 521380
rect 181013 521346 181071 521380
rect 181105 521346 181163 521380
rect 181197 521346 181255 521380
rect 181289 521346 181347 521380
rect 181381 521346 181439 521380
rect 181473 521346 181531 521380
rect 181565 521346 181623 521380
rect 181657 521346 181715 521380
rect 181749 521346 181807 521380
rect 181841 521346 181899 521380
rect 181933 521346 181991 521380
rect 182025 521346 182083 521380
rect 182117 521346 182175 521380
rect 182209 521346 182267 521380
rect 182301 521346 182359 521380
rect 182393 521346 182451 521380
rect 182485 521346 182543 521380
rect 182577 521346 182635 521380
rect 182669 521346 182727 521380
rect 182761 521346 182819 521380
rect 182853 521346 182911 521380
rect 182945 521346 183003 521380
rect 183037 521346 183095 521380
rect 183129 521346 183187 521380
rect 183221 521346 183279 521380
rect 183313 521346 183371 521380
rect 183405 521346 183463 521380
rect 183497 521346 183555 521380
rect 183589 521346 183647 521380
rect 183681 521346 183739 521380
rect 183773 521346 183831 521380
rect 183865 521346 183923 521380
rect 183957 521346 184015 521380
rect 184049 521346 184107 521380
rect 184141 521346 184199 521380
rect 184233 521346 184291 521380
rect 184325 521346 184383 521380
rect 184417 521346 184475 521380
rect 184509 521346 184567 521380
rect 184601 521346 184659 521380
rect 184693 521346 184751 521380
rect 184785 521346 184843 521380
rect 184877 521346 184935 521380
rect 184969 521346 185027 521380
rect 185061 521346 185119 521380
rect 185153 521346 185211 521380
rect 185245 521346 185303 521380
rect 185337 521346 185395 521380
rect 185429 521346 185487 521380
rect 185521 521346 185579 521380
rect 185613 521346 185671 521380
rect 185705 521346 185763 521380
rect 185797 521346 185855 521380
rect 185889 521346 185947 521380
rect 185981 521346 186039 521380
rect 186073 521346 186131 521380
rect 186165 521346 186223 521380
rect 186257 521346 186315 521380
rect 186349 521346 186407 521380
rect 186441 521346 186499 521380
rect 186533 521346 186591 521380
rect 186625 521346 186683 521380
rect 186717 521346 186775 521380
rect 186809 521346 186867 521380
rect 186901 521346 186959 521380
rect 186993 521346 187051 521380
rect 187085 521346 187143 521380
rect 187177 521346 187235 521380
rect 187269 521346 187327 521380
rect 187361 521346 187419 521380
rect 187453 521346 187482 521380
rect 172227 521304 172469 521346
rect 172227 521270 172245 521304
rect 172279 521270 172417 521304
rect 172451 521270 172469 521304
rect 172227 521209 172469 521270
rect 172503 521304 173572 521346
rect 172503 521270 172521 521304
rect 172555 521270 173521 521304
rect 173555 521270 173572 521304
rect 172503 521259 173572 521270
rect 173607 521304 174676 521346
rect 173607 521270 173625 521304
rect 173659 521270 174625 521304
rect 174659 521270 174676 521304
rect 173607 521259 174676 521270
rect 174711 521304 175780 521346
rect 174711 521270 174729 521304
rect 174763 521270 175729 521304
rect 175763 521270 175780 521304
rect 174711 521259 175780 521270
rect 175815 521304 176884 521346
rect 175815 521270 175833 521304
rect 175867 521270 176833 521304
rect 176867 521270 176884 521304
rect 175815 521259 176884 521270
rect 176919 521304 177253 521346
rect 176919 521270 176937 521304
rect 176971 521270 177201 521304
rect 177235 521270 177253 521304
rect 172227 521175 172245 521209
rect 172279 521175 172417 521209
rect 172451 521175 172469 521209
rect 172227 521128 172469 521175
rect 172227 521060 172277 521094
rect 172311 521060 172331 521094
rect 172227 520986 172331 521060
rect 172365 521054 172469 521128
rect 172365 521020 172385 521054
rect 172419 521020 172469 521054
rect 172820 521094 172888 521111
rect 172820 521060 172837 521094
rect 172871 521060 172888 521094
rect 172227 520933 172469 520986
rect 172820 520945 172888 521060
rect 173184 521058 173254 521259
rect 173184 521024 173201 521058
rect 173235 521024 173254 521058
rect 173184 521009 173254 521024
rect 173924 521094 173992 521111
rect 173924 521060 173941 521094
rect 173975 521060 173992 521094
rect 173924 520945 173992 521060
rect 174288 521058 174358 521259
rect 174288 521024 174305 521058
rect 174339 521024 174358 521058
rect 174288 521009 174358 521024
rect 175028 521094 175096 521111
rect 175028 521060 175045 521094
rect 175079 521060 175096 521094
rect 175028 520945 175096 521060
rect 175392 521058 175462 521259
rect 175392 521024 175409 521058
rect 175443 521024 175462 521058
rect 175392 521009 175462 521024
rect 176132 521094 176200 521111
rect 176132 521060 176149 521094
rect 176183 521060 176200 521094
rect 176132 520945 176200 521060
rect 176496 521058 176566 521259
rect 176919 521202 177253 521270
rect 176919 521168 176937 521202
rect 176971 521168 177201 521202
rect 177235 521168 177253 521202
rect 176919 521128 177253 521168
rect 176496 521024 176513 521058
rect 176547 521024 176566 521058
rect 176496 521009 176566 521024
rect 176919 521060 176939 521094
rect 176973 521060 177069 521094
rect 176919 520990 177069 521060
rect 177103 521058 177253 521128
rect 177379 521275 177437 521346
rect 177379 521241 177391 521275
rect 177425 521241 177437 521275
rect 177471 521304 178540 521346
rect 177471 521270 177489 521304
rect 177523 521270 178489 521304
rect 178523 521270 178540 521304
rect 177471 521259 178540 521270
rect 178575 521304 179644 521346
rect 178575 521270 178593 521304
rect 178627 521270 179593 521304
rect 179627 521270 179644 521304
rect 178575 521259 179644 521270
rect 179679 521304 180748 521346
rect 179679 521270 179697 521304
rect 179731 521270 180697 521304
rect 180731 521270 180748 521304
rect 179679 521259 180748 521270
rect 180783 521304 181852 521346
rect 180783 521270 180801 521304
rect 180835 521270 181801 521304
rect 181835 521270 181852 521304
rect 180783 521259 181852 521270
rect 181887 521304 182405 521346
rect 181887 521270 181905 521304
rect 181939 521270 182353 521304
rect 182387 521270 182405 521304
rect 177379 521182 177437 521241
rect 177379 521148 177391 521182
rect 177425 521148 177437 521182
rect 177379 521113 177437 521148
rect 177103 521024 177199 521058
rect 177233 521024 177253 521058
rect 177788 521094 177856 521111
rect 177788 521060 177805 521094
rect 177839 521060 177856 521094
rect 172227 520899 172245 520933
rect 172279 520899 172417 520933
rect 172451 520899 172469 520933
rect 172227 520836 172469 520899
rect 172503 520931 173572 520945
rect 172503 520897 172521 520931
rect 172555 520897 173521 520931
rect 173555 520897 173572 520931
rect 172503 520836 173572 520897
rect 173607 520931 174676 520945
rect 173607 520897 173625 520931
rect 173659 520897 174625 520931
rect 174659 520897 174676 520931
rect 173607 520836 174676 520897
rect 174711 520931 175780 520945
rect 174711 520897 174729 520931
rect 174763 520897 175729 520931
rect 175763 520897 175780 520931
rect 174711 520836 175780 520897
rect 175815 520931 176884 520945
rect 175815 520897 175833 520931
rect 175867 520897 176833 520931
rect 176867 520897 176884 520931
rect 175815 520836 176884 520897
rect 176919 520938 177253 520990
rect 176919 520904 176937 520938
rect 176971 520904 177201 520938
rect 177235 520904 177253 520938
rect 176919 520836 177253 520904
rect 177379 520964 177437 520981
rect 177379 520930 177391 520964
rect 177425 520930 177437 520964
rect 177788 520945 177856 521060
rect 178152 521058 178222 521259
rect 178152 521024 178169 521058
rect 178203 521024 178222 521058
rect 178152 521009 178222 521024
rect 178892 521094 178960 521111
rect 178892 521060 178909 521094
rect 178943 521060 178960 521094
rect 178892 520945 178960 521060
rect 179256 521058 179326 521259
rect 179256 521024 179273 521058
rect 179307 521024 179326 521058
rect 179256 521009 179326 521024
rect 179996 521094 180064 521111
rect 179996 521060 180013 521094
rect 180047 521060 180064 521094
rect 179996 520945 180064 521060
rect 180360 521058 180430 521259
rect 180360 521024 180377 521058
rect 180411 521024 180430 521058
rect 180360 521009 180430 521024
rect 181100 521094 181168 521111
rect 181100 521060 181117 521094
rect 181151 521060 181168 521094
rect 181100 520945 181168 521060
rect 181464 521058 181534 521259
rect 181887 521202 182405 521270
rect 181887 521168 181905 521202
rect 181939 521168 182353 521202
rect 182387 521168 182405 521202
rect 181887 521128 182405 521168
rect 181464 521024 181481 521058
rect 181515 521024 181534 521058
rect 181464 521009 181534 521024
rect 181887 521060 181965 521094
rect 181999 521060 182075 521094
rect 182109 521060 182129 521094
rect 181887 520990 182129 521060
rect 182163 521058 182405 521128
rect 182531 521275 182589 521346
rect 182531 521241 182543 521275
rect 182577 521241 182589 521275
rect 182623 521304 183692 521346
rect 182623 521270 182641 521304
rect 182675 521270 183641 521304
rect 183675 521270 183692 521304
rect 182623 521259 183692 521270
rect 183727 521304 184796 521346
rect 183727 521270 183745 521304
rect 183779 521270 184745 521304
rect 184779 521270 184796 521304
rect 183727 521259 184796 521270
rect 184831 521304 185900 521346
rect 184831 521270 184849 521304
rect 184883 521270 185849 521304
rect 185883 521270 185900 521304
rect 184831 521259 185900 521270
rect 185935 521304 187004 521346
rect 185935 521270 185953 521304
rect 185987 521270 186953 521304
rect 186987 521270 187004 521304
rect 185935 521259 187004 521270
rect 187223 521304 187465 521346
rect 187223 521270 187241 521304
rect 187275 521270 187413 521304
rect 187447 521270 187465 521304
rect 182531 521182 182589 521241
rect 182531 521148 182543 521182
rect 182577 521148 182589 521182
rect 182531 521113 182589 521148
rect 182163 521024 182183 521058
rect 182217 521024 182293 521058
rect 182327 521024 182405 521058
rect 182940 521094 183008 521111
rect 182940 521060 182957 521094
rect 182991 521060 183008 521094
rect 177379 520836 177437 520930
rect 177471 520931 178540 520945
rect 177471 520897 177489 520931
rect 177523 520897 178489 520931
rect 178523 520897 178540 520931
rect 177471 520836 178540 520897
rect 178575 520931 179644 520945
rect 178575 520897 178593 520931
rect 178627 520897 179593 520931
rect 179627 520897 179644 520931
rect 178575 520836 179644 520897
rect 179679 520931 180748 520945
rect 179679 520897 179697 520931
rect 179731 520897 180697 520931
rect 180731 520897 180748 520931
rect 179679 520836 180748 520897
rect 180783 520931 181852 520945
rect 180783 520897 180801 520931
rect 180835 520897 181801 520931
rect 181835 520897 181852 520931
rect 180783 520836 181852 520897
rect 181887 520931 182405 520990
rect 181887 520897 181905 520931
rect 181939 520897 182353 520931
rect 182387 520897 182405 520931
rect 181887 520836 182405 520897
rect 182531 520964 182589 520981
rect 182531 520930 182543 520964
rect 182577 520930 182589 520964
rect 182940 520945 183008 521060
rect 183304 521058 183374 521259
rect 183304 521024 183321 521058
rect 183355 521024 183374 521058
rect 183304 521009 183374 521024
rect 184044 521094 184112 521111
rect 184044 521060 184061 521094
rect 184095 521060 184112 521094
rect 184044 520945 184112 521060
rect 184408 521058 184478 521259
rect 184408 521024 184425 521058
rect 184459 521024 184478 521058
rect 184408 521009 184478 521024
rect 185148 521094 185216 521111
rect 185148 521060 185165 521094
rect 185199 521060 185216 521094
rect 185148 520945 185216 521060
rect 185512 521058 185582 521259
rect 185512 521024 185529 521058
rect 185563 521024 185582 521058
rect 185512 521009 185582 521024
rect 186252 521094 186320 521111
rect 186252 521060 186269 521094
rect 186303 521060 186320 521094
rect 186252 520945 186320 521060
rect 186616 521058 186686 521259
rect 186616 521024 186633 521058
rect 186667 521024 186686 521058
rect 186616 521009 186686 521024
rect 187223 521209 187465 521270
rect 187223 521175 187241 521209
rect 187275 521175 187413 521209
rect 187447 521175 187465 521209
rect 187223 521128 187465 521175
rect 187223 521054 187327 521128
rect 187223 521020 187273 521054
rect 187307 521020 187327 521054
rect 187361 521060 187381 521094
rect 187415 521060 187465 521094
rect 187361 520986 187465 521060
rect 182531 520836 182589 520930
rect 182623 520931 183692 520945
rect 182623 520897 182641 520931
rect 182675 520897 183641 520931
rect 183675 520897 183692 520931
rect 182623 520836 183692 520897
rect 183727 520931 184796 520945
rect 183727 520897 183745 520931
rect 183779 520897 184745 520931
rect 184779 520897 184796 520931
rect 183727 520836 184796 520897
rect 184831 520931 185900 520945
rect 184831 520897 184849 520931
rect 184883 520897 185849 520931
rect 185883 520897 185900 520931
rect 184831 520836 185900 520897
rect 185935 520931 187004 520945
rect 185935 520897 185953 520931
rect 185987 520897 186953 520931
rect 186987 520897 187004 520931
rect 185935 520836 187004 520897
rect 187223 520933 187465 520986
rect 187223 520899 187241 520933
rect 187275 520899 187413 520933
rect 187447 520899 187465 520933
rect 187223 520836 187465 520899
rect 172210 520802 172239 520836
rect 172273 520802 172331 520836
rect 172365 520802 172423 520836
rect 172457 520802 172515 520836
rect 172549 520802 172607 520836
rect 172641 520802 172699 520836
rect 172733 520802 172791 520836
rect 172825 520802 172883 520836
rect 172917 520802 172975 520836
rect 173009 520802 173067 520836
rect 173101 520802 173159 520836
rect 173193 520802 173251 520836
rect 173285 520802 173343 520836
rect 173377 520802 173435 520836
rect 173469 520802 173527 520836
rect 173561 520802 173619 520836
rect 173653 520802 173711 520836
rect 173745 520802 173803 520836
rect 173837 520802 173895 520836
rect 173929 520802 173987 520836
rect 174021 520802 174079 520836
rect 174113 520802 174171 520836
rect 174205 520802 174263 520836
rect 174297 520802 174355 520836
rect 174389 520802 174447 520836
rect 174481 520802 174539 520836
rect 174573 520802 174631 520836
rect 174665 520802 174723 520836
rect 174757 520802 174815 520836
rect 174849 520802 174907 520836
rect 174941 520802 174999 520836
rect 175033 520802 175091 520836
rect 175125 520802 175183 520836
rect 175217 520802 175275 520836
rect 175309 520802 175367 520836
rect 175401 520802 175459 520836
rect 175493 520802 175551 520836
rect 175585 520802 175643 520836
rect 175677 520802 175735 520836
rect 175769 520802 175827 520836
rect 175861 520802 175919 520836
rect 175953 520802 176011 520836
rect 176045 520802 176103 520836
rect 176137 520802 176195 520836
rect 176229 520802 176287 520836
rect 176321 520802 176379 520836
rect 176413 520802 176471 520836
rect 176505 520802 176563 520836
rect 176597 520802 176655 520836
rect 176689 520802 176747 520836
rect 176781 520802 176839 520836
rect 176873 520802 176931 520836
rect 176965 520802 177023 520836
rect 177057 520802 177115 520836
rect 177149 520802 177207 520836
rect 177241 520802 177299 520836
rect 177333 520802 177391 520836
rect 177425 520802 177483 520836
rect 177517 520802 177575 520836
rect 177609 520802 177667 520836
rect 177701 520802 177759 520836
rect 177793 520802 177851 520836
rect 177885 520802 177943 520836
rect 177977 520802 178035 520836
rect 178069 520802 178127 520836
rect 178161 520802 178219 520836
rect 178253 520802 178311 520836
rect 178345 520802 178403 520836
rect 178437 520802 178495 520836
rect 178529 520802 178587 520836
rect 178621 520802 178679 520836
rect 178713 520802 178771 520836
rect 178805 520802 178863 520836
rect 178897 520802 178955 520836
rect 178989 520802 179047 520836
rect 179081 520802 179139 520836
rect 179173 520802 179231 520836
rect 179265 520802 179323 520836
rect 179357 520802 179415 520836
rect 179449 520802 179507 520836
rect 179541 520802 179599 520836
rect 179633 520802 179691 520836
rect 179725 520802 179783 520836
rect 179817 520802 179875 520836
rect 179909 520802 179967 520836
rect 180001 520802 180059 520836
rect 180093 520802 180151 520836
rect 180185 520802 180243 520836
rect 180277 520802 180335 520836
rect 180369 520802 180427 520836
rect 180461 520802 180519 520836
rect 180553 520802 180611 520836
rect 180645 520802 180703 520836
rect 180737 520802 180795 520836
rect 180829 520802 180887 520836
rect 180921 520802 180979 520836
rect 181013 520802 181071 520836
rect 181105 520802 181163 520836
rect 181197 520802 181255 520836
rect 181289 520802 181347 520836
rect 181381 520802 181439 520836
rect 181473 520802 181531 520836
rect 181565 520802 181623 520836
rect 181657 520802 181715 520836
rect 181749 520802 181807 520836
rect 181841 520802 181899 520836
rect 181933 520802 181991 520836
rect 182025 520802 182083 520836
rect 182117 520802 182175 520836
rect 182209 520802 182267 520836
rect 182301 520802 182359 520836
rect 182393 520802 182451 520836
rect 182485 520802 182543 520836
rect 182577 520802 182635 520836
rect 182669 520802 182727 520836
rect 182761 520802 182819 520836
rect 182853 520802 182911 520836
rect 182945 520802 183003 520836
rect 183037 520802 183095 520836
rect 183129 520802 183187 520836
rect 183221 520802 183279 520836
rect 183313 520802 183371 520836
rect 183405 520802 183463 520836
rect 183497 520802 183555 520836
rect 183589 520802 183647 520836
rect 183681 520802 183739 520836
rect 183773 520802 183831 520836
rect 183865 520802 183923 520836
rect 183957 520802 184015 520836
rect 184049 520802 184107 520836
rect 184141 520802 184199 520836
rect 184233 520802 184291 520836
rect 184325 520802 184383 520836
rect 184417 520802 184475 520836
rect 184509 520802 184567 520836
rect 184601 520802 184659 520836
rect 184693 520802 184751 520836
rect 184785 520802 184843 520836
rect 184877 520802 184935 520836
rect 184969 520802 185027 520836
rect 185061 520802 185119 520836
rect 185153 520802 185211 520836
rect 185245 520802 185303 520836
rect 185337 520802 185395 520836
rect 185429 520802 185487 520836
rect 185521 520802 185579 520836
rect 185613 520802 185671 520836
rect 185705 520802 185763 520836
rect 185797 520802 185855 520836
rect 185889 520802 185947 520836
rect 185981 520802 186039 520836
rect 186073 520802 186131 520836
rect 186165 520802 186223 520836
rect 186257 520802 186315 520836
rect 186349 520802 186407 520836
rect 186441 520802 186499 520836
rect 186533 520802 186591 520836
rect 186625 520802 186683 520836
rect 186717 520802 186775 520836
rect 186809 520802 186867 520836
rect 186901 520802 186959 520836
rect 186993 520802 187051 520836
rect 187085 520802 187143 520836
rect 187177 520802 187235 520836
rect 187269 520802 187327 520836
rect 187361 520802 187419 520836
rect 187453 520802 187482 520836
rect 172227 520739 172469 520802
rect 172227 520705 172245 520739
rect 172279 520705 172417 520739
rect 172451 520705 172469 520739
rect 172227 520652 172469 520705
rect 172503 520741 173572 520802
rect 172503 520707 172521 520741
rect 172555 520707 173521 520741
rect 173555 520707 173572 520741
rect 172503 520693 173572 520707
rect 173607 520741 174676 520802
rect 173607 520707 173625 520741
rect 173659 520707 174625 520741
rect 174659 520707 174676 520741
rect 173607 520693 174676 520707
rect 174803 520708 174861 520802
rect 172227 520578 172331 520652
rect 172227 520544 172277 520578
rect 172311 520544 172331 520578
rect 172365 520584 172385 520618
rect 172419 520584 172469 520618
rect 172365 520510 172469 520584
rect 172820 520578 172888 520693
rect 172820 520544 172837 520578
rect 172871 520544 172888 520578
rect 172820 520527 172888 520544
rect 173184 520614 173254 520629
rect 173184 520580 173201 520614
rect 173235 520580 173254 520614
rect 172227 520463 172469 520510
rect 172227 520429 172245 520463
rect 172279 520429 172417 520463
rect 172451 520429 172469 520463
rect 172227 520368 172469 520429
rect 173184 520379 173254 520580
rect 173924 520578 173992 520693
rect 174803 520674 174815 520708
rect 174849 520674 174861 520708
rect 174895 520741 175964 520802
rect 174895 520707 174913 520741
rect 174947 520707 175913 520741
rect 175947 520707 175964 520741
rect 174895 520693 175964 520707
rect 175999 520741 177068 520802
rect 175999 520707 176017 520741
rect 176051 520707 177017 520741
rect 177051 520707 177068 520741
rect 175999 520693 177068 520707
rect 177103 520741 178172 520802
rect 177103 520707 177121 520741
rect 177155 520707 178121 520741
rect 178155 520707 178172 520741
rect 177103 520693 178172 520707
rect 178207 520741 179276 520802
rect 178207 520707 178225 520741
rect 178259 520707 179225 520741
rect 179259 520707 179276 520741
rect 178207 520693 179276 520707
rect 179311 520741 179829 520802
rect 179311 520707 179329 520741
rect 179363 520707 179777 520741
rect 179811 520707 179829 520741
rect 174803 520657 174861 520674
rect 173924 520544 173941 520578
rect 173975 520544 173992 520578
rect 173924 520527 173992 520544
rect 174288 520614 174358 520629
rect 174288 520580 174305 520614
rect 174339 520580 174358 520614
rect 174288 520379 174358 520580
rect 175212 520578 175280 520693
rect 175212 520544 175229 520578
rect 175263 520544 175280 520578
rect 175212 520527 175280 520544
rect 175576 520614 175646 520629
rect 175576 520580 175593 520614
rect 175627 520580 175646 520614
rect 174803 520490 174861 520525
rect 174803 520456 174815 520490
rect 174849 520456 174861 520490
rect 174803 520397 174861 520456
rect 172227 520334 172245 520368
rect 172279 520334 172417 520368
rect 172451 520334 172469 520368
rect 172227 520292 172469 520334
rect 172503 520368 173572 520379
rect 172503 520334 172521 520368
rect 172555 520334 173521 520368
rect 173555 520334 173572 520368
rect 172503 520292 173572 520334
rect 173607 520368 174676 520379
rect 173607 520334 173625 520368
rect 173659 520334 174625 520368
rect 174659 520334 174676 520368
rect 173607 520292 174676 520334
rect 174803 520363 174815 520397
rect 174849 520363 174861 520397
rect 175576 520379 175646 520580
rect 176316 520578 176384 520693
rect 176316 520544 176333 520578
rect 176367 520544 176384 520578
rect 176316 520527 176384 520544
rect 176680 520614 176750 520629
rect 176680 520580 176697 520614
rect 176731 520580 176750 520614
rect 176680 520379 176750 520580
rect 177420 520578 177488 520693
rect 177420 520544 177437 520578
rect 177471 520544 177488 520578
rect 177420 520527 177488 520544
rect 177784 520614 177854 520629
rect 177784 520580 177801 520614
rect 177835 520580 177854 520614
rect 177784 520379 177854 520580
rect 178524 520578 178592 520693
rect 179311 520648 179829 520707
rect 179955 520708 180013 520802
rect 179955 520674 179967 520708
rect 180001 520674 180013 520708
rect 180047 520741 181116 520802
rect 180047 520707 180065 520741
rect 180099 520707 181065 520741
rect 181099 520707 181116 520741
rect 180047 520693 181116 520707
rect 181151 520741 182220 520802
rect 181151 520707 181169 520741
rect 181203 520707 182169 520741
rect 182203 520707 182220 520741
rect 181151 520693 182220 520707
rect 182255 520741 183324 520802
rect 182255 520707 182273 520741
rect 182307 520707 183273 520741
rect 183307 520707 183324 520741
rect 182255 520693 183324 520707
rect 183359 520741 184428 520802
rect 183359 520707 183377 520741
rect 183411 520707 184377 520741
rect 184411 520707 184428 520741
rect 183359 520693 184428 520707
rect 184463 520741 184981 520802
rect 184463 520707 184481 520741
rect 184515 520707 184929 520741
rect 184963 520707 184981 520741
rect 179955 520657 180013 520674
rect 178524 520544 178541 520578
rect 178575 520544 178592 520578
rect 178524 520527 178592 520544
rect 178888 520614 178958 520629
rect 178888 520580 178905 520614
rect 178939 520580 178958 520614
rect 178888 520379 178958 520580
rect 179311 520578 179553 520648
rect 179311 520544 179389 520578
rect 179423 520544 179499 520578
rect 179533 520544 179553 520578
rect 179587 520580 179607 520614
rect 179641 520580 179717 520614
rect 179751 520580 179829 520614
rect 179587 520510 179829 520580
rect 180364 520578 180432 520693
rect 180364 520544 180381 520578
rect 180415 520544 180432 520578
rect 180364 520527 180432 520544
rect 180728 520614 180798 520629
rect 180728 520580 180745 520614
rect 180779 520580 180798 520614
rect 179311 520470 179829 520510
rect 179311 520436 179329 520470
rect 179363 520436 179777 520470
rect 179811 520436 179829 520470
rect 174803 520292 174861 520363
rect 174895 520368 175964 520379
rect 174895 520334 174913 520368
rect 174947 520334 175913 520368
rect 175947 520334 175964 520368
rect 174895 520292 175964 520334
rect 175999 520368 177068 520379
rect 175999 520334 176017 520368
rect 176051 520334 177017 520368
rect 177051 520334 177068 520368
rect 175999 520292 177068 520334
rect 177103 520368 178172 520379
rect 177103 520334 177121 520368
rect 177155 520334 178121 520368
rect 178155 520334 178172 520368
rect 177103 520292 178172 520334
rect 178207 520368 179276 520379
rect 178207 520334 178225 520368
rect 178259 520334 179225 520368
rect 179259 520334 179276 520368
rect 178207 520292 179276 520334
rect 179311 520368 179829 520436
rect 179311 520334 179329 520368
rect 179363 520334 179777 520368
rect 179811 520334 179829 520368
rect 179311 520292 179829 520334
rect 179955 520490 180013 520525
rect 179955 520456 179967 520490
rect 180001 520456 180013 520490
rect 179955 520397 180013 520456
rect 179955 520363 179967 520397
rect 180001 520363 180013 520397
rect 180728 520379 180798 520580
rect 181468 520578 181536 520693
rect 181468 520544 181485 520578
rect 181519 520544 181536 520578
rect 181468 520527 181536 520544
rect 181832 520614 181902 520629
rect 181832 520580 181849 520614
rect 181883 520580 181902 520614
rect 181832 520379 181902 520580
rect 182572 520578 182640 520693
rect 182572 520544 182589 520578
rect 182623 520544 182640 520578
rect 182572 520527 182640 520544
rect 182936 520614 183006 520629
rect 182936 520580 182953 520614
rect 182987 520580 183006 520614
rect 182936 520379 183006 520580
rect 183676 520578 183744 520693
rect 184463 520648 184981 520707
rect 185107 520708 185165 520802
rect 185107 520674 185119 520708
rect 185153 520674 185165 520708
rect 185199 520741 186268 520802
rect 185199 520707 185217 520741
rect 185251 520707 186217 520741
rect 186251 520707 186268 520741
rect 185199 520693 186268 520707
rect 186303 520741 187005 520802
rect 186303 520707 186321 520741
rect 186355 520707 186953 520741
rect 186987 520707 187005 520741
rect 185107 520657 185165 520674
rect 183676 520544 183693 520578
rect 183727 520544 183744 520578
rect 183676 520527 183744 520544
rect 184040 520614 184110 520629
rect 184040 520580 184057 520614
rect 184091 520580 184110 520614
rect 184040 520379 184110 520580
rect 184463 520578 184705 520648
rect 184463 520544 184541 520578
rect 184575 520544 184651 520578
rect 184685 520544 184705 520578
rect 184739 520580 184759 520614
rect 184793 520580 184869 520614
rect 184903 520580 184981 520614
rect 184739 520510 184981 520580
rect 185516 520578 185584 520693
rect 186303 520648 187005 520707
rect 187223 520739 187465 520802
rect 187223 520705 187241 520739
rect 187275 520705 187413 520739
rect 187447 520705 187465 520739
rect 187223 520652 187465 520705
rect 185516 520544 185533 520578
rect 185567 520544 185584 520578
rect 185516 520527 185584 520544
rect 185880 520614 185950 520629
rect 185880 520580 185897 520614
rect 185931 520580 185950 520614
rect 184463 520470 184981 520510
rect 184463 520436 184481 520470
rect 184515 520436 184929 520470
rect 184963 520436 184981 520470
rect 179955 520292 180013 520363
rect 180047 520368 181116 520379
rect 180047 520334 180065 520368
rect 180099 520334 181065 520368
rect 181099 520334 181116 520368
rect 180047 520292 181116 520334
rect 181151 520368 182220 520379
rect 181151 520334 181169 520368
rect 181203 520334 182169 520368
rect 182203 520334 182220 520368
rect 181151 520292 182220 520334
rect 182255 520368 183324 520379
rect 182255 520334 182273 520368
rect 182307 520334 183273 520368
rect 183307 520334 183324 520368
rect 182255 520292 183324 520334
rect 183359 520368 184428 520379
rect 183359 520334 183377 520368
rect 183411 520334 184377 520368
rect 184411 520334 184428 520368
rect 183359 520292 184428 520334
rect 184463 520368 184981 520436
rect 184463 520334 184481 520368
rect 184515 520334 184929 520368
rect 184963 520334 184981 520368
rect 184463 520292 184981 520334
rect 185107 520490 185165 520525
rect 185107 520456 185119 520490
rect 185153 520456 185165 520490
rect 185107 520397 185165 520456
rect 185107 520363 185119 520397
rect 185153 520363 185165 520397
rect 185880 520379 185950 520580
rect 186303 520578 186633 520648
rect 186303 520544 186381 520578
rect 186415 520544 186480 520578
rect 186514 520544 186579 520578
rect 186613 520544 186633 520578
rect 186667 520580 186687 520614
rect 186721 520580 186790 520614
rect 186824 520580 186893 520614
rect 186927 520580 187005 520614
rect 186667 520510 187005 520580
rect 186303 520470 187005 520510
rect 186303 520436 186321 520470
rect 186355 520436 186953 520470
rect 186987 520436 187005 520470
rect 185107 520292 185165 520363
rect 185199 520368 186268 520379
rect 185199 520334 185217 520368
rect 185251 520334 186217 520368
rect 186251 520334 186268 520368
rect 185199 520292 186268 520334
rect 186303 520368 187005 520436
rect 186303 520334 186321 520368
rect 186355 520334 186953 520368
rect 186987 520334 187005 520368
rect 186303 520292 187005 520334
rect 187223 520584 187273 520618
rect 187307 520584 187327 520618
rect 187223 520510 187327 520584
rect 187361 520578 187465 520652
rect 187361 520544 187381 520578
rect 187415 520544 187465 520578
rect 187223 520463 187465 520510
rect 187223 520429 187241 520463
rect 187275 520429 187413 520463
rect 187447 520429 187465 520463
rect 187223 520368 187465 520429
rect 187223 520334 187241 520368
rect 187275 520334 187413 520368
rect 187447 520334 187465 520368
rect 187223 520292 187465 520334
rect 172210 520258 172239 520292
rect 172273 520258 172331 520292
rect 172365 520258 172423 520292
rect 172457 520258 172515 520292
rect 172549 520258 172607 520292
rect 172641 520258 172699 520292
rect 172733 520258 172791 520292
rect 172825 520258 172883 520292
rect 172917 520258 172975 520292
rect 173009 520258 173067 520292
rect 173101 520258 173159 520292
rect 173193 520258 173251 520292
rect 173285 520258 173343 520292
rect 173377 520258 173435 520292
rect 173469 520258 173527 520292
rect 173561 520258 173619 520292
rect 173653 520258 173711 520292
rect 173745 520258 173803 520292
rect 173837 520258 173895 520292
rect 173929 520258 173987 520292
rect 174021 520258 174079 520292
rect 174113 520258 174171 520292
rect 174205 520258 174263 520292
rect 174297 520258 174355 520292
rect 174389 520258 174447 520292
rect 174481 520258 174539 520292
rect 174573 520258 174631 520292
rect 174665 520258 174723 520292
rect 174757 520258 174815 520292
rect 174849 520258 174907 520292
rect 174941 520258 174999 520292
rect 175033 520258 175091 520292
rect 175125 520258 175183 520292
rect 175217 520258 175275 520292
rect 175309 520258 175367 520292
rect 175401 520258 175459 520292
rect 175493 520258 175551 520292
rect 175585 520258 175643 520292
rect 175677 520258 175735 520292
rect 175769 520258 175827 520292
rect 175861 520258 175919 520292
rect 175953 520258 176011 520292
rect 176045 520258 176103 520292
rect 176137 520258 176195 520292
rect 176229 520258 176287 520292
rect 176321 520258 176379 520292
rect 176413 520258 176471 520292
rect 176505 520258 176563 520292
rect 176597 520258 176655 520292
rect 176689 520258 176747 520292
rect 176781 520258 176839 520292
rect 176873 520258 176931 520292
rect 176965 520258 177023 520292
rect 177057 520258 177115 520292
rect 177149 520258 177207 520292
rect 177241 520258 177299 520292
rect 177333 520258 177391 520292
rect 177425 520258 177483 520292
rect 177517 520258 177575 520292
rect 177609 520258 177667 520292
rect 177701 520258 177759 520292
rect 177793 520258 177851 520292
rect 177885 520258 177943 520292
rect 177977 520258 178035 520292
rect 178069 520258 178127 520292
rect 178161 520258 178219 520292
rect 178253 520258 178311 520292
rect 178345 520258 178403 520292
rect 178437 520258 178495 520292
rect 178529 520258 178587 520292
rect 178621 520258 178679 520292
rect 178713 520258 178771 520292
rect 178805 520258 178863 520292
rect 178897 520258 178955 520292
rect 178989 520258 179047 520292
rect 179081 520258 179139 520292
rect 179173 520258 179231 520292
rect 179265 520258 179323 520292
rect 179357 520258 179415 520292
rect 179449 520258 179507 520292
rect 179541 520258 179599 520292
rect 179633 520258 179691 520292
rect 179725 520258 179783 520292
rect 179817 520258 179875 520292
rect 179909 520258 179967 520292
rect 180001 520258 180059 520292
rect 180093 520258 180151 520292
rect 180185 520258 180243 520292
rect 180277 520258 180335 520292
rect 180369 520258 180427 520292
rect 180461 520258 180519 520292
rect 180553 520258 180611 520292
rect 180645 520258 180703 520292
rect 180737 520258 180795 520292
rect 180829 520258 180887 520292
rect 180921 520258 180979 520292
rect 181013 520258 181071 520292
rect 181105 520258 181163 520292
rect 181197 520258 181255 520292
rect 181289 520258 181347 520292
rect 181381 520258 181439 520292
rect 181473 520258 181531 520292
rect 181565 520258 181623 520292
rect 181657 520258 181715 520292
rect 181749 520258 181807 520292
rect 181841 520258 181899 520292
rect 181933 520258 181991 520292
rect 182025 520258 182083 520292
rect 182117 520258 182175 520292
rect 182209 520258 182267 520292
rect 182301 520258 182359 520292
rect 182393 520258 182451 520292
rect 182485 520258 182543 520292
rect 182577 520258 182635 520292
rect 182669 520258 182727 520292
rect 182761 520258 182819 520292
rect 182853 520258 182911 520292
rect 182945 520258 183003 520292
rect 183037 520258 183095 520292
rect 183129 520258 183187 520292
rect 183221 520258 183279 520292
rect 183313 520258 183371 520292
rect 183405 520258 183463 520292
rect 183497 520258 183555 520292
rect 183589 520258 183647 520292
rect 183681 520258 183739 520292
rect 183773 520258 183831 520292
rect 183865 520258 183923 520292
rect 183957 520258 184015 520292
rect 184049 520258 184107 520292
rect 184141 520258 184199 520292
rect 184233 520258 184291 520292
rect 184325 520258 184383 520292
rect 184417 520258 184475 520292
rect 184509 520258 184567 520292
rect 184601 520258 184659 520292
rect 184693 520258 184751 520292
rect 184785 520258 184843 520292
rect 184877 520258 184935 520292
rect 184969 520258 185027 520292
rect 185061 520258 185119 520292
rect 185153 520258 185211 520292
rect 185245 520258 185303 520292
rect 185337 520258 185395 520292
rect 185429 520258 185487 520292
rect 185521 520258 185579 520292
rect 185613 520258 185671 520292
rect 185705 520258 185763 520292
rect 185797 520258 185855 520292
rect 185889 520258 185947 520292
rect 185981 520258 186039 520292
rect 186073 520258 186131 520292
rect 186165 520258 186223 520292
rect 186257 520258 186315 520292
rect 186349 520258 186407 520292
rect 186441 520258 186499 520292
rect 186533 520258 186591 520292
rect 186625 520258 186683 520292
rect 186717 520258 186775 520292
rect 186809 520258 186867 520292
rect 186901 520258 186959 520292
rect 186993 520258 187051 520292
rect 187085 520258 187143 520292
rect 187177 520258 187235 520292
rect 187269 520258 187327 520292
rect 187361 520258 187419 520292
rect 187453 520258 187482 520292
rect 172227 520216 172469 520258
rect 172227 520182 172245 520216
rect 172279 520182 172417 520216
rect 172451 520182 172469 520216
rect 172227 520121 172469 520182
rect 172503 520216 173572 520258
rect 172503 520182 172521 520216
rect 172555 520182 173521 520216
rect 173555 520182 173572 520216
rect 172503 520171 173572 520182
rect 173607 520216 174676 520258
rect 173607 520182 173625 520216
rect 173659 520182 174625 520216
rect 174659 520182 174676 520216
rect 173607 520171 174676 520182
rect 174711 520216 175780 520258
rect 174711 520182 174729 520216
rect 174763 520182 175729 520216
rect 175763 520182 175780 520216
rect 174711 520171 175780 520182
rect 175815 520216 176884 520258
rect 175815 520182 175833 520216
rect 175867 520182 176833 520216
rect 176867 520182 176884 520216
rect 175815 520171 176884 520182
rect 176919 520216 177253 520258
rect 176919 520182 176937 520216
rect 176971 520182 177201 520216
rect 177235 520182 177253 520216
rect 172227 520087 172245 520121
rect 172279 520087 172417 520121
rect 172451 520087 172469 520121
rect 172227 520040 172469 520087
rect 172227 519972 172277 520006
rect 172311 519972 172331 520006
rect 172227 519898 172331 519972
rect 172365 519966 172469 520040
rect 172365 519932 172385 519966
rect 172419 519932 172469 519966
rect 172820 520006 172888 520023
rect 172820 519972 172837 520006
rect 172871 519972 172888 520006
rect 172227 519845 172469 519898
rect 172820 519857 172888 519972
rect 173184 519970 173254 520171
rect 173184 519936 173201 519970
rect 173235 519936 173254 519970
rect 173184 519921 173254 519936
rect 173924 520006 173992 520023
rect 173924 519972 173941 520006
rect 173975 519972 173992 520006
rect 173924 519857 173992 519972
rect 174288 519970 174358 520171
rect 174288 519936 174305 519970
rect 174339 519936 174358 519970
rect 174288 519921 174358 519936
rect 175028 520006 175096 520023
rect 175028 519972 175045 520006
rect 175079 519972 175096 520006
rect 175028 519857 175096 519972
rect 175392 519970 175462 520171
rect 175392 519936 175409 519970
rect 175443 519936 175462 519970
rect 175392 519921 175462 519936
rect 176132 520006 176200 520023
rect 176132 519972 176149 520006
rect 176183 519972 176200 520006
rect 176132 519857 176200 519972
rect 176496 519970 176566 520171
rect 176919 520114 177253 520182
rect 176919 520080 176937 520114
rect 176971 520080 177201 520114
rect 177235 520080 177253 520114
rect 176919 520040 177253 520080
rect 176496 519936 176513 519970
rect 176547 519936 176566 519970
rect 176496 519921 176566 519936
rect 176919 519972 176939 520006
rect 176973 519972 177069 520006
rect 176919 519902 177069 519972
rect 177103 519970 177253 520040
rect 177379 520187 177437 520258
rect 177379 520153 177391 520187
rect 177425 520153 177437 520187
rect 177471 520216 178540 520258
rect 177471 520182 177489 520216
rect 177523 520182 178489 520216
rect 178523 520182 178540 520216
rect 177471 520171 178540 520182
rect 178575 520216 179644 520258
rect 178575 520182 178593 520216
rect 178627 520182 179593 520216
rect 179627 520182 179644 520216
rect 178575 520171 179644 520182
rect 179679 520216 180748 520258
rect 179679 520182 179697 520216
rect 179731 520182 180697 520216
rect 180731 520182 180748 520216
rect 179679 520171 180748 520182
rect 180783 520216 181852 520258
rect 180783 520182 180801 520216
rect 180835 520182 181801 520216
rect 181835 520182 181852 520216
rect 180783 520171 181852 520182
rect 181887 520216 182405 520258
rect 181887 520182 181905 520216
rect 181939 520182 182353 520216
rect 182387 520182 182405 520216
rect 177379 520094 177437 520153
rect 177379 520060 177391 520094
rect 177425 520060 177437 520094
rect 177379 520025 177437 520060
rect 177103 519936 177199 519970
rect 177233 519936 177253 519970
rect 177788 520006 177856 520023
rect 177788 519972 177805 520006
rect 177839 519972 177856 520006
rect 172227 519811 172245 519845
rect 172279 519811 172417 519845
rect 172451 519811 172469 519845
rect 172227 519748 172469 519811
rect 172503 519843 173572 519857
rect 172503 519809 172521 519843
rect 172555 519809 173521 519843
rect 173555 519809 173572 519843
rect 172503 519748 173572 519809
rect 173607 519843 174676 519857
rect 173607 519809 173625 519843
rect 173659 519809 174625 519843
rect 174659 519809 174676 519843
rect 173607 519748 174676 519809
rect 174711 519843 175780 519857
rect 174711 519809 174729 519843
rect 174763 519809 175729 519843
rect 175763 519809 175780 519843
rect 174711 519748 175780 519809
rect 175815 519843 176884 519857
rect 175815 519809 175833 519843
rect 175867 519809 176833 519843
rect 176867 519809 176884 519843
rect 175815 519748 176884 519809
rect 176919 519850 177253 519902
rect 176919 519816 176937 519850
rect 176971 519816 177201 519850
rect 177235 519816 177253 519850
rect 176919 519748 177253 519816
rect 177379 519876 177437 519893
rect 177379 519842 177391 519876
rect 177425 519842 177437 519876
rect 177788 519857 177856 519972
rect 178152 519970 178222 520171
rect 178152 519936 178169 519970
rect 178203 519936 178222 519970
rect 178152 519921 178222 519936
rect 178892 520006 178960 520023
rect 178892 519972 178909 520006
rect 178943 519972 178960 520006
rect 178892 519857 178960 519972
rect 179256 519970 179326 520171
rect 179256 519936 179273 519970
rect 179307 519936 179326 519970
rect 179256 519921 179326 519936
rect 179996 520006 180064 520023
rect 179996 519972 180013 520006
rect 180047 519972 180064 520006
rect 179996 519857 180064 519972
rect 180360 519970 180430 520171
rect 180360 519936 180377 519970
rect 180411 519936 180430 519970
rect 180360 519921 180430 519936
rect 181100 520006 181168 520023
rect 181100 519972 181117 520006
rect 181151 519972 181168 520006
rect 181100 519857 181168 519972
rect 181464 519970 181534 520171
rect 181887 520114 182405 520182
rect 181887 520080 181905 520114
rect 181939 520080 182353 520114
rect 182387 520080 182405 520114
rect 181887 520040 182405 520080
rect 181464 519936 181481 519970
rect 181515 519936 181534 519970
rect 181464 519921 181534 519936
rect 181887 519972 181965 520006
rect 181999 519972 182075 520006
rect 182109 519972 182129 520006
rect 181887 519902 182129 519972
rect 182163 519970 182405 520040
rect 182531 520187 182589 520258
rect 182531 520153 182543 520187
rect 182577 520153 182589 520187
rect 182623 520216 183692 520258
rect 182623 520182 182641 520216
rect 182675 520182 183641 520216
rect 183675 520182 183692 520216
rect 182623 520171 183692 520182
rect 183727 520216 184796 520258
rect 183727 520182 183745 520216
rect 183779 520182 184745 520216
rect 184779 520182 184796 520216
rect 183727 520171 184796 520182
rect 184831 520216 185900 520258
rect 184831 520182 184849 520216
rect 184883 520182 185849 520216
rect 185883 520182 185900 520216
rect 184831 520171 185900 520182
rect 185935 520216 187004 520258
rect 185935 520182 185953 520216
rect 185987 520182 186953 520216
rect 186987 520182 187004 520216
rect 185935 520171 187004 520182
rect 187223 520216 187465 520258
rect 187223 520182 187241 520216
rect 187275 520182 187413 520216
rect 187447 520182 187465 520216
rect 182531 520094 182589 520153
rect 182531 520060 182543 520094
rect 182577 520060 182589 520094
rect 182531 520025 182589 520060
rect 182163 519936 182183 519970
rect 182217 519936 182293 519970
rect 182327 519936 182405 519970
rect 182940 520006 183008 520023
rect 182940 519972 182957 520006
rect 182991 519972 183008 520006
rect 177379 519748 177437 519842
rect 177471 519843 178540 519857
rect 177471 519809 177489 519843
rect 177523 519809 178489 519843
rect 178523 519809 178540 519843
rect 177471 519748 178540 519809
rect 178575 519843 179644 519857
rect 178575 519809 178593 519843
rect 178627 519809 179593 519843
rect 179627 519809 179644 519843
rect 178575 519748 179644 519809
rect 179679 519843 180748 519857
rect 179679 519809 179697 519843
rect 179731 519809 180697 519843
rect 180731 519809 180748 519843
rect 179679 519748 180748 519809
rect 180783 519843 181852 519857
rect 180783 519809 180801 519843
rect 180835 519809 181801 519843
rect 181835 519809 181852 519843
rect 180783 519748 181852 519809
rect 181887 519843 182405 519902
rect 181887 519809 181905 519843
rect 181939 519809 182353 519843
rect 182387 519809 182405 519843
rect 181887 519748 182405 519809
rect 182531 519876 182589 519893
rect 182531 519842 182543 519876
rect 182577 519842 182589 519876
rect 182940 519857 183008 519972
rect 183304 519970 183374 520171
rect 183304 519936 183321 519970
rect 183355 519936 183374 519970
rect 183304 519921 183374 519936
rect 184044 520006 184112 520023
rect 184044 519972 184061 520006
rect 184095 519972 184112 520006
rect 184044 519857 184112 519972
rect 184408 519970 184478 520171
rect 184408 519936 184425 519970
rect 184459 519936 184478 519970
rect 184408 519921 184478 519936
rect 185148 520006 185216 520023
rect 185148 519972 185165 520006
rect 185199 519972 185216 520006
rect 185148 519857 185216 519972
rect 185512 519970 185582 520171
rect 185512 519936 185529 519970
rect 185563 519936 185582 519970
rect 185512 519921 185582 519936
rect 186252 520006 186320 520023
rect 186252 519972 186269 520006
rect 186303 519972 186320 520006
rect 186252 519857 186320 519972
rect 186616 519970 186686 520171
rect 186616 519936 186633 519970
rect 186667 519936 186686 519970
rect 186616 519921 186686 519936
rect 187223 520121 187465 520182
rect 187223 520087 187241 520121
rect 187275 520087 187413 520121
rect 187447 520087 187465 520121
rect 187223 520040 187465 520087
rect 187223 519966 187327 520040
rect 187223 519932 187273 519966
rect 187307 519932 187327 519966
rect 187361 519972 187381 520006
rect 187415 519972 187465 520006
rect 187361 519898 187465 519972
rect 182531 519748 182589 519842
rect 182623 519843 183692 519857
rect 182623 519809 182641 519843
rect 182675 519809 183641 519843
rect 183675 519809 183692 519843
rect 182623 519748 183692 519809
rect 183727 519843 184796 519857
rect 183727 519809 183745 519843
rect 183779 519809 184745 519843
rect 184779 519809 184796 519843
rect 183727 519748 184796 519809
rect 184831 519843 185900 519857
rect 184831 519809 184849 519843
rect 184883 519809 185849 519843
rect 185883 519809 185900 519843
rect 184831 519748 185900 519809
rect 185935 519843 187004 519857
rect 185935 519809 185953 519843
rect 185987 519809 186953 519843
rect 186987 519809 187004 519843
rect 185935 519748 187004 519809
rect 187223 519845 187465 519898
rect 187223 519811 187241 519845
rect 187275 519811 187413 519845
rect 187447 519811 187465 519845
rect 187223 519748 187465 519811
rect 172210 519714 172239 519748
rect 172273 519714 172331 519748
rect 172365 519714 172423 519748
rect 172457 519714 172515 519748
rect 172549 519714 172607 519748
rect 172641 519714 172699 519748
rect 172733 519714 172791 519748
rect 172825 519714 172883 519748
rect 172917 519714 172975 519748
rect 173009 519714 173067 519748
rect 173101 519714 173159 519748
rect 173193 519714 173251 519748
rect 173285 519714 173343 519748
rect 173377 519714 173435 519748
rect 173469 519714 173527 519748
rect 173561 519714 173619 519748
rect 173653 519714 173711 519748
rect 173745 519714 173803 519748
rect 173837 519714 173895 519748
rect 173929 519714 173987 519748
rect 174021 519714 174079 519748
rect 174113 519714 174171 519748
rect 174205 519714 174263 519748
rect 174297 519714 174355 519748
rect 174389 519714 174447 519748
rect 174481 519714 174539 519748
rect 174573 519714 174631 519748
rect 174665 519714 174723 519748
rect 174757 519714 174815 519748
rect 174849 519714 174907 519748
rect 174941 519714 174999 519748
rect 175033 519714 175091 519748
rect 175125 519714 175183 519748
rect 175217 519714 175275 519748
rect 175309 519714 175367 519748
rect 175401 519714 175459 519748
rect 175493 519714 175551 519748
rect 175585 519714 175643 519748
rect 175677 519714 175735 519748
rect 175769 519714 175827 519748
rect 175861 519714 175919 519748
rect 175953 519714 176011 519748
rect 176045 519714 176103 519748
rect 176137 519714 176195 519748
rect 176229 519714 176287 519748
rect 176321 519714 176379 519748
rect 176413 519714 176471 519748
rect 176505 519714 176563 519748
rect 176597 519714 176655 519748
rect 176689 519714 176747 519748
rect 176781 519714 176839 519748
rect 176873 519714 176931 519748
rect 176965 519714 177023 519748
rect 177057 519714 177115 519748
rect 177149 519714 177207 519748
rect 177241 519714 177299 519748
rect 177333 519714 177391 519748
rect 177425 519714 177483 519748
rect 177517 519714 177575 519748
rect 177609 519714 177667 519748
rect 177701 519714 177759 519748
rect 177793 519714 177851 519748
rect 177885 519714 177943 519748
rect 177977 519714 178035 519748
rect 178069 519714 178127 519748
rect 178161 519714 178219 519748
rect 178253 519714 178311 519748
rect 178345 519714 178403 519748
rect 178437 519714 178495 519748
rect 178529 519714 178587 519748
rect 178621 519714 178679 519748
rect 178713 519714 178771 519748
rect 178805 519714 178863 519748
rect 178897 519714 178955 519748
rect 178989 519714 179047 519748
rect 179081 519714 179139 519748
rect 179173 519714 179231 519748
rect 179265 519714 179323 519748
rect 179357 519714 179415 519748
rect 179449 519714 179507 519748
rect 179541 519714 179599 519748
rect 179633 519714 179691 519748
rect 179725 519714 179783 519748
rect 179817 519714 179875 519748
rect 179909 519714 179967 519748
rect 180001 519714 180059 519748
rect 180093 519714 180151 519748
rect 180185 519714 180243 519748
rect 180277 519714 180335 519748
rect 180369 519714 180427 519748
rect 180461 519714 180519 519748
rect 180553 519714 180611 519748
rect 180645 519714 180703 519748
rect 180737 519714 180795 519748
rect 180829 519714 180887 519748
rect 180921 519714 180979 519748
rect 181013 519714 181071 519748
rect 181105 519714 181163 519748
rect 181197 519714 181255 519748
rect 181289 519714 181347 519748
rect 181381 519714 181439 519748
rect 181473 519714 181531 519748
rect 181565 519714 181623 519748
rect 181657 519714 181715 519748
rect 181749 519714 181807 519748
rect 181841 519714 181899 519748
rect 181933 519714 181991 519748
rect 182025 519714 182083 519748
rect 182117 519714 182175 519748
rect 182209 519714 182267 519748
rect 182301 519714 182359 519748
rect 182393 519714 182451 519748
rect 182485 519714 182543 519748
rect 182577 519714 182635 519748
rect 182669 519714 182727 519748
rect 182761 519714 182819 519748
rect 182853 519714 182911 519748
rect 182945 519714 183003 519748
rect 183037 519714 183095 519748
rect 183129 519714 183187 519748
rect 183221 519714 183279 519748
rect 183313 519714 183371 519748
rect 183405 519714 183463 519748
rect 183497 519714 183555 519748
rect 183589 519714 183647 519748
rect 183681 519714 183739 519748
rect 183773 519714 183831 519748
rect 183865 519714 183923 519748
rect 183957 519714 184015 519748
rect 184049 519714 184107 519748
rect 184141 519714 184199 519748
rect 184233 519714 184291 519748
rect 184325 519714 184383 519748
rect 184417 519714 184475 519748
rect 184509 519714 184567 519748
rect 184601 519714 184659 519748
rect 184693 519714 184751 519748
rect 184785 519714 184843 519748
rect 184877 519714 184935 519748
rect 184969 519714 185027 519748
rect 185061 519714 185119 519748
rect 185153 519714 185211 519748
rect 185245 519714 185303 519748
rect 185337 519714 185395 519748
rect 185429 519714 185487 519748
rect 185521 519714 185579 519748
rect 185613 519714 185671 519748
rect 185705 519714 185763 519748
rect 185797 519714 185855 519748
rect 185889 519714 185947 519748
rect 185981 519714 186039 519748
rect 186073 519714 186131 519748
rect 186165 519714 186223 519748
rect 186257 519714 186315 519748
rect 186349 519714 186407 519748
rect 186441 519714 186499 519748
rect 186533 519714 186591 519748
rect 186625 519714 186683 519748
rect 186717 519714 186775 519748
rect 186809 519714 186867 519748
rect 186901 519714 186959 519748
rect 186993 519714 187051 519748
rect 187085 519714 187143 519748
rect 187177 519714 187235 519748
rect 187269 519714 187327 519748
rect 187361 519714 187419 519748
rect 187453 519714 187482 519748
rect 172227 519651 172469 519714
rect 172227 519617 172245 519651
rect 172279 519617 172417 519651
rect 172451 519617 172469 519651
rect 172227 519564 172469 519617
rect 172503 519653 173572 519714
rect 172503 519619 172521 519653
rect 172555 519619 173521 519653
rect 173555 519619 173572 519653
rect 172503 519605 173572 519619
rect 173607 519653 174676 519714
rect 173607 519619 173625 519653
rect 173659 519619 174625 519653
rect 174659 519619 174676 519653
rect 173607 519605 174676 519619
rect 174803 519620 174861 519714
rect 172227 519490 172331 519564
rect 172227 519456 172277 519490
rect 172311 519456 172331 519490
rect 172365 519496 172385 519530
rect 172419 519496 172469 519530
rect 172365 519422 172469 519496
rect 172820 519490 172888 519605
rect 172820 519456 172837 519490
rect 172871 519456 172888 519490
rect 172820 519439 172888 519456
rect 173184 519526 173254 519541
rect 173184 519492 173201 519526
rect 173235 519492 173254 519526
rect 172227 519375 172469 519422
rect 172227 519341 172245 519375
rect 172279 519341 172417 519375
rect 172451 519341 172469 519375
rect 172227 519280 172469 519341
rect 173184 519291 173254 519492
rect 173924 519490 173992 519605
rect 174803 519586 174815 519620
rect 174849 519586 174861 519620
rect 174895 519653 175964 519714
rect 174895 519619 174913 519653
rect 174947 519619 175913 519653
rect 175947 519619 175964 519653
rect 174895 519605 175964 519619
rect 175999 519653 177068 519714
rect 175999 519619 176017 519653
rect 176051 519619 177017 519653
rect 177051 519619 177068 519653
rect 175999 519605 177068 519619
rect 177103 519653 178172 519714
rect 177103 519619 177121 519653
rect 177155 519619 178121 519653
rect 178155 519619 178172 519653
rect 177103 519605 178172 519619
rect 178207 519653 179276 519714
rect 178207 519619 178225 519653
rect 178259 519619 179225 519653
rect 179259 519619 179276 519653
rect 178207 519605 179276 519619
rect 179311 519653 179829 519714
rect 179311 519619 179329 519653
rect 179363 519619 179777 519653
rect 179811 519619 179829 519653
rect 174803 519569 174861 519586
rect 173924 519456 173941 519490
rect 173975 519456 173992 519490
rect 173924 519439 173992 519456
rect 174288 519526 174358 519541
rect 174288 519492 174305 519526
rect 174339 519492 174358 519526
rect 174288 519291 174358 519492
rect 175212 519490 175280 519605
rect 175212 519456 175229 519490
rect 175263 519456 175280 519490
rect 175212 519439 175280 519456
rect 175576 519526 175646 519541
rect 175576 519492 175593 519526
rect 175627 519492 175646 519526
rect 174803 519402 174861 519437
rect 174803 519368 174815 519402
rect 174849 519368 174861 519402
rect 174803 519309 174861 519368
rect 172227 519246 172245 519280
rect 172279 519246 172417 519280
rect 172451 519246 172469 519280
rect 172227 519204 172469 519246
rect 172503 519280 173572 519291
rect 172503 519246 172521 519280
rect 172555 519246 173521 519280
rect 173555 519246 173572 519280
rect 172503 519204 173572 519246
rect 173607 519280 174676 519291
rect 173607 519246 173625 519280
rect 173659 519246 174625 519280
rect 174659 519246 174676 519280
rect 173607 519204 174676 519246
rect 174803 519275 174815 519309
rect 174849 519275 174861 519309
rect 175576 519291 175646 519492
rect 176316 519490 176384 519605
rect 176316 519456 176333 519490
rect 176367 519456 176384 519490
rect 176316 519439 176384 519456
rect 176680 519526 176750 519541
rect 176680 519492 176697 519526
rect 176731 519492 176750 519526
rect 176680 519291 176750 519492
rect 177420 519490 177488 519605
rect 177420 519456 177437 519490
rect 177471 519456 177488 519490
rect 177420 519439 177488 519456
rect 177784 519526 177854 519541
rect 177784 519492 177801 519526
rect 177835 519492 177854 519526
rect 177784 519291 177854 519492
rect 178524 519490 178592 519605
rect 179311 519560 179829 519619
rect 179955 519620 180013 519714
rect 179955 519586 179967 519620
rect 180001 519586 180013 519620
rect 180047 519653 181116 519714
rect 180047 519619 180065 519653
rect 180099 519619 181065 519653
rect 181099 519619 181116 519653
rect 180047 519605 181116 519619
rect 181151 519653 182220 519714
rect 181151 519619 181169 519653
rect 181203 519619 182169 519653
rect 182203 519619 182220 519653
rect 181151 519605 182220 519619
rect 182255 519653 183324 519714
rect 182255 519619 182273 519653
rect 182307 519619 183273 519653
rect 183307 519619 183324 519653
rect 182255 519605 183324 519619
rect 183359 519653 184428 519714
rect 183359 519619 183377 519653
rect 183411 519619 184377 519653
rect 184411 519619 184428 519653
rect 183359 519605 184428 519619
rect 184463 519653 184981 519714
rect 184463 519619 184481 519653
rect 184515 519619 184929 519653
rect 184963 519619 184981 519653
rect 179955 519569 180013 519586
rect 178524 519456 178541 519490
rect 178575 519456 178592 519490
rect 178524 519439 178592 519456
rect 178888 519526 178958 519541
rect 178888 519492 178905 519526
rect 178939 519492 178958 519526
rect 178888 519291 178958 519492
rect 179311 519490 179553 519560
rect 179311 519456 179389 519490
rect 179423 519456 179499 519490
rect 179533 519456 179553 519490
rect 179587 519492 179607 519526
rect 179641 519492 179717 519526
rect 179751 519492 179829 519526
rect 179587 519422 179829 519492
rect 180364 519490 180432 519605
rect 180364 519456 180381 519490
rect 180415 519456 180432 519490
rect 180364 519439 180432 519456
rect 180728 519526 180798 519541
rect 180728 519492 180745 519526
rect 180779 519492 180798 519526
rect 179311 519382 179829 519422
rect 179311 519348 179329 519382
rect 179363 519348 179777 519382
rect 179811 519348 179829 519382
rect 174803 519204 174861 519275
rect 174895 519280 175964 519291
rect 174895 519246 174913 519280
rect 174947 519246 175913 519280
rect 175947 519246 175964 519280
rect 174895 519204 175964 519246
rect 175999 519280 177068 519291
rect 175999 519246 176017 519280
rect 176051 519246 177017 519280
rect 177051 519246 177068 519280
rect 175999 519204 177068 519246
rect 177103 519280 178172 519291
rect 177103 519246 177121 519280
rect 177155 519246 178121 519280
rect 178155 519246 178172 519280
rect 177103 519204 178172 519246
rect 178207 519280 179276 519291
rect 178207 519246 178225 519280
rect 178259 519246 179225 519280
rect 179259 519246 179276 519280
rect 178207 519204 179276 519246
rect 179311 519280 179829 519348
rect 179311 519246 179329 519280
rect 179363 519246 179777 519280
rect 179811 519246 179829 519280
rect 179311 519204 179829 519246
rect 179955 519402 180013 519437
rect 179955 519368 179967 519402
rect 180001 519368 180013 519402
rect 179955 519309 180013 519368
rect 179955 519275 179967 519309
rect 180001 519275 180013 519309
rect 180728 519291 180798 519492
rect 181468 519490 181536 519605
rect 181468 519456 181485 519490
rect 181519 519456 181536 519490
rect 181468 519439 181536 519456
rect 181832 519526 181902 519541
rect 181832 519492 181849 519526
rect 181883 519492 181902 519526
rect 181832 519291 181902 519492
rect 182572 519490 182640 519605
rect 182572 519456 182589 519490
rect 182623 519456 182640 519490
rect 182572 519439 182640 519456
rect 182936 519526 183006 519541
rect 182936 519492 182953 519526
rect 182987 519492 183006 519526
rect 182936 519291 183006 519492
rect 183676 519490 183744 519605
rect 184463 519560 184981 519619
rect 185107 519620 185165 519714
rect 185107 519586 185119 519620
rect 185153 519586 185165 519620
rect 185199 519653 186268 519714
rect 185199 519619 185217 519653
rect 185251 519619 186217 519653
rect 186251 519619 186268 519653
rect 185199 519605 186268 519619
rect 186303 519653 187005 519714
rect 186303 519619 186321 519653
rect 186355 519619 186953 519653
rect 186987 519619 187005 519653
rect 185107 519569 185165 519586
rect 183676 519456 183693 519490
rect 183727 519456 183744 519490
rect 183676 519439 183744 519456
rect 184040 519526 184110 519541
rect 184040 519492 184057 519526
rect 184091 519492 184110 519526
rect 184040 519291 184110 519492
rect 184463 519490 184705 519560
rect 184463 519456 184541 519490
rect 184575 519456 184651 519490
rect 184685 519456 184705 519490
rect 184739 519492 184759 519526
rect 184793 519492 184869 519526
rect 184903 519492 184981 519526
rect 184739 519422 184981 519492
rect 185516 519490 185584 519605
rect 186303 519560 187005 519619
rect 187223 519651 187465 519714
rect 187223 519617 187241 519651
rect 187275 519617 187413 519651
rect 187447 519617 187465 519651
rect 187223 519564 187465 519617
rect 185516 519456 185533 519490
rect 185567 519456 185584 519490
rect 185516 519439 185584 519456
rect 185880 519526 185950 519541
rect 185880 519492 185897 519526
rect 185931 519492 185950 519526
rect 184463 519382 184981 519422
rect 184463 519348 184481 519382
rect 184515 519348 184929 519382
rect 184963 519348 184981 519382
rect 179955 519204 180013 519275
rect 180047 519280 181116 519291
rect 180047 519246 180065 519280
rect 180099 519246 181065 519280
rect 181099 519246 181116 519280
rect 180047 519204 181116 519246
rect 181151 519280 182220 519291
rect 181151 519246 181169 519280
rect 181203 519246 182169 519280
rect 182203 519246 182220 519280
rect 181151 519204 182220 519246
rect 182255 519280 183324 519291
rect 182255 519246 182273 519280
rect 182307 519246 183273 519280
rect 183307 519246 183324 519280
rect 182255 519204 183324 519246
rect 183359 519280 184428 519291
rect 183359 519246 183377 519280
rect 183411 519246 184377 519280
rect 184411 519246 184428 519280
rect 183359 519204 184428 519246
rect 184463 519280 184981 519348
rect 184463 519246 184481 519280
rect 184515 519246 184929 519280
rect 184963 519246 184981 519280
rect 184463 519204 184981 519246
rect 185107 519402 185165 519437
rect 185107 519368 185119 519402
rect 185153 519368 185165 519402
rect 185107 519309 185165 519368
rect 185107 519275 185119 519309
rect 185153 519275 185165 519309
rect 185880 519291 185950 519492
rect 186303 519490 186633 519560
rect 186303 519456 186381 519490
rect 186415 519456 186480 519490
rect 186514 519456 186579 519490
rect 186613 519456 186633 519490
rect 186667 519492 186687 519526
rect 186721 519492 186790 519526
rect 186824 519492 186893 519526
rect 186927 519492 187005 519526
rect 186667 519422 187005 519492
rect 186303 519382 187005 519422
rect 186303 519348 186321 519382
rect 186355 519348 186953 519382
rect 186987 519348 187005 519382
rect 185107 519204 185165 519275
rect 185199 519280 186268 519291
rect 185199 519246 185217 519280
rect 185251 519246 186217 519280
rect 186251 519246 186268 519280
rect 185199 519204 186268 519246
rect 186303 519280 187005 519348
rect 186303 519246 186321 519280
rect 186355 519246 186953 519280
rect 186987 519246 187005 519280
rect 186303 519204 187005 519246
rect 187223 519496 187273 519530
rect 187307 519496 187327 519530
rect 187223 519422 187327 519496
rect 187361 519490 187465 519564
rect 187361 519456 187381 519490
rect 187415 519456 187465 519490
rect 187223 519375 187465 519422
rect 187223 519341 187241 519375
rect 187275 519341 187413 519375
rect 187447 519341 187465 519375
rect 187223 519280 187465 519341
rect 187223 519246 187241 519280
rect 187275 519246 187413 519280
rect 187447 519246 187465 519280
rect 187223 519204 187465 519246
rect 172210 519170 172239 519204
rect 172273 519170 172331 519204
rect 172365 519170 172423 519204
rect 172457 519170 172515 519204
rect 172549 519170 172607 519204
rect 172641 519170 172699 519204
rect 172733 519170 172791 519204
rect 172825 519170 172883 519204
rect 172917 519170 172975 519204
rect 173009 519170 173067 519204
rect 173101 519170 173159 519204
rect 173193 519170 173251 519204
rect 173285 519170 173343 519204
rect 173377 519170 173435 519204
rect 173469 519170 173527 519204
rect 173561 519170 173619 519204
rect 173653 519170 173711 519204
rect 173745 519170 173803 519204
rect 173837 519170 173895 519204
rect 173929 519170 173987 519204
rect 174021 519170 174079 519204
rect 174113 519170 174171 519204
rect 174205 519170 174263 519204
rect 174297 519170 174355 519204
rect 174389 519170 174447 519204
rect 174481 519170 174539 519204
rect 174573 519170 174631 519204
rect 174665 519170 174723 519204
rect 174757 519170 174815 519204
rect 174849 519170 174907 519204
rect 174941 519170 174999 519204
rect 175033 519170 175091 519204
rect 175125 519170 175183 519204
rect 175217 519170 175275 519204
rect 175309 519170 175367 519204
rect 175401 519170 175459 519204
rect 175493 519170 175551 519204
rect 175585 519170 175643 519204
rect 175677 519170 175735 519204
rect 175769 519170 175827 519204
rect 175861 519170 175919 519204
rect 175953 519170 176011 519204
rect 176045 519170 176103 519204
rect 176137 519170 176195 519204
rect 176229 519170 176287 519204
rect 176321 519170 176379 519204
rect 176413 519170 176471 519204
rect 176505 519170 176563 519204
rect 176597 519170 176655 519204
rect 176689 519170 176747 519204
rect 176781 519170 176839 519204
rect 176873 519170 176931 519204
rect 176965 519170 177023 519204
rect 177057 519170 177115 519204
rect 177149 519170 177207 519204
rect 177241 519170 177299 519204
rect 177333 519170 177391 519204
rect 177425 519170 177483 519204
rect 177517 519170 177575 519204
rect 177609 519170 177667 519204
rect 177701 519170 177759 519204
rect 177793 519170 177851 519204
rect 177885 519170 177943 519204
rect 177977 519170 178035 519204
rect 178069 519170 178127 519204
rect 178161 519170 178219 519204
rect 178253 519170 178311 519204
rect 178345 519170 178403 519204
rect 178437 519170 178495 519204
rect 178529 519170 178587 519204
rect 178621 519170 178679 519204
rect 178713 519170 178771 519204
rect 178805 519170 178863 519204
rect 178897 519170 178955 519204
rect 178989 519170 179047 519204
rect 179081 519170 179139 519204
rect 179173 519170 179231 519204
rect 179265 519170 179323 519204
rect 179357 519170 179415 519204
rect 179449 519170 179507 519204
rect 179541 519170 179599 519204
rect 179633 519170 179691 519204
rect 179725 519170 179783 519204
rect 179817 519170 179875 519204
rect 179909 519170 179967 519204
rect 180001 519170 180059 519204
rect 180093 519170 180151 519204
rect 180185 519170 180243 519204
rect 180277 519170 180335 519204
rect 180369 519170 180427 519204
rect 180461 519170 180519 519204
rect 180553 519170 180611 519204
rect 180645 519170 180703 519204
rect 180737 519170 180795 519204
rect 180829 519170 180887 519204
rect 180921 519170 180979 519204
rect 181013 519170 181071 519204
rect 181105 519170 181163 519204
rect 181197 519170 181255 519204
rect 181289 519170 181347 519204
rect 181381 519170 181439 519204
rect 181473 519170 181531 519204
rect 181565 519170 181623 519204
rect 181657 519170 181715 519204
rect 181749 519170 181807 519204
rect 181841 519170 181899 519204
rect 181933 519170 181991 519204
rect 182025 519170 182083 519204
rect 182117 519170 182175 519204
rect 182209 519170 182267 519204
rect 182301 519170 182359 519204
rect 182393 519170 182451 519204
rect 182485 519170 182543 519204
rect 182577 519170 182635 519204
rect 182669 519170 182727 519204
rect 182761 519170 182819 519204
rect 182853 519170 182911 519204
rect 182945 519170 183003 519204
rect 183037 519170 183095 519204
rect 183129 519170 183187 519204
rect 183221 519170 183279 519204
rect 183313 519170 183371 519204
rect 183405 519170 183463 519204
rect 183497 519170 183555 519204
rect 183589 519170 183647 519204
rect 183681 519170 183739 519204
rect 183773 519170 183831 519204
rect 183865 519170 183923 519204
rect 183957 519170 184015 519204
rect 184049 519170 184107 519204
rect 184141 519170 184199 519204
rect 184233 519170 184291 519204
rect 184325 519170 184383 519204
rect 184417 519170 184475 519204
rect 184509 519170 184567 519204
rect 184601 519170 184659 519204
rect 184693 519170 184751 519204
rect 184785 519170 184843 519204
rect 184877 519170 184935 519204
rect 184969 519170 185027 519204
rect 185061 519170 185119 519204
rect 185153 519170 185211 519204
rect 185245 519170 185303 519204
rect 185337 519170 185395 519204
rect 185429 519170 185487 519204
rect 185521 519170 185579 519204
rect 185613 519170 185671 519204
rect 185705 519170 185763 519204
rect 185797 519170 185855 519204
rect 185889 519170 185947 519204
rect 185981 519170 186039 519204
rect 186073 519170 186131 519204
rect 186165 519170 186223 519204
rect 186257 519170 186315 519204
rect 186349 519170 186407 519204
rect 186441 519170 186499 519204
rect 186533 519170 186591 519204
rect 186625 519170 186683 519204
rect 186717 519170 186775 519204
rect 186809 519170 186867 519204
rect 186901 519170 186959 519204
rect 186993 519170 187051 519204
rect 187085 519170 187143 519204
rect 187177 519170 187235 519204
rect 187269 519170 187327 519204
rect 187361 519170 187419 519204
rect 187453 519170 187482 519204
rect 172227 519128 172469 519170
rect 172227 519094 172245 519128
rect 172279 519094 172417 519128
rect 172451 519094 172469 519128
rect 172227 519033 172469 519094
rect 172503 519128 173572 519170
rect 172503 519094 172521 519128
rect 172555 519094 173521 519128
rect 173555 519094 173572 519128
rect 172503 519083 173572 519094
rect 173607 519128 174676 519170
rect 173607 519094 173625 519128
rect 173659 519094 174625 519128
rect 174659 519094 174676 519128
rect 173607 519083 174676 519094
rect 174711 519128 175780 519170
rect 174711 519094 174729 519128
rect 174763 519094 175729 519128
rect 175763 519094 175780 519128
rect 174711 519083 175780 519094
rect 175815 519128 176884 519170
rect 175815 519094 175833 519128
rect 175867 519094 176833 519128
rect 176867 519094 176884 519128
rect 175815 519083 176884 519094
rect 176919 519128 177253 519170
rect 176919 519094 176937 519128
rect 176971 519094 177201 519128
rect 177235 519094 177253 519128
rect 172227 518999 172245 519033
rect 172279 518999 172417 519033
rect 172451 518999 172469 519033
rect 172227 518952 172469 518999
rect 172227 518884 172277 518918
rect 172311 518884 172331 518918
rect 172227 518810 172331 518884
rect 172365 518878 172469 518952
rect 172365 518844 172385 518878
rect 172419 518844 172469 518878
rect 172820 518918 172888 518935
rect 172820 518884 172837 518918
rect 172871 518884 172888 518918
rect 172227 518757 172469 518810
rect 172820 518769 172888 518884
rect 173184 518882 173254 519083
rect 173184 518848 173201 518882
rect 173235 518848 173254 518882
rect 173184 518833 173254 518848
rect 173924 518918 173992 518935
rect 173924 518884 173941 518918
rect 173975 518884 173992 518918
rect 173924 518769 173992 518884
rect 174288 518882 174358 519083
rect 174288 518848 174305 518882
rect 174339 518848 174358 518882
rect 174288 518833 174358 518848
rect 175028 518918 175096 518935
rect 175028 518884 175045 518918
rect 175079 518884 175096 518918
rect 175028 518769 175096 518884
rect 175392 518882 175462 519083
rect 175392 518848 175409 518882
rect 175443 518848 175462 518882
rect 175392 518833 175462 518848
rect 176132 518918 176200 518935
rect 176132 518884 176149 518918
rect 176183 518884 176200 518918
rect 176132 518769 176200 518884
rect 176496 518882 176566 519083
rect 176919 519026 177253 519094
rect 176919 518992 176937 519026
rect 176971 518992 177201 519026
rect 177235 518992 177253 519026
rect 176919 518952 177253 518992
rect 176496 518848 176513 518882
rect 176547 518848 176566 518882
rect 176496 518833 176566 518848
rect 176919 518884 176939 518918
rect 176973 518884 177069 518918
rect 176919 518814 177069 518884
rect 177103 518882 177253 518952
rect 177379 519099 177437 519170
rect 177379 519065 177391 519099
rect 177425 519065 177437 519099
rect 177471 519128 178540 519170
rect 177471 519094 177489 519128
rect 177523 519094 178489 519128
rect 178523 519094 178540 519128
rect 177471 519083 178540 519094
rect 178575 519128 179644 519170
rect 178575 519094 178593 519128
rect 178627 519094 179593 519128
rect 179627 519094 179644 519128
rect 178575 519083 179644 519094
rect 179679 519128 180748 519170
rect 179679 519094 179697 519128
rect 179731 519094 180697 519128
rect 180731 519094 180748 519128
rect 179679 519083 180748 519094
rect 180783 519128 181852 519170
rect 180783 519094 180801 519128
rect 180835 519094 181801 519128
rect 181835 519094 181852 519128
rect 180783 519083 181852 519094
rect 181887 519128 182405 519170
rect 181887 519094 181905 519128
rect 181939 519094 182353 519128
rect 182387 519094 182405 519128
rect 177379 519006 177437 519065
rect 177379 518972 177391 519006
rect 177425 518972 177437 519006
rect 177379 518937 177437 518972
rect 177103 518848 177199 518882
rect 177233 518848 177253 518882
rect 177788 518918 177856 518935
rect 177788 518884 177805 518918
rect 177839 518884 177856 518918
rect 172227 518723 172245 518757
rect 172279 518723 172417 518757
rect 172451 518723 172469 518757
rect 172227 518660 172469 518723
rect 172503 518755 173572 518769
rect 172503 518721 172521 518755
rect 172555 518721 173521 518755
rect 173555 518721 173572 518755
rect 172503 518660 173572 518721
rect 173607 518755 174676 518769
rect 173607 518721 173625 518755
rect 173659 518721 174625 518755
rect 174659 518721 174676 518755
rect 173607 518660 174676 518721
rect 174711 518755 175780 518769
rect 174711 518721 174729 518755
rect 174763 518721 175729 518755
rect 175763 518721 175780 518755
rect 174711 518660 175780 518721
rect 175815 518755 176884 518769
rect 175815 518721 175833 518755
rect 175867 518721 176833 518755
rect 176867 518721 176884 518755
rect 175815 518660 176884 518721
rect 176919 518762 177253 518814
rect 176919 518728 176937 518762
rect 176971 518728 177201 518762
rect 177235 518728 177253 518762
rect 176919 518660 177253 518728
rect 177379 518788 177437 518805
rect 177379 518754 177391 518788
rect 177425 518754 177437 518788
rect 177788 518769 177856 518884
rect 178152 518882 178222 519083
rect 178152 518848 178169 518882
rect 178203 518848 178222 518882
rect 178152 518833 178222 518848
rect 178892 518918 178960 518935
rect 178892 518884 178909 518918
rect 178943 518884 178960 518918
rect 178892 518769 178960 518884
rect 179256 518882 179326 519083
rect 179256 518848 179273 518882
rect 179307 518848 179326 518882
rect 179256 518833 179326 518848
rect 179996 518918 180064 518935
rect 179996 518884 180013 518918
rect 180047 518884 180064 518918
rect 179996 518769 180064 518884
rect 180360 518882 180430 519083
rect 180360 518848 180377 518882
rect 180411 518848 180430 518882
rect 180360 518833 180430 518848
rect 181100 518918 181168 518935
rect 181100 518884 181117 518918
rect 181151 518884 181168 518918
rect 181100 518769 181168 518884
rect 181464 518882 181534 519083
rect 181887 519026 182405 519094
rect 181887 518992 181905 519026
rect 181939 518992 182353 519026
rect 182387 518992 182405 519026
rect 181887 518952 182405 518992
rect 181464 518848 181481 518882
rect 181515 518848 181534 518882
rect 181464 518833 181534 518848
rect 181887 518884 181965 518918
rect 181999 518884 182075 518918
rect 182109 518884 182129 518918
rect 181887 518814 182129 518884
rect 182163 518882 182405 518952
rect 182531 519099 182589 519170
rect 182531 519065 182543 519099
rect 182577 519065 182589 519099
rect 182623 519128 183692 519170
rect 182623 519094 182641 519128
rect 182675 519094 183641 519128
rect 183675 519094 183692 519128
rect 182623 519083 183692 519094
rect 183727 519128 184796 519170
rect 183727 519094 183745 519128
rect 183779 519094 184745 519128
rect 184779 519094 184796 519128
rect 183727 519083 184796 519094
rect 184831 519128 185900 519170
rect 184831 519094 184849 519128
rect 184883 519094 185849 519128
rect 185883 519094 185900 519128
rect 184831 519083 185900 519094
rect 185935 519128 187004 519170
rect 185935 519094 185953 519128
rect 185987 519094 186953 519128
rect 186987 519094 187004 519128
rect 185935 519083 187004 519094
rect 187223 519128 187465 519170
rect 187223 519094 187241 519128
rect 187275 519094 187413 519128
rect 187447 519094 187465 519128
rect 182531 519006 182589 519065
rect 182531 518972 182543 519006
rect 182577 518972 182589 519006
rect 182531 518937 182589 518972
rect 182163 518848 182183 518882
rect 182217 518848 182293 518882
rect 182327 518848 182405 518882
rect 182940 518918 183008 518935
rect 182940 518884 182957 518918
rect 182991 518884 183008 518918
rect 177379 518660 177437 518754
rect 177471 518755 178540 518769
rect 177471 518721 177489 518755
rect 177523 518721 178489 518755
rect 178523 518721 178540 518755
rect 177471 518660 178540 518721
rect 178575 518755 179644 518769
rect 178575 518721 178593 518755
rect 178627 518721 179593 518755
rect 179627 518721 179644 518755
rect 178575 518660 179644 518721
rect 179679 518755 180748 518769
rect 179679 518721 179697 518755
rect 179731 518721 180697 518755
rect 180731 518721 180748 518755
rect 179679 518660 180748 518721
rect 180783 518755 181852 518769
rect 180783 518721 180801 518755
rect 180835 518721 181801 518755
rect 181835 518721 181852 518755
rect 180783 518660 181852 518721
rect 181887 518755 182405 518814
rect 181887 518721 181905 518755
rect 181939 518721 182353 518755
rect 182387 518721 182405 518755
rect 181887 518660 182405 518721
rect 182531 518788 182589 518805
rect 182531 518754 182543 518788
rect 182577 518754 182589 518788
rect 182940 518769 183008 518884
rect 183304 518882 183374 519083
rect 183304 518848 183321 518882
rect 183355 518848 183374 518882
rect 183304 518833 183374 518848
rect 184044 518918 184112 518935
rect 184044 518884 184061 518918
rect 184095 518884 184112 518918
rect 184044 518769 184112 518884
rect 184408 518882 184478 519083
rect 184408 518848 184425 518882
rect 184459 518848 184478 518882
rect 184408 518833 184478 518848
rect 185148 518918 185216 518935
rect 185148 518884 185165 518918
rect 185199 518884 185216 518918
rect 185148 518769 185216 518884
rect 185512 518882 185582 519083
rect 185512 518848 185529 518882
rect 185563 518848 185582 518882
rect 185512 518833 185582 518848
rect 186252 518918 186320 518935
rect 186252 518884 186269 518918
rect 186303 518884 186320 518918
rect 186252 518769 186320 518884
rect 186616 518882 186686 519083
rect 186616 518848 186633 518882
rect 186667 518848 186686 518882
rect 186616 518833 186686 518848
rect 187223 519033 187465 519094
rect 187223 518999 187241 519033
rect 187275 518999 187413 519033
rect 187447 518999 187465 519033
rect 187223 518952 187465 518999
rect 187223 518878 187327 518952
rect 187223 518844 187273 518878
rect 187307 518844 187327 518878
rect 187361 518884 187381 518918
rect 187415 518884 187465 518918
rect 187361 518810 187465 518884
rect 182531 518660 182589 518754
rect 182623 518755 183692 518769
rect 182623 518721 182641 518755
rect 182675 518721 183641 518755
rect 183675 518721 183692 518755
rect 182623 518660 183692 518721
rect 183727 518755 184796 518769
rect 183727 518721 183745 518755
rect 183779 518721 184745 518755
rect 184779 518721 184796 518755
rect 183727 518660 184796 518721
rect 184831 518755 185900 518769
rect 184831 518721 184849 518755
rect 184883 518721 185849 518755
rect 185883 518721 185900 518755
rect 184831 518660 185900 518721
rect 185935 518755 187004 518769
rect 185935 518721 185953 518755
rect 185987 518721 186953 518755
rect 186987 518721 187004 518755
rect 185935 518660 187004 518721
rect 187223 518757 187465 518810
rect 187223 518723 187241 518757
rect 187275 518723 187413 518757
rect 187447 518723 187465 518757
rect 187223 518660 187465 518723
rect 172210 518626 172239 518660
rect 172273 518626 172331 518660
rect 172365 518626 172423 518660
rect 172457 518626 172515 518660
rect 172549 518626 172607 518660
rect 172641 518626 172699 518660
rect 172733 518626 172791 518660
rect 172825 518626 172883 518660
rect 172917 518626 172975 518660
rect 173009 518626 173067 518660
rect 173101 518626 173159 518660
rect 173193 518626 173251 518660
rect 173285 518626 173343 518660
rect 173377 518626 173435 518660
rect 173469 518626 173527 518660
rect 173561 518626 173619 518660
rect 173653 518626 173711 518660
rect 173745 518626 173803 518660
rect 173837 518626 173895 518660
rect 173929 518626 173987 518660
rect 174021 518626 174079 518660
rect 174113 518626 174171 518660
rect 174205 518626 174263 518660
rect 174297 518626 174355 518660
rect 174389 518626 174447 518660
rect 174481 518626 174539 518660
rect 174573 518626 174631 518660
rect 174665 518626 174723 518660
rect 174757 518626 174815 518660
rect 174849 518626 174907 518660
rect 174941 518626 174999 518660
rect 175033 518626 175091 518660
rect 175125 518626 175183 518660
rect 175217 518626 175275 518660
rect 175309 518626 175367 518660
rect 175401 518626 175459 518660
rect 175493 518626 175551 518660
rect 175585 518626 175643 518660
rect 175677 518626 175735 518660
rect 175769 518626 175827 518660
rect 175861 518626 175919 518660
rect 175953 518626 176011 518660
rect 176045 518626 176103 518660
rect 176137 518626 176195 518660
rect 176229 518626 176287 518660
rect 176321 518626 176379 518660
rect 176413 518626 176471 518660
rect 176505 518626 176563 518660
rect 176597 518626 176655 518660
rect 176689 518626 176747 518660
rect 176781 518626 176839 518660
rect 176873 518626 176931 518660
rect 176965 518626 177023 518660
rect 177057 518626 177115 518660
rect 177149 518626 177207 518660
rect 177241 518626 177299 518660
rect 177333 518626 177391 518660
rect 177425 518626 177483 518660
rect 177517 518626 177575 518660
rect 177609 518626 177667 518660
rect 177701 518626 177759 518660
rect 177793 518626 177851 518660
rect 177885 518626 177943 518660
rect 177977 518626 178035 518660
rect 178069 518626 178127 518660
rect 178161 518626 178219 518660
rect 178253 518626 178311 518660
rect 178345 518626 178403 518660
rect 178437 518626 178495 518660
rect 178529 518626 178587 518660
rect 178621 518626 178679 518660
rect 178713 518626 178771 518660
rect 178805 518626 178863 518660
rect 178897 518626 178955 518660
rect 178989 518626 179047 518660
rect 179081 518626 179139 518660
rect 179173 518626 179231 518660
rect 179265 518626 179323 518660
rect 179357 518626 179415 518660
rect 179449 518626 179507 518660
rect 179541 518626 179599 518660
rect 179633 518626 179691 518660
rect 179725 518626 179783 518660
rect 179817 518626 179875 518660
rect 179909 518626 179967 518660
rect 180001 518626 180059 518660
rect 180093 518626 180151 518660
rect 180185 518626 180243 518660
rect 180277 518626 180335 518660
rect 180369 518626 180427 518660
rect 180461 518626 180519 518660
rect 180553 518626 180611 518660
rect 180645 518626 180703 518660
rect 180737 518626 180795 518660
rect 180829 518626 180887 518660
rect 180921 518626 180979 518660
rect 181013 518626 181071 518660
rect 181105 518626 181163 518660
rect 181197 518626 181255 518660
rect 181289 518626 181347 518660
rect 181381 518626 181439 518660
rect 181473 518626 181531 518660
rect 181565 518626 181623 518660
rect 181657 518626 181715 518660
rect 181749 518626 181807 518660
rect 181841 518626 181899 518660
rect 181933 518626 181991 518660
rect 182025 518626 182083 518660
rect 182117 518626 182175 518660
rect 182209 518626 182267 518660
rect 182301 518626 182359 518660
rect 182393 518626 182451 518660
rect 182485 518626 182543 518660
rect 182577 518626 182635 518660
rect 182669 518626 182727 518660
rect 182761 518626 182819 518660
rect 182853 518626 182911 518660
rect 182945 518626 183003 518660
rect 183037 518626 183095 518660
rect 183129 518626 183187 518660
rect 183221 518626 183279 518660
rect 183313 518626 183371 518660
rect 183405 518626 183463 518660
rect 183497 518626 183555 518660
rect 183589 518626 183647 518660
rect 183681 518626 183739 518660
rect 183773 518626 183831 518660
rect 183865 518626 183923 518660
rect 183957 518626 184015 518660
rect 184049 518626 184107 518660
rect 184141 518626 184199 518660
rect 184233 518626 184291 518660
rect 184325 518626 184383 518660
rect 184417 518626 184475 518660
rect 184509 518626 184567 518660
rect 184601 518626 184659 518660
rect 184693 518626 184751 518660
rect 184785 518626 184843 518660
rect 184877 518626 184935 518660
rect 184969 518626 185027 518660
rect 185061 518626 185119 518660
rect 185153 518626 185211 518660
rect 185245 518626 185303 518660
rect 185337 518626 185395 518660
rect 185429 518626 185487 518660
rect 185521 518626 185579 518660
rect 185613 518626 185671 518660
rect 185705 518626 185763 518660
rect 185797 518626 185855 518660
rect 185889 518626 185947 518660
rect 185981 518626 186039 518660
rect 186073 518626 186131 518660
rect 186165 518626 186223 518660
rect 186257 518626 186315 518660
rect 186349 518626 186407 518660
rect 186441 518626 186499 518660
rect 186533 518626 186591 518660
rect 186625 518626 186683 518660
rect 186717 518626 186775 518660
rect 186809 518626 186867 518660
rect 186901 518626 186959 518660
rect 186993 518626 187051 518660
rect 187085 518626 187143 518660
rect 187177 518626 187235 518660
rect 187269 518626 187327 518660
rect 187361 518626 187419 518660
rect 187453 518626 187482 518660
rect 172227 518563 172469 518626
rect 172227 518529 172245 518563
rect 172279 518529 172417 518563
rect 172451 518529 172469 518563
rect 172227 518476 172469 518529
rect 172503 518565 173572 518626
rect 172503 518531 172521 518565
rect 172555 518531 173521 518565
rect 173555 518531 173572 518565
rect 172503 518517 173572 518531
rect 173607 518565 174676 518626
rect 173607 518531 173625 518565
rect 173659 518531 174625 518565
rect 174659 518531 174676 518565
rect 173607 518517 174676 518531
rect 174803 518532 174861 518626
rect 172227 518402 172331 518476
rect 172227 518368 172277 518402
rect 172311 518368 172331 518402
rect 172365 518408 172385 518442
rect 172419 518408 172469 518442
rect 172365 518334 172469 518408
rect 172820 518402 172888 518517
rect 172820 518368 172837 518402
rect 172871 518368 172888 518402
rect 172820 518351 172888 518368
rect 173184 518438 173254 518453
rect 173184 518404 173201 518438
rect 173235 518404 173254 518438
rect 172227 518287 172469 518334
rect 172227 518253 172245 518287
rect 172279 518253 172417 518287
rect 172451 518253 172469 518287
rect 172227 518192 172469 518253
rect 173184 518203 173254 518404
rect 173924 518402 173992 518517
rect 174803 518498 174815 518532
rect 174849 518498 174861 518532
rect 174895 518565 175964 518626
rect 174895 518531 174913 518565
rect 174947 518531 175913 518565
rect 175947 518531 175964 518565
rect 174895 518517 175964 518531
rect 175999 518565 177068 518626
rect 175999 518531 176017 518565
rect 176051 518531 177017 518565
rect 177051 518531 177068 518565
rect 175999 518517 177068 518531
rect 177103 518565 178172 518626
rect 177103 518531 177121 518565
rect 177155 518531 178121 518565
rect 178155 518531 178172 518565
rect 177103 518517 178172 518531
rect 178207 518565 179276 518626
rect 178207 518531 178225 518565
rect 178259 518531 179225 518565
rect 179259 518531 179276 518565
rect 178207 518517 179276 518531
rect 179311 518565 179829 518626
rect 179311 518531 179329 518565
rect 179363 518531 179777 518565
rect 179811 518531 179829 518565
rect 174803 518481 174861 518498
rect 173924 518368 173941 518402
rect 173975 518368 173992 518402
rect 173924 518351 173992 518368
rect 174288 518438 174358 518453
rect 174288 518404 174305 518438
rect 174339 518404 174358 518438
rect 174288 518203 174358 518404
rect 175212 518402 175280 518517
rect 175212 518368 175229 518402
rect 175263 518368 175280 518402
rect 175212 518351 175280 518368
rect 175576 518438 175646 518453
rect 175576 518404 175593 518438
rect 175627 518404 175646 518438
rect 174803 518314 174861 518349
rect 174803 518280 174815 518314
rect 174849 518280 174861 518314
rect 174803 518221 174861 518280
rect 172227 518158 172245 518192
rect 172279 518158 172417 518192
rect 172451 518158 172469 518192
rect 172227 518116 172469 518158
rect 172503 518192 173572 518203
rect 172503 518158 172521 518192
rect 172555 518158 173521 518192
rect 173555 518158 173572 518192
rect 172503 518116 173572 518158
rect 173607 518192 174676 518203
rect 173607 518158 173625 518192
rect 173659 518158 174625 518192
rect 174659 518158 174676 518192
rect 173607 518116 174676 518158
rect 174803 518187 174815 518221
rect 174849 518187 174861 518221
rect 175576 518203 175646 518404
rect 176316 518402 176384 518517
rect 176316 518368 176333 518402
rect 176367 518368 176384 518402
rect 176316 518351 176384 518368
rect 176680 518438 176750 518453
rect 176680 518404 176697 518438
rect 176731 518404 176750 518438
rect 176680 518203 176750 518404
rect 177420 518402 177488 518517
rect 177420 518368 177437 518402
rect 177471 518368 177488 518402
rect 177420 518351 177488 518368
rect 177784 518438 177854 518453
rect 177784 518404 177801 518438
rect 177835 518404 177854 518438
rect 177784 518203 177854 518404
rect 178524 518402 178592 518517
rect 179311 518472 179829 518531
rect 179955 518532 180013 518626
rect 179955 518498 179967 518532
rect 180001 518498 180013 518532
rect 180047 518565 181116 518626
rect 180047 518531 180065 518565
rect 180099 518531 181065 518565
rect 181099 518531 181116 518565
rect 180047 518517 181116 518531
rect 181151 518565 182220 518626
rect 181151 518531 181169 518565
rect 181203 518531 182169 518565
rect 182203 518531 182220 518565
rect 181151 518517 182220 518531
rect 182255 518565 183324 518626
rect 182255 518531 182273 518565
rect 182307 518531 183273 518565
rect 183307 518531 183324 518565
rect 182255 518517 183324 518531
rect 183359 518565 184428 518626
rect 183359 518531 183377 518565
rect 183411 518531 184377 518565
rect 184411 518531 184428 518565
rect 183359 518517 184428 518531
rect 184463 518565 184981 518626
rect 184463 518531 184481 518565
rect 184515 518531 184929 518565
rect 184963 518531 184981 518565
rect 179955 518481 180013 518498
rect 178524 518368 178541 518402
rect 178575 518368 178592 518402
rect 178524 518351 178592 518368
rect 178888 518438 178958 518453
rect 178888 518404 178905 518438
rect 178939 518404 178958 518438
rect 178888 518203 178958 518404
rect 179311 518402 179553 518472
rect 179311 518368 179389 518402
rect 179423 518368 179499 518402
rect 179533 518368 179553 518402
rect 179587 518404 179607 518438
rect 179641 518404 179717 518438
rect 179751 518404 179829 518438
rect 179587 518334 179829 518404
rect 180364 518402 180432 518517
rect 180364 518368 180381 518402
rect 180415 518368 180432 518402
rect 180364 518351 180432 518368
rect 180728 518438 180798 518453
rect 180728 518404 180745 518438
rect 180779 518404 180798 518438
rect 179311 518294 179829 518334
rect 179311 518260 179329 518294
rect 179363 518260 179777 518294
rect 179811 518260 179829 518294
rect 174803 518116 174861 518187
rect 174895 518192 175964 518203
rect 174895 518158 174913 518192
rect 174947 518158 175913 518192
rect 175947 518158 175964 518192
rect 174895 518116 175964 518158
rect 175999 518192 177068 518203
rect 175999 518158 176017 518192
rect 176051 518158 177017 518192
rect 177051 518158 177068 518192
rect 175999 518116 177068 518158
rect 177103 518192 178172 518203
rect 177103 518158 177121 518192
rect 177155 518158 178121 518192
rect 178155 518158 178172 518192
rect 177103 518116 178172 518158
rect 178207 518192 179276 518203
rect 178207 518158 178225 518192
rect 178259 518158 179225 518192
rect 179259 518158 179276 518192
rect 178207 518116 179276 518158
rect 179311 518192 179829 518260
rect 179311 518158 179329 518192
rect 179363 518158 179777 518192
rect 179811 518158 179829 518192
rect 179311 518116 179829 518158
rect 179955 518314 180013 518349
rect 179955 518280 179967 518314
rect 180001 518280 180013 518314
rect 179955 518221 180013 518280
rect 179955 518187 179967 518221
rect 180001 518187 180013 518221
rect 180728 518203 180798 518404
rect 181468 518402 181536 518517
rect 181468 518368 181485 518402
rect 181519 518368 181536 518402
rect 181468 518351 181536 518368
rect 181832 518438 181902 518453
rect 181832 518404 181849 518438
rect 181883 518404 181902 518438
rect 181832 518203 181902 518404
rect 182572 518402 182640 518517
rect 182572 518368 182589 518402
rect 182623 518368 182640 518402
rect 182572 518351 182640 518368
rect 182936 518438 183006 518453
rect 182936 518404 182953 518438
rect 182987 518404 183006 518438
rect 182936 518203 183006 518404
rect 183676 518402 183744 518517
rect 184463 518472 184981 518531
rect 185107 518532 185165 518626
rect 185107 518498 185119 518532
rect 185153 518498 185165 518532
rect 185199 518565 186268 518626
rect 185199 518531 185217 518565
rect 185251 518531 186217 518565
rect 186251 518531 186268 518565
rect 185199 518517 186268 518531
rect 186303 518565 187005 518626
rect 186303 518531 186321 518565
rect 186355 518531 186953 518565
rect 186987 518531 187005 518565
rect 185107 518481 185165 518498
rect 183676 518368 183693 518402
rect 183727 518368 183744 518402
rect 183676 518351 183744 518368
rect 184040 518438 184110 518453
rect 184040 518404 184057 518438
rect 184091 518404 184110 518438
rect 184040 518203 184110 518404
rect 184463 518402 184705 518472
rect 184463 518368 184541 518402
rect 184575 518368 184651 518402
rect 184685 518368 184705 518402
rect 184739 518404 184759 518438
rect 184793 518404 184869 518438
rect 184903 518404 184981 518438
rect 184739 518334 184981 518404
rect 185516 518402 185584 518517
rect 186303 518472 187005 518531
rect 187223 518563 187465 518626
rect 187223 518529 187241 518563
rect 187275 518529 187413 518563
rect 187447 518529 187465 518563
rect 187223 518476 187465 518529
rect 185516 518368 185533 518402
rect 185567 518368 185584 518402
rect 185516 518351 185584 518368
rect 185880 518438 185950 518453
rect 185880 518404 185897 518438
rect 185931 518404 185950 518438
rect 184463 518294 184981 518334
rect 184463 518260 184481 518294
rect 184515 518260 184929 518294
rect 184963 518260 184981 518294
rect 179955 518116 180013 518187
rect 180047 518192 181116 518203
rect 180047 518158 180065 518192
rect 180099 518158 181065 518192
rect 181099 518158 181116 518192
rect 180047 518116 181116 518158
rect 181151 518192 182220 518203
rect 181151 518158 181169 518192
rect 181203 518158 182169 518192
rect 182203 518158 182220 518192
rect 181151 518116 182220 518158
rect 182255 518192 183324 518203
rect 182255 518158 182273 518192
rect 182307 518158 183273 518192
rect 183307 518158 183324 518192
rect 182255 518116 183324 518158
rect 183359 518192 184428 518203
rect 183359 518158 183377 518192
rect 183411 518158 184377 518192
rect 184411 518158 184428 518192
rect 183359 518116 184428 518158
rect 184463 518192 184981 518260
rect 184463 518158 184481 518192
rect 184515 518158 184929 518192
rect 184963 518158 184981 518192
rect 184463 518116 184981 518158
rect 185107 518314 185165 518349
rect 185107 518280 185119 518314
rect 185153 518280 185165 518314
rect 185107 518221 185165 518280
rect 185107 518187 185119 518221
rect 185153 518187 185165 518221
rect 185880 518203 185950 518404
rect 186303 518402 186633 518472
rect 186303 518368 186381 518402
rect 186415 518368 186480 518402
rect 186514 518368 186579 518402
rect 186613 518368 186633 518402
rect 186667 518404 186687 518438
rect 186721 518404 186790 518438
rect 186824 518404 186893 518438
rect 186927 518404 187005 518438
rect 186667 518334 187005 518404
rect 186303 518294 187005 518334
rect 186303 518260 186321 518294
rect 186355 518260 186953 518294
rect 186987 518260 187005 518294
rect 185107 518116 185165 518187
rect 185199 518192 186268 518203
rect 185199 518158 185217 518192
rect 185251 518158 186217 518192
rect 186251 518158 186268 518192
rect 185199 518116 186268 518158
rect 186303 518192 187005 518260
rect 186303 518158 186321 518192
rect 186355 518158 186953 518192
rect 186987 518158 187005 518192
rect 186303 518116 187005 518158
rect 187223 518408 187273 518442
rect 187307 518408 187327 518442
rect 187223 518334 187327 518408
rect 187361 518402 187465 518476
rect 187361 518368 187381 518402
rect 187415 518368 187465 518402
rect 187223 518287 187465 518334
rect 187223 518253 187241 518287
rect 187275 518253 187413 518287
rect 187447 518253 187465 518287
rect 187223 518192 187465 518253
rect 187223 518158 187241 518192
rect 187275 518158 187413 518192
rect 187447 518158 187465 518192
rect 187223 518116 187465 518158
rect 172210 518082 172239 518116
rect 172273 518082 172331 518116
rect 172365 518082 172423 518116
rect 172457 518082 172515 518116
rect 172549 518082 172607 518116
rect 172641 518082 172699 518116
rect 172733 518082 172791 518116
rect 172825 518082 172883 518116
rect 172917 518082 172975 518116
rect 173009 518082 173067 518116
rect 173101 518082 173159 518116
rect 173193 518082 173251 518116
rect 173285 518082 173343 518116
rect 173377 518082 173435 518116
rect 173469 518082 173527 518116
rect 173561 518082 173619 518116
rect 173653 518082 173711 518116
rect 173745 518082 173803 518116
rect 173837 518082 173895 518116
rect 173929 518082 173987 518116
rect 174021 518082 174079 518116
rect 174113 518082 174171 518116
rect 174205 518082 174263 518116
rect 174297 518082 174355 518116
rect 174389 518082 174447 518116
rect 174481 518082 174539 518116
rect 174573 518082 174631 518116
rect 174665 518082 174723 518116
rect 174757 518082 174815 518116
rect 174849 518082 174907 518116
rect 174941 518082 174999 518116
rect 175033 518082 175091 518116
rect 175125 518082 175183 518116
rect 175217 518082 175275 518116
rect 175309 518082 175367 518116
rect 175401 518082 175459 518116
rect 175493 518082 175551 518116
rect 175585 518082 175643 518116
rect 175677 518082 175735 518116
rect 175769 518082 175827 518116
rect 175861 518082 175919 518116
rect 175953 518082 176011 518116
rect 176045 518082 176103 518116
rect 176137 518082 176195 518116
rect 176229 518082 176287 518116
rect 176321 518082 176379 518116
rect 176413 518082 176471 518116
rect 176505 518082 176563 518116
rect 176597 518082 176655 518116
rect 176689 518082 176747 518116
rect 176781 518082 176839 518116
rect 176873 518082 176931 518116
rect 176965 518082 177023 518116
rect 177057 518082 177115 518116
rect 177149 518082 177207 518116
rect 177241 518082 177299 518116
rect 177333 518082 177391 518116
rect 177425 518082 177483 518116
rect 177517 518082 177575 518116
rect 177609 518082 177667 518116
rect 177701 518082 177759 518116
rect 177793 518082 177851 518116
rect 177885 518082 177943 518116
rect 177977 518082 178035 518116
rect 178069 518082 178127 518116
rect 178161 518082 178219 518116
rect 178253 518082 178311 518116
rect 178345 518082 178403 518116
rect 178437 518082 178495 518116
rect 178529 518082 178587 518116
rect 178621 518082 178679 518116
rect 178713 518082 178771 518116
rect 178805 518082 178863 518116
rect 178897 518082 178955 518116
rect 178989 518082 179047 518116
rect 179081 518082 179139 518116
rect 179173 518082 179231 518116
rect 179265 518082 179323 518116
rect 179357 518082 179415 518116
rect 179449 518082 179507 518116
rect 179541 518082 179599 518116
rect 179633 518082 179691 518116
rect 179725 518082 179783 518116
rect 179817 518082 179875 518116
rect 179909 518082 179967 518116
rect 180001 518082 180059 518116
rect 180093 518082 180151 518116
rect 180185 518082 180243 518116
rect 180277 518082 180335 518116
rect 180369 518082 180427 518116
rect 180461 518082 180519 518116
rect 180553 518082 180611 518116
rect 180645 518082 180703 518116
rect 180737 518082 180795 518116
rect 180829 518082 180887 518116
rect 180921 518082 180979 518116
rect 181013 518082 181071 518116
rect 181105 518082 181163 518116
rect 181197 518082 181255 518116
rect 181289 518082 181347 518116
rect 181381 518082 181439 518116
rect 181473 518082 181531 518116
rect 181565 518082 181623 518116
rect 181657 518082 181715 518116
rect 181749 518082 181807 518116
rect 181841 518082 181899 518116
rect 181933 518082 181991 518116
rect 182025 518082 182083 518116
rect 182117 518082 182175 518116
rect 182209 518082 182267 518116
rect 182301 518082 182359 518116
rect 182393 518082 182451 518116
rect 182485 518082 182543 518116
rect 182577 518082 182635 518116
rect 182669 518082 182727 518116
rect 182761 518082 182819 518116
rect 182853 518082 182911 518116
rect 182945 518082 183003 518116
rect 183037 518082 183095 518116
rect 183129 518082 183187 518116
rect 183221 518082 183279 518116
rect 183313 518082 183371 518116
rect 183405 518082 183463 518116
rect 183497 518082 183555 518116
rect 183589 518082 183647 518116
rect 183681 518082 183739 518116
rect 183773 518082 183831 518116
rect 183865 518082 183923 518116
rect 183957 518082 184015 518116
rect 184049 518082 184107 518116
rect 184141 518082 184199 518116
rect 184233 518082 184291 518116
rect 184325 518082 184383 518116
rect 184417 518082 184475 518116
rect 184509 518082 184567 518116
rect 184601 518082 184659 518116
rect 184693 518082 184751 518116
rect 184785 518082 184843 518116
rect 184877 518082 184935 518116
rect 184969 518082 185027 518116
rect 185061 518082 185119 518116
rect 185153 518082 185211 518116
rect 185245 518082 185303 518116
rect 185337 518082 185395 518116
rect 185429 518082 185487 518116
rect 185521 518082 185579 518116
rect 185613 518082 185671 518116
rect 185705 518082 185763 518116
rect 185797 518082 185855 518116
rect 185889 518082 185947 518116
rect 185981 518082 186039 518116
rect 186073 518082 186131 518116
rect 186165 518082 186223 518116
rect 186257 518082 186315 518116
rect 186349 518082 186407 518116
rect 186441 518082 186499 518116
rect 186533 518082 186591 518116
rect 186625 518082 186683 518116
rect 186717 518082 186775 518116
rect 186809 518082 186867 518116
rect 186901 518082 186959 518116
rect 186993 518082 187051 518116
rect 187085 518082 187143 518116
rect 187177 518082 187235 518116
rect 187269 518082 187327 518116
rect 187361 518082 187419 518116
rect 187453 518082 187482 518116
rect 172227 518040 172469 518082
rect 172227 518006 172245 518040
rect 172279 518006 172417 518040
rect 172451 518006 172469 518040
rect 172227 517945 172469 518006
rect 172503 518040 173572 518082
rect 172503 518006 172521 518040
rect 172555 518006 173521 518040
rect 173555 518006 173572 518040
rect 172503 517995 173572 518006
rect 173607 518040 174676 518082
rect 173607 518006 173625 518040
rect 173659 518006 174625 518040
rect 174659 518006 174676 518040
rect 173607 517995 174676 518006
rect 174711 518040 175780 518082
rect 174711 518006 174729 518040
rect 174763 518006 175729 518040
rect 175763 518006 175780 518040
rect 174711 517995 175780 518006
rect 175815 518040 176884 518082
rect 175815 518006 175833 518040
rect 175867 518006 176833 518040
rect 176867 518006 176884 518040
rect 175815 517995 176884 518006
rect 176919 518040 177253 518082
rect 176919 518006 176937 518040
rect 176971 518006 177201 518040
rect 177235 518006 177253 518040
rect 172227 517911 172245 517945
rect 172279 517911 172417 517945
rect 172451 517911 172469 517945
rect 172227 517864 172469 517911
rect 172227 517796 172277 517830
rect 172311 517796 172331 517830
rect 172227 517722 172331 517796
rect 172365 517790 172469 517864
rect 172365 517756 172385 517790
rect 172419 517756 172469 517790
rect 172820 517830 172888 517847
rect 172820 517796 172837 517830
rect 172871 517796 172888 517830
rect 172227 517669 172469 517722
rect 172820 517681 172888 517796
rect 173184 517794 173254 517995
rect 173184 517760 173201 517794
rect 173235 517760 173254 517794
rect 173184 517745 173254 517760
rect 173924 517830 173992 517847
rect 173924 517796 173941 517830
rect 173975 517796 173992 517830
rect 173924 517681 173992 517796
rect 174288 517794 174358 517995
rect 174288 517760 174305 517794
rect 174339 517760 174358 517794
rect 174288 517745 174358 517760
rect 175028 517830 175096 517847
rect 175028 517796 175045 517830
rect 175079 517796 175096 517830
rect 175028 517681 175096 517796
rect 175392 517794 175462 517995
rect 175392 517760 175409 517794
rect 175443 517760 175462 517794
rect 175392 517745 175462 517760
rect 176132 517830 176200 517847
rect 176132 517796 176149 517830
rect 176183 517796 176200 517830
rect 176132 517681 176200 517796
rect 176496 517794 176566 517995
rect 176919 517938 177253 518006
rect 176919 517904 176937 517938
rect 176971 517904 177201 517938
rect 177235 517904 177253 517938
rect 176919 517864 177253 517904
rect 176496 517760 176513 517794
rect 176547 517760 176566 517794
rect 176496 517745 176566 517760
rect 176919 517796 176939 517830
rect 176973 517796 177069 517830
rect 176919 517726 177069 517796
rect 177103 517794 177253 517864
rect 177379 518011 177437 518082
rect 177379 517977 177391 518011
rect 177425 517977 177437 518011
rect 177471 518040 178540 518082
rect 177471 518006 177489 518040
rect 177523 518006 178489 518040
rect 178523 518006 178540 518040
rect 177471 517995 178540 518006
rect 178575 518040 179644 518082
rect 178575 518006 178593 518040
rect 178627 518006 179593 518040
rect 179627 518006 179644 518040
rect 178575 517995 179644 518006
rect 179679 518040 180748 518082
rect 179679 518006 179697 518040
rect 179731 518006 180697 518040
rect 180731 518006 180748 518040
rect 179679 517995 180748 518006
rect 180783 518040 181852 518082
rect 180783 518006 180801 518040
rect 180835 518006 181801 518040
rect 181835 518006 181852 518040
rect 180783 517995 181852 518006
rect 181887 518040 182405 518082
rect 181887 518006 181905 518040
rect 181939 518006 182353 518040
rect 182387 518006 182405 518040
rect 177379 517918 177437 517977
rect 177379 517884 177391 517918
rect 177425 517884 177437 517918
rect 177379 517849 177437 517884
rect 177103 517760 177199 517794
rect 177233 517760 177253 517794
rect 177788 517830 177856 517847
rect 177788 517796 177805 517830
rect 177839 517796 177856 517830
rect 172227 517635 172245 517669
rect 172279 517635 172417 517669
rect 172451 517635 172469 517669
rect 172227 517572 172469 517635
rect 172503 517667 173572 517681
rect 172503 517633 172521 517667
rect 172555 517633 173521 517667
rect 173555 517633 173572 517667
rect 172503 517572 173572 517633
rect 173607 517667 174676 517681
rect 173607 517633 173625 517667
rect 173659 517633 174625 517667
rect 174659 517633 174676 517667
rect 173607 517572 174676 517633
rect 174711 517667 175780 517681
rect 174711 517633 174729 517667
rect 174763 517633 175729 517667
rect 175763 517633 175780 517667
rect 174711 517572 175780 517633
rect 175815 517667 176884 517681
rect 175815 517633 175833 517667
rect 175867 517633 176833 517667
rect 176867 517633 176884 517667
rect 175815 517572 176884 517633
rect 176919 517674 177253 517726
rect 176919 517640 176937 517674
rect 176971 517640 177201 517674
rect 177235 517640 177253 517674
rect 176919 517572 177253 517640
rect 177379 517700 177437 517717
rect 177379 517666 177391 517700
rect 177425 517666 177437 517700
rect 177788 517681 177856 517796
rect 178152 517794 178222 517995
rect 178152 517760 178169 517794
rect 178203 517760 178222 517794
rect 178152 517745 178222 517760
rect 178892 517830 178960 517847
rect 178892 517796 178909 517830
rect 178943 517796 178960 517830
rect 178892 517681 178960 517796
rect 179256 517794 179326 517995
rect 179256 517760 179273 517794
rect 179307 517760 179326 517794
rect 179256 517745 179326 517760
rect 179996 517830 180064 517847
rect 179996 517796 180013 517830
rect 180047 517796 180064 517830
rect 179996 517681 180064 517796
rect 180360 517794 180430 517995
rect 180360 517760 180377 517794
rect 180411 517760 180430 517794
rect 180360 517745 180430 517760
rect 181100 517830 181168 517847
rect 181100 517796 181117 517830
rect 181151 517796 181168 517830
rect 181100 517681 181168 517796
rect 181464 517794 181534 517995
rect 181887 517938 182405 518006
rect 181887 517904 181905 517938
rect 181939 517904 182353 517938
rect 182387 517904 182405 517938
rect 181887 517864 182405 517904
rect 181464 517760 181481 517794
rect 181515 517760 181534 517794
rect 181464 517745 181534 517760
rect 181887 517796 181965 517830
rect 181999 517796 182075 517830
rect 182109 517796 182129 517830
rect 181887 517726 182129 517796
rect 182163 517794 182405 517864
rect 182531 518011 182589 518082
rect 182531 517977 182543 518011
rect 182577 517977 182589 518011
rect 182623 518040 183692 518082
rect 182623 518006 182641 518040
rect 182675 518006 183641 518040
rect 183675 518006 183692 518040
rect 182623 517995 183692 518006
rect 183727 518040 184796 518082
rect 183727 518006 183745 518040
rect 183779 518006 184745 518040
rect 184779 518006 184796 518040
rect 183727 517995 184796 518006
rect 184831 518040 185900 518082
rect 184831 518006 184849 518040
rect 184883 518006 185849 518040
rect 185883 518006 185900 518040
rect 184831 517995 185900 518006
rect 185935 518040 187004 518082
rect 185935 518006 185953 518040
rect 185987 518006 186953 518040
rect 186987 518006 187004 518040
rect 185935 517995 187004 518006
rect 187223 518040 187465 518082
rect 187223 518006 187241 518040
rect 187275 518006 187413 518040
rect 187447 518006 187465 518040
rect 182531 517918 182589 517977
rect 182531 517884 182543 517918
rect 182577 517884 182589 517918
rect 182531 517849 182589 517884
rect 182163 517760 182183 517794
rect 182217 517760 182293 517794
rect 182327 517760 182405 517794
rect 182940 517830 183008 517847
rect 182940 517796 182957 517830
rect 182991 517796 183008 517830
rect 177379 517572 177437 517666
rect 177471 517667 178540 517681
rect 177471 517633 177489 517667
rect 177523 517633 178489 517667
rect 178523 517633 178540 517667
rect 177471 517572 178540 517633
rect 178575 517667 179644 517681
rect 178575 517633 178593 517667
rect 178627 517633 179593 517667
rect 179627 517633 179644 517667
rect 178575 517572 179644 517633
rect 179679 517667 180748 517681
rect 179679 517633 179697 517667
rect 179731 517633 180697 517667
rect 180731 517633 180748 517667
rect 179679 517572 180748 517633
rect 180783 517667 181852 517681
rect 180783 517633 180801 517667
rect 180835 517633 181801 517667
rect 181835 517633 181852 517667
rect 180783 517572 181852 517633
rect 181887 517667 182405 517726
rect 181887 517633 181905 517667
rect 181939 517633 182353 517667
rect 182387 517633 182405 517667
rect 181887 517572 182405 517633
rect 182531 517700 182589 517717
rect 182531 517666 182543 517700
rect 182577 517666 182589 517700
rect 182940 517681 183008 517796
rect 183304 517794 183374 517995
rect 183304 517760 183321 517794
rect 183355 517760 183374 517794
rect 183304 517745 183374 517760
rect 184044 517830 184112 517847
rect 184044 517796 184061 517830
rect 184095 517796 184112 517830
rect 184044 517681 184112 517796
rect 184408 517794 184478 517995
rect 184408 517760 184425 517794
rect 184459 517760 184478 517794
rect 184408 517745 184478 517760
rect 185148 517830 185216 517847
rect 185148 517796 185165 517830
rect 185199 517796 185216 517830
rect 185148 517681 185216 517796
rect 185512 517794 185582 517995
rect 185512 517760 185529 517794
rect 185563 517760 185582 517794
rect 185512 517745 185582 517760
rect 186252 517830 186320 517847
rect 186252 517796 186269 517830
rect 186303 517796 186320 517830
rect 186252 517681 186320 517796
rect 186616 517794 186686 517995
rect 186616 517760 186633 517794
rect 186667 517760 186686 517794
rect 186616 517745 186686 517760
rect 187223 517945 187465 518006
rect 187223 517911 187241 517945
rect 187275 517911 187413 517945
rect 187447 517911 187465 517945
rect 187223 517864 187465 517911
rect 187223 517790 187327 517864
rect 187223 517756 187273 517790
rect 187307 517756 187327 517790
rect 187361 517796 187381 517830
rect 187415 517796 187465 517830
rect 187361 517722 187465 517796
rect 182531 517572 182589 517666
rect 182623 517667 183692 517681
rect 182623 517633 182641 517667
rect 182675 517633 183641 517667
rect 183675 517633 183692 517667
rect 182623 517572 183692 517633
rect 183727 517667 184796 517681
rect 183727 517633 183745 517667
rect 183779 517633 184745 517667
rect 184779 517633 184796 517667
rect 183727 517572 184796 517633
rect 184831 517667 185900 517681
rect 184831 517633 184849 517667
rect 184883 517633 185849 517667
rect 185883 517633 185900 517667
rect 184831 517572 185900 517633
rect 185935 517667 187004 517681
rect 185935 517633 185953 517667
rect 185987 517633 186953 517667
rect 186987 517633 187004 517667
rect 185935 517572 187004 517633
rect 187223 517669 187465 517722
rect 187223 517635 187241 517669
rect 187275 517635 187413 517669
rect 187447 517635 187465 517669
rect 187223 517572 187465 517635
rect 172210 517538 172239 517572
rect 172273 517538 172331 517572
rect 172365 517538 172423 517572
rect 172457 517538 172515 517572
rect 172549 517538 172607 517572
rect 172641 517538 172699 517572
rect 172733 517538 172791 517572
rect 172825 517538 172883 517572
rect 172917 517538 172975 517572
rect 173009 517538 173067 517572
rect 173101 517538 173159 517572
rect 173193 517538 173251 517572
rect 173285 517538 173343 517572
rect 173377 517538 173435 517572
rect 173469 517538 173527 517572
rect 173561 517538 173619 517572
rect 173653 517538 173711 517572
rect 173745 517538 173803 517572
rect 173837 517538 173895 517572
rect 173929 517538 173987 517572
rect 174021 517538 174079 517572
rect 174113 517538 174171 517572
rect 174205 517538 174263 517572
rect 174297 517538 174355 517572
rect 174389 517538 174447 517572
rect 174481 517538 174539 517572
rect 174573 517538 174631 517572
rect 174665 517538 174723 517572
rect 174757 517538 174815 517572
rect 174849 517538 174907 517572
rect 174941 517538 174999 517572
rect 175033 517538 175091 517572
rect 175125 517538 175183 517572
rect 175217 517538 175275 517572
rect 175309 517538 175367 517572
rect 175401 517538 175459 517572
rect 175493 517538 175551 517572
rect 175585 517538 175643 517572
rect 175677 517538 175735 517572
rect 175769 517538 175827 517572
rect 175861 517538 175919 517572
rect 175953 517538 176011 517572
rect 176045 517538 176103 517572
rect 176137 517538 176195 517572
rect 176229 517538 176287 517572
rect 176321 517538 176379 517572
rect 176413 517538 176471 517572
rect 176505 517538 176563 517572
rect 176597 517538 176655 517572
rect 176689 517538 176747 517572
rect 176781 517538 176839 517572
rect 176873 517538 176931 517572
rect 176965 517538 177023 517572
rect 177057 517538 177115 517572
rect 177149 517538 177207 517572
rect 177241 517538 177299 517572
rect 177333 517538 177391 517572
rect 177425 517538 177483 517572
rect 177517 517538 177575 517572
rect 177609 517538 177667 517572
rect 177701 517538 177759 517572
rect 177793 517538 177851 517572
rect 177885 517538 177943 517572
rect 177977 517538 178035 517572
rect 178069 517538 178127 517572
rect 178161 517538 178219 517572
rect 178253 517538 178311 517572
rect 178345 517538 178403 517572
rect 178437 517538 178495 517572
rect 178529 517538 178587 517572
rect 178621 517538 178679 517572
rect 178713 517538 178771 517572
rect 178805 517538 178863 517572
rect 178897 517538 178955 517572
rect 178989 517538 179047 517572
rect 179081 517538 179139 517572
rect 179173 517538 179231 517572
rect 179265 517538 179323 517572
rect 179357 517538 179415 517572
rect 179449 517538 179507 517572
rect 179541 517538 179599 517572
rect 179633 517538 179691 517572
rect 179725 517538 179783 517572
rect 179817 517538 179875 517572
rect 179909 517538 179967 517572
rect 180001 517538 180059 517572
rect 180093 517538 180151 517572
rect 180185 517538 180243 517572
rect 180277 517538 180335 517572
rect 180369 517538 180427 517572
rect 180461 517538 180519 517572
rect 180553 517538 180611 517572
rect 180645 517538 180703 517572
rect 180737 517538 180795 517572
rect 180829 517538 180887 517572
rect 180921 517538 180979 517572
rect 181013 517538 181071 517572
rect 181105 517538 181163 517572
rect 181197 517538 181255 517572
rect 181289 517538 181347 517572
rect 181381 517538 181439 517572
rect 181473 517538 181531 517572
rect 181565 517538 181623 517572
rect 181657 517538 181715 517572
rect 181749 517538 181807 517572
rect 181841 517538 181899 517572
rect 181933 517538 181991 517572
rect 182025 517538 182083 517572
rect 182117 517538 182175 517572
rect 182209 517538 182267 517572
rect 182301 517538 182359 517572
rect 182393 517538 182451 517572
rect 182485 517538 182543 517572
rect 182577 517538 182635 517572
rect 182669 517538 182727 517572
rect 182761 517538 182819 517572
rect 182853 517538 182911 517572
rect 182945 517538 183003 517572
rect 183037 517538 183095 517572
rect 183129 517538 183187 517572
rect 183221 517538 183279 517572
rect 183313 517538 183371 517572
rect 183405 517538 183463 517572
rect 183497 517538 183555 517572
rect 183589 517538 183647 517572
rect 183681 517538 183739 517572
rect 183773 517538 183831 517572
rect 183865 517538 183923 517572
rect 183957 517538 184015 517572
rect 184049 517538 184107 517572
rect 184141 517538 184199 517572
rect 184233 517538 184291 517572
rect 184325 517538 184383 517572
rect 184417 517538 184475 517572
rect 184509 517538 184567 517572
rect 184601 517538 184659 517572
rect 184693 517538 184751 517572
rect 184785 517538 184843 517572
rect 184877 517538 184935 517572
rect 184969 517538 185027 517572
rect 185061 517538 185119 517572
rect 185153 517538 185211 517572
rect 185245 517538 185303 517572
rect 185337 517538 185395 517572
rect 185429 517538 185487 517572
rect 185521 517538 185579 517572
rect 185613 517538 185671 517572
rect 185705 517538 185763 517572
rect 185797 517538 185855 517572
rect 185889 517538 185947 517572
rect 185981 517538 186039 517572
rect 186073 517538 186131 517572
rect 186165 517538 186223 517572
rect 186257 517538 186315 517572
rect 186349 517538 186407 517572
rect 186441 517538 186499 517572
rect 186533 517538 186591 517572
rect 186625 517538 186683 517572
rect 186717 517538 186775 517572
rect 186809 517538 186867 517572
rect 186901 517538 186959 517572
rect 186993 517538 187051 517572
rect 187085 517538 187143 517572
rect 187177 517538 187235 517572
rect 187269 517538 187327 517572
rect 187361 517538 187419 517572
rect 187453 517538 187482 517572
rect 172227 517475 172469 517538
rect 172227 517441 172245 517475
rect 172279 517441 172417 517475
rect 172451 517441 172469 517475
rect 172227 517388 172469 517441
rect 172503 517477 173572 517538
rect 172503 517443 172521 517477
rect 172555 517443 173521 517477
rect 173555 517443 173572 517477
rect 172503 517429 173572 517443
rect 173607 517477 174676 517538
rect 173607 517443 173625 517477
rect 173659 517443 174625 517477
rect 174659 517443 174676 517477
rect 173607 517429 174676 517443
rect 174803 517444 174861 517538
rect 172227 517314 172331 517388
rect 172227 517280 172277 517314
rect 172311 517280 172331 517314
rect 172365 517320 172385 517354
rect 172419 517320 172469 517354
rect 172365 517246 172469 517320
rect 172820 517314 172888 517429
rect 172820 517280 172837 517314
rect 172871 517280 172888 517314
rect 172820 517263 172888 517280
rect 173184 517350 173254 517365
rect 173184 517316 173201 517350
rect 173235 517316 173254 517350
rect 172227 517199 172469 517246
rect 172227 517165 172245 517199
rect 172279 517165 172417 517199
rect 172451 517165 172469 517199
rect 172227 517104 172469 517165
rect 173184 517115 173254 517316
rect 173924 517314 173992 517429
rect 174803 517410 174815 517444
rect 174849 517410 174861 517444
rect 174895 517477 175964 517538
rect 174895 517443 174913 517477
rect 174947 517443 175913 517477
rect 175947 517443 175964 517477
rect 174895 517429 175964 517443
rect 175999 517477 177068 517538
rect 175999 517443 176017 517477
rect 176051 517443 177017 517477
rect 177051 517443 177068 517477
rect 175999 517429 177068 517443
rect 177103 517477 178172 517538
rect 177103 517443 177121 517477
rect 177155 517443 178121 517477
rect 178155 517443 178172 517477
rect 177103 517429 178172 517443
rect 178207 517477 179276 517538
rect 178207 517443 178225 517477
rect 178259 517443 179225 517477
rect 179259 517443 179276 517477
rect 178207 517429 179276 517443
rect 179311 517477 179829 517538
rect 179311 517443 179329 517477
rect 179363 517443 179777 517477
rect 179811 517443 179829 517477
rect 174803 517393 174861 517410
rect 173924 517280 173941 517314
rect 173975 517280 173992 517314
rect 173924 517263 173992 517280
rect 174288 517350 174358 517365
rect 174288 517316 174305 517350
rect 174339 517316 174358 517350
rect 174288 517115 174358 517316
rect 175212 517314 175280 517429
rect 175212 517280 175229 517314
rect 175263 517280 175280 517314
rect 175212 517263 175280 517280
rect 175576 517350 175646 517365
rect 175576 517316 175593 517350
rect 175627 517316 175646 517350
rect 174803 517226 174861 517261
rect 174803 517192 174815 517226
rect 174849 517192 174861 517226
rect 174803 517133 174861 517192
rect 172227 517070 172245 517104
rect 172279 517070 172417 517104
rect 172451 517070 172469 517104
rect 172227 517028 172469 517070
rect 172503 517104 173572 517115
rect 172503 517070 172521 517104
rect 172555 517070 173521 517104
rect 173555 517070 173572 517104
rect 172503 517028 173572 517070
rect 173607 517104 174676 517115
rect 173607 517070 173625 517104
rect 173659 517070 174625 517104
rect 174659 517070 174676 517104
rect 173607 517028 174676 517070
rect 174803 517099 174815 517133
rect 174849 517099 174861 517133
rect 175576 517115 175646 517316
rect 176316 517314 176384 517429
rect 176316 517280 176333 517314
rect 176367 517280 176384 517314
rect 176316 517263 176384 517280
rect 176680 517350 176750 517365
rect 176680 517316 176697 517350
rect 176731 517316 176750 517350
rect 176680 517115 176750 517316
rect 177420 517314 177488 517429
rect 177420 517280 177437 517314
rect 177471 517280 177488 517314
rect 177420 517263 177488 517280
rect 177784 517350 177854 517365
rect 177784 517316 177801 517350
rect 177835 517316 177854 517350
rect 177784 517115 177854 517316
rect 178524 517314 178592 517429
rect 179311 517384 179829 517443
rect 179955 517444 180013 517538
rect 179955 517410 179967 517444
rect 180001 517410 180013 517444
rect 180047 517477 181116 517538
rect 180047 517443 180065 517477
rect 180099 517443 181065 517477
rect 181099 517443 181116 517477
rect 180047 517429 181116 517443
rect 181151 517477 182220 517538
rect 181151 517443 181169 517477
rect 181203 517443 182169 517477
rect 182203 517443 182220 517477
rect 181151 517429 182220 517443
rect 182255 517477 183324 517538
rect 182255 517443 182273 517477
rect 182307 517443 183273 517477
rect 183307 517443 183324 517477
rect 182255 517429 183324 517443
rect 183359 517477 184428 517538
rect 183359 517443 183377 517477
rect 183411 517443 184377 517477
rect 184411 517443 184428 517477
rect 183359 517429 184428 517443
rect 184463 517477 184981 517538
rect 184463 517443 184481 517477
rect 184515 517443 184929 517477
rect 184963 517443 184981 517477
rect 179955 517393 180013 517410
rect 178524 517280 178541 517314
rect 178575 517280 178592 517314
rect 178524 517263 178592 517280
rect 178888 517350 178958 517365
rect 178888 517316 178905 517350
rect 178939 517316 178958 517350
rect 178888 517115 178958 517316
rect 179311 517314 179553 517384
rect 179311 517280 179389 517314
rect 179423 517280 179499 517314
rect 179533 517280 179553 517314
rect 179587 517316 179607 517350
rect 179641 517316 179717 517350
rect 179751 517316 179829 517350
rect 179587 517246 179829 517316
rect 180364 517314 180432 517429
rect 180364 517280 180381 517314
rect 180415 517280 180432 517314
rect 180364 517263 180432 517280
rect 180728 517350 180798 517365
rect 180728 517316 180745 517350
rect 180779 517316 180798 517350
rect 179311 517206 179829 517246
rect 179311 517172 179329 517206
rect 179363 517172 179777 517206
rect 179811 517172 179829 517206
rect 174803 517028 174861 517099
rect 174895 517104 175964 517115
rect 174895 517070 174913 517104
rect 174947 517070 175913 517104
rect 175947 517070 175964 517104
rect 174895 517028 175964 517070
rect 175999 517104 177068 517115
rect 175999 517070 176017 517104
rect 176051 517070 177017 517104
rect 177051 517070 177068 517104
rect 175999 517028 177068 517070
rect 177103 517104 178172 517115
rect 177103 517070 177121 517104
rect 177155 517070 178121 517104
rect 178155 517070 178172 517104
rect 177103 517028 178172 517070
rect 178207 517104 179276 517115
rect 178207 517070 178225 517104
rect 178259 517070 179225 517104
rect 179259 517070 179276 517104
rect 178207 517028 179276 517070
rect 179311 517104 179829 517172
rect 179311 517070 179329 517104
rect 179363 517070 179777 517104
rect 179811 517070 179829 517104
rect 179311 517028 179829 517070
rect 179955 517226 180013 517261
rect 179955 517192 179967 517226
rect 180001 517192 180013 517226
rect 179955 517133 180013 517192
rect 179955 517099 179967 517133
rect 180001 517099 180013 517133
rect 180728 517115 180798 517316
rect 181468 517314 181536 517429
rect 181468 517280 181485 517314
rect 181519 517280 181536 517314
rect 181468 517263 181536 517280
rect 181832 517350 181902 517365
rect 181832 517316 181849 517350
rect 181883 517316 181902 517350
rect 181832 517115 181902 517316
rect 182572 517314 182640 517429
rect 182572 517280 182589 517314
rect 182623 517280 182640 517314
rect 182572 517263 182640 517280
rect 182936 517350 183006 517365
rect 182936 517316 182953 517350
rect 182987 517316 183006 517350
rect 182936 517115 183006 517316
rect 183676 517314 183744 517429
rect 184463 517384 184981 517443
rect 185107 517444 185165 517538
rect 185107 517410 185119 517444
rect 185153 517410 185165 517444
rect 185199 517477 186268 517538
rect 185199 517443 185217 517477
rect 185251 517443 186217 517477
rect 186251 517443 186268 517477
rect 185199 517429 186268 517443
rect 186303 517477 187005 517538
rect 186303 517443 186321 517477
rect 186355 517443 186953 517477
rect 186987 517443 187005 517477
rect 185107 517393 185165 517410
rect 183676 517280 183693 517314
rect 183727 517280 183744 517314
rect 183676 517263 183744 517280
rect 184040 517350 184110 517365
rect 184040 517316 184057 517350
rect 184091 517316 184110 517350
rect 184040 517115 184110 517316
rect 184463 517314 184705 517384
rect 184463 517280 184541 517314
rect 184575 517280 184651 517314
rect 184685 517280 184705 517314
rect 184739 517316 184759 517350
rect 184793 517316 184869 517350
rect 184903 517316 184981 517350
rect 184739 517246 184981 517316
rect 185516 517314 185584 517429
rect 186303 517384 187005 517443
rect 187223 517475 187465 517538
rect 187223 517441 187241 517475
rect 187275 517441 187413 517475
rect 187447 517441 187465 517475
rect 187223 517388 187465 517441
rect 185516 517280 185533 517314
rect 185567 517280 185584 517314
rect 185516 517263 185584 517280
rect 185880 517350 185950 517365
rect 185880 517316 185897 517350
rect 185931 517316 185950 517350
rect 184463 517206 184981 517246
rect 184463 517172 184481 517206
rect 184515 517172 184929 517206
rect 184963 517172 184981 517206
rect 179955 517028 180013 517099
rect 180047 517104 181116 517115
rect 180047 517070 180065 517104
rect 180099 517070 181065 517104
rect 181099 517070 181116 517104
rect 180047 517028 181116 517070
rect 181151 517104 182220 517115
rect 181151 517070 181169 517104
rect 181203 517070 182169 517104
rect 182203 517070 182220 517104
rect 181151 517028 182220 517070
rect 182255 517104 183324 517115
rect 182255 517070 182273 517104
rect 182307 517070 183273 517104
rect 183307 517070 183324 517104
rect 182255 517028 183324 517070
rect 183359 517104 184428 517115
rect 183359 517070 183377 517104
rect 183411 517070 184377 517104
rect 184411 517070 184428 517104
rect 183359 517028 184428 517070
rect 184463 517104 184981 517172
rect 184463 517070 184481 517104
rect 184515 517070 184929 517104
rect 184963 517070 184981 517104
rect 184463 517028 184981 517070
rect 185107 517226 185165 517261
rect 185107 517192 185119 517226
rect 185153 517192 185165 517226
rect 185107 517133 185165 517192
rect 185107 517099 185119 517133
rect 185153 517099 185165 517133
rect 185880 517115 185950 517316
rect 186303 517314 186633 517384
rect 186303 517280 186381 517314
rect 186415 517280 186480 517314
rect 186514 517280 186579 517314
rect 186613 517280 186633 517314
rect 186667 517316 186687 517350
rect 186721 517316 186790 517350
rect 186824 517316 186893 517350
rect 186927 517316 187005 517350
rect 186667 517246 187005 517316
rect 186303 517206 187005 517246
rect 186303 517172 186321 517206
rect 186355 517172 186953 517206
rect 186987 517172 187005 517206
rect 185107 517028 185165 517099
rect 185199 517104 186268 517115
rect 185199 517070 185217 517104
rect 185251 517070 186217 517104
rect 186251 517070 186268 517104
rect 185199 517028 186268 517070
rect 186303 517104 187005 517172
rect 186303 517070 186321 517104
rect 186355 517070 186953 517104
rect 186987 517070 187005 517104
rect 186303 517028 187005 517070
rect 187223 517320 187273 517354
rect 187307 517320 187327 517354
rect 187223 517246 187327 517320
rect 187361 517314 187465 517388
rect 187361 517280 187381 517314
rect 187415 517280 187465 517314
rect 187223 517199 187465 517246
rect 187223 517165 187241 517199
rect 187275 517165 187413 517199
rect 187447 517165 187465 517199
rect 187223 517104 187465 517165
rect 187223 517070 187241 517104
rect 187275 517070 187413 517104
rect 187447 517070 187465 517104
rect 187223 517028 187465 517070
rect 172210 516994 172239 517028
rect 172273 516994 172331 517028
rect 172365 516994 172423 517028
rect 172457 516994 172515 517028
rect 172549 516994 172607 517028
rect 172641 516994 172699 517028
rect 172733 516994 172791 517028
rect 172825 516994 172883 517028
rect 172917 516994 172975 517028
rect 173009 516994 173067 517028
rect 173101 516994 173159 517028
rect 173193 516994 173251 517028
rect 173285 516994 173343 517028
rect 173377 516994 173435 517028
rect 173469 516994 173527 517028
rect 173561 516994 173619 517028
rect 173653 516994 173711 517028
rect 173745 516994 173803 517028
rect 173837 516994 173895 517028
rect 173929 516994 173987 517028
rect 174021 516994 174079 517028
rect 174113 516994 174171 517028
rect 174205 516994 174263 517028
rect 174297 516994 174355 517028
rect 174389 516994 174447 517028
rect 174481 516994 174539 517028
rect 174573 516994 174631 517028
rect 174665 516994 174723 517028
rect 174757 516994 174815 517028
rect 174849 516994 174907 517028
rect 174941 516994 174999 517028
rect 175033 516994 175091 517028
rect 175125 516994 175183 517028
rect 175217 516994 175275 517028
rect 175309 516994 175367 517028
rect 175401 516994 175459 517028
rect 175493 516994 175551 517028
rect 175585 516994 175643 517028
rect 175677 516994 175735 517028
rect 175769 516994 175827 517028
rect 175861 516994 175919 517028
rect 175953 516994 176011 517028
rect 176045 516994 176103 517028
rect 176137 516994 176195 517028
rect 176229 516994 176287 517028
rect 176321 516994 176379 517028
rect 176413 516994 176471 517028
rect 176505 516994 176563 517028
rect 176597 516994 176655 517028
rect 176689 516994 176747 517028
rect 176781 516994 176839 517028
rect 176873 516994 176931 517028
rect 176965 516994 177023 517028
rect 177057 516994 177115 517028
rect 177149 516994 177207 517028
rect 177241 516994 177299 517028
rect 177333 516994 177391 517028
rect 177425 516994 177483 517028
rect 177517 516994 177575 517028
rect 177609 516994 177667 517028
rect 177701 516994 177759 517028
rect 177793 516994 177851 517028
rect 177885 516994 177943 517028
rect 177977 516994 178035 517028
rect 178069 516994 178127 517028
rect 178161 516994 178219 517028
rect 178253 516994 178311 517028
rect 178345 516994 178403 517028
rect 178437 516994 178495 517028
rect 178529 516994 178587 517028
rect 178621 516994 178679 517028
rect 178713 516994 178771 517028
rect 178805 516994 178863 517028
rect 178897 516994 178955 517028
rect 178989 516994 179047 517028
rect 179081 516994 179139 517028
rect 179173 516994 179231 517028
rect 179265 516994 179323 517028
rect 179357 516994 179415 517028
rect 179449 516994 179507 517028
rect 179541 516994 179599 517028
rect 179633 516994 179691 517028
rect 179725 516994 179783 517028
rect 179817 516994 179875 517028
rect 179909 516994 179967 517028
rect 180001 516994 180059 517028
rect 180093 516994 180151 517028
rect 180185 516994 180243 517028
rect 180277 516994 180335 517028
rect 180369 516994 180427 517028
rect 180461 516994 180519 517028
rect 180553 516994 180611 517028
rect 180645 516994 180703 517028
rect 180737 516994 180795 517028
rect 180829 516994 180887 517028
rect 180921 516994 180979 517028
rect 181013 516994 181071 517028
rect 181105 516994 181163 517028
rect 181197 516994 181255 517028
rect 181289 516994 181347 517028
rect 181381 516994 181439 517028
rect 181473 516994 181531 517028
rect 181565 516994 181623 517028
rect 181657 516994 181715 517028
rect 181749 516994 181807 517028
rect 181841 516994 181899 517028
rect 181933 516994 181991 517028
rect 182025 516994 182083 517028
rect 182117 516994 182175 517028
rect 182209 516994 182267 517028
rect 182301 516994 182359 517028
rect 182393 516994 182451 517028
rect 182485 516994 182543 517028
rect 182577 516994 182635 517028
rect 182669 516994 182727 517028
rect 182761 516994 182819 517028
rect 182853 516994 182911 517028
rect 182945 516994 183003 517028
rect 183037 516994 183095 517028
rect 183129 516994 183187 517028
rect 183221 516994 183279 517028
rect 183313 516994 183371 517028
rect 183405 516994 183463 517028
rect 183497 516994 183555 517028
rect 183589 516994 183647 517028
rect 183681 516994 183739 517028
rect 183773 516994 183831 517028
rect 183865 516994 183923 517028
rect 183957 516994 184015 517028
rect 184049 516994 184107 517028
rect 184141 516994 184199 517028
rect 184233 516994 184291 517028
rect 184325 516994 184383 517028
rect 184417 516994 184475 517028
rect 184509 516994 184567 517028
rect 184601 516994 184659 517028
rect 184693 516994 184751 517028
rect 184785 516994 184843 517028
rect 184877 516994 184935 517028
rect 184969 516994 185027 517028
rect 185061 516994 185119 517028
rect 185153 516994 185211 517028
rect 185245 516994 185303 517028
rect 185337 516994 185395 517028
rect 185429 516994 185487 517028
rect 185521 516994 185579 517028
rect 185613 516994 185671 517028
rect 185705 516994 185763 517028
rect 185797 516994 185855 517028
rect 185889 516994 185947 517028
rect 185981 516994 186039 517028
rect 186073 516994 186131 517028
rect 186165 516994 186223 517028
rect 186257 516994 186315 517028
rect 186349 516994 186407 517028
rect 186441 516994 186499 517028
rect 186533 516994 186591 517028
rect 186625 516994 186683 517028
rect 186717 516994 186775 517028
rect 186809 516994 186867 517028
rect 186901 516994 186959 517028
rect 186993 516994 187051 517028
rect 187085 516994 187143 517028
rect 187177 516994 187235 517028
rect 187269 516994 187327 517028
rect 187361 516994 187419 517028
rect 187453 516994 187482 517028
rect 172227 516952 172469 516994
rect 172227 516918 172245 516952
rect 172279 516918 172417 516952
rect 172451 516918 172469 516952
rect 172227 516857 172469 516918
rect 172503 516952 173572 516994
rect 172503 516918 172521 516952
rect 172555 516918 173521 516952
rect 173555 516918 173572 516952
rect 172503 516907 173572 516918
rect 173607 516952 174676 516994
rect 173607 516918 173625 516952
rect 173659 516918 174625 516952
rect 174659 516918 174676 516952
rect 173607 516907 174676 516918
rect 174711 516952 175780 516994
rect 174711 516918 174729 516952
rect 174763 516918 175729 516952
rect 175763 516918 175780 516952
rect 174711 516907 175780 516918
rect 175815 516952 176884 516994
rect 175815 516918 175833 516952
rect 175867 516918 176833 516952
rect 176867 516918 176884 516952
rect 175815 516907 176884 516918
rect 176919 516952 177253 516994
rect 176919 516918 176937 516952
rect 176971 516918 177201 516952
rect 177235 516918 177253 516952
rect 172227 516823 172245 516857
rect 172279 516823 172417 516857
rect 172451 516823 172469 516857
rect 172227 516776 172469 516823
rect 172227 516708 172277 516742
rect 172311 516708 172331 516742
rect 172227 516634 172331 516708
rect 172365 516702 172469 516776
rect 172365 516668 172385 516702
rect 172419 516668 172469 516702
rect 172820 516742 172888 516759
rect 172820 516708 172837 516742
rect 172871 516708 172888 516742
rect 172227 516581 172469 516634
rect 172820 516593 172888 516708
rect 173184 516706 173254 516907
rect 173184 516672 173201 516706
rect 173235 516672 173254 516706
rect 173184 516657 173254 516672
rect 173924 516742 173992 516759
rect 173924 516708 173941 516742
rect 173975 516708 173992 516742
rect 173924 516593 173992 516708
rect 174288 516706 174358 516907
rect 174288 516672 174305 516706
rect 174339 516672 174358 516706
rect 174288 516657 174358 516672
rect 175028 516742 175096 516759
rect 175028 516708 175045 516742
rect 175079 516708 175096 516742
rect 175028 516593 175096 516708
rect 175392 516706 175462 516907
rect 175392 516672 175409 516706
rect 175443 516672 175462 516706
rect 175392 516657 175462 516672
rect 176132 516742 176200 516759
rect 176132 516708 176149 516742
rect 176183 516708 176200 516742
rect 176132 516593 176200 516708
rect 176496 516706 176566 516907
rect 176919 516850 177253 516918
rect 176919 516816 176937 516850
rect 176971 516816 177201 516850
rect 177235 516816 177253 516850
rect 176919 516776 177253 516816
rect 176496 516672 176513 516706
rect 176547 516672 176566 516706
rect 176496 516657 176566 516672
rect 176919 516708 176939 516742
rect 176973 516708 177069 516742
rect 176919 516638 177069 516708
rect 177103 516706 177253 516776
rect 177379 516923 177437 516994
rect 177379 516889 177391 516923
rect 177425 516889 177437 516923
rect 177471 516952 178540 516994
rect 177471 516918 177489 516952
rect 177523 516918 178489 516952
rect 178523 516918 178540 516952
rect 177471 516907 178540 516918
rect 178575 516952 179644 516994
rect 178575 516918 178593 516952
rect 178627 516918 179593 516952
rect 179627 516918 179644 516952
rect 178575 516907 179644 516918
rect 179679 516952 180748 516994
rect 179679 516918 179697 516952
rect 179731 516918 180697 516952
rect 180731 516918 180748 516952
rect 179679 516907 180748 516918
rect 180783 516952 181852 516994
rect 180783 516918 180801 516952
rect 180835 516918 181801 516952
rect 181835 516918 181852 516952
rect 180783 516907 181852 516918
rect 181887 516952 182405 516994
rect 181887 516918 181905 516952
rect 181939 516918 182353 516952
rect 182387 516918 182405 516952
rect 177379 516830 177437 516889
rect 177379 516796 177391 516830
rect 177425 516796 177437 516830
rect 177379 516761 177437 516796
rect 177103 516672 177199 516706
rect 177233 516672 177253 516706
rect 177788 516742 177856 516759
rect 177788 516708 177805 516742
rect 177839 516708 177856 516742
rect 172227 516547 172245 516581
rect 172279 516547 172417 516581
rect 172451 516547 172469 516581
rect 172227 516484 172469 516547
rect 172503 516579 173572 516593
rect 172503 516545 172521 516579
rect 172555 516545 173521 516579
rect 173555 516545 173572 516579
rect 172503 516484 173572 516545
rect 173607 516579 174676 516593
rect 173607 516545 173625 516579
rect 173659 516545 174625 516579
rect 174659 516545 174676 516579
rect 173607 516484 174676 516545
rect 174711 516579 175780 516593
rect 174711 516545 174729 516579
rect 174763 516545 175729 516579
rect 175763 516545 175780 516579
rect 174711 516484 175780 516545
rect 175815 516579 176884 516593
rect 175815 516545 175833 516579
rect 175867 516545 176833 516579
rect 176867 516545 176884 516579
rect 175815 516484 176884 516545
rect 176919 516586 177253 516638
rect 176919 516552 176937 516586
rect 176971 516552 177201 516586
rect 177235 516552 177253 516586
rect 176919 516484 177253 516552
rect 177379 516612 177437 516629
rect 177379 516578 177391 516612
rect 177425 516578 177437 516612
rect 177788 516593 177856 516708
rect 178152 516706 178222 516907
rect 178152 516672 178169 516706
rect 178203 516672 178222 516706
rect 178152 516657 178222 516672
rect 178892 516742 178960 516759
rect 178892 516708 178909 516742
rect 178943 516708 178960 516742
rect 178892 516593 178960 516708
rect 179256 516706 179326 516907
rect 179256 516672 179273 516706
rect 179307 516672 179326 516706
rect 179256 516657 179326 516672
rect 179996 516742 180064 516759
rect 179996 516708 180013 516742
rect 180047 516708 180064 516742
rect 179996 516593 180064 516708
rect 180360 516706 180430 516907
rect 180360 516672 180377 516706
rect 180411 516672 180430 516706
rect 180360 516657 180430 516672
rect 181100 516742 181168 516759
rect 181100 516708 181117 516742
rect 181151 516708 181168 516742
rect 181100 516593 181168 516708
rect 181464 516706 181534 516907
rect 181887 516850 182405 516918
rect 181887 516816 181905 516850
rect 181939 516816 182353 516850
rect 182387 516816 182405 516850
rect 181887 516776 182405 516816
rect 181464 516672 181481 516706
rect 181515 516672 181534 516706
rect 181464 516657 181534 516672
rect 181887 516708 181965 516742
rect 181999 516708 182075 516742
rect 182109 516708 182129 516742
rect 181887 516638 182129 516708
rect 182163 516706 182405 516776
rect 182531 516923 182589 516994
rect 182531 516889 182543 516923
rect 182577 516889 182589 516923
rect 182623 516952 183692 516994
rect 182623 516918 182641 516952
rect 182675 516918 183641 516952
rect 183675 516918 183692 516952
rect 182623 516907 183692 516918
rect 183727 516952 184796 516994
rect 183727 516918 183745 516952
rect 183779 516918 184745 516952
rect 184779 516918 184796 516952
rect 183727 516907 184796 516918
rect 184831 516952 185900 516994
rect 184831 516918 184849 516952
rect 184883 516918 185849 516952
rect 185883 516918 185900 516952
rect 184831 516907 185900 516918
rect 185935 516952 187004 516994
rect 185935 516918 185953 516952
rect 185987 516918 186953 516952
rect 186987 516918 187004 516952
rect 185935 516907 187004 516918
rect 187223 516952 187465 516994
rect 187223 516918 187241 516952
rect 187275 516918 187413 516952
rect 187447 516918 187465 516952
rect 182531 516830 182589 516889
rect 182531 516796 182543 516830
rect 182577 516796 182589 516830
rect 182531 516761 182589 516796
rect 182163 516672 182183 516706
rect 182217 516672 182293 516706
rect 182327 516672 182405 516706
rect 182940 516742 183008 516759
rect 182940 516708 182957 516742
rect 182991 516708 183008 516742
rect 177379 516484 177437 516578
rect 177471 516579 178540 516593
rect 177471 516545 177489 516579
rect 177523 516545 178489 516579
rect 178523 516545 178540 516579
rect 177471 516484 178540 516545
rect 178575 516579 179644 516593
rect 178575 516545 178593 516579
rect 178627 516545 179593 516579
rect 179627 516545 179644 516579
rect 178575 516484 179644 516545
rect 179679 516579 180748 516593
rect 179679 516545 179697 516579
rect 179731 516545 180697 516579
rect 180731 516545 180748 516579
rect 179679 516484 180748 516545
rect 180783 516579 181852 516593
rect 180783 516545 180801 516579
rect 180835 516545 181801 516579
rect 181835 516545 181852 516579
rect 180783 516484 181852 516545
rect 181887 516579 182405 516638
rect 181887 516545 181905 516579
rect 181939 516545 182353 516579
rect 182387 516545 182405 516579
rect 181887 516484 182405 516545
rect 182531 516612 182589 516629
rect 182531 516578 182543 516612
rect 182577 516578 182589 516612
rect 182940 516593 183008 516708
rect 183304 516706 183374 516907
rect 183304 516672 183321 516706
rect 183355 516672 183374 516706
rect 183304 516657 183374 516672
rect 184044 516742 184112 516759
rect 184044 516708 184061 516742
rect 184095 516708 184112 516742
rect 184044 516593 184112 516708
rect 184408 516706 184478 516907
rect 184408 516672 184425 516706
rect 184459 516672 184478 516706
rect 184408 516657 184478 516672
rect 185148 516742 185216 516759
rect 185148 516708 185165 516742
rect 185199 516708 185216 516742
rect 185148 516593 185216 516708
rect 185512 516706 185582 516907
rect 185512 516672 185529 516706
rect 185563 516672 185582 516706
rect 185512 516657 185582 516672
rect 186252 516742 186320 516759
rect 186252 516708 186269 516742
rect 186303 516708 186320 516742
rect 186252 516593 186320 516708
rect 186616 516706 186686 516907
rect 186616 516672 186633 516706
rect 186667 516672 186686 516706
rect 186616 516657 186686 516672
rect 187223 516857 187465 516918
rect 187223 516823 187241 516857
rect 187275 516823 187413 516857
rect 187447 516823 187465 516857
rect 187223 516776 187465 516823
rect 187223 516702 187327 516776
rect 187223 516668 187273 516702
rect 187307 516668 187327 516702
rect 187361 516708 187381 516742
rect 187415 516708 187465 516742
rect 187361 516634 187465 516708
rect 182531 516484 182589 516578
rect 182623 516579 183692 516593
rect 182623 516545 182641 516579
rect 182675 516545 183641 516579
rect 183675 516545 183692 516579
rect 182623 516484 183692 516545
rect 183727 516579 184796 516593
rect 183727 516545 183745 516579
rect 183779 516545 184745 516579
rect 184779 516545 184796 516579
rect 183727 516484 184796 516545
rect 184831 516579 185900 516593
rect 184831 516545 184849 516579
rect 184883 516545 185849 516579
rect 185883 516545 185900 516579
rect 184831 516484 185900 516545
rect 185935 516579 187004 516593
rect 185935 516545 185953 516579
rect 185987 516545 186953 516579
rect 186987 516545 187004 516579
rect 185935 516484 187004 516545
rect 187223 516581 187465 516634
rect 187223 516547 187241 516581
rect 187275 516547 187413 516581
rect 187447 516547 187465 516581
rect 187223 516484 187465 516547
rect 172210 516450 172239 516484
rect 172273 516450 172331 516484
rect 172365 516450 172423 516484
rect 172457 516450 172515 516484
rect 172549 516450 172607 516484
rect 172641 516450 172699 516484
rect 172733 516450 172791 516484
rect 172825 516450 172883 516484
rect 172917 516450 172975 516484
rect 173009 516450 173067 516484
rect 173101 516450 173159 516484
rect 173193 516450 173251 516484
rect 173285 516450 173343 516484
rect 173377 516450 173435 516484
rect 173469 516450 173527 516484
rect 173561 516450 173619 516484
rect 173653 516450 173711 516484
rect 173745 516450 173803 516484
rect 173837 516450 173895 516484
rect 173929 516450 173987 516484
rect 174021 516450 174079 516484
rect 174113 516450 174171 516484
rect 174205 516450 174263 516484
rect 174297 516450 174355 516484
rect 174389 516450 174447 516484
rect 174481 516450 174539 516484
rect 174573 516450 174631 516484
rect 174665 516450 174723 516484
rect 174757 516450 174815 516484
rect 174849 516450 174907 516484
rect 174941 516450 174999 516484
rect 175033 516450 175091 516484
rect 175125 516450 175183 516484
rect 175217 516450 175275 516484
rect 175309 516450 175367 516484
rect 175401 516450 175459 516484
rect 175493 516450 175551 516484
rect 175585 516450 175643 516484
rect 175677 516450 175735 516484
rect 175769 516450 175827 516484
rect 175861 516450 175919 516484
rect 175953 516450 176011 516484
rect 176045 516450 176103 516484
rect 176137 516450 176195 516484
rect 176229 516450 176287 516484
rect 176321 516450 176379 516484
rect 176413 516450 176471 516484
rect 176505 516450 176563 516484
rect 176597 516450 176655 516484
rect 176689 516450 176747 516484
rect 176781 516450 176839 516484
rect 176873 516450 176931 516484
rect 176965 516450 177023 516484
rect 177057 516450 177115 516484
rect 177149 516450 177207 516484
rect 177241 516450 177299 516484
rect 177333 516450 177391 516484
rect 177425 516450 177483 516484
rect 177517 516450 177575 516484
rect 177609 516450 177667 516484
rect 177701 516450 177759 516484
rect 177793 516450 177851 516484
rect 177885 516450 177943 516484
rect 177977 516450 178035 516484
rect 178069 516450 178127 516484
rect 178161 516450 178219 516484
rect 178253 516450 178311 516484
rect 178345 516450 178403 516484
rect 178437 516450 178495 516484
rect 178529 516450 178587 516484
rect 178621 516450 178679 516484
rect 178713 516450 178771 516484
rect 178805 516450 178863 516484
rect 178897 516450 178955 516484
rect 178989 516450 179047 516484
rect 179081 516450 179139 516484
rect 179173 516450 179231 516484
rect 179265 516450 179323 516484
rect 179357 516450 179415 516484
rect 179449 516450 179507 516484
rect 179541 516450 179599 516484
rect 179633 516450 179691 516484
rect 179725 516450 179783 516484
rect 179817 516450 179875 516484
rect 179909 516450 179967 516484
rect 180001 516450 180059 516484
rect 180093 516450 180151 516484
rect 180185 516450 180243 516484
rect 180277 516450 180335 516484
rect 180369 516450 180427 516484
rect 180461 516450 180519 516484
rect 180553 516450 180611 516484
rect 180645 516450 180703 516484
rect 180737 516450 180795 516484
rect 180829 516450 180887 516484
rect 180921 516450 180979 516484
rect 181013 516450 181071 516484
rect 181105 516450 181163 516484
rect 181197 516450 181255 516484
rect 181289 516450 181347 516484
rect 181381 516450 181439 516484
rect 181473 516450 181531 516484
rect 181565 516450 181623 516484
rect 181657 516450 181715 516484
rect 181749 516450 181807 516484
rect 181841 516450 181899 516484
rect 181933 516450 181991 516484
rect 182025 516450 182083 516484
rect 182117 516450 182175 516484
rect 182209 516450 182267 516484
rect 182301 516450 182359 516484
rect 182393 516450 182451 516484
rect 182485 516450 182543 516484
rect 182577 516450 182635 516484
rect 182669 516450 182727 516484
rect 182761 516450 182819 516484
rect 182853 516450 182911 516484
rect 182945 516450 183003 516484
rect 183037 516450 183095 516484
rect 183129 516450 183187 516484
rect 183221 516450 183279 516484
rect 183313 516450 183371 516484
rect 183405 516450 183463 516484
rect 183497 516450 183555 516484
rect 183589 516450 183647 516484
rect 183681 516450 183739 516484
rect 183773 516450 183831 516484
rect 183865 516450 183923 516484
rect 183957 516450 184015 516484
rect 184049 516450 184107 516484
rect 184141 516450 184199 516484
rect 184233 516450 184291 516484
rect 184325 516450 184383 516484
rect 184417 516450 184475 516484
rect 184509 516450 184567 516484
rect 184601 516450 184659 516484
rect 184693 516450 184751 516484
rect 184785 516450 184843 516484
rect 184877 516450 184935 516484
rect 184969 516450 185027 516484
rect 185061 516450 185119 516484
rect 185153 516450 185211 516484
rect 185245 516450 185303 516484
rect 185337 516450 185395 516484
rect 185429 516450 185487 516484
rect 185521 516450 185579 516484
rect 185613 516450 185671 516484
rect 185705 516450 185763 516484
rect 185797 516450 185855 516484
rect 185889 516450 185947 516484
rect 185981 516450 186039 516484
rect 186073 516450 186131 516484
rect 186165 516450 186223 516484
rect 186257 516450 186315 516484
rect 186349 516450 186407 516484
rect 186441 516450 186499 516484
rect 186533 516450 186591 516484
rect 186625 516450 186683 516484
rect 186717 516450 186775 516484
rect 186809 516450 186867 516484
rect 186901 516450 186959 516484
rect 186993 516450 187051 516484
rect 187085 516450 187143 516484
rect 187177 516450 187235 516484
rect 187269 516450 187327 516484
rect 187361 516450 187419 516484
rect 187453 516450 187482 516484
rect 172227 516387 172469 516450
rect 172227 516353 172245 516387
rect 172279 516353 172417 516387
rect 172451 516353 172469 516387
rect 172227 516300 172469 516353
rect 172503 516389 173572 516450
rect 172503 516355 172521 516389
rect 172555 516355 173521 516389
rect 173555 516355 173572 516389
rect 172503 516341 173572 516355
rect 173607 516389 174676 516450
rect 173607 516355 173625 516389
rect 173659 516355 174625 516389
rect 174659 516355 174676 516389
rect 173607 516341 174676 516355
rect 174803 516356 174861 516450
rect 172227 516226 172331 516300
rect 172227 516192 172277 516226
rect 172311 516192 172331 516226
rect 172365 516232 172385 516266
rect 172419 516232 172469 516266
rect 172365 516158 172469 516232
rect 172820 516226 172888 516341
rect 172820 516192 172837 516226
rect 172871 516192 172888 516226
rect 172820 516175 172888 516192
rect 173184 516262 173254 516277
rect 173184 516228 173201 516262
rect 173235 516228 173254 516262
rect 172227 516111 172469 516158
rect 172227 516077 172245 516111
rect 172279 516077 172417 516111
rect 172451 516077 172469 516111
rect 172227 516016 172469 516077
rect 173184 516027 173254 516228
rect 173924 516226 173992 516341
rect 174803 516322 174815 516356
rect 174849 516322 174861 516356
rect 174895 516389 175964 516450
rect 174895 516355 174913 516389
rect 174947 516355 175913 516389
rect 175947 516355 175964 516389
rect 174895 516341 175964 516355
rect 175999 516389 177068 516450
rect 175999 516355 176017 516389
rect 176051 516355 177017 516389
rect 177051 516355 177068 516389
rect 175999 516341 177068 516355
rect 177103 516389 178172 516450
rect 177103 516355 177121 516389
rect 177155 516355 178121 516389
rect 178155 516355 178172 516389
rect 177103 516341 178172 516355
rect 178207 516389 179276 516450
rect 178207 516355 178225 516389
rect 178259 516355 179225 516389
rect 179259 516355 179276 516389
rect 178207 516341 179276 516355
rect 179311 516389 179829 516450
rect 179311 516355 179329 516389
rect 179363 516355 179777 516389
rect 179811 516355 179829 516389
rect 174803 516305 174861 516322
rect 173924 516192 173941 516226
rect 173975 516192 173992 516226
rect 173924 516175 173992 516192
rect 174288 516262 174358 516277
rect 174288 516228 174305 516262
rect 174339 516228 174358 516262
rect 174288 516027 174358 516228
rect 175212 516226 175280 516341
rect 175212 516192 175229 516226
rect 175263 516192 175280 516226
rect 175212 516175 175280 516192
rect 175576 516262 175646 516277
rect 175576 516228 175593 516262
rect 175627 516228 175646 516262
rect 174803 516138 174861 516173
rect 174803 516104 174815 516138
rect 174849 516104 174861 516138
rect 174803 516045 174861 516104
rect 172227 515982 172245 516016
rect 172279 515982 172417 516016
rect 172451 515982 172469 516016
rect 172227 515940 172469 515982
rect 172503 516016 173572 516027
rect 172503 515982 172521 516016
rect 172555 515982 173521 516016
rect 173555 515982 173572 516016
rect 172503 515940 173572 515982
rect 173607 516016 174676 516027
rect 173607 515982 173625 516016
rect 173659 515982 174625 516016
rect 174659 515982 174676 516016
rect 173607 515940 174676 515982
rect 174803 516011 174815 516045
rect 174849 516011 174861 516045
rect 175576 516027 175646 516228
rect 176316 516226 176384 516341
rect 176316 516192 176333 516226
rect 176367 516192 176384 516226
rect 176316 516175 176384 516192
rect 176680 516262 176750 516277
rect 176680 516228 176697 516262
rect 176731 516228 176750 516262
rect 176680 516027 176750 516228
rect 177420 516226 177488 516341
rect 177420 516192 177437 516226
rect 177471 516192 177488 516226
rect 177420 516175 177488 516192
rect 177784 516262 177854 516277
rect 177784 516228 177801 516262
rect 177835 516228 177854 516262
rect 177784 516027 177854 516228
rect 178524 516226 178592 516341
rect 179311 516296 179829 516355
rect 179955 516356 180013 516450
rect 179955 516322 179967 516356
rect 180001 516322 180013 516356
rect 180047 516389 181116 516450
rect 180047 516355 180065 516389
rect 180099 516355 181065 516389
rect 181099 516355 181116 516389
rect 180047 516341 181116 516355
rect 181151 516389 182220 516450
rect 181151 516355 181169 516389
rect 181203 516355 182169 516389
rect 182203 516355 182220 516389
rect 181151 516341 182220 516355
rect 182255 516389 183324 516450
rect 182255 516355 182273 516389
rect 182307 516355 183273 516389
rect 183307 516355 183324 516389
rect 182255 516341 183324 516355
rect 183359 516389 184428 516450
rect 183359 516355 183377 516389
rect 183411 516355 184377 516389
rect 184411 516355 184428 516389
rect 183359 516341 184428 516355
rect 184463 516389 184981 516450
rect 184463 516355 184481 516389
rect 184515 516355 184929 516389
rect 184963 516355 184981 516389
rect 179955 516305 180013 516322
rect 178524 516192 178541 516226
rect 178575 516192 178592 516226
rect 178524 516175 178592 516192
rect 178888 516262 178958 516277
rect 178888 516228 178905 516262
rect 178939 516228 178958 516262
rect 178888 516027 178958 516228
rect 179311 516226 179553 516296
rect 179311 516192 179389 516226
rect 179423 516192 179499 516226
rect 179533 516192 179553 516226
rect 179587 516228 179607 516262
rect 179641 516228 179717 516262
rect 179751 516228 179829 516262
rect 179587 516158 179829 516228
rect 180364 516226 180432 516341
rect 180364 516192 180381 516226
rect 180415 516192 180432 516226
rect 180364 516175 180432 516192
rect 180728 516262 180798 516277
rect 180728 516228 180745 516262
rect 180779 516228 180798 516262
rect 179311 516118 179829 516158
rect 179311 516084 179329 516118
rect 179363 516084 179777 516118
rect 179811 516084 179829 516118
rect 174803 515940 174861 516011
rect 174895 516016 175964 516027
rect 174895 515982 174913 516016
rect 174947 515982 175913 516016
rect 175947 515982 175964 516016
rect 174895 515940 175964 515982
rect 175999 516016 177068 516027
rect 175999 515982 176017 516016
rect 176051 515982 177017 516016
rect 177051 515982 177068 516016
rect 175999 515940 177068 515982
rect 177103 516016 178172 516027
rect 177103 515982 177121 516016
rect 177155 515982 178121 516016
rect 178155 515982 178172 516016
rect 177103 515940 178172 515982
rect 178207 516016 179276 516027
rect 178207 515982 178225 516016
rect 178259 515982 179225 516016
rect 179259 515982 179276 516016
rect 178207 515940 179276 515982
rect 179311 516016 179829 516084
rect 179311 515982 179329 516016
rect 179363 515982 179777 516016
rect 179811 515982 179829 516016
rect 179311 515940 179829 515982
rect 179955 516138 180013 516173
rect 179955 516104 179967 516138
rect 180001 516104 180013 516138
rect 179955 516045 180013 516104
rect 179955 516011 179967 516045
rect 180001 516011 180013 516045
rect 180728 516027 180798 516228
rect 181468 516226 181536 516341
rect 181468 516192 181485 516226
rect 181519 516192 181536 516226
rect 181468 516175 181536 516192
rect 181832 516262 181902 516277
rect 181832 516228 181849 516262
rect 181883 516228 181902 516262
rect 181832 516027 181902 516228
rect 182572 516226 182640 516341
rect 182572 516192 182589 516226
rect 182623 516192 182640 516226
rect 182572 516175 182640 516192
rect 182936 516262 183006 516277
rect 182936 516228 182953 516262
rect 182987 516228 183006 516262
rect 182936 516027 183006 516228
rect 183676 516226 183744 516341
rect 184463 516296 184981 516355
rect 185107 516356 185165 516450
rect 185107 516322 185119 516356
rect 185153 516322 185165 516356
rect 185199 516389 186268 516450
rect 185199 516355 185217 516389
rect 185251 516355 186217 516389
rect 186251 516355 186268 516389
rect 185199 516341 186268 516355
rect 186303 516389 187005 516450
rect 186303 516355 186321 516389
rect 186355 516355 186953 516389
rect 186987 516355 187005 516389
rect 185107 516305 185165 516322
rect 183676 516192 183693 516226
rect 183727 516192 183744 516226
rect 183676 516175 183744 516192
rect 184040 516262 184110 516277
rect 184040 516228 184057 516262
rect 184091 516228 184110 516262
rect 184040 516027 184110 516228
rect 184463 516226 184705 516296
rect 184463 516192 184541 516226
rect 184575 516192 184651 516226
rect 184685 516192 184705 516226
rect 184739 516228 184759 516262
rect 184793 516228 184869 516262
rect 184903 516228 184981 516262
rect 184739 516158 184981 516228
rect 185516 516226 185584 516341
rect 186303 516296 187005 516355
rect 187223 516387 187465 516450
rect 187223 516353 187241 516387
rect 187275 516353 187413 516387
rect 187447 516353 187465 516387
rect 187223 516300 187465 516353
rect 185516 516192 185533 516226
rect 185567 516192 185584 516226
rect 185516 516175 185584 516192
rect 185880 516262 185950 516277
rect 185880 516228 185897 516262
rect 185931 516228 185950 516262
rect 184463 516118 184981 516158
rect 184463 516084 184481 516118
rect 184515 516084 184929 516118
rect 184963 516084 184981 516118
rect 179955 515940 180013 516011
rect 180047 516016 181116 516027
rect 180047 515982 180065 516016
rect 180099 515982 181065 516016
rect 181099 515982 181116 516016
rect 180047 515940 181116 515982
rect 181151 516016 182220 516027
rect 181151 515982 181169 516016
rect 181203 515982 182169 516016
rect 182203 515982 182220 516016
rect 181151 515940 182220 515982
rect 182255 516016 183324 516027
rect 182255 515982 182273 516016
rect 182307 515982 183273 516016
rect 183307 515982 183324 516016
rect 182255 515940 183324 515982
rect 183359 516016 184428 516027
rect 183359 515982 183377 516016
rect 183411 515982 184377 516016
rect 184411 515982 184428 516016
rect 183359 515940 184428 515982
rect 184463 516016 184981 516084
rect 184463 515982 184481 516016
rect 184515 515982 184929 516016
rect 184963 515982 184981 516016
rect 184463 515940 184981 515982
rect 185107 516138 185165 516173
rect 185107 516104 185119 516138
rect 185153 516104 185165 516138
rect 185107 516045 185165 516104
rect 185107 516011 185119 516045
rect 185153 516011 185165 516045
rect 185880 516027 185950 516228
rect 186303 516226 186633 516296
rect 186303 516192 186381 516226
rect 186415 516192 186480 516226
rect 186514 516192 186579 516226
rect 186613 516192 186633 516226
rect 186667 516228 186687 516262
rect 186721 516228 186790 516262
rect 186824 516228 186893 516262
rect 186927 516228 187005 516262
rect 186667 516158 187005 516228
rect 186303 516118 187005 516158
rect 186303 516084 186321 516118
rect 186355 516084 186953 516118
rect 186987 516084 187005 516118
rect 185107 515940 185165 516011
rect 185199 516016 186268 516027
rect 185199 515982 185217 516016
rect 185251 515982 186217 516016
rect 186251 515982 186268 516016
rect 185199 515940 186268 515982
rect 186303 516016 187005 516084
rect 186303 515982 186321 516016
rect 186355 515982 186953 516016
rect 186987 515982 187005 516016
rect 186303 515940 187005 515982
rect 187223 516232 187273 516266
rect 187307 516232 187327 516266
rect 187223 516158 187327 516232
rect 187361 516226 187465 516300
rect 187361 516192 187381 516226
rect 187415 516192 187465 516226
rect 187223 516111 187465 516158
rect 187223 516077 187241 516111
rect 187275 516077 187413 516111
rect 187447 516077 187465 516111
rect 187223 516016 187465 516077
rect 187223 515982 187241 516016
rect 187275 515982 187413 516016
rect 187447 515982 187465 516016
rect 187223 515940 187465 515982
rect 172210 515906 172239 515940
rect 172273 515906 172331 515940
rect 172365 515906 172423 515940
rect 172457 515906 172515 515940
rect 172549 515906 172607 515940
rect 172641 515906 172699 515940
rect 172733 515906 172791 515940
rect 172825 515906 172883 515940
rect 172917 515906 172975 515940
rect 173009 515906 173067 515940
rect 173101 515906 173159 515940
rect 173193 515906 173251 515940
rect 173285 515906 173343 515940
rect 173377 515906 173435 515940
rect 173469 515906 173527 515940
rect 173561 515906 173619 515940
rect 173653 515906 173711 515940
rect 173745 515906 173803 515940
rect 173837 515906 173895 515940
rect 173929 515906 173987 515940
rect 174021 515906 174079 515940
rect 174113 515906 174171 515940
rect 174205 515906 174263 515940
rect 174297 515906 174355 515940
rect 174389 515906 174447 515940
rect 174481 515906 174539 515940
rect 174573 515906 174631 515940
rect 174665 515906 174723 515940
rect 174757 515906 174815 515940
rect 174849 515906 174907 515940
rect 174941 515906 174999 515940
rect 175033 515906 175091 515940
rect 175125 515906 175183 515940
rect 175217 515906 175275 515940
rect 175309 515906 175367 515940
rect 175401 515906 175459 515940
rect 175493 515906 175551 515940
rect 175585 515906 175643 515940
rect 175677 515906 175735 515940
rect 175769 515906 175827 515940
rect 175861 515906 175919 515940
rect 175953 515906 176011 515940
rect 176045 515906 176103 515940
rect 176137 515906 176195 515940
rect 176229 515906 176287 515940
rect 176321 515906 176379 515940
rect 176413 515906 176471 515940
rect 176505 515906 176563 515940
rect 176597 515906 176655 515940
rect 176689 515906 176747 515940
rect 176781 515906 176839 515940
rect 176873 515906 176931 515940
rect 176965 515906 177023 515940
rect 177057 515906 177115 515940
rect 177149 515906 177207 515940
rect 177241 515906 177299 515940
rect 177333 515906 177391 515940
rect 177425 515906 177483 515940
rect 177517 515906 177575 515940
rect 177609 515906 177667 515940
rect 177701 515906 177759 515940
rect 177793 515906 177851 515940
rect 177885 515906 177943 515940
rect 177977 515906 178035 515940
rect 178069 515906 178127 515940
rect 178161 515906 178219 515940
rect 178253 515906 178311 515940
rect 178345 515906 178403 515940
rect 178437 515906 178495 515940
rect 178529 515906 178587 515940
rect 178621 515906 178679 515940
rect 178713 515906 178771 515940
rect 178805 515906 178863 515940
rect 178897 515906 178955 515940
rect 178989 515906 179047 515940
rect 179081 515906 179139 515940
rect 179173 515906 179231 515940
rect 179265 515906 179323 515940
rect 179357 515906 179415 515940
rect 179449 515906 179507 515940
rect 179541 515906 179599 515940
rect 179633 515906 179691 515940
rect 179725 515906 179783 515940
rect 179817 515906 179875 515940
rect 179909 515906 179967 515940
rect 180001 515906 180059 515940
rect 180093 515906 180151 515940
rect 180185 515906 180243 515940
rect 180277 515906 180335 515940
rect 180369 515906 180427 515940
rect 180461 515906 180519 515940
rect 180553 515906 180611 515940
rect 180645 515906 180703 515940
rect 180737 515906 180795 515940
rect 180829 515906 180887 515940
rect 180921 515906 180979 515940
rect 181013 515906 181071 515940
rect 181105 515906 181163 515940
rect 181197 515906 181255 515940
rect 181289 515906 181347 515940
rect 181381 515906 181439 515940
rect 181473 515906 181531 515940
rect 181565 515906 181623 515940
rect 181657 515906 181715 515940
rect 181749 515906 181807 515940
rect 181841 515906 181899 515940
rect 181933 515906 181991 515940
rect 182025 515906 182083 515940
rect 182117 515906 182175 515940
rect 182209 515906 182267 515940
rect 182301 515906 182359 515940
rect 182393 515906 182451 515940
rect 182485 515906 182543 515940
rect 182577 515906 182635 515940
rect 182669 515906 182727 515940
rect 182761 515906 182819 515940
rect 182853 515906 182911 515940
rect 182945 515906 183003 515940
rect 183037 515906 183095 515940
rect 183129 515906 183187 515940
rect 183221 515906 183279 515940
rect 183313 515906 183371 515940
rect 183405 515906 183463 515940
rect 183497 515906 183555 515940
rect 183589 515906 183647 515940
rect 183681 515906 183739 515940
rect 183773 515906 183831 515940
rect 183865 515906 183923 515940
rect 183957 515906 184015 515940
rect 184049 515906 184107 515940
rect 184141 515906 184199 515940
rect 184233 515906 184291 515940
rect 184325 515906 184383 515940
rect 184417 515906 184475 515940
rect 184509 515906 184567 515940
rect 184601 515906 184659 515940
rect 184693 515906 184751 515940
rect 184785 515906 184843 515940
rect 184877 515906 184935 515940
rect 184969 515906 185027 515940
rect 185061 515906 185119 515940
rect 185153 515906 185211 515940
rect 185245 515906 185303 515940
rect 185337 515906 185395 515940
rect 185429 515906 185487 515940
rect 185521 515906 185579 515940
rect 185613 515906 185671 515940
rect 185705 515906 185763 515940
rect 185797 515906 185855 515940
rect 185889 515906 185947 515940
rect 185981 515906 186039 515940
rect 186073 515906 186131 515940
rect 186165 515906 186223 515940
rect 186257 515906 186315 515940
rect 186349 515906 186407 515940
rect 186441 515906 186499 515940
rect 186533 515906 186591 515940
rect 186625 515906 186683 515940
rect 186717 515906 186775 515940
rect 186809 515906 186867 515940
rect 186901 515906 186959 515940
rect 186993 515906 187051 515940
rect 187085 515906 187143 515940
rect 187177 515906 187235 515940
rect 187269 515906 187327 515940
rect 187361 515906 187419 515940
rect 187453 515906 187482 515940
rect 172227 515864 172469 515906
rect 172227 515830 172245 515864
rect 172279 515830 172417 515864
rect 172451 515830 172469 515864
rect 172227 515769 172469 515830
rect 172227 515735 172245 515769
rect 172279 515735 172417 515769
rect 172451 515735 172469 515769
rect 172227 515688 172469 515735
rect 172503 515864 173205 515906
rect 172503 515830 172521 515864
rect 172555 515830 173153 515864
rect 173187 515830 173205 515864
rect 172503 515762 173205 515830
rect 172503 515728 172521 515762
rect 172555 515728 173153 515762
rect 173187 515728 173205 515762
rect 172503 515688 173205 515728
rect 172227 515620 172277 515654
rect 172311 515620 172331 515654
rect 172227 515546 172331 515620
rect 172365 515614 172469 515688
rect 172365 515580 172385 515614
rect 172419 515580 172469 515614
rect 172503 515620 172581 515654
rect 172615 515620 172680 515654
rect 172714 515620 172779 515654
rect 172813 515620 172833 515654
rect 172503 515550 172833 515620
rect 172867 515618 173205 515688
rect 172867 515584 172887 515618
rect 172921 515584 172990 515618
rect 173024 515584 173093 515618
rect 173127 515584 173205 515618
rect 173423 515856 173485 515872
rect 173423 515822 173441 515856
rect 173475 515822 173485 515856
rect 173423 515734 173485 515822
rect 173519 515864 173581 515906
rect 173519 515830 173527 515864
rect 173561 515830 173581 515864
rect 173519 515796 173581 515830
rect 173519 515762 173527 515796
rect 173561 515762 173581 515796
rect 173519 515746 173581 515762
rect 173615 515838 173667 515872
rect 173615 515804 173619 515838
rect 173653 515829 173667 515838
rect 173615 515795 173623 515804
rect 173657 515795 173667 515829
rect 173701 515864 173752 515906
rect 173701 515830 173709 515864
rect 173743 515830 173752 515864
rect 173701 515814 173752 515830
rect 173787 515856 173839 515872
rect 173787 515822 173795 515856
rect 173829 515822 173839 515856
rect 173615 515780 173667 515795
rect 173787 515788 173839 515822
rect 173787 515780 173795 515788
rect 173615 515754 173795 515780
rect 173829 515754 173839 515788
rect 173615 515746 173839 515754
rect 173423 515700 173441 515734
rect 173475 515712 173485 515734
rect 173787 515720 173839 515746
rect 173873 515850 173930 515906
rect 173873 515816 173881 515850
rect 173915 515816 173930 515850
rect 173873 515782 173930 515816
rect 173873 515748 173881 515782
rect 173915 515748 173930 515782
rect 173873 515732 173930 515748
rect 173975 515864 174677 515906
rect 173975 515830 173993 515864
rect 174027 515830 174625 515864
rect 174659 515830 174677 515864
rect 173975 515762 174677 515830
rect 173475 515700 173629 515712
rect 173423 515678 173629 515700
rect 172227 515493 172469 515546
rect 172227 515459 172245 515493
rect 172279 515459 172417 515493
rect 172451 515459 172469 515493
rect 172227 515396 172469 515459
rect 172503 515491 173205 515550
rect 172503 515457 172521 515491
rect 172555 515457 173153 515491
rect 173187 515457 173205 515491
rect 172503 515396 173205 515457
rect 173423 515496 173457 515678
rect 173491 515628 173561 515644
rect 173525 515594 173561 515628
rect 173595 515628 173629 515678
rect 173787 515686 173795 515720
rect 173829 515696 173839 515720
rect 173975 515728 173993 515762
rect 174027 515728 174625 515762
rect 174659 515728 174677 515762
rect 173829 515686 173938 515696
rect 173975 515688 174677 515728
rect 173787 515662 173938 515686
rect 173595 515594 173637 515628
rect 173671 515594 173705 515628
rect 173739 515594 173773 515628
rect 173807 515594 173823 515628
rect 173491 515566 173561 515594
rect 173491 515532 173527 515566
rect 173857 515560 173938 515662
rect 173491 515530 173561 515532
rect 173608 515526 173938 515560
rect 173975 515620 174053 515654
rect 174087 515620 174152 515654
rect 174186 515620 174251 515654
rect 174285 515620 174305 515654
rect 173975 515550 174305 515620
rect 174339 515618 174677 515688
rect 174803 515835 174861 515906
rect 174803 515801 174815 515835
rect 174849 515801 174861 515835
rect 174895 515864 175964 515906
rect 174895 515830 174913 515864
rect 174947 515830 175913 515864
rect 175947 515830 175964 515864
rect 174895 515819 175964 515830
rect 175999 515864 177068 515906
rect 175999 515830 176017 515864
rect 176051 515830 177017 515864
rect 177051 515830 177068 515864
rect 175999 515819 177068 515830
rect 177103 515864 177345 515906
rect 177103 515830 177121 515864
rect 177155 515830 177293 515864
rect 177327 515830 177345 515864
rect 174803 515742 174861 515801
rect 174803 515708 174815 515742
rect 174849 515708 174861 515742
rect 174803 515673 174861 515708
rect 174339 515584 174359 515618
rect 174393 515584 174462 515618
rect 174496 515584 174565 515618
rect 174599 515584 174677 515618
rect 175212 515654 175280 515671
rect 175212 515620 175229 515654
rect 175263 515620 175280 515654
rect 173608 515498 173667 515526
rect 173423 515480 173483 515496
rect 173423 515446 173441 515480
rect 173475 515446 173483 515480
rect 173423 515430 173483 515446
rect 173517 515476 173572 515492
rect 173517 515442 173527 515476
rect 173561 515442 173572 515476
rect 173608 515464 173624 515498
rect 173658 515464 173667 515498
rect 173787 515498 173839 515526
rect 173608 515448 173667 515464
rect 173701 515476 173752 515492
rect 173517 515396 173572 515442
rect 173701 515442 173710 515476
rect 173744 515442 173752 515476
rect 173787 515464 173796 515498
rect 173830 515464 173839 515498
rect 173787 515448 173839 515464
rect 173873 515476 173929 515492
rect 173701 515396 173752 515442
rect 173873 515442 173882 515476
rect 173916 515442 173929 515476
rect 173873 515396 173929 515442
rect 173975 515491 174677 515550
rect 173975 515457 173993 515491
rect 174027 515457 174625 515491
rect 174659 515457 174677 515491
rect 173975 515396 174677 515457
rect 174803 515524 174861 515541
rect 174803 515490 174815 515524
rect 174849 515490 174861 515524
rect 175212 515505 175280 515620
rect 175576 515618 175646 515819
rect 175576 515584 175593 515618
rect 175627 515584 175646 515618
rect 175576 515569 175646 515584
rect 176316 515654 176384 515671
rect 176316 515620 176333 515654
rect 176367 515620 176384 515654
rect 176316 515505 176384 515620
rect 176680 515618 176750 515819
rect 177103 515769 177345 515830
rect 177103 515735 177121 515769
rect 177155 515735 177293 515769
rect 177327 515735 177345 515769
rect 177103 515688 177345 515735
rect 176680 515584 176697 515618
rect 176731 515584 176750 515618
rect 176680 515569 176750 515584
rect 177103 515620 177153 515654
rect 177187 515620 177207 515654
rect 177103 515546 177207 515620
rect 177241 515614 177345 515688
rect 177379 515835 177437 515906
rect 177379 515801 177391 515835
rect 177425 515801 177437 515835
rect 177471 515864 178540 515906
rect 177471 515830 177489 515864
rect 177523 515830 178489 515864
rect 178523 515830 178540 515864
rect 177471 515819 178540 515830
rect 178575 515864 179644 515906
rect 178575 515830 178593 515864
rect 178627 515830 179593 515864
rect 179627 515830 179644 515864
rect 178575 515819 179644 515830
rect 179679 515864 179921 515906
rect 179679 515830 179697 515864
rect 179731 515830 179869 515864
rect 179903 515830 179921 515864
rect 177379 515742 177437 515801
rect 177379 515708 177391 515742
rect 177425 515708 177437 515742
rect 177379 515673 177437 515708
rect 177241 515580 177261 515614
rect 177295 515580 177345 515614
rect 177788 515654 177856 515671
rect 177788 515620 177805 515654
rect 177839 515620 177856 515654
rect 174803 515396 174861 515490
rect 174895 515491 175964 515505
rect 174895 515457 174913 515491
rect 174947 515457 175913 515491
rect 175947 515457 175964 515491
rect 174895 515396 175964 515457
rect 175999 515491 177068 515505
rect 175999 515457 176017 515491
rect 176051 515457 177017 515491
rect 177051 515457 177068 515491
rect 175999 515396 177068 515457
rect 177103 515493 177345 515546
rect 177103 515459 177121 515493
rect 177155 515459 177293 515493
rect 177327 515459 177345 515493
rect 177103 515396 177345 515459
rect 177379 515524 177437 515541
rect 177379 515490 177391 515524
rect 177425 515490 177437 515524
rect 177788 515505 177856 515620
rect 178152 515618 178222 515819
rect 178152 515584 178169 515618
rect 178203 515584 178222 515618
rect 178152 515569 178222 515584
rect 178892 515654 178960 515671
rect 178892 515620 178909 515654
rect 178943 515620 178960 515654
rect 178892 515505 178960 515620
rect 179256 515618 179326 515819
rect 179679 515769 179921 515830
rect 179679 515735 179697 515769
rect 179731 515735 179869 515769
rect 179903 515735 179921 515769
rect 179679 515688 179921 515735
rect 179256 515584 179273 515618
rect 179307 515584 179326 515618
rect 179256 515569 179326 515584
rect 179679 515620 179729 515654
rect 179763 515620 179783 515654
rect 179679 515546 179783 515620
rect 179817 515614 179921 515688
rect 179955 515835 180013 515906
rect 179955 515801 179967 515835
rect 180001 515801 180013 515835
rect 180047 515864 181116 515906
rect 180047 515830 180065 515864
rect 180099 515830 181065 515864
rect 181099 515830 181116 515864
rect 180047 515819 181116 515830
rect 181151 515864 181853 515906
rect 181151 515830 181169 515864
rect 181203 515830 181801 515864
rect 181835 515830 181853 515864
rect 179955 515742 180013 515801
rect 179955 515708 179967 515742
rect 180001 515708 180013 515742
rect 179955 515673 180013 515708
rect 179817 515580 179837 515614
rect 179871 515580 179921 515614
rect 180364 515654 180432 515671
rect 180364 515620 180381 515654
rect 180415 515620 180432 515654
rect 177379 515396 177437 515490
rect 177471 515491 178540 515505
rect 177471 515457 177489 515491
rect 177523 515457 178489 515491
rect 178523 515457 178540 515491
rect 177471 515396 178540 515457
rect 178575 515491 179644 515505
rect 178575 515457 178593 515491
rect 178627 515457 179593 515491
rect 179627 515457 179644 515491
rect 178575 515396 179644 515457
rect 179679 515493 179921 515546
rect 179679 515459 179697 515493
rect 179731 515459 179869 515493
rect 179903 515459 179921 515493
rect 179679 515396 179921 515459
rect 179955 515524 180013 515541
rect 179955 515490 179967 515524
rect 180001 515490 180013 515524
rect 180364 515505 180432 515620
rect 180728 515618 180798 515819
rect 181151 515762 181853 515830
rect 181151 515728 181169 515762
rect 181203 515728 181801 515762
rect 181835 515728 181853 515762
rect 181151 515688 181853 515728
rect 180728 515584 180745 515618
rect 180779 515584 180798 515618
rect 180728 515569 180798 515584
rect 181151 515620 181229 515654
rect 181263 515620 181328 515654
rect 181362 515620 181427 515654
rect 181461 515620 181481 515654
rect 181151 515550 181481 515620
rect 181515 515618 181853 515688
rect 181515 515584 181535 515618
rect 181569 515584 181638 515618
rect 181672 515584 181741 515618
rect 181775 515584 181853 515618
rect 182071 515856 182125 515872
rect 182071 515838 182089 515856
rect 182071 515804 182083 515838
rect 182123 515822 182125 515856
rect 182117 515804 182125 515822
rect 182071 515775 182125 515804
rect 182071 515741 182089 515775
rect 182123 515741 182125 515775
rect 182159 515856 182225 515906
rect 182159 515822 182175 515856
rect 182209 515822 182225 515856
rect 182159 515788 182225 515822
rect 182159 515754 182175 515788
rect 182209 515754 182225 515788
rect 182261 515856 182297 515872
rect 182295 515822 182297 515856
rect 182261 515788 182297 515822
rect 182295 515754 182297 515788
rect 182071 515691 182125 515741
rect 182261 515720 182297 515754
rect 179955 515396 180013 515490
rect 180047 515491 181116 515505
rect 180047 515457 180065 515491
rect 180099 515457 181065 515491
rect 181099 515457 181116 515491
rect 180047 515396 181116 515457
rect 181151 515491 181853 515550
rect 181151 515457 181169 515491
rect 181203 515457 181801 515491
rect 181835 515457 181853 515491
rect 181151 515396 181853 515457
rect 182071 515531 182107 515691
rect 182162 515686 182297 515720
rect 182531 515835 182589 515906
rect 182531 515801 182543 515835
rect 182577 515801 182589 515835
rect 182623 515864 183692 515906
rect 182623 515830 182641 515864
rect 182675 515830 183641 515864
rect 183675 515830 183692 515864
rect 182623 515819 183692 515830
rect 183727 515864 184796 515906
rect 183727 515830 183745 515864
rect 183779 515830 184745 515864
rect 184779 515830 184796 515864
rect 183727 515819 184796 515830
rect 184831 515864 185073 515906
rect 184831 515830 184849 515864
rect 184883 515830 185021 515864
rect 185055 515830 185073 515864
rect 182531 515742 182589 515801
rect 182531 515708 182543 515742
rect 182577 515708 182589 515742
rect 182162 515657 182196 515686
rect 182531 515673 182589 515708
rect 182141 515641 182196 515657
rect 182940 515654 183008 515671
rect 182175 515607 182196 515641
rect 182141 515591 182196 515607
rect 182162 515540 182196 515591
rect 182241 515634 182309 515650
rect 182241 515628 182267 515634
rect 182241 515594 182259 515628
rect 182301 515600 182309 515634
rect 182293 515594 182309 515600
rect 182241 515576 182309 515594
rect 182940 515620 182957 515654
rect 182991 515620 183008 515654
rect 182071 515502 182123 515531
rect 182162 515506 182295 515540
rect 182071 515468 182089 515502
rect 182261 515485 182295 515506
rect 182071 515430 182123 515468
rect 182159 515438 182175 515472
rect 182209 515438 182225 515472
rect 182159 515396 182225 515438
rect 182261 515430 182295 515451
rect 182531 515524 182589 515541
rect 182531 515490 182543 515524
rect 182577 515490 182589 515524
rect 182940 515505 183008 515620
rect 183304 515618 183374 515819
rect 183304 515584 183321 515618
rect 183355 515584 183374 515618
rect 183304 515569 183374 515584
rect 184044 515654 184112 515671
rect 184044 515620 184061 515654
rect 184095 515620 184112 515654
rect 184044 515505 184112 515620
rect 184408 515618 184478 515819
rect 184831 515769 185073 515830
rect 184831 515735 184849 515769
rect 184883 515735 185021 515769
rect 185055 515735 185073 515769
rect 184831 515688 185073 515735
rect 184408 515584 184425 515618
rect 184459 515584 184478 515618
rect 184408 515569 184478 515584
rect 184831 515620 184881 515654
rect 184915 515620 184935 515654
rect 184831 515546 184935 515620
rect 184969 515614 185073 515688
rect 185107 515835 185165 515906
rect 185107 515801 185119 515835
rect 185153 515801 185165 515835
rect 185199 515864 186268 515906
rect 185199 515830 185217 515864
rect 185251 515830 186217 515864
rect 186251 515830 186268 515864
rect 185199 515819 186268 515830
rect 186395 515856 186457 515872
rect 186395 515822 186413 515856
rect 186447 515822 186457 515856
rect 185107 515742 185165 515801
rect 185107 515708 185119 515742
rect 185153 515708 185165 515742
rect 185107 515673 185165 515708
rect 184969 515580 184989 515614
rect 185023 515580 185073 515614
rect 185516 515654 185584 515671
rect 185516 515620 185533 515654
rect 185567 515620 185584 515654
rect 182531 515396 182589 515490
rect 182623 515491 183692 515505
rect 182623 515457 182641 515491
rect 182675 515457 183641 515491
rect 183675 515457 183692 515491
rect 182623 515396 183692 515457
rect 183727 515491 184796 515505
rect 183727 515457 183745 515491
rect 183779 515457 184745 515491
rect 184779 515457 184796 515491
rect 183727 515396 184796 515457
rect 184831 515493 185073 515546
rect 184831 515459 184849 515493
rect 184883 515459 185021 515493
rect 185055 515459 185073 515493
rect 184831 515396 185073 515459
rect 185107 515524 185165 515541
rect 185107 515490 185119 515524
rect 185153 515490 185165 515524
rect 185516 515505 185584 515620
rect 185880 515618 185950 515819
rect 185880 515584 185897 515618
rect 185931 515584 185950 515618
rect 185880 515569 185950 515584
rect 186395 515734 186457 515822
rect 186491 515864 186553 515906
rect 186491 515830 186499 515864
rect 186533 515830 186553 515864
rect 186491 515796 186553 515830
rect 186491 515762 186499 515796
rect 186533 515762 186553 515796
rect 186491 515746 186553 515762
rect 186587 515838 186639 515872
rect 186587 515804 186591 515838
rect 186625 515829 186639 515838
rect 186587 515795 186595 515804
rect 186629 515795 186639 515829
rect 186673 515864 186724 515906
rect 186673 515830 186681 515864
rect 186715 515830 186724 515864
rect 186673 515814 186724 515830
rect 186759 515856 186811 515872
rect 186759 515822 186767 515856
rect 186801 515822 186811 515856
rect 186587 515780 186639 515795
rect 186759 515788 186811 515822
rect 186759 515780 186767 515788
rect 186587 515754 186767 515780
rect 186801 515754 186811 515788
rect 186587 515746 186811 515754
rect 186395 515700 186413 515734
rect 186447 515712 186457 515734
rect 186759 515720 186811 515746
rect 186845 515850 186902 515906
rect 186845 515816 186853 515850
rect 186887 515816 186902 515850
rect 186845 515782 186902 515816
rect 186845 515748 186853 515782
rect 186887 515748 186902 515782
rect 186845 515732 186902 515748
rect 186947 515864 187189 515906
rect 186947 515830 186965 515864
rect 186999 515830 187137 515864
rect 187171 515830 187189 515864
rect 186947 515769 187189 515830
rect 186947 515735 186965 515769
rect 186999 515735 187137 515769
rect 187171 515735 187189 515769
rect 186447 515700 186601 515712
rect 186395 515678 186601 515700
rect 185107 515396 185165 515490
rect 185199 515491 186268 515505
rect 185199 515457 185217 515491
rect 185251 515457 186217 515491
rect 186251 515457 186268 515491
rect 185199 515396 186268 515457
rect 186395 515496 186429 515678
rect 186463 515628 186533 515644
rect 186497 515594 186533 515628
rect 186567 515628 186601 515678
rect 186759 515686 186767 515720
rect 186801 515696 186811 515720
rect 186801 515686 186910 515696
rect 186947 515688 187189 515735
rect 186759 515662 186910 515686
rect 186567 515594 186609 515628
rect 186643 515594 186677 515628
rect 186711 515594 186745 515628
rect 186779 515594 186795 515628
rect 186463 515566 186533 515594
rect 186463 515532 186499 515566
rect 186829 515560 186910 515662
rect 186463 515530 186533 515532
rect 186580 515526 186910 515560
rect 186947 515620 186997 515654
rect 187031 515620 187051 515654
rect 186947 515546 187051 515620
rect 187085 515614 187189 515688
rect 187085 515580 187105 515614
rect 187139 515580 187189 515614
rect 187223 515864 187465 515906
rect 187223 515830 187241 515864
rect 187275 515830 187413 515864
rect 187447 515830 187465 515864
rect 187223 515769 187465 515830
rect 187223 515735 187241 515769
rect 187275 515735 187413 515769
rect 187447 515735 187465 515769
rect 187223 515688 187465 515735
rect 187223 515614 187327 515688
rect 187223 515580 187273 515614
rect 187307 515580 187327 515614
rect 187361 515620 187381 515654
rect 187415 515620 187465 515654
rect 187361 515546 187465 515620
rect 186580 515498 186639 515526
rect 186395 515480 186455 515496
rect 186395 515446 186413 515480
rect 186447 515446 186455 515480
rect 186395 515430 186455 515446
rect 186489 515476 186544 515492
rect 186489 515442 186499 515476
rect 186533 515442 186544 515476
rect 186580 515464 186596 515498
rect 186630 515464 186639 515498
rect 186759 515498 186811 515526
rect 186580 515448 186639 515464
rect 186673 515476 186724 515492
rect 186489 515396 186544 515442
rect 186673 515442 186682 515476
rect 186716 515442 186724 515476
rect 186759 515464 186768 515498
rect 186802 515464 186811 515498
rect 186947 515493 187189 515546
rect 186759 515448 186811 515464
rect 186845 515476 186901 515492
rect 186673 515396 186724 515442
rect 186845 515442 186854 515476
rect 186888 515442 186901 515476
rect 186845 515396 186901 515442
rect 186947 515459 186965 515493
rect 186999 515459 187137 515493
rect 187171 515459 187189 515493
rect 186947 515396 187189 515459
rect 187223 515493 187465 515546
rect 187223 515459 187241 515493
rect 187275 515459 187413 515493
rect 187447 515459 187465 515493
rect 187223 515396 187465 515459
rect 172210 515362 172239 515396
rect 172273 515362 172331 515396
rect 172365 515362 172423 515396
rect 172457 515362 172515 515396
rect 172549 515362 172607 515396
rect 172641 515362 172699 515396
rect 172733 515362 172791 515396
rect 172825 515362 172883 515396
rect 172917 515362 172975 515396
rect 173009 515362 173067 515396
rect 173101 515362 173159 515396
rect 173193 515362 173251 515396
rect 173285 515362 173343 515396
rect 173377 515362 173435 515396
rect 173469 515362 173527 515396
rect 173561 515362 173619 515396
rect 173653 515362 173711 515396
rect 173745 515362 173803 515396
rect 173837 515362 173895 515396
rect 173929 515362 173987 515396
rect 174021 515362 174079 515396
rect 174113 515362 174171 515396
rect 174205 515362 174263 515396
rect 174297 515362 174355 515396
rect 174389 515362 174447 515396
rect 174481 515362 174539 515396
rect 174573 515362 174631 515396
rect 174665 515362 174723 515396
rect 174757 515362 174815 515396
rect 174849 515362 174907 515396
rect 174941 515362 174999 515396
rect 175033 515362 175091 515396
rect 175125 515362 175183 515396
rect 175217 515362 175275 515396
rect 175309 515362 175367 515396
rect 175401 515362 175459 515396
rect 175493 515362 175551 515396
rect 175585 515362 175643 515396
rect 175677 515362 175735 515396
rect 175769 515362 175827 515396
rect 175861 515362 175919 515396
rect 175953 515362 176011 515396
rect 176045 515362 176103 515396
rect 176137 515362 176195 515396
rect 176229 515362 176287 515396
rect 176321 515362 176379 515396
rect 176413 515362 176471 515396
rect 176505 515362 176563 515396
rect 176597 515362 176655 515396
rect 176689 515362 176747 515396
rect 176781 515362 176839 515396
rect 176873 515362 176931 515396
rect 176965 515362 177023 515396
rect 177057 515362 177115 515396
rect 177149 515362 177207 515396
rect 177241 515362 177299 515396
rect 177333 515362 177391 515396
rect 177425 515362 177483 515396
rect 177517 515362 177575 515396
rect 177609 515362 177667 515396
rect 177701 515362 177759 515396
rect 177793 515362 177851 515396
rect 177885 515362 177943 515396
rect 177977 515362 178035 515396
rect 178069 515362 178127 515396
rect 178161 515362 178219 515396
rect 178253 515362 178311 515396
rect 178345 515362 178403 515396
rect 178437 515362 178495 515396
rect 178529 515362 178587 515396
rect 178621 515362 178679 515396
rect 178713 515362 178771 515396
rect 178805 515362 178863 515396
rect 178897 515362 178955 515396
rect 178989 515362 179047 515396
rect 179081 515362 179139 515396
rect 179173 515362 179231 515396
rect 179265 515362 179323 515396
rect 179357 515362 179415 515396
rect 179449 515362 179507 515396
rect 179541 515362 179599 515396
rect 179633 515362 179691 515396
rect 179725 515362 179783 515396
rect 179817 515362 179875 515396
rect 179909 515362 179967 515396
rect 180001 515362 180059 515396
rect 180093 515362 180151 515396
rect 180185 515362 180243 515396
rect 180277 515362 180335 515396
rect 180369 515362 180427 515396
rect 180461 515362 180519 515396
rect 180553 515362 180611 515396
rect 180645 515362 180703 515396
rect 180737 515362 180795 515396
rect 180829 515362 180887 515396
rect 180921 515362 180979 515396
rect 181013 515362 181071 515396
rect 181105 515362 181163 515396
rect 181197 515362 181255 515396
rect 181289 515362 181347 515396
rect 181381 515362 181439 515396
rect 181473 515362 181531 515396
rect 181565 515362 181623 515396
rect 181657 515362 181715 515396
rect 181749 515362 181807 515396
rect 181841 515362 181899 515396
rect 181933 515362 181991 515396
rect 182025 515362 182083 515396
rect 182117 515362 182175 515396
rect 182209 515362 182267 515396
rect 182301 515362 182359 515396
rect 182393 515362 182451 515396
rect 182485 515362 182543 515396
rect 182577 515362 182635 515396
rect 182669 515362 182727 515396
rect 182761 515362 182819 515396
rect 182853 515362 182911 515396
rect 182945 515362 183003 515396
rect 183037 515362 183095 515396
rect 183129 515362 183187 515396
rect 183221 515362 183279 515396
rect 183313 515362 183371 515396
rect 183405 515362 183463 515396
rect 183497 515362 183555 515396
rect 183589 515362 183647 515396
rect 183681 515362 183739 515396
rect 183773 515362 183831 515396
rect 183865 515362 183923 515396
rect 183957 515362 184015 515396
rect 184049 515362 184107 515396
rect 184141 515362 184199 515396
rect 184233 515362 184291 515396
rect 184325 515362 184383 515396
rect 184417 515362 184475 515396
rect 184509 515362 184567 515396
rect 184601 515362 184659 515396
rect 184693 515362 184751 515396
rect 184785 515362 184843 515396
rect 184877 515362 184935 515396
rect 184969 515362 185027 515396
rect 185061 515362 185119 515396
rect 185153 515362 185211 515396
rect 185245 515362 185303 515396
rect 185337 515362 185395 515396
rect 185429 515362 185487 515396
rect 185521 515362 185579 515396
rect 185613 515362 185671 515396
rect 185705 515362 185763 515396
rect 185797 515362 185855 515396
rect 185889 515362 185947 515396
rect 185981 515362 186039 515396
rect 186073 515362 186131 515396
rect 186165 515362 186223 515396
rect 186257 515362 186315 515396
rect 186349 515362 186407 515396
rect 186441 515362 186499 515396
rect 186533 515362 186591 515396
rect 186625 515362 186683 515396
rect 186717 515362 186775 515396
rect 186809 515362 186867 515396
rect 186901 515362 186959 515396
rect 186993 515362 187051 515396
rect 187085 515362 187143 515396
rect 187177 515362 187235 515396
rect 187269 515362 187327 515396
rect 187361 515362 187419 515396
rect 187453 515362 187482 515396
<< viali >>
rect 164730 541117 164764 541151
rect 165033 541124 165067 541158
rect 165225 541124 165259 541158
rect 165417 541124 165451 541158
rect 165609 541124 165643 541158
rect 165801 541124 165835 541158
rect 165993 541124 166027 541158
rect 166410 541117 166444 541151
rect 164686 540562 164720 541050
rect 164774 540562 164808 541050
rect 164889 540115 164923 540603
rect 164985 540569 165019 541057
rect 165081 540115 165115 540603
rect 165177 540569 165211 541057
rect 165273 540115 165307 540603
rect 165369 540569 165403 541057
rect 165465 540115 165499 540603
rect 165561 540569 165595 541057
rect 165657 540115 165691 540603
rect 165753 540569 165787 541057
rect 165849 540115 165883 540603
rect 165945 540569 165979 541057
rect 166041 540115 166075 540603
rect 166210 540317 166244 540351
rect 166166 540091 166200 540267
rect 166254 540091 166288 540267
rect 166366 540108 166400 540596
rect 166454 540108 166488 540596
rect 166570 540117 166580 540247
rect 166580 540117 166620 540247
rect 166620 540117 166630 540247
rect 164730 540007 164764 540041
rect 164937 540014 164971 540048
rect 165129 540014 165163 540048
rect 165321 540014 165355 540048
rect 165513 540014 165547 540048
rect 165705 540014 165739 540048
rect 165897 540014 165931 540048
rect 166210 540007 166244 540041
rect 166410 540007 166444 540041
rect 168530 541117 168564 541151
rect 168833 541124 168867 541158
rect 169025 541124 169059 541158
rect 169217 541124 169251 541158
rect 169409 541124 169443 541158
rect 169601 541124 169635 541158
rect 169793 541124 169827 541158
rect 170210 541117 170244 541151
rect 168486 540562 168520 541050
rect 168574 540562 168608 541050
rect 168689 540115 168723 540603
rect 168785 540569 168819 541057
rect 168881 540115 168915 540603
rect 168977 540569 169011 541057
rect 169073 540115 169107 540603
rect 169169 540569 169203 541057
rect 169265 540115 169299 540603
rect 169361 540569 169395 541057
rect 169457 540115 169491 540603
rect 169553 540569 169587 541057
rect 169649 540115 169683 540603
rect 169745 540569 169779 541057
rect 169841 540115 169875 540603
rect 170010 540317 170044 540351
rect 169966 540091 170000 540267
rect 170054 540091 170088 540267
rect 170166 540108 170200 540596
rect 170254 540108 170288 540596
rect 170370 540117 170380 540247
rect 170380 540117 170420 540247
rect 170420 540117 170430 540247
rect 168530 540007 168564 540041
rect 168737 540014 168771 540048
rect 168929 540014 168963 540048
rect 169121 540014 169155 540048
rect 169313 540014 169347 540048
rect 169505 540014 169539 540048
rect 169697 540014 169731 540048
rect 170010 540007 170044 540041
rect 170210 540007 170244 540041
rect 172230 541117 172264 541151
rect 172533 541124 172567 541158
rect 172725 541124 172759 541158
rect 172917 541124 172951 541158
rect 173109 541124 173143 541158
rect 173301 541124 173335 541158
rect 173493 541124 173527 541158
rect 173910 541117 173944 541151
rect 172186 540562 172220 541050
rect 172274 540562 172308 541050
rect 172389 540115 172423 540603
rect 172485 540569 172519 541057
rect 172581 540115 172615 540603
rect 172677 540569 172711 541057
rect 172773 540115 172807 540603
rect 172869 540569 172903 541057
rect 172965 540115 172999 540603
rect 173061 540569 173095 541057
rect 173157 540115 173191 540603
rect 173253 540569 173287 541057
rect 173349 540115 173383 540603
rect 173445 540569 173479 541057
rect 173541 540115 173575 540603
rect 173710 540317 173744 540351
rect 173666 540091 173700 540267
rect 173754 540091 173788 540267
rect 173866 540108 173900 540596
rect 173954 540108 173988 540596
rect 174070 540117 174080 540247
rect 174080 540117 174120 540247
rect 174120 540117 174130 540247
rect 172230 540007 172264 540041
rect 172437 540014 172471 540048
rect 172629 540014 172663 540048
rect 172821 540014 172855 540048
rect 173013 540014 173047 540048
rect 173205 540014 173239 540048
rect 173397 540014 173431 540048
rect 173710 540007 173744 540041
rect 173910 540007 173944 540041
rect 175730 541117 175764 541151
rect 176033 541124 176067 541158
rect 176225 541124 176259 541158
rect 176417 541124 176451 541158
rect 176609 541124 176643 541158
rect 176801 541124 176835 541158
rect 176993 541124 177027 541158
rect 177410 541117 177444 541151
rect 175686 540562 175720 541050
rect 175774 540562 175808 541050
rect 175889 540115 175923 540603
rect 175985 540569 176019 541057
rect 176081 540115 176115 540603
rect 176177 540569 176211 541057
rect 176273 540115 176307 540603
rect 176369 540569 176403 541057
rect 176465 540115 176499 540603
rect 176561 540569 176595 541057
rect 176657 540115 176691 540603
rect 176753 540569 176787 541057
rect 176849 540115 176883 540603
rect 176945 540569 176979 541057
rect 177041 540115 177075 540603
rect 177210 540317 177244 540351
rect 177166 540091 177200 540267
rect 177254 540091 177288 540267
rect 177366 540108 177400 540596
rect 177454 540108 177488 540596
rect 177570 540117 177580 540247
rect 177580 540117 177620 540247
rect 177620 540117 177630 540247
rect 175730 540007 175764 540041
rect 175937 540014 175971 540048
rect 176129 540014 176163 540048
rect 176321 540014 176355 540048
rect 176513 540014 176547 540048
rect 176705 540014 176739 540048
rect 176897 540014 176931 540048
rect 177210 540007 177244 540041
rect 177410 540007 177444 540041
rect 179330 541117 179364 541151
rect 179633 541124 179667 541158
rect 179825 541124 179859 541158
rect 180017 541124 180051 541158
rect 180209 541124 180243 541158
rect 180401 541124 180435 541158
rect 180593 541124 180627 541158
rect 181010 541117 181044 541151
rect 179286 540562 179320 541050
rect 179374 540562 179408 541050
rect 179489 540115 179523 540603
rect 179585 540569 179619 541057
rect 179681 540115 179715 540603
rect 179777 540569 179811 541057
rect 179873 540115 179907 540603
rect 179969 540569 180003 541057
rect 180065 540115 180099 540603
rect 180161 540569 180195 541057
rect 180257 540115 180291 540603
rect 180353 540569 180387 541057
rect 180449 540115 180483 540603
rect 180545 540569 180579 541057
rect 180641 540115 180675 540603
rect 180810 540317 180844 540351
rect 180766 540091 180800 540267
rect 180854 540091 180888 540267
rect 180966 540108 181000 540596
rect 181054 540108 181088 540596
rect 181170 540117 181180 540247
rect 181180 540117 181220 540247
rect 181220 540117 181230 540247
rect 179330 540007 179364 540041
rect 179537 540014 179571 540048
rect 179729 540014 179763 540048
rect 179921 540014 179955 540048
rect 180113 540014 180147 540048
rect 180305 540014 180339 540048
rect 180497 540014 180531 540048
rect 180810 540007 180844 540041
rect 181010 540007 181044 540041
rect 182630 541117 182664 541151
rect 182933 541124 182967 541158
rect 183125 541124 183159 541158
rect 183317 541124 183351 541158
rect 183509 541124 183543 541158
rect 183701 541124 183735 541158
rect 183893 541124 183927 541158
rect 184310 541117 184344 541151
rect 182586 540562 182620 541050
rect 182674 540562 182708 541050
rect 182789 540115 182823 540603
rect 182885 540569 182919 541057
rect 182981 540115 183015 540603
rect 183077 540569 183111 541057
rect 183173 540115 183207 540603
rect 183269 540569 183303 541057
rect 183365 540115 183399 540603
rect 183461 540569 183495 541057
rect 183557 540115 183591 540603
rect 183653 540569 183687 541057
rect 183749 540115 183783 540603
rect 183845 540569 183879 541057
rect 183941 540115 183975 540603
rect 184110 540317 184144 540351
rect 184066 540091 184100 540267
rect 184154 540091 184188 540267
rect 184266 540108 184300 540596
rect 184354 540108 184388 540596
rect 184470 540117 184480 540247
rect 184480 540117 184520 540247
rect 184520 540117 184530 540247
rect 182630 540007 182664 540041
rect 182837 540014 182871 540048
rect 183029 540014 183063 540048
rect 183221 540014 183255 540048
rect 183413 540014 183447 540048
rect 183605 540014 183639 540048
rect 183797 540014 183831 540048
rect 184110 540007 184144 540041
rect 184310 540007 184344 540041
rect 185930 541117 185964 541151
rect 186233 541124 186267 541158
rect 186425 541124 186459 541158
rect 186617 541124 186651 541158
rect 186809 541124 186843 541158
rect 187001 541124 187035 541158
rect 187193 541124 187227 541158
rect 187610 541117 187644 541151
rect 185886 540562 185920 541050
rect 185974 540562 186008 541050
rect 186089 540115 186123 540603
rect 186185 540569 186219 541057
rect 186281 540115 186315 540603
rect 186377 540569 186411 541057
rect 186473 540115 186507 540603
rect 186569 540569 186603 541057
rect 186665 540115 186699 540603
rect 186761 540569 186795 541057
rect 186857 540115 186891 540603
rect 186953 540569 186987 541057
rect 187049 540115 187083 540603
rect 187145 540569 187179 541057
rect 187241 540115 187275 540603
rect 187410 540317 187444 540351
rect 187366 540091 187400 540267
rect 187454 540091 187488 540267
rect 187566 540108 187600 540596
rect 187654 540108 187688 540596
rect 187770 540117 187780 540247
rect 187780 540117 187820 540247
rect 187820 540117 187830 540247
rect 185930 540007 185964 540041
rect 186137 540014 186171 540048
rect 186329 540014 186363 540048
rect 186521 540014 186555 540048
rect 186713 540014 186747 540048
rect 186905 540014 186939 540048
rect 187097 540014 187131 540048
rect 187410 540007 187444 540041
rect 187610 540007 187644 540041
rect 189230 541117 189264 541151
rect 189533 541124 189567 541158
rect 189725 541124 189759 541158
rect 189917 541124 189951 541158
rect 190109 541124 190143 541158
rect 190301 541124 190335 541158
rect 190493 541124 190527 541158
rect 190910 541117 190944 541151
rect 189186 540562 189220 541050
rect 189274 540562 189308 541050
rect 189389 540115 189423 540603
rect 189485 540569 189519 541057
rect 189581 540115 189615 540603
rect 189677 540569 189711 541057
rect 189773 540115 189807 540603
rect 189869 540569 189903 541057
rect 189965 540115 189999 540603
rect 190061 540569 190095 541057
rect 190157 540115 190191 540603
rect 190253 540569 190287 541057
rect 190349 540115 190383 540603
rect 190445 540569 190479 541057
rect 190541 540115 190575 540603
rect 190710 540317 190744 540351
rect 190666 540091 190700 540267
rect 190754 540091 190788 540267
rect 190866 540108 190900 540596
rect 190954 540108 190988 540596
rect 191070 540117 191080 540247
rect 191080 540117 191120 540247
rect 191120 540117 191130 540247
rect 189230 540007 189264 540041
rect 189437 540014 189471 540048
rect 189629 540014 189663 540048
rect 189821 540014 189855 540048
rect 190013 540014 190047 540048
rect 190205 540014 190239 540048
rect 190397 540014 190431 540048
rect 190710 540007 190744 540041
rect 190910 540007 190944 540041
rect 191810 540097 191990 540277
rect 162270 538697 162530 538737
rect 158728 538467 158896 538501
rect 159104 538467 159272 538501
rect 159362 538467 159530 538501
rect 159620 538467 159788 538501
rect 159878 538467 160046 538501
rect 160136 538467 160304 538501
rect 160394 538467 160562 538501
rect 160652 538467 160820 538501
rect 160910 538467 161078 538501
rect 161168 538467 161336 538501
rect 161548 538467 161716 538501
rect 161948 538467 162116 538501
rect 162328 538467 162496 538501
rect 158666 538241 158700 538417
rect 158924 538241 158958 538417
rect 159042 538312 159076 538400
rect 159300 538258 159334 538346
rect 159558 538312 159592 538400
rect 159816 538258 159850 538346
rect 160074 538312 160108 538400
rect 160332 538258 160366 538346
rect 160590 538312 160624 538400
rect 160848 538258 160882 538346
rect 161106 538312 161140 538400
rect 161364 538258 161398 538346
rect 161486 538241 161520 538417
rect 161744 538241 161778 538417
rect 161886 538241 161920 538417
rect 162144 538241 162178 538417
rect 162266 538241 162300 538417
rect 162524 538241 162558 538417
rect 158728 538157 158896 538191
rect 159104 538157 159272 538191
rect 159362 538157 159530 538191
rect 159620 538157 159788 538191
rect 159878 538157 160046 538191
rect 160136 538157 160304 538191
rect 160394 538157 160562 538191
rect 160652 538157 160820 538191
rect 160910 538157 161078 538191
rect 161168 538157 161336 538191
rect 161548 538157 161716 538191
rect 161948 538157 162116 538191
rect 162328 538157 162496 538191
rect 164714 539604 164748 539638
rect 165037 539611 165071 539645
rect 165229 539611 165263 539645
rect 165421 539611 165455 539645
rect 165613 539611 165647 539645
rect 165805 539611 165839 539645
rect 165997 539611 166031 539645
rect 166214 539604 166248 539638
rect 166414 539604 166448 539638
rect 164670 538569 164704 539545
rect 164758 538569 164792 539545
rect 164893 538593 164927 539081
rect 164989 539047 165023 539535
rect 165085 538593 165119 539081
rect 165181 539047 165215 539535
rect 165277 538593 165311 539081
rect 165373 539047 165407 539535
rect 165469 538593 165503 539081
rect 165565 539047 165599 539535
rect 165661 538593 165695 539081
rect 165757 539047 165791 539535
rect 165853 538593 165887 539081
rect 165949 539047 165983 539535
rect 166045 538593 166079 539081
rect 166170 538969 166204 539545
rect 166258 538969 166292 539545
rect 166214 538876 166248 538910
rect 166370 538586 166404 539074
rect 166458 538586 166492 539074
rect 166570 539207 166580 539297
rect 166580 539207 166620 539297
rect 164714 538476 164748 538510
rect 164941 538483 164975 538517
rect 165133 538483 165167 538517
rect 165325 538483 165359 538517
rect 165517 538483 165551 538517
rect 165709 538483 165743 538517
rect 165901 538483 165935 538517
rect 166414 538476 166448 538510
rect 168514 539604 168548 539638
rect 168837 539611 168871 539645
rect 169029 539611 169063 539645
rect 169221 539611 169255 539645
rect 169413 539611 169447 539645
rect 169605 539611 169639 539645
rect 169797 539611 169831 539645
rect 170014 539604 170048 539638
rect 170214 539604 170248 539638
rect 168470 538569 168504 539545
rect 168558 538569 168592 539545
rect 168693 538593 168727 539081
rect 168789 539047 168823 539535
rect 168885 538593 168919 539081
rect 168981 539047 169015 539535
rect 169077 538593 169111 539081
rect 169173 539047 169207 539535
rect 169269 538593 169303 539081
rect 169365 539047 169399 539535
rect 169461 538593 169495 539081
rect 169557 539047 169591 539535
rect 169653 538593 169687 539081
rect 169749 539047 169783 539535
rect 169845 538593 169879 539081
rect 169970 538969 170004 539545
rect 170058 538969 170092 539545
rect 170014 538876 170048 538910
rect 170170 538586 170204 539074
rect 170258 538586 170292 539074
rect 170370 539207 170380 539297
rect 170380 539207 170420 539297
rect 168514 538476 168548 538510
rect 168741 538483 168775 538517
rect 168933 538483 168967 538517
rect 169125 538483 169159 538517
rect 169317 538483 169351 538517
rect 169509 538483 169543 538517
rect 169701 538483 169735 538517
rect 170214 538476 170248 538510
rect 172214 539604 172248 539638
rect 172537 539611 172571 539645
rect 172729 539611 172763 539645
rect 172921 539611 172955 539645
rect 173113 539611 173147 539645
rect 173305 539611 173339 539645
rect 173497 539611 173531 539645
rect 173714 539604 173748 539638
rect 173914 539604 173948 539638
rect 172170 538569 172204 539545
rect 172258 538569 172292 539545
rect 172393 538593 172427 539081
rect 172489 539047 172523 539535
rect 172585 538593 172619 539081
rect 172681 539047 172715 539535
rect 172777 538593 172811 539081
rect 172873 539047 172907 539535
rect 172969 538593 173003 539081
rect 173065 539047 173099 539535
rect 173161 538593 173195 539081
rect 173257 539047 173291 539535
rect 173353 538593 173387 539081
rect 173449 539047 173483 539535
rect 173545 538593 173579 539081
rect 173670 538969 173704 539545
rect 173758 538969 173792 539545
rect 173714 538876 173748 538910
rect 173870 538586 173904 539074
rect 173958 538586 173992 539074
rect 174070 539207 174080 539297
rect 174080 539207 174120 539297
rect 172214 538476 172248 538510
rect 172441 538483 172475 538517
rect 172633 538483 172667 538517
rect 172825 538483 172859 538517
rect 173017 538483 173051 538517
rect 173209 538483 173243 538517
rect 173401 538483 173435 538517
rect 173914 538476 173948 538510
rect 175714 539604 175748 539638
rect 176037 539611 176071 539645
rect 176229 539611 176263 539645
rect 176421 539611 176455 539645
rect 176613 539611 176647 539645
rect 176805 539611 176839 539645
rect 176997 539611 177031 539645
rect 177214 539604 177248 539638
rect 177414 539604 177448 539638
rect 175670 538569 175704 539545
rect 175758 538569 175792 539545
rect 175893 538593 175927 539081
rect 175989 539047 176023 539535
rect 176085 538593 176119 539081
rect 176181 539047 176215 539535
rect 176277 538593 176311 539081
rect 176373 539047 176407 539535
rect 176469 538593 176503 539081
rect 176565 539047 176599 539535
rect 176661 538593 176695 539081
rect 176757 539047 176791 539535
rect 176853 538593 176887 539081
rect 176949 539047 176983 539535
rect 177045 538593 177079 539081
rect 177170 538969 177204 539545
rect 177258 538969 177292 539545
rect 177214 538876 177248 538910
rect 177370 538586 177404 539074
rect 177458 538586 177492 539074
rect 177570 539207 177580 539297
rect 177580 539207 177620 539297
rect 175714 538476 175748 538510
rect 175941 538483 175975 538517
rect 176133 538483 176167 538517
rect 176325 538483 176359 538517
rect 176517 538483 176551 538517
rect 176709 538483 176743 538517
rect 176901 538483 176935 538517
rect 177414 538476 177448 538510
rect 179314 539604 179348 539638
rect 179637 539611 179671 539645
rect 179829 539611 179863 539645
rect 180021 539611 180055 539645
rect 180213 539611 180247 539645
rect 180405 539611 180439 539645
rect 180597 539611 180631 539645
rect 180814 539604 180848 539638
rect 181014 539604 181048 539638
rect 179270 538569 179304 539545
rect 179358 538569 179392 539545
rect 179493 538593 179527 539081
rect 179589 539047 179623 539535
rect 179685 538593 179719 539081
rect 179781 539047 179815 539535
rect 179877 538593 179911 539081
rect 179973 539047 180007 539535
rect 180069 538593 180103 539081
rect 180165 539047 180199 539535
rect 180261 538593 180295 539081
rect 180357 539047 180391 539535
rect 180453 538593 180487 539081
rect 180549 539047 180583 539535
rect 180645 538593 180679 539081
rect 180770 538969 180804 539545
rect 180858 538969 180892 539545
rect 180814 538876 180848 538910
rect 180970 538586 181004 539074
rect 181058 538586 181092 539074
rect 181170 539207 181180 539297
rect 181180 539207 181220 539297
rect 179314 538476 179348 538510
rect 179541 538483 179575 538517
rect 179733 538483 179767 538517
rect 179925 538483 179959 538517
rect 180117 538483 180151 538517
rect 180309 538483 180343 538517
rect 180501 538483 180535 538517
rect 181014 538476 181048 538510
rect 182614 539604 182648 539638
rect 182937 539611 182971 539645
rect 183129 539611 183163 539645
rect 183321 539611 183355 539645
rect 183513 539611 183547 539645
rect 183705 539611 183739 539645
rect 183897 539611 183931 539645
rect 184114 539604 184148 539638
rect 184314 539604 184348 539638
rect 182570 538569 182604 539545
rect 182658 538569 182692 539545
rect 182793 538593 182827 539081
rect 182889 539047 182923 539535
rect 182985 538593 183019 539081
rect 183081 539047 183115 539535
rect 183177 538593 183211 539081
rect 183273 539047 183307 539535
rect 183369 538593 183403 539081
rect 183465 539047 183499 539535
rect 183561 538593 183595 539081
rect 183657 539047 183691 539535
rect 183753 538593 183787 539081
rect 183849 539047 183883 539535
rect 183945 538593 183979 539081
rect 184070 538969 184104 539545
rect 184158 538969 184192 539545
rect 184114 538876 184148 538910
rect 184270 538586 184304 539074
rect 184358 538586 184392 539074
rect 184470 539207 184480 539297
rect 184480 539207 184520 539297
rect 182614 538476 182648 538510
rect 182841 538483 182875 538517
rect 183033 538483 183067 538517
rect 183225 538483 183259 538517
rect 183417 538483 183451 538517
rect 183609 538483 183643 538517
rect 183801 538483 183835 538517
rect 184314 538476 184348 538510
rect 185914 539604 185948 539638
rect 186237 539611 186271 539645
rect 186429 539611 186463 539645
rect 186621 539611 186655 539645
rect 186813 539611 186847 539645
rect 187005 539611 187039 539645
rect 187197 539611 187231 539645
rect 187414 539604 187448 539638
rect 187614 539604 187648 539638
rect 185870 538569 185904 539545
rect 185958 538569 185992 539545
rect 186093 538593 186127 539081
rect 186189 539047 186223 539535
rect 186285 538593 186319 539081
rect 186381 539047 186415 539535
rect 186477 538593 186511 539081
rect 186573 539047 186607 539535
rect 186669 538593 186703 539081
rect 186765 539047 186799 539535
rect 186861 538593 186895 539081
rect 186957 539047 186991 539535
rect 187053 538593 187087 539081
rect 187149 539047 187183 539535
rect 187245 538593 187279 539081
rect 187370 538969 187404 539545
rect 187458 538969 187492 539545
rect 187414 538876 187448 538910
rect 187570 538586 187604 539074
rect 187658 538586 187692 539074
rect 187770 539207 187780 539297
rect 187780 539207 187820 539297
rect 185914 538476 185948 538510
rect 186141 538483 186175 538517
rect 186333 538483 186367 538517
rect 186525 538483 186559 538517
rect 186717 538483 186751 538517
rect 186909 538483 186943 538517
rect 187101 538483 187135 538517
rect 187614 538476 187648 538510
rect 189214 539604 189248 539638
rect 189537 539611 189571 539645
rect 189729 539611 189763 539645
rect 189921 539611 189955 539645
rect 190113 539611 190147 539645
rect 190305 539611 190339 539645
rect 190497 539611 190531 539645
rect 190714 539604 190748 539638
rect 190914 539604 190948 539638
rect 189170 538569 189204 539545
rect 189258 538569 189292 539545
rect 189393 538593 189427 539081
rect 189489 539047 189523 539535
rect 189585 538593 189619 539081
rect 189681 539047 189715 539535
rect 189777 538593 189811 539081
rect 189873 539047 189907 539535
rect 189969 538593 190003 539081
rect 190065 539047 190099 539535
rect 190161 538593 190195 539081
rect 190257 539047 190291 539535
rect 190353 538593 190387 539081
rect 190449 539047 190483 539535
rect 190545 538593 190579 539081
rect 190670 538969 190704 539545
rect 190758 538969 190792 539545
rect 190714 538876 190748 538910
rect 190870 538586 190904 539074
rect 190958 538586 190992 539074
rect 191070 539207 191080 539297
rect 191080 539207 191120 539297
rect 189214 538476 189248 538510
rect 189441 538483 189475 538517
rect 189633 538483 189667 538517
rect 189825 538483 189859 538517
rect 190017 538483 190051 538517
rect 190209 538483 190243 538517
rect 190401 538483 190435 538517
rect 190914 538476 190948 538510
rect 161304 537704 161338 537738
rect 161508 537704 161542 537738
rect 161700 537704 161734 537738
rect 161908 537704 161942 537738
rect 162100 537704 162134 537738
rect 162324 537704 162358 537738
rect 161260 537086 161294 537374
rect 161348 537086 161382 537374
rect 161460 537086 161494 537374
rect 161556 537340 161590 537628
rect 161652 537086 161686 537374
rect 161748 537340 161782 537628
rect 161860 537340 161894 537628
rect 161956 537086 161990 537374
rect 162052 537340 162086 537628
rect 162148 537086 162182 537374
rect 162280 537086 162314 537374
rect 162368 537086 162402 537374
rect 161304 536976 161338 537010
rect 161604 536976 161638 537010
rect 162004 536976 162038 537010
rect 162324 536976 162358 537010
rect 157812 536684 157980 536718
rect 158190 536684 158358 536718
rect 158448 536684 158616 536718
rect 158706 536684 158874 536718
rect 158964 536684 159132 536718
rect 159222 536684 159390 536718
rect 159480 536684 159648 536718
rect 159738 536684 159906 536718
rect 159996 536684 160164 536718
rect 160254 536684 160422 536718
rect 160512 536684 160680 536718
rect 160896 536684 161064 536718
rect 161154 536684 161322 536718
rect 161412 536684 161580 536718
rect 161794 536684 161962 536718
rect 162052 536684 162220 536718
rect 162432 536684 162600 536718
rect 157750 536049 157784 536625
rect 158008 536049 158042 536625
rect 158128 536066 158162 536354
rect 158386 536320 158420 536608
rect 158644 536066 158678 536354
rect 158902 536320 158936 536608
rect 159160 536066 159194 536354
rect 159418 536320 159452 536608
rect 159676 536066 159710 536354
rect 159934 536320 159968 536608
rect 160192 536066 160226 536354
rect 160450 536320 160484 536608
rect 160708 536066 160742 536354
rect 160834 536320 160868 536608
rect 161092 536066 161126 536354
rect 161350 536320 161384 536608
rect 161608 536066 161642 536354
rect 161732 536066 161766 536354
rect 161990 536320 162024 536608
rect 162248 536066 162282 536354
rect 162370 536049 162404 536625
rect 162628 536049 162662 536625
rect 157812 535956 157980 535990
rect 158190 535956 158358 535990
rect 158448 535956 158616 535990
rect 158706 535956 158874 535990
rect 158964 535956 159132 535990
rect 159222 535956 159390 535990
rect 159480 535956 159648 535990
rect 159738 535956 159906 535990
rect 159996 535956 160164 535990
rect 160254 535956 160422 535990
rect 160512 535956 160680 535990
rect 160896 535956 161064 535990
rect 161154 535956 161322 535990
rect 161412 535956 161580 535990
rect 161794 535956 161962 535990
rect 162052 535956 162220 535990
rect 162432 535956 162600 535990
rect 164334 537566 164372 537963
rect 164652 537566 164690 537963
rect 164970 537566 165008 537963
rect 165288 537566 165326 537963
rect 165606 537566 165644 537963
rect 165924 537566 165962 537963
rect 166242 537566 166280 537963
rect 166560 537566 166598 537963
rect 164334 536051 164372 536448
rect 164652 536051 164690 536448
rect 164970 536051 165008 536448
rect 165288 536051 165326 536448
rect 165606 536051 165644 536448
rect 165924 536051 165962 536448
rect 166242 536051 166280 536448
rect 166560 536051 166598 536448
rect 168106 537566 168144 537963
rect 168424 537566 168462 537963
rect 168742 537566 168780 537963
rect 169060 537566 169098 537963
rect 168106 536051 168144 536448
rect 168424 536051 168462 536448
rect 168742 536051 168780 536448
rect 169060 536051 169098 536448
rect 171842 537566 171880 537963
rect 172160 537566 172198 537963
rect 171842 536051 171880 536448
rect 172160 536051 172198 536448
rect 175360 537566 175398 537963
rect 175360 536051 175398 536448
rect 178960 537566 178998 537963
rect 178960 536611 178998 537008
rect 182260 537566 182298 537963
rect 182260 536891 182298 537288
rect 185560 537566 185598 537963
rect 185560 537031 185598 537428
rect 188860 537566 188898 537963
rect 188860 536935 188898 537332
rect 162050 535737 162650 535777
rect 164304 535226 164342 535623
rect 164622 535226 164660 535623
rect 164940 535226 164978 535623
rect 165258 535226 165296 535623
rect 165576 535226 165614 535623
rect 165894 535226 165932 535623
rect 166212 535226 166250 535623
rect 166530 535226 166568 535623
rect 164304 533711 164342 534108
rect 164622 533711 164660 534108
rect 164940 533711 164978 534108
rect 165258 533711 165296 534108
rect 165576 533711 165614 534108
rect 165894 533711 165932 534108
rect 166212 533711 166250 534108
rect 166530 533711 166568 534108
rect 172239 530594 172273 530628
rect 172331 530594 172365 530628
rect 172423 530594 172457 530628
rect 172515 530594 172549 530628
rect 172607 530594 172641 530628
rect 172699 530594 172733 530628
rect 172791 530594 172825 530628
rect 172883 530594 172917 530628
rect 172975 530594 173009 530628
rect 173067 530594 173101 530628
rect 173159 530594 173193 530628
rect 173251 530594 173285 530628
rect 173343 530594 173377 530628
rect 173435 530594 173469 530628
rect 173527 530594 173561 530628
rect 173619 530594 173653 530628
rect 173711 530594 173745 530628
rect 173803 530594 173837 530628
rect 173895 530594 173929 530628
rect 173987 530594 174021 530628
rect 174079 530594 174113 530628
rect 174171 530594 174205 530628
rect 174263 530594 174297 530628
rect 174355 530594 174389 530628
rect 174447 530594 174481 530628
rect 174539 530594 174573 530628
rect 174631 530594 174665 530628
rect 174723 530594 174757 530628
rect 174815 530594 174849 530628
rect 174907 530594 174941 530628
rect 174999 530594 175033 530628
rect 175091 530594 175125 530628
rect 175183 530594 175217 530628
rect 175275 530594 175309 530628
rect 175367 530594 175401 530628
rect 175459 530594 175493 530628
rect 175551 530594 175585 530628
rect 175643 530594 175677 530628
rect 175735 530594 175769 530628
rect 175827 530594 175861 530628
rect 175919 530594 175953 530628
rect 176011 530594 176045 530628
rect 176103 530594 176137 530628
rect 176195 530594 176229 530628
rect 176287 530594 176321 530628
rect 176379 530594 176413 530628
rect 176471 530594 176505 530628
rect 176563 530594 176597 530628
rect 176655 530594 176689 530628
rect 176747 530594 176781 530628
rect 176839 530594 176873 530628
rect 176931 530594 176965 530628
rect 177023 530594 177057 530628
rect 177115 530594 177149 530628
rect 177207 530594 177241 530628
rect 177299 530594 177333 530628
rect 177391 530594 177425 530628
rect 177483 530594 177517 530628
rect 177575 530594 177609 530628
rect 177667 530594 177701 530628
rect 177759 530594 177793 530628
rect 177851 530594 177885 530628
rect 177943 530594 177977 530628
rect 178035 530594 178069 530628
rect 178127 530594 178161 530628
rect 178219 530594 178253 530628
rect 178311 530594 178345 530628
rect 178403 530594 178437 530628
rect 178495 530594 178529 530628
rect 178587 530594 178621 530628
rect 178679 530594 178713 530628
rect 178771 530594 178805 530628
rect 178863 530594 178897 530628
rect 178955 530594 178989 530628
rect 179047 530594 179081 530628
rect 179139 530594 179173 530628
rect 179231 530594 179265 530628
rect 179323 530594 179357 530628
rect 179415 530594 179449 530628
rect 179507 530594 179541 530628
rect 179599 530594 179633 530628
rect 179691 530594 179725 530628
rect 179783 530594 179817 530628
rect 179875 530594 179909 530628
rect 179967 530594 180001 530628
rect 180059 530594 180093 530628
rect 180151 530594 180185 530628
rect 180243 530594 180277 530628
rect 180335 530594 180369 530628
rect 180427 530594 180461 530628
rect 180519 530594 180553 530628
rect 180611 530594 180645 530628
rect 180703 530594 180737 530628
rect 180795 530594 180829 530628
rect 180887 530594 180921 530628
rect 180979 530594 181013 530628
rect 181071 530594 181105 530628
rect 181163 530594 181197 530628
rect 181255 530594 181289 530628
rect 181347 530594 181381 530628
rect 181439 530594 181473 530628
rect 181531 530594 181565 530628
rect 181623 530594 181657 530628
rect 181715 530594 181749 530628
rect 181807 530594 181841 530628
rect 181899 530594 181933 530628
rect 181991 530594 182025 530628
rect 182083 530594 182117 530628
rect 182175 530594 182209 530628
rect 182267 530594 182301 530628
rect 182359 530594 182393 530628
rect 182451 530594 182485 530628
rect 182543 530594 182577 530628
rect 182635 530594 182669 530628
rect 182727 530594 182761 530628
rect 182819 530594 182853 530628
rect 182911 530594 182945 530628
rect 183003 530594 183037 530628
rect 183095 530594 183129 530628
rect 183187 530594 183221 530628
rect 183279 530594 183313 530628
rect 183371 530594 183405 530628
rect 183463 530594 183497 530628
rect 183555 530594 183589 530628
rect 183647 530594 183681 530628
rect 183739 530594 183773 530628
rect 183831 530594 183865 530628
rect 183923 530594 183957 530628
rect 184015 530594 184049 530628
rect 184107 530594 184141 530628
rect 184199 530594 184233 530628
rect 184291 530594 184325 530628
rect 184383 530594 184417 530628
rect 184475 530594 184509 530628
rect 184567 530594 184601 530628
rect 184659 530594 184693 530628
rect 184751 530594 184785 530628
rect 184843 530594 184877 530628
rect 184935 530594 184969 530628
rect 185027 530594 185061 530628
rect 185119 530594 185153 530628
rect 185211 530594 185245 530628
rect 185303 530594 185337 530628
rect 185395 530594 185429 530628
rect 185487 530594 185521 530628
rect 185579 530594 185613 530628
rect 185671 530594 185705 530628
rect 185763 530594 185797 530628
rect 185855 530594 185889 530628
rect 185947 530594 185981 530628
rect 186039 530594 186073 530628
rect 186131 530594 186165 530628
rect 186223 530594 186257 530628
rect 186315 530594 186349 530628
rect 186407 530594 186441 530628
rect 186499 530594 186533 530628
rect 186591 530594 186625 530628
rect 186683 530594 186717 530628
rect 186775 530594 186809 530628
rect 186867 530594 186901 530628
rect 186959 530594 186993 530628
rect 187051 530594 187085 530628
rect 187143 530594 187177 530628
rect 187235 530594 187269 530628
rect 187327 530594 187361 530628
rect 187419 530594 187453 530628
rect 172515 530424 172549 530458
rect 172883 530356 172917 530390
rect 174907 530424 174941 530458
rect 175275 530356 175309 530390
rect 175847 530424 175881 530458
rect 175907 530370 175925 530395
rect 175925 530370 175941 530395
rect 175907 530361 175941 530370
rect 175551 530288 175585 530322
rect 176123 530372 176131 530390
rect 176131 530372 176157 530390
rect 176123 530356 176157 530372
rect 176495 530442 176529 530458
rect 176495 530424 176505 530442
rect 176505 530424 176529 530442
rect 176567 530424 176601 530458
rect 176123 530246 176126 530254
rect 176126 530246 176157 530254
rect 176123 530220 176157 530246
rect 176839 530356 176873 530390
rect 176747 530220 176781 530254
rect 177023 530288 177057 530322
rect 177125 530236 177159 530254
rect 177125 530220 177159 530236
rect 177206 530381 177240 530390
rect 177206 530356 177228 530381
rect 177228 530356 177240 530381
rect 177299 530288 177333 530322
rect 177667 530152 177692 530186
rect 177692 530152 177701 530186
rect 178219 530288 178253 530322
rect 178771 530492 178778 530526
rect 178778 530492 178805 530526
rect 178587 530362 178613 530390
rect 178613 530362 178621 530390
rect 178587 530356 178621 530362
rect 179047 530356 179081 530390
rect 178403 530168 178437 530186
rect 178403 530152 178409 530168
rect 178409 530152 178437 530168
rect 179415 530492 179420 530526
rect 179420 530492 179449 530526
rect 179323 530356 179357 530390
rect 180243 530160 180277 530186
rect 180243 530152 180249 530160
rect 180249 530152 180277 530160
rect 180611 530356 180645 530390
rect 180703 530492 180737 530526
rect 180795 530288 180829 530322
rect 181255 530319 181289 530322
rect 181255 530288 181269 530319
rect 181269 530288 181289 530319
rect 181531 530356 181565 530390
rect 181439 530319 181473 530322
rect 181439 530288 181471 530319
rect 181471 530288 181473 530319
rect 181899 530228 181933 530254
rect 181899 530220 181927 530228
rect 181927 530220 181933 530228
rect 182083 530424 182117 530458
rect 182175 530161 182179 530186
rect 182179 530161 182209 530186
rect 182175 530152 182209 530161
rect 183279 530492 183284 530526
rect 183284 530492 183313 530526
rect 183187 530356 183221 530390
rect 185395 530492 185400 530526
rect 185400 530492 185429 530526
rect 185303 530424 185337 530458
rect 187143 530356 187177 530390
rect 172239 530050 172273 530084
rect 172331 530050 172365 530084
rect 172423 530050 172457 530084
rect 172515 530050 172549 530084
rect 172607 530050 172641 530084
rect 172699 530050 172733 530084
rect 172791 530050 172825 530084
rect 172883 530050 172917 530084
rect 172975 530050 173009 530084
rect 173067 530050 173101 530084
rect 173159 530050 173193 530084
rect 173251 530050 173285 530084
rect 173343 530050 173377 530084
rect 173435 530050 173469 530084
rect 173527 530050 173561 530084
rect 173619 530050 173653 530084
rect 173711 530050 173745 530084
rect 173803 530050 173837 530084
rect 173895 530050 173929 530084
rect 173987 530050 174021 530084
rect 174079 530050 174113 530084
rect 174171 530050 174205 530084
rect 174263 530050 174297 530084
rect 174355 530050 174389 530084
rect 174447 530050 174481 530084
rect 174539 530050 174573 530084
rect 174631 530050 174665 530084
rect 174723 530050 174757 530084
rect 174815 530050 174849 530084
rect 174907 530050 174941 530084
rect 174999 530050 175033 530084
rect 175091 530050 175125 530084
rect 175183 530050 175217 530084
rect 175275 530050 175309 530084
rect 175367 530050 175401 530084
rect 175459 530050 175493 530084
rect 175551 530050 175585 530084
rect 175643 530050 175677 530084
rect 175735 530050 175769 530084
rect 175827 530050 175861 530084
rect 175919 530050 175953 530084
rect 176011 530050 176045 530084
rect 176103 530050 176137 530084
rect 176195 530050 176229 530084
rect 176287 530050 176321 530084
rect 176379 530050 176413 530084
rect 176471 530050 176505 530084
rect 176563 530050 176597 530084
rect 176655 530050 176689 530084
rect 176747 530050 176781 530084
rect 176839 530050 176873 530084
rect 176931 530050 176965 530084
rect 177023 530050 177057 530084
rect 177115 530050 177149 530084
rect 177207 530050 177241 530084
rect 177299 530050 177333 530084
rect 177391 530050 177425 530084
rect 177483 530050 177517 530084
rect 177575 530050 177609 530084
rect 177667 530050 177701 530084
rect 177759 530050 177793 530084
rect 177851 530050 177885 530084
rect 177943 530050 177977 530084
rect 178035 530050 178069 530084
rect 178127 530050 178161 530084
rect 178219 530050 178253 530084
rect 178311 530050 178345 530084
rect 178403 530050 178437 530084
rect 178495 530050 178529 530084
rect 178587 530050 178621 530084
rect 178679 530050 178713 530084
rect 178771 530050 178805 530084
rect 178863 530050 178897 530084
rect 178955 530050 178989 530084
rect 179047 530050 179081 530084
rect 179139 530050 179173 530084
rect 179231 530050 179265 530084
rect 179323 530050 179357 530084
rect 179415 530050 179449 530084
rect 179507 530050 179541 530084
rect 179599 530050 179633 530084
rect 179691 530050 179725 530084
rect 179783 530050 179817 530084
rect 179875 530050 179909 530084
rect 179967 530050 180001 530084
rect 180059 530050 180093 530084
rect 180151 530050 180185 530084
rect 180243 530050 180277 530084
rect 180335 530050 180369 530084
rect 180427 530050 180461 530084
rect 180519 530050 180553 530084
rect 180611 530050 180645 530084
rect 180703 530050 180737 530084
rect 180795 530050 180829 530084
rect 180887 530050 180921 530084
rect 180979 530050 181013 530084
rect 181071 530050 181105 530084
rect 181163 530050 181197 530084
rect 181255 530050 181289 530084
rect 181347 530050 181381 530084
rect 181439 530050 181473 530084
rect 181531 530050 181565 530084
rect 181623 530050 181657 530084
rect 181715 530050 181749 530084
rect 181807 530050 181841 530084
rect 181899 530050 181933 530084
rect 181991 530050 182025 530084
rect 182083 530050 182117 530084
rect 182175 530050 182209 530084
rect 182267 530050 182301 530084
rect 182359 530050 182393 530084
rect 182451 530050 182485 530084
rect 182543 530050 182577 530084
rect 182635 530050 182669 530084
rect 182727 530050 182761 530084
rect 182819 530050 182853 530084
rect 182911 530050 182945 530084
rect 183003 530050 183037 530084
rect 183095 530050 183129 530084
rect 183187 530050 183221 530084
rect 183279 530050 183313 530084
rect 183371 530050 183405 530084
rect 183463 530050 183497 530084
rect 183555 530050 183589 530084
rect 183647 530050 183681 530084
rect 183739 530050 183773 530084
rect 183831 530050 183865 530084
rect 183923 530050 183957 530084
rect 184015 530050 184049 530084
rect 184107 530050 184141 530084
rect 184199 530050 184233 530084
rect 184291 530050 184325 530084
rect 184383 530050 184417 530084
rect 184475 530050 184509 530084
rect 184567 530050 184601 530084
rect 184659 530050 184693 530084
rect 184751 530050 184785 530084
rect 184843 530050 184877 530084
rect 184935 530050 184969 530084
rect 185027 530050 185061 530084
rect 185119 530050 185153 530084
rect 185211 530050 185245 530084
rect 185303 530050 185337 530084
rect 185395 530050 185429 530084
rect 185487 530050 185521 530084
rect 185579 530050 185613 530084
rect 185671 530050 185705 530084
rect 185763 530050 185797 530084
rect 185855 530050 185889 530084
rect 185947 530050 185981 530084
rect 186039 530050 186073 530084
rect 186131 530050 186165 530084
rect 186223 530050 186257 530084
rect 186315 530050 186349 530084
rect 186407 530050 186441 530084
rect 186499 530050 186533 530084
rect 186591 530050 186625 530084
rect 186683 530050 186717 530084
rect 186775 530050 186809 530084
rect 186867 530050 186901 530084
rect 186959 530050 186993 530084
rect 187051 530050 187085 530084
rect 187143 530050 187177 530084
rect 187235 530050 187269 530084
rect 187327 530050 187361 530084
rect 187419 530050 187453 530084
rect 174815 529812 174849 529846
rect 175551 529772 175585 529778
rect 175551 529744 175554 529772
rect 175554 529744 175585 529772
rect 175644 529753 175656 529778
rect 175656 529753 175678 529778
rect 175644 529744 175678 529753
rect 175459 529608 175468 529642
rect 175468 529608 175493 529642
rect 175725 529898 175759 529914
rect 175725 529880 175759 529898
rect 175827 529812 175861 529846
rect 176103 529880 176137 529914
rect 176011 529744 176045 529778
rect 176727 529888 176761 529914
rect 176727 529880 176758 529888
rect 176758 529880 176761 529888
rect 176283 529676 176317 529710
rect 176355 529692 176379 529710
rect 176379 529692 176389 529710
rect 176355 529676 176389 529692
rect 176727 529762 176761 529778
rect 176727 529744 176753 529762
rect 176753 529744 176761 529762
rect 177299 529972 177333 529982
rect 177299 529948 177327 529972
rect 177327 529948 177333 529972
rect 176943 529764 176977 529773
rect 176943 529739 176959 529764
rect 176959 529739 176977 529764
rect 177003 529676 177037 529710
rect 177667 529815 177681 529846
rect 177681 529815 177701 529846
rect 177667 529812 177701 529815
rect 177851 529676 177885 529710
rect 177943 529744 177977 529778
rect 178311 529906 178339 529914
rect 178339 529906 178345 529914
rect 178311 529880 178345 529906
rect 178403 529972 178437 529982
rect 178403 529948 178409 529972
rect 178409 529948 178437 529972
rect 178975 529888 179009 529914
rect 178975 529880 178978 529888
rect 178978 529880 179009 529888
rect 178759 529764 178793 529773
rect 178759 529739 178777 529764
rect 178777 529739 178793 529764
rect 178699 529676 178733 529710
rect 178975 529762 179009 529778
rect 178975 529744 178983 529762
rect 178983 529744 179009 529762
rect 179599 529880 179633 529914
rect 179347 529692 179357 529710
rect 179357 529692 179381 529710
rect 179347 529676 179381 529692
rect 179419 529676 179453 529710
rect 179691 529744 179725 529778
rect 179977 529898 180011 529914
rect 179977 529880 180011 529898
rect 179875 529812 179909 529846
rect 180058 529753 180080 529778
rect 180080 529753 180092 529778
rect 180058 529744 180092 529753
rect 180151 529772 180185 529778
rect 180151 529744 180182 529772
rect 180182 529744 180185 529772
rect 180243 529772 180277 529778
rect 180243 529744 180246 529772
rect 180246 529744 180277 529772
rect 180336 529753 180348 529778
rect 180348 529753 180370 529778
rect 180336 529744 180370 529753
rect 180417 529898 180451 529914
rect 180417 529880 180451 529898
rect 180519 529812 180553 529846
rect 180795 529880 180829 529914
rect 180703 529744 180737 529778
rect 181419 529888 181453 529914
rect 181419 529880 181450 529888
rect 181450 529880 181453 529888
rect 180975 529676 181009 529710
rect 181047 529692 181071 529710
rect 181071 529692 181081 529710
rect 181047 529676 181081 529692
rect 181419 529762 181453 529778
rect 181419 529744 181445 529762
rect 181445 529744 181453 529762
rect 181991 529812 182025 529846
rect 181635 529764 181669 529773
rect 181635 529739 181651 529764
rect 181651 529739 181669 529764
rect 181695 529676 181729 529710
rect 182635 529948 182660 529982
rect 182660 529948 182669 529982
rect 183187 529812 183221 529846
rect 172239 529506 172273 529540
rect 172331 529506 172365 529540
rect 172423 529506 172457 529540
rect 172515 529506 172549 529540
rect 172607 529506 172641 529540
rect 172699 529506 172733 529540
rect 172791 529506 172825 529540
rect 172883 529506 172917 529540
rect 172975 529506 173009 529540
rect 173067 529506 173101 529540
rect 173159 529506 173193 529540
rect 173251 529506 173285 529540
rect 173343 529506 173377 529540
rect 173435 529506 173469 529540
rect 173527 529506 173561 529540
rect 173619 529506 173653 529540
rect 173711 529506 173745 529540
rect 173803 529506 173837 529540
rect 173895 529506 173929 529540
rect 173987 529506 174021 529540
rect 174079 529506 174113 529540
rect 174171 529506 174205 529540
rect 174263 529506 174297 529540
rect 174355 529506 174389 529540
rect 174447 529506 174481 529540
rect 174539 529506 174573 529540
rect 174631 529506 174665 529540
rect 174723 529506 174757 529540
rect 174815 529506 174849 529540
rect 174907 529506 174941 529540
rect 174999 529506 175033 529540
rect 175091 529506 175125 529540
rect 175183 529506 175217 529540
rect 175275 529506 175309 529540
rect 175367 529506 175401 529540
rect 175459 529506 175493 529540
rect 175551 529506 175585 529540
rect 175643 529506 175677 529540
rect 175735 529506 175769 529540
rect 175827 529506 175861 529540
rect 175919 529506 175953 529540
rect 176011 529506 176045 529540
rect 176103 529506 176137 529540
rect 176195 529506 176229 529540
rect 176287 529506 176321 529540
rect 176379 529506 176413 529540
rect 176471 529506 176505 529540
rect 176563 529506 176597 529540
rect 176655 529506 176689 529540
rect 176747 529506 176781 529540
rect 176839 529506 176873 529540
rect 176931 529506 176965 529540
rect 177023 529506 177057 529540
rect 177115 529506 177149 529540
rect 177207 529506 177241 529540
rect 177299 529506 177333 529540
rect 177391 529506 177425 529540
rect 177483 529506 177517 529540
rect 177575 529506 177609 529540
rect 177667 529506 177701 529540
rect 177759 529506 177793 529540
rect 177851 529506 177885 529540
rect 177943 529506 177977 529540
rect 178035 529506 178069 529540
rect 178127 529506 178161 529540
rect 178219 529506 178253 529540
rect 178311 529506 178345 529540
rect 178403 529506 178437 529540
rect 178495 529506 178529 529540
rect 178587 529506 178621 529540
rect 178679 529506 178713 529540
rect 178771 529506 178805 529540
rect 178863 529506 178897 529540
rect 178955 529506 178989 529540
rect 179047 529506 179081 529540
rect 179139 529506 179173 529540
rect 179231 529506 179265 529540
rect 179323 529506 179357 529540
rect 179415 529506 179449 529540
rect 179507 529506 179541 529540
rect 179599 529506 179633 529540
rect 179691 529506 179725 529540
rect 179783 529506 179817 529540
rect 179875 529506 179909 529540
rect 179967 529506 180001 529540
rect 180059 529506 180093 529540
rect 180151 529506 180185 529540
rect 180243 529506 180277 529540
rect 180335 529506 180369 529540
rect 180427 529506 180461 529540
rect 180519 529506 180553 529540
rect 180611 529506 180645 529540
rect 180703 529506 180737 529540
rect 180795 529506 180829 529540
rect 180887 529506 180921 529540
rect 180979 529506 181013 529540
rect 181071 529506 181105 529540
rect 181163 529506 181197 529540
rect 181255 529506 181289 529540
rect 181347 529506 181381 529540
rect 181439 529506 181473 529540
rect 181531 529506 181565 529540
rect 181623 529506 181657 529540
rect 181715 529506 181749 529540
rect 181807 529506 181841 529540
rect 181899 529506 181933 529540
rect 181991 529506 182025 529540
rect 182083 529506 182117 529540
rect 182175 529506 182209 529540
rect 182267 529506 182301 529540
rect 182359 529506 182393 529540
rect 182451 529506 182485 529540
rect 182543 529506 182577 529540
rect 182635 529506 182669 529540
rect 182727 529506 182761 529540
rect 182819 529506 182853 529540
rect 182911 529506 182945 529540
rect 183003 529506 183037 529540
rect 183095 529506 183129 529540
rect 183187 529506 183221 529540
rect 183279 529506 183313 529540
rect 183371 529506 183405 529540
rect 183463 529506 183497 529540
rect 183555 529506 183589 529540
rect 183647 529506 183681 529540
rect 183739 529506 183773 529540
rect 183831 529506 183865 529540
rect 183923 529506 183957 529540
rect 184015 529506 184049 529540
rect 184107 529506 184141 529540
rect 184199 529506 184233 529540
rect 184291 529506 184325 529540
rect 184383 529506 184417 529540
rect 184475 529506 184509 529540
rect 184567 529506 184601 529540
rect 184659 529506 184693 529540
rect 184751 529506 184785 529540
rect 184843 529506 184877 529540
rect 184935 529506 184969 529540
rect 185027 529506 185061 529540
rect 185119 529506 185153 529540
rect 185211 529506 185245 529540
rect 185303 529506 185337 529540
rect 185395 529506 185429 529540
rect 185487 529506 185521 529540
rect 185579 529506 185613 529540
rect 185671 529506 185705 529540
rect 185763 529506 185797 529540
rect 185855 529506 185889 529540
rect 185947 529506 185981 529540
rect 186039 529506 186073 529540
rect 186131 529506 186165 529540
rect 186223 529506 186257 529540
rect 186315 529506 186349 529540
rect 186407 529506 186441 529540
rect 186499 529506 186533 529540
rect 186591 529506 186625 529540
rect 186683 529506 186717 529540
rect 186775 529506 186809 529540
rect 186867 529506 186901 529540
rect 186959 529506 186993 529540
rect 187051 529506 187085 529540
rect 187143 529506 187177 529540
rect 187235 529506 187269 529540
rect 187327 529506 187361 529540
rect 187419 529506 187453 529540
rect 175367 529404 175401 529438
rect 175275 529200 175309 529234
rect 175459 529268 175493 529302
rect 177667 529274 177693 529302
rect 177693 529274 177701 529302
rect 177667 529268 177701 529274
rect 175827 529072 175861 529098
rect 175827 529064 175855 529072
rect 175855 529064 175861 529072
rect 176195 529082 176200 529098
rect 176200 529082 176229 529098
rect 176195 529064 176229 529082
rect 177759 529200 177793 529234
rect 177852 529293 177886 529302
rect 177852 529268 177864 529293
rect 177864 529268 177886 529293
rect 178035 529336 178069 529370
rect 177933 529148 177967 529166
rect 177933 529132 177967 529148
rect 178219 529268 178253 529302
rect 178491 529336 178525 529370
rect 178563 529354 178597 529370
rect 178563 529336 178587 529354
rect 178587 529336 178597 529354
rect 178311 529132 178345 529166
rect 178935 529284 178961 529302
rect 178961 529284 178969 529302
rect 178935 529268 178969 529284
rect 179211 529336 179245 529370
rect 179151 529282 179167 529307
rect 179167 529282 179185 529307
rect 179151 529273 179185 529282
rect 178935 529158 178966 529166
rect 178966 529158 178969 529166
rect 178935 529132 178969 529158
rect 179875 529434 179909 529438
rect 179875 529404 179903 529434
rect 179903 529404 179909 529434
rect 179691 529274 179699 529302
rect 179699 529274 179725 529302
rect 179691 529268 179725 529274
rect 179507 529074 179535 529098
rect 179535 529074 179541 529098
rect 179507 529064 179541 529074
rect 180703 529274 180711 529302
rect 180711 529274 180737 529302
rect 180703 529268 180737 529274
rect 182543 529434 182577 529438
rect 182543 529404 182549 529434
rect 182549 529404 182577 529434
rect 181991 529082 181998 529098
rect 181998 529082 182025 529098
rect 181991 529064 182025 529082
rect 182727 529274 182753 529302
rect 182753 529274 182761 529302
rect 182727 529268 182761 529274
rect 172239 528962 172273 528996
rect 172331 528962 172365 528996
rect 172423 528962 172457 528996
rect 172515 528962 172549 528996
rect 172607 528962 172641 528996
rect 172699 528962 172733 528996
rect 172791 528962 172825 528996
rect 172883 528962 172917 528996
rect 172975 528962 173009 528996
rect 173067 528962 173101 528996
rect 173159 528962 173193 528996
rect 173251 528962 173285 528996
rect 173343 528962 173377 528996
rect 173435 528962 173469 528996
rect 173527 528962 173561 528996
rect 173619 528962 173653 528996
rect 173711 528962 173745 528996
rect 173803 528962 173837 528996
rect 173895 528962 173929 528996
rect 173987 528962 174021 528996
rect 174079 528962 174113 528996
rect 174171 528962 174205 528996
rect 174263 528962 174297 528996
rect 174355 528962 174389 528996
rect 174447 528962 174481 528996
rect 174539 528962 174573 528996
rect 174631 528962 174665 528996
rect 174723 528962 174757 528996
rect 174815 528962 174849 528996
rect 174907 528962 174941 528996
rect 174999 528962 175033 528996
rect 175091 528962 175125 528996
rect 175183 528962 175217 528996
rect 175275 528962 175309 528996
rect 175367 528962 175401 528996
rect 175459 528962 175493 528996
rect 175551 528962 175585 528996
rect 175643 528962 175677 528996
rect 175735 528962 175769 528996
rect 175827 528962 175861 528996
rect 175919 528962 175953 528996
rect 176011 528962 176045 528996
rect 176103 528962 176137 528996
rect 176195 528962 176229 528996
rect 176287 528962 176321 528996
rect 176379 528962 176413 528996
rect 176471 528962 176505 528996
rect 176563 528962 176597 528996
rect 176655 528962 176689 528996
rect 176747 528962 176781 528996
rect 176839 528962 176873 528996
rect 176931 528962 176965 528996
rect 177023 528962 177057 528996
rect 177115 528962 177149 528996
rect 177207 528962 177241 528996
rect 177299 528962 177333 528996
rect 177391 528962 177425 528996
rect 177483 528962 177517 528996
rect 177575 528962 177609 528996
rect 177667 528962 177701 528996
rect 177759 528962 177793 528996
rect 177851 528962 177885 528996
rect 177943 528962 177977 528996
rect 178035 528962 178069 528996
rect 178127 528962 178161 528996
rect 178219 528962 178253 528996
rect 178311 528962 178345 528996
rect 178403 528962 178437 528996
rect 178495 528962 178529 528996
rect 178587 528962 178621 528996
rect 178679 528962 178713 528996
rect 178771 528962 178805 528996
rect 178863 528962 178897 528996
rect 178955 528962 178989 528996
rect 179047 528962 179081 528996
rect 179139 528962 179173 528996
rect 179231 528962 179265 528996
rect 179323 528962 179357 528996
rect 179415 528962 179449 528996
rect 179507 528962 179541 528996
rect 179599 528962 179633 528996
rect 179691 528962 179725 528996
rect 179783 528962 179817 528996
rect 179875 528962 179909 528996
rect 179967 528962 180001 528996
rect 180059 528962 180093 528996
rect 180151 528962 180185 528996
rect 180243 528962 180277 528996
rect 180335 528962 180369 528996
rect 180427 528962 180461 528996
rect 180519 528962 180553 528996
rect 180611 528962 180645 528996
rect 180703 528962 180737 528996
rect 180795 528962 180829 528996
rect 180887 528962 180921 528996
rect 180979 528962 181013 528996
rect 181071 528962 181105 528996
rect 181163 528962 181197 528996
rect 181255 528962 181289 528996
rect 181347 528962 181381 528996
rect 181439 528962 181473 528996
rect 181531 528962 181565 528996
rect 181623 528962 181657 528996
rect 181715 528962 181749 528996
rect 181807 528962 181841 528996
rect 181899 528962 181933 528996
rect 181991 528962 182025 528996
rect 182083 528962 182117 528996
rect 182175 528962 182209 528996
rect 182267 528962 182301 528996
rect 182359 528962 182393 528996
rect 182451 528962 182485 528996
rect 182543 528962 182577 528996
rect 182635 528962 182669 528996
rect 182727 528962 182761 528996
rect 182819 528962 182853 528996
rect 182911 528962 182945 528996
rect 183003 528962 183037 528996
rect 183095 528962 183129 528996
rect 183187 528962 183221 528996
rect 183279 528962 183313 528996
rect 183371 528962 183405 528996
rect 183463 528962 183497 528996
rect 183555 528962 183589 528996
rect 183647 528962 183681 528996
rect 183739 528962 183773 528996
rect 183831 528962 183865 528996
rect 183923 528962 183957 528996
rect 184015 528962 184049 528996
rect 184107 528962 184141 528996
rect 184199 528962 184233 528996
rect 184291 528962 184325 528996
rect 184383 528962 184417 528996
rect 184475 528962 184509 528996
rect 184567 528962 184601 528996
rect 184659 528962 184693 528996
rect 184751 528962 184785 528996
rect 184843 528962 184877 528996
rect 184935 528962 184969 528996
rect 185027 528962 185061 528996
rect 185119 528962 185153 528996
rect 185211 528962 185245 528996
rect 185303 528962 185337 528996
rect 185395 528962 185429 528996
rect 185487 528962 185521 528996
rect 185579 528962 185613 528996
rect 185671 528962 185705 528996
rect 185763 528962 185797 528996
rect 185855 528962 185889 528996
rect 185947 528962 185981 528996
rect 186039 528962 186073 528996
rect 186131 528962 186165 528996
rect 186223 528962 186257 528996
rect 186315 528962 186349 528996
rect 186407 528962 186441 528996
rect 186499 528962 186533 528996
rect 186591 528962 186625 528996
rect 186683 528962 186717 528996
rect 186775 528962 186809 528996
rect 186867 528962 186901 528996
rect 186959 528962 186993 528996
rect 187051 528962 187085 528996
rect 187143 528962 187177 528996
rect 187235 528962 187269 528996
rect 187327 528962 187361 528996
rect 187419 528962 187453 528996
rect 176103 528878 176131 528894
rect 176131 528878 176137 528894
rect 176103 528860 176137 528878
rect 175919 528684 175953 528690
rect 175919 528656 175927 528684
rect 175927 528656 175953 528684
rect 176195 528684 176229 528690
rect 176195 528656 176203 528684
rect 176203 528656 176229 528684
rect 176563 528727 176577 528758
rect 176577 528727 176597 528758
rect 176563 528724 176597 528727
rect 176379 528524 176407 528554
rect 176407 528524 176413 528554
rect 176379 528520 176413 528524
rect 176747 528520 176781 528554
rect 176839 528656 176873 528690
rect 177483 528656 177517 528690
rect 177207 528547 177241 528554
rect 177207 528520 177235 528547
rect 177235 528520 177241 528547
rect 178127 528724 178161 528758
rect 179691 528876 179725 528894
rect 179691 528860 179698 528876
rect 179698 528860 179725 528876
rect 180427 528797 180455 528826
rect 180455 528797 180461 528826
rect 180427 528792 180461 528797
rect 178403 528588 178437 528622
rect 180243 528684 180277 528690
rect 180243 528656 180251 528684
rect 180251 528656 180277 528684
rect 180519 528724 180553 528758
rect 180612 528665 180624 528690
rect 180624 528665 180646 528690
rect 180612 528656 180646 528665
rect 180693 528810 180727 528826
rect 180693 528792 180727 528810
rect 180795 528724 180829 528758
rect 181071 528792 181105 528826
rect 180979 528656 181013 528690
rect 181695 528800 181729 528826
rect 181695 528792 181726 528800
rect 181726 528792 181729 528800
rect 181251 528588 181285 528622
rect 181323 528604 181347 528622
rect 181347 528604 181357 528622
rect 181323 528588 181357 528604
rect 181695 528674 181729 528690
rect 181695 528656 181721 528674
rect 181721 528656 181729 528674
rect 182267 528884 182301 528894
rect 182267 528860 182295 528884
rect 182295 528860 182301 528884
rect 181911 528676 181945 528685
rect 181911 528651 181927 528676
rect 181927 528651 181945 528676
rect 181971 528588 182005 528622
rect 172239 528418 172273 528452
rect 172331 528418 172365 528452
rect 172423 528418 172457 528452
rect 172515 528418 172549 528452
rect 172607 528418 172641 528452
rect 172699 528418 172733 528452
rect 172791 528418 172825 528452
rect 172883 528418 172917 528452
rect 172975 528418 173009 528452
rect 173067 528418 173101 528452
rect 173159 528418 173193 528452
rect 173251 528418 173285 528452
rect 173343 528418 173377 528452
rect 173435 528418 173469 528452
rect 173527 528418 173561 528452
rect 173619 528418 173653 528452
rect 173711 528418 173745 528452
rect 173803 528418 173837 528452
rect 173895 528418 173929 528452
rect 173987 528418 174021 528452
rect 174079 528418 174113 528452
rect 174171 528418 174205 528452
rect 174263 528418 174297 528452
rect 174355 528418 174389 528452
rect 174447 528418 174481 528452
rect 174539 528418 174573 528452
rect 174631 528418 174665 528452
rect 174723 528418 174757 528452
rect 174815 528418 174849 528452
rect 174907 528418 174941 528452
rect 174999 528418 175033 528452
rect 175091 528418 175125 528452
rect 175183 528418 175217 528452
rect 175275 528418 175309 528452
rect 175367 528418 175401 528452
rect 175459 528418 175493 528452
rect 175551 528418 175585 528452
rect 175643 528418 175677 528452
rect 175735 528418 175769 528452
rect 175827 528418 175861 528452
rect 175919 528418 175953 528452
rect 176011 528418 176045 528452
rect 176103 528418 176137 528452
rect 176195 528418 176229 528452
rect 176287 528418 176321 528452
rect 176379 528418 176413 528452
rect 176471 528418 176505 528452
rect 176563 528418 176597 528452
rect 176655 528418 176689 528452
rect 176747 528418 176781 528452
rect 176839 528418 176873 528452
rect 176931 528418 176965 528452
rect 177023 528418 177057 528452
rect 177115 528418 177149 528452
rect 177207 528418 177241 528452
rect 177299 528418 177333 528452
rect 177391 528418 177425 528452
rect 177483 528418 177517 528452
rect 177575 528418 177609 528452
rect 177667 528418 177701 528452
rect 177759 528418 177793 528452
rect 177851 528418 177885 528452
rect 177943 528418 177977 528452
rect 178035 528418 178069 528452
rect 178127 528418 178161 528452
rect 178219 528418 178253 528452
rect 178311 528418 178345 528452
rect 178403 528418 178437 528452
rect 178495 528418 178529 528452
rect 178587 528418 178621 528452
rect 178679 528418 178713 528452
rect 178771 528418 178805 528452
rect 178863 528418 178897 528452
rect 178955 528418 178989 528452
rect 179047 528418 179081 528452
rect 179139 528418 179173 528452
rect 179231 528418 179265 528452
rect 179323 528418 179357 528452
rect 179415 528418 179449 528452
rect 179507 528418 179541 528452
rect 179599 528418 179633 528452
rect 179691 528418 179725 528452
rect 179783 528418 179817 528452
rect 179875 528418 179909 528452
rect 179967 528418 180001 528452
rect 180059 528418 180093 528452
rect 180151 528418 180185 528452
rect 180243 528418 180277 528452
rect 180335 528418 180369 528452
rect 180427 528418 180461 528452
rect 180519 528418 180553 528452
rect 180611 528418 180645 528452
rect 180703 528418 180737 528452
rect 180795 528418 180829 528452
rect 180887 528418 180921 528452
rect 180979 528418 181013 528452
rect 181071 528418 181105 528452
rect 181163 528418 181197 528452
rect 181255 528418 181289 528452
rect 181347 528418 181381 528452
rect 181439 528418 181473 528452
rect 181531 528418 181565 528452
rect 181623 528418 181657 528452
rect 181715 528418 181749 528452
rect 181807 528418 181841 528452
rect 181899 528418 181933 528452
rect 181991 528418 182025 528452
rect 182083 528418 182117 528452
rect 182175 528418 182209 528452
rect 182267 528418 182301 528452
rect 182359 528418 182393 528452
rect 182451 528418 182485 528452
rect 182543 528418 182577 528452
rect 182635 528418 182669 528452
rect 182727 528418 182761 528452
rect 182819 528418 182853 528452
rect 182911 528418 182945 528452
rect 183003 528418 183037 528452
rect 183095 528418 183129 528452
rect 183187 528418 183221 528452
rect 183279 528418 183313 528452
rect 183371 528418 183405 528452
rect 183463 528418 183497 528452
rect 183555 528418 183589 528452
rect 183647 528418 183681 528452
rect 183739 528418 183773 528452
rect 183831 528418 183865 528452
rect 183923 528418 183957 528452
rect 184015 528418 184049 528452
rect 184107 528418 184141 528452
rect 184199 528418 184233 528452
rect 184291 528418 184325 528452
rect 184383 528418 184417 528452
rect 184475 528418 184509 528452
rect 184567 528418 184601 528452
rect 184659 528418 184693 528452
rect 184751 528418 184785 528452
rect 184843 528418 184877 528452
rect 184935 528418 184969 528452
rect 185027 528418 185061 528452
rect 185119 528418 185153 528452
rect 185211 528418 185245 528452
rect 185303 528418 185337 528452
rect 185395 528418 185429 528452
rect 185487 528418 185521 528452
rect 185579 528418 185613 528452
rect 185671 528418 185705 528452
rect 185763 528418 185797 528452
rect 185855 528418 185889 528452
rect 185947 528418 185981 528452
rect 186039 528418 186073 528452
rect 186131 528418 186165 528452
rect 186223 528418 186257 528452
rect 186315 528418 186349 528452
rect 186407 528418 186441 528452
rect 186499 528418 186533 528452
rect 186591 528418 186625 528452
rect 186683 528418 186717 528452
rect 186775 528418 186809 528452
rect 186867 528418 186901 528452
rect 186959 528418 186993 528452
rect 187051 528418 187085 528452
rect 187143 528418 187177 528452
rect 187235 528418 187269 528452
rect 187327 528418 187361 528452
rect 187419 528418 187453 528452
rect 176103 528186 176106 528214
rect 176106 528186 176137 528214
rect 176103 528180 176137 528186
rect 176196 528205 176230 528214
rect 176196 528180 176208 528205
rect 176208 528180 176230 528205
rect 176379 528248 176413 528282
rect 176277 528060 176311 528078
rect 176277 528044 176311 528060
rect 176563 528180 176597 528214
rect 176835 528248 176869 528282
rect 176907 528266 176941 528282
rect 176907 528248 176931 528266
rect 176931 528248 176941 528266
rect 176655 528044 176689 528078
rect 177279 528196 177305 528214
rect 177305 528196 177313 528214
rect 177279 528180 177313 528196
rect 177851 528326 177885 528350
rect 177555 528248 177589 528282
rect 177495 528194 177511 528219
rect 177511 528194 177529 528219
rect 177495 528185 177529 528194
rect 177851 528316 177879 528326
rect 177879 528316 177885 528326
rect 177279 528070 177310 528078
rect 177310 528070 177313 528078
rect 177279 528044 177313 528070
rect 178955 528323 178961 528350
rect 178961 528323 178989 528350
rect 178955 528316 178989 528323
rect 178127 528186 178153 528214
rect 178153 528186 178161 528214
rect 178127 528180 178161 528186
rect 177943 528073 177977 528078
rect 177943 528044 177949 528073
rect 177949 528044 177977 528073
rect 179323 528180 179357 528214
rect 179415 528316 179449 528350
rect 180979 528323 180985 528350
rect 180985 528323 181013 528350
rect 180979 528316 181013 528323
rect 179507 528112 179541 528146
rect 181347 528180 181381 528214
rect 181439 528316 181473 528350
rect 181531 528112 181565 528146
rect 172239 527874 172273 527908
rect 172331 527874 172365 527908
rect 172423 527874 172457 527908
rect 172515 527874 172549 527908
rect 172607 527874 172641 527908
rect 172699 527874 172733 527908
rect 172791 527874 172825 527908
rect 172883 527874 172917 527908
rect 172975 527874 173009 527908
rect 173067 527874 173101 527908
rect 173159 527874 173193 527908
rect 173251 527874 173285 527908
rect 173343 527874 173377 527908
rect 173435 527874 173469 527908
rect 173527 527874 173561 527908
rect 173619 527874 173653 527908
rect 173711 527874 173745 527908
rect 173803 527874 173837 527908
rect 173895 527874 173929 527908
rect 173987 527874 174021 527908
rect 174079 527874 174113 527908
rect 174171 527874 174205 527908
rect 174263 527874 174297 527908
rect 174355 527874 174389 527908
rect 174447 527874 174481 527908
rect 174539 527874 174573 527908
rect 174631 527874 174665 527908
rect 174723 527874 174757 527908
rect 174815 527874 174849 527908
rect 174907 527874 174941 527908
rect 174999 527874 175033 527908
rect 175091 527874 175125 527908
rect 175183 527874 175217 527908
rect 175275 527874 175309 527908
rect 175367 527874 175401 527908
rect 175459 527874 175493 527908
rect 175551 527874 175585 527908
rect 175643 527874 175677 527908
rect 175735 527874 175769 527908
rect 175827 527874 175861 527908
rect 175919 527874 175953 527908
rect 176011 527874 176045 527908
rect 176103 527874 176137 527908
rect 176195 527874 176229 527908
rect 176287 527874 176321 527908
rect 176379 527874 176413 527908
rect 176471 527874 176505 527908
rect 176563 527874 176597 527908
rect 176655 527874 176689 527908
rect 176747 527874 176781 527908
rect 176839 527874 176873 527908
rect 176931 527874 176965 527908
rect 177023 527874 177057 527908
rect 177115 527874 177149 527908
rect 177207 527874 177241 527908
rect 177299 527874 177333 527908
rect 177391 527874 177425 527908
rect 177483 527874 177517 527908
rect 177575 527874 177609 527908
rect 177667 527874 177701 527908
rect 177759 527874 177793 527908
rect 177851 527874 177885 527908
rect 177943 527874 177977 527908
rect 178035 527874 178069 527908
rect 178127 527874 178161 527908
rect 178219 527874 178253 527908
rect 178311 527874 178345 527908
rect 178403 527874 178437 527908
rect 178495 527874 178529 527908
rect 178587 527874 178621 527908
rect 178679 527874 178713 527908
rect 178771 527874 178805 527908
rect 178863 527874 178897 527908
rect 178955 527874 178989 527908
rect 179047 527874 179081 527908
rect 179139 527874 179173 527908
rect 179231 527874 179265 527908
rect 179323 527874 179357 527908
rect 179415 527874 179449 527908
rect 179507 527874 179541 527908
rect 179599 527874 179633 527908
rect 179691 527874 179725 527908
rect 179783 527874 179817 527908
rect 179875 527874 179909 527908
rect 179967 527874 180001 527908
rect 180059 527874 180093 527908
rect 180151 527874 180185 527908
rect 180243 527874 180277 527908
rect 180335 527874 180369 527908
rect 180427 527874 180461 527908
rect 180519 527874 180553 527908
rect 180611 527874 180645 527908
rect 180703 527874 180737 527908
rect 180795 527874 180829 527908
rect 180887 527874 180921 527908
rect 180979 527874 181013 527908
rect 181071 527874 181105 527908
rect 181163 527874 181197 527908
rect 181255 527874 181289 527908
rect 181347 527874 181381 527908
rect 181439 527874 181473 527908
rect 181531 527874 181565 527908
rect 181623 527874 181657 527908
rect 181715 527874 181749 527908
rect 181807 527874 181841 527908
rect 181899 527874 181933 527908
rect 181991 527874 182025 527908
rect 182083 527874 182117 527908
rect 182175 527874 182209 527908
rect 182267 527874 182301 527908
rect 182359 527874 182393 527908
rect 182451 527874 182485 527908
rect 182543 527874 182577 527908
rect 182635 527874 182669 527908
rect 182727 527874 182761 527908
rect 182819 527874 182853 527908
rect 182911 527874 182945 527908
rect 183003 527874 183037 527908
rect 183095 527874 183129 527908
rect 183187 527874 183221 527908
rect 183279 527874 183313 527908
rect 183371 527874 183405 527908
rect 183463 527874 183497 527908
rect 183555 527874 183589 527908
rect 183647 527874 183681 527908
rect 183739 527874 183773 527908
rect 183831 527874 183865 527908
rect 183923 527874 183957 527908
rect 184015 527874 184049 527908
rect 184107 527874 184141 527908
rect 184199 527874 184233 527908
rect 184291 527874 184325 527908
rect 184383 527874 184417 527908
rect 184475 527874 184509 527908
rect 184567 527874 184601 527908
rect 184659 527874 184693 527908
rect 184751 527874 184785 527908
rect 184843 527874 184877 527908
rect 184935 527874 184969 527908
rect 185027 527874 185061 527908
rect 185119 527874 185153 527908
rect 185211 527874 185245 527908
rect 185303 527874 185337 527908
rect 185395 527874 185429 527908
rect 185487 527874 185521 527908
rect 185579 527874 185613 527908
rect 185671 527874 185705 527908
rect 185763 527874 185797 527908
rect 185855 527874 185889 527908
rect 185947 527874 185981 527908
rect 186039 527874 186073 527908
rect 186131 527874 186165 527908
rect 186223 527874 186257 527908
rect 186315 527874 186349 527908
rect 186407 527874 186441 527908
rect 186499 527874 186533 527908
rect 186591 527874 186625 527908
rect 186683 527874 186717 527908
rect 186775 527874 186809 527908
rect 186867 527874 186901 527908
rect 186959 527874 186993 527908
rect 187051 527874 187085 527908
rect 187143 527874 187177 527908
rect 187235 527874 187269 527908
rect 187327 527874 187361 527908
rect 187419 527874 187453 527908
rect 176379 527772 176404 527806
rect 176404 527772 176413 527806
rect 177023 527636 177057 527670
rect 178955 527772 178980 527806
rect 178980 527772 178989 527806
rect 179507 527636 179541 527670
rect 172239 527330 172273 527364
rect 172331 527330 172365 527364
rect 172423 527330 172457 527364
rect 172515 527330 172549 527364
rect 172607 527330 172641 527364
rect 172699 527330 172733 527364
rect 172791 527330 172825 527364
rect 172883 527330 172917 527364
rect 172975 527330 173009 527364
rect 173067 527330 173101 527364
rect 173159 527330 173193 527364
rect 173251 527330 173285 527364
rect 173343 527330 173377 527364
rect 173435 527330 173469 527364
rect 173527 527330 173561 527364
rect 173619 527330 173653 527364
rect 173711 527330 173745 527364
rect 173803 527330 173837 527364
rect 173895 527330 173929 527364
rect 173987 527330 174021 527364
rect 174079 527330 174113 527364
rect 174171 527330 174205 527364
rect 174263 527330 174297 527364
rect 174355 527330 174389 527364
rect 174447 527330 174481 527364
rect 174539 527330 174573 527364
rect 174631 527330 174665 527364
rect 174723 527330 174757 527364
rect 174815 527330 174849 527364
rect 174907 527330 174941 527364
rect 174999 527330 175033 527364
rect 175091 527330 175125 527364
rect 175183 527330 175217 527364
rect 175275 527330 175309 527364
rect 175367 527330 175401 527364
rect 175459 527330 175493 527364
rect 175551 527330 175585 527364
rect 175643 527330 175677 527364
rect 175735 527330 175769 527364
rect 175827 527330 175861 527364
rect 175919 527330 175953 527364
rect 176011 527330 176045 527364
rect 176103 527330 176137 527364
rect 176195 527330 176229 527364
rect 176287 527330 176321 527364
rect 176379 527330 176413 527364
rect 176471 527330 176505 527364
rect 176563 527330 176597 527364
rect 176655 527330 176689 527364
rect 176747 527330 176781 527364
rect 176839 527330 176873 527364
rect 176931 527330 176965 527364
rect 177023 527330 177057 527364
rect 177115 527330 177149 527364
rect 177207 527330 177241 527364
rect 177299 527330 177333 527364
rect 177391 527330 177425 527364
rect 177483 527330 177517 527364
rect 177575 527330 177609 527364
rect 177667 527330 177701 527364
rect 177759 527330 177793 527364
rect 177851 527330 177885 527364
rect 177943 527330 177977 527364
rect 178035 527330 178069 527364
rect 178127 527330 178161 527364
rect 178219 527330 178253 527364
rect 178311 527330 178345 527364
rect 178403 527330 178437 527364
rect 178495 527330 178529 527364
rect 178587 527330 178621 527364
rect 178679 527330 178713 527364
rect 178771 527330 178805 527364
rect 178863 527330 178897 527364
rect 178955 527330 178989 527364
rect 179047 527330 179081 527364
rect 179139 527330 179173 527364
rect 179231 527330 179265 527364
rect 179323 527330 179357 527364
rect 179415 527330 179449 527364
rect 179507 527330 179541 527364
rect 179599 527330 179633 527364
rect 179691 527330 179725 527364
rect 179783 527330 179817 527364
rect 179875 527330 179909 527364
rect 179967 527330 180001 527364
rect 180059 527330 180093 527364
rect 180151 527330 180185 527364
rect 180243 527330 180277 527364
rect 180335 527330 180369 527364
rect 180427 527330 180461 527364
rect 180519 527330 180553 527364
rect 180611 527330 180645 527364
rect 180703 527330 180737 527364
rect 180795 527330 180829 527364
rect 180887 527330 180921 527364
rect 180979 527330 181013 527364
rect 181071 527330 181105 527364
rect 181163 527330 181197 527364
rect 181255 527330 181289 527364
rect 181347 527330 181381 527364
rect 181439 527330 181473 527364
rect 181531 527330 181565 527364
rect 181623 527330 181657 527364
rect 181715 527330 181749 527364
rect 181807 527330 181841 527364
rect 181899 527330 181933 527364
rect 181991 527330 182025 527364
rect 182083 527330 182117 527364
rect 182175 527330 182209 527364
rect 182267 527330 182301 527364
rect 182359 527330 182393 527364
rect 182451 527330 182485 527364
rect 182543 527330 182577 527364
rect 182635 527330 182669 527364
rect 182727 527330 182761 527364
rect 182819 527330 182853 527364
rect 182911 527330 182945 527364
rect 183003 527330 183037 527364
rect 183095 527330 183129 527364
rect 183187 527330 183221 527364
rect 183279 527330 183313 527364
rect 183371 527330 183405 527364
rect 183463 527330 183497 527364
rect 183555 527330 183589 527364
rect 183647 527330 183681 527364
rect 183739 527330 183773 527364
rect 183831 527330 183865 527364
rect 183923 527330 183957 527364
rect 184015 527330 184049 527364
rect 184107 527330 184141 527364
rect 184199 527330 184233 527364
rect 184291 527330 184325 527364
rect 184383 527330 184417 527364
rect 184475 527330 184509 527364
rect 184567 527330 184601 527364
rect 184659 527330 184693 527364
rect 184751 527330 184785 527364
rect 184843 527330 184877 527364
rect 184935 527330 184969 527364
rect 185027 527330 185061 527364
rect 185119 527330 185153 527364
rect 185211 527330 185245 527364
rect 185303 527330 185337 527364
rect 185395 527330 185429 527364
rect 185487 527330 185521 527364
rect 185579 527330 185613 527364
rect 185671 527330 185705 527364
rect 185763 527330 185797 527364
rect 185855 527330 185889 527364
rect 185947 527330 185981 527364
rect 186039 527330 186073 527364
rect 186131 527330 186165 527364
rect 186223 527330 186257 527364
rect 186315 527330 186349 527364
rect 186407 527330 186441 527364
rect 186499 527330 186533 527364
rect 186591 527330 186625 527364
rect 186683 527330 186717 527364
rect 186775 527330 186809 527364
rect 186867 527330 186901 527364
rect 186959 527330 186993 527364
rect 187051 527330 187085 527364
rect 187143 527330 187177 527364
rect 187235 527330 187269 527364
rect 187327 527330 187361 527364
rect 187419 527330 187453 527364
rect 172239 526786 172273 526820
rect 172331 526786 172365 526820
rect 172423 526786 172457 526820
rect 172515 526786 172549 526820
rect 172607 526786 172641 526820
rect 172699 526786 172733 526820
rect 172791 526786 172825 526820
rect 172883 526786 172917 526820
rect 172975 526786 173009 526820
rect 173067 526786 173101 526820
rect 173159 526786 173193 526820
rect 173251 526786 173285 526820
rect 173343 526786 173377 526820
rect 173435 526786 173469 526820
rect 173527 526786 173561 526820
rect 173619 526786 173653 526820
rect 173711 526786 173745 526820
rect 173803 526786 173837 526820
rect 173895 526786 173929 526820
rect 173987 526786 174021 526820
rect 174079 526786 174113 526820
rect 174171 526786 174205 526820
rect 174263 526786 174297 526820
rect 174355 526786 174389 526820
rect 174447 526786 174481 526820
rect 174539 526786 174573 526820
rect 174631 526786 174665 526820
rect 174723 526786 174757 526820
rect 174815 526786 174849 526820
rect 174907 526786 174941 526820
rect 174999 526786 175033 526820
rect 175091 526786 175125 526820
rect 175183 526786 175217 526820
rect 175275 526786 175309 526820
rect 175367 526786 175401 526820
rect 175459 526786 175493 526820
rect 175551 526786 175585 526820
rect 175643 526786 175677 526820
rect 175735 526786 175769 526820
rect 175827 526786 175861 526820
rect 175919 526786 175953 526820
rect 176011 526786 176045 526820
rect 176103 526786 176137 526820
rect 176195 526786 176229 526820
rect 176287 526786 176321 526820
rect 176379 526786 176413 526820
rect 176471 526786 176505 526820
rect 176563 526786 176597 526820
rect 176655 526786 176689 526820
rect 176747 526786 176781 526820
rect 176839 526786 176873 526820
rect 176931 526786 176965 526820
rect 177023 526786 177057 526820
rect 177115 526786 177149 526820
rect 177207 526786 177241 526820
rect 177299 526786 177333 526820
rect 177391 526786 177425 526820
rect 177483 526786 177517 526820
rect 177575 526786 177609 526820
rect 177667 526786 177701 526820
rect 177759 526786 177793 526820
rect 177851 526786 177885 526820
rect 177943 526786 177977 526820
rect 178035 526786 178069 526820
rect 178127 526786 178161 526820
rect 178219 526786 178253 526820
rect 178311 526786 178345 526820
rect 178403 526786 178437 526820
rect 178495 526786 178529 526820
rect 178587 526786 178621 526820
rect 178679 526786 178713 526820
rect 178771 526786 178805 526820
rect 178863 526786 178897 526820
rect 178955 526786 178989 526820
rect 179047 526786 179081 526820
rect 179139 526786 179173 526820
rect 179231 526786 179265 526820
rect 179323 526786 179357 526820
rect 179415 526786 179449 526820
rect 179507 526786 179541 526820
rect 179599 526786 179633 526820
rect 179691 526786 179725 526820
rect 179783 526786 179817 526820
rect 179875 526786 179909 526820
rect 179967 526786 180001 526820
rect 180059 526786 180093 526820
rect 180151 526786 180185 526820
rect 180243 526786 180277 526820
rect 180335 526786 180369 526820
rect 180427 526786 180461 526820
rect 180519 526786 180553 526820
rect 180611 526786 180645 526820
rect 180703 526786 180737 526820
rect 180795 526786 180829 526820
rect 180887 526786 180921 526820
rect 180979 526786 181013 526820
rect 181071 526786 181105 526820
rect 181163 526786 181197 526820
rect 181255 526786 181289 526820
rect 181347 526786 181381 526820
rect 181439 526786 181473 526820
rect 181531 526786 181565 526820
rect 181623 526786 181657 526820
rect 181715 526786 181749 526820
rect 181807 526786 181841 526820
rect 181899 526786 181933 526820
rect 181991 526786 182025 526820
rect 182083 526786 182117 526820
rect 182175 526786 182209 526820
rect 182267 526786 182301 526820
rect 182359 526786 182393 526820
rect 182451 526786 182485 526820
rect 182543 526786 182577 526820
rect 182635 526786 182669 526820
rect 182727 526786 182761 526820
rect 182819 526786 182853 526820
rect 182911 526786 182945 526820
rect 183003 526786 183037 526820
rect 183095 526786 183129 526820
rect 183187 526786 183221 526820
rect 183279 526786 183313 526820
rect 183371 526786 183405 526820
rect 183463 526786 183497 526820
rect 183555 526786 183589 526820
rect 183647 526786 183681 526820
rect 183739 526786 183773 526820
rect 183831 526786 183865 526820
rect 183923 526786 183957 526820
rect 184015 526786 184049 526820
rect 184107 526786 184141 526820
rect 184199 526786 184233 526820
rect 184291 526786 184325 526820
rect 184383 526786 184417 526820
rect 184475 526786 184509 526820
rect 184567 526786 184601 526820
rect 184659 526786 184693 526820
rect 184751 526786 184785 526820
rect 184843 526786 184877 526820
rect 184935 526786 184969 526820
rect 185027 526786 185061 526820
rect 185119 526786 185153 526820
rect 185211 526786 185245 526820
rect 185303 526786 185337 526820
rect 185395 526786 185429 526820
rect 185487 526786 185521 526820
rect 185579 526786 185613 526820
rect 185671 526786 185705 526820
rect 185763 526786 185797 526820
rect 185855 526786 185889 526820
rect 185947 526786 185981 526820
rect 186039 526786 186073 526820
rect 186131 526786 186165 526820
rect 186223 526786 186257 526820
rect 186315 526786 186349 526820
rect 186407 526786 186441 526820
rect 186499 526786 186533 526820
rect 186591 526786 186625 526820
rect 186683 526786 186717 526820
rect 186775 526786 186809 526820
rect 186867 526786 186901 526820
rect 186959 526786 186993 526820
rect 187051 526786 187085 526820
rect 187143 526786 187177 526820
rect 187235 526786 187269 526820
rect 187327 526786 187361 526820
rect 187419 526786 187453 526820
rect 172239 526242 172273 526276
rect 172331 526242 172365 526276
rect 172423 526242 172457 526276
rect 172515 526242 172549 526276
rect 172607 526242 172641 526276
rect 172699 526242 172733 526276
rect 172791 526242 172825 526276
rect 172883 526242 172917 526276
rect 172975 526242 173009 526276
rect 173067 526242 173101 526276
rect 173159 526242 173193 526276
rect 173251 526242 173285 526276
rect 173343 526242 173377 526276
rect 173435 526242 173469 526276
rect 173527 526242 173561 526276
rect 173619 526242 173653 526276
rect 173711 526242 173745 526276
rect 173803 526242 173837 526276
rect 173895 526242 173929 526276
rect 173987 526242 174021 526276
rect 174079 526242 174113 526276
rect 174171 526242 174205 526276
rect 174263 526242 174297 526276
rect 174355 526242 174389 526276
rect 174447 526242 174481 526276
rect 174539 526242 174573 526276
rect 174631 526242 174665 526276
rect 174723 526242 174757 526276
rect 174815 526242 174849 526276
rect 174907 526242 174941 526276
rect 174999 526242 175033 526276
rect 175091 526242 175125 526276
rect 175183 526242 175217 526276
rect 175275 526242 175309 526276
rect 175367 526242 175401 526276
rect 175459 526242 175493 526276
rect 175551 526242 175585 526276
rect 175643 526242 175677 526276
rect 175735 526242 175769 526276
rect 175827 526242 175861 526276
rect 175919 526242 175953 526276
rect 176011 526242 176045 526276
rect 176103 526242 176137 526276
rect 176195 526242 176229 526276
rect 176287 526242 176321 526276
rect 176379 526242 176413 526276
rect 176471 526242 176505 526276
rect 176563 526242 176597 526276
rect 176655 526242 176689 526276
rect 176747 526242 176781 526276
rect 176839 526242 176873 526276
rect 176931 526242 176965 526276
rect 177023 526242 177057 526276
rect 177115 526242 177149 526276
rect 177207 526242 177241 526276
rect 177299 526242 177333 526276
rect 177391 526242 177425 526276
rect 177483 526242 177517 526276
rect 177575 526242 177609 526276
rect 177667 526242 177701 526276
rect 177759 526242 177793 526276
rect 177851 526242 177885 526276
rect 177943 526242 177977 526276
rect 178035 526242 178069 526276
rect 178127 526242 178161 526276
rect 178219 526242 178253 526276
rect 178311 526242 178345 526276
rect 178403 526242 178437 526276
rect 178495 526242 178529 526276
rect 178587 526242 178621 526276
rect 178679 526242 178713 526276
rect 178771 526242 178805 526276
rect 178863 526242 178897 526276
rect 178955 526242 178989 526276
rect 179047 526242 179081 526276
rect 179139 526242 179173 526276
rect 179231 526242 179265 526276
rect 179323 526242 179357 526276
rect 179415 526242 179449 526276
rect 179507 526242 179541 526276
rect 179599 526242 179633 526276
rect 179691 526242 179725 526276
rect 179783 526242 179817 526276
rect 179875 526242 179909 526276
rect 179967 526242 180001 526276
rect 180059 526242 180093 526276
rect 180151 526242 180185 526276
rect 180243 526242 180277 526276
rect 180335 526242 180369 526276
rect 180427 526242 180461 526276
rect 180519 526242 180553 526276
rect 180611 526242 180645 526276
rect 180703 526242 180737 526276
rect 180795 526242 180829 526276
rect 180887 526242 180921 526276
rect 180979 526242 181013 526276
rect 181071 526242 181105 526276
rect 181163 526242 181197 526276
rect 181255 526242 181289 526276
rect 181347 526242 181381 526276
rect 181439 526242 181473 526276
rect 181531 526242 181565 526276
rect 181623 526242 181657 526276
rect 181715 526242 181749 526276
rect 181807 526242 181841 526276
rect 181899 526242 181933 526276
rect 181991 526242 182025 526276
rect 182083 526242 182117 526276
rect 182175 526242 182209 526276
rect 182267 526242 182301 526276
rect 182359 526242 182393 526276
rect 182451 526242 182485 526276
rect 182543 526242 182577 526276
rect 182635 526242 182669 526276
rect 182727 526242 182761 526276
rect 182819 526242 182853 526276
rect 182911 526242 182945 526276
rect 183003 526242 183037 526276
rect 183095 526242 183129 526276
rect 183187 526242 183221 526276
rect 183279 526242 183313 526276
rect 183371 526242 183405 526276
rect 183463 526242 183497 526276
rect 183555 526242 183589 526276
rect 183647 526242 183681 526276
rect 183739 526242 183773 526276
rect 183831 526242 183865 526276
rect 183923 526242 183957 526276
rect 184015 526242 184049 526276
rect 184107 526242 184141 526276
rect 184199 526242 184233 526276
rect 184291 526242 184325 526276
rect 184383 526242 184417 526276
rect 184475 526242 184509 526276
rect 184567 526242 184601 526276
rect 184659 526242 184693 526276
rect 184751 526242 184785 526276
rect 184843 526242 184877 526276
rect 184935 526242 184969 526276
rect 185027 526242 185061 526276
rect 185119 526242 185153 526276
rect 185211 526242 185245 526276
rect 185303 526242 185337 526276
rect 185395 526242 185429 526276
rect 185487 526242 185521 526276
rect 185579 526242 185613 526276
rect 185671 526242 185705 526276
rect 185763 526242 185797 526276
rect 185855 526242 185889 526276
rect 185947 526242 185981 526276
rect 186039 526242 186073 526276
rect 186131 526242 186165 526276
rect 186223 526242 186257 526276
rect 186315 526242 186349 526276
rect 186407 526242 186441 526276
rect 186499 526242 186533 526276
rect 186591 526242 186625 526276
rect 186683 526242 186717 526276
rect 186775 526242 186809 526276
rect 186867 526242 186901 526276
rect 186959 526242 186993 526276
rect 187051 526242 187085 526276
rect 187143 526242 187177 526276
rect 187235 526242 187269 526276
rect 187327 526242 187361 526276
rect 187419 526242 187453 526276
rect 172239 525698 172273 525732
rect 172331 525698 172365 525732
rect 172423 525698 172457 525732
rect 172515 525698 172549 525732
rect 172607 525698 172641 525732
rect 172699 525698 172733 525732
rect 172791 525698 172825 525732
rect 172883 525698 172917 525732
rect 172975 525698 173009 525732
rect 173067 525698 173101 525732
rect 173159 525698 173193 525732
rect 173251 525698 173285 525732
rect 173343 525698 173377 525732
rect 173435 525698 173469 525732
rect 173527 525698 173561 525732
rect 173619 525698 173653 525732
rect 173711 525698 173745 525732
rect 173803 525698 173837 525732
rect 173895 525698 173929 525732
rect 173987 525698 174021 525732
rect 174079 525698 174113 525732
rect 174171 525698 174205 525732
rect 174263 525698 174297 525732
rect 174355 525698 174389 525732
rect 174447 525698 174481 525732
rect 174539 525698 174573 525732
rect 174631 525698 174665 525732
rect 174723 525698 174757 525732
rect 174815 525698 174849 525732
rect 174907 525698 174941 525732
rect 174999 525698 175033 525732
rect 175091 525698 175125 525732
rect 175183 525698 175217 525732
rect 175275 525698 175309 525732
rect 175367 525698 175401 525732
rect 175459 525698 175493 525732
rect 175551 525698 175585 525732
rect 175643 525698 175677 525732
rect 175735 525698 175769 525732
rect 175827 525698 175861 525732
rect 175919 525698 175953 525732
rect 176011 525698 176045 525732
rect 176103 525698 176137 525732
rect 176195 525698 176229 525732
rect 176287 525698 176321 525732
rect 176379 525698 176413 525732
rect 176471 525698 176505 525732
rect 176563 525698 176597 525732
rect 176655 525698 176689 525732
rect 176747 525698 176781 525732
rect 176839 525698 176873 525732
rect 176931 525698 176965 525732
rect 177023 525698 177057 525732
rect 177115 525698 177149 525732
rect 177207 525698 177241 525732
rect 177299 525698 177333 525732
rect 177391 525698 177425 525732
rect 177483 525698 177517 525732
rect 177575 525698 177609 525732
rect 177667 525698 177701 525732
rect 177759 525698 177793 525732
rect 177851 525698 177885 525732
rect 177943 525698 177977 525732
rect 178035 525698 178069 525732
rect 178127 525698 178161 525732
rect 178219 525698 178253 525732
rect 178311 525698 178345 525732
rect 178403 525698 178437 525732
rect 178495 525698 178529 525732
rect 178587 525698 178621 525732
rect 178679 525698 178713 525732
rect 178771 525698 178805 525732
rect 178863 525698 178897 525732
rect 178955 525698 178989 525732
rect 179047 525698 179081 525732
rect 179139 525698 179173 525732
rect 179231 525698 179265 525732
rect 179323 525698 179357 525732
rect 179415 525698 179449 525732
rect 179507 525698 179541 525732
rect 179599 525698 179633 525732
rect 179691 525698 179725 525732
rect 179783 525698 179817 525732
rect 179875 525698 179909 525732
rect 179967 525698 180001 525732
rect 180059 525698 180093 525732
rect 180151 525698 180185 525732
rect 180243 525698 180277 525732
rect 180335 525698 180369 525732
rect 180427 525698 180461 525732
rect 180519 525698 180553 525732
rect 180611 525698 180645 525732
rect 180703 525698 180737 525732
rect 180795 525698 180829 525732
rect 180887 525698 180921 525732
rect 180979 525698 181013 525732
rect 181071 525698 181105 525732
rect 181163 525698 181197 525732
rect 181255 525698 181289 525732
rect 181347 525698 181381 525732
rect 181439 525698 181473 525732
rect 181531 525698 181565 525732
rect 181623 525698 181657 525732
rect 181715 525698 181749 525732
rect 181807 525698 181841 525732
rect 181899 525698 181933 525732
rect 181991 525698 182025 525732
rect 182083 525698 182117 525732
rect 182175 525698 182209 525732
rect 182267 525698 182301 525732
rect 182359 525698 182393 525732
rect 182451 525698 182485 525732
rect 182543 525698 182577 525732
rect 182635 525698 182669 525732
rect 182727 525698 182761 525732
rect 182819 525698 182853 525732
rect 182911 525698 182945 525732
rect 183003 525698 183037 525732
rect 183095 525698 183129 525732
rect 183187 525698 183221 525732
rect 183279 525698 183313 525732
rect 183371 525698 183405 525732
rect 183463 525698 183497 525732
rect 183555 525698 183589 525732
rect 183647 525698 183681 525732
rect 183739 525698 183773 525732
rect 183831 525698 183865 525732
rect 183923 525698 183957 525732
rect 184015 525698 184049 525732
rect 184107 525698 184141 525732
rect 184199 525698 184233 525732
rect 184291 525698 184325 525732
rect 184383 525698 184417 525732
rect 184475 525698 184509 525732
rect 184567 525698 184601 525732
rect 184659 525698 184693 525732
rect 184751 525698 184785 525732
rect 184843 525698 184877 525732
rect 184935 525698 184969 525732
rect 185027 525698 185061 525732
rect 185119 525698 185153 525732
rect 185211 525698 185245 525732
rect 185303 525698 185337 525732
rect 185395 525698 185429 525732
rect 185487 525698 185521 525732
rect 185579 525698 185613 525732
rect 185671 525698 185705 525732
rect 185763 525698 185797 525732
rect 185855 525698 185889 525732
rect 185947 525698 185981 525732
rect 186039 525698 186073 525732
rect 186131 525698 186165 525732
rect 186223 525698 186257 525732
rect 186315 525698 186349 525732
rect 186407 525698 186441 525732
rect 186499 525698 186533 525732
rect 186591 525698 186625 525732
rect 186683 525698 186717 525732
rect 186775 525698 186809 525732
rect 186867 525698 186901 525732
rect 186959 525698 186993 525732
rect 187051 525698 187085 525732
rect 187143 525698 187177 525732
rect 187235 525698 187269 525732
rect 187327 525698 187361 525732
rect 187419 525698 187453 525732
rect 172239 525154 172273 525188
rect 172331 525154 172365 525188
rect 172423 525154 172457 525188
rect 172515 525154 172549 525188
rect 172607 525154 172641 525188
rect 172699 525154 172733 525188
rect 172791 525154 172825 525188
rect 172883 525154 172917 525188
rect 172975 525154 173009 525188
rect 173067 525154 173101 525188
rect 173159 525154 173193 525188
rect 173251 525154 173285 525188
rect 173343 525154 173377 525188
rect 173435 525154 173469 525188
rect 173527 525154 173561 525188
rect 173619 525154 173653 525188
rect 173711 525154 173745 525188
rect 173803 525154 173837 525188
rect 173895 525154 173929 525188
rect 173987 525154 174021 525188
rect 174079 525154 174113 525188
rect 174171 525154 174205 525188
rect 174263 525154 174297 525188
rect 174355 525154 174389 525188
rect 174447 525154 174481 525188
rect 174539 525154 174573 525188
rect 174631 525154 174665 525188
rect 174723 525154 174757 525188
rect 174815 525154 174849 525188
rect 174907 525154 174941 525188
rect 174999 525154 175033 525188
rect 175091 525154 175125 525188
rect 175183 525154 175217 525188
rect 175275 525154 175309 525188
rect 175367 525154 175401 525188
rect 175459 525154 175493 525188
rect 175551 525154 175585 525188
rect 175643 525154 175677 525188
rect 175735 525154 175769 525188
rect 175827 525154 175861 525188
rect 175919 525154 175953 525188
rect 176011 525154 176045 525188
rect 176103 525154 176137 525188
rect 176195 525154 176229 525188
rect 176287 525154 176321 525188
rect 176379 525154 176413 525188
rect 176471 525154 176505 525188
rect 176563 525154 176597 525188
rect 176655 525154 176689 525188
rect 176747 525154 176781 525188
rect 176839 525154 176873 525188
rect 176931 525154 176965 525188
rect 177023 525154 177057 525188
rect 177115 525154 177149 525188
rect 177207 525154 177241 525188
rect 177299 525154 177333 525188
rect 177391 525154 177425 525188
rect 177483 525154 177517 525188
rect 177575 525154 177609 525188
rect 177667 525154 177701 525188
rect 177759 525154 177793 525188
rect 177851 525154 177885 525188
rect 177943 525154 177977 525188
rect 178035 525154 178069 525188
rect 178127 525154 178161 525188
rect 178219 525154 178253 525188
rect 178311 525154 178345 525188
rect 178403 525154 178437 525188
rect 178495 525154 178529 525188
rect 178587 525154 178621 525188
rect 178679 525154 178713 525188
rect 178771 525154 178805 525188
rect 178863 525154 178897 525188
rect 178955 525154 178989 525188
rect 179047 525154 179081 525188
rect 179139 525154 179173 525188
rect 179231 525154 179265 525188
rect 179323 525154 179357 525188
rect 179415 525154 179449 525188
rect 179507 525154 179541 525188
rect 179599 525154 179633 525188
rect 179691 525154 179725 525188
rect 179783 525154 179817 525188
rect 179875 525154 179909 525188
rect 179967 525154 180001 525188
rect 180059 525154 180093 525188
rect 180151 525154 180185 525188
rect 180243 525154 180277 525188
rect 180335 525154 180369 525188
rect 180427 525154 180461 525188
rect 180519 525154 180553 525188
rect 180611 525154 180645 525188
rect 180703 525154 180737 525188
rect 180795 525154 180829 525188
rect 180887 525154 180921 525188
rect 180979 525154 181013 525188
rect 181071 525154 181105 525188
rect 181163 525154 181197 525188
rect 181255 525154 181289 525188
rect 181347 525154 181381 525188
rect 181439 525154 181473 525188
rect 181531 525154 181565 525188
rect 181623 525154 181657 525188
rect 181715 525154 181749 525188
rect 181807 525154 181841 525188
rect 181899 525154 181933 525188
rect 181991 525154 182025 525188
rect 182083 525154 182117 525188
rect 182175 525154 182209 525188
rect 182267 525154 182301 525188
rect 182359 525154 182393 525188
rect 182451 525154 182485 525188
rect 182543 525154 182577 525188
rect 182635 525154 182669 525188
rect 182727 525154 182761 525188
rect 182819 525154 182853 525188
rect 182911 525154 182945 525188
rect 183003 525154 183037 525188
rect 183095 525154 183129 525188
rect 183187 525154 183221 525188
rect 183279 525154 183313 525188
rect 183371 525154 183405 525188
rect 183463 525154 183497 525188
rect 183555 525154 183589 525188
rect 183647 525154 183681 525188
rect 183739 525154 183773 525188
rect 183831 525154 183865 525188
rect 183923 525154 183957 525188
rect 184015 525154 184049 525188
rect 184107 525154 184141 525188
rect 184199 525154 184233 525188
rect 184291 525154 184325 525188
rect 184383 525154 184417 525188
rect 184475 525154 184509 525188
rect 184567 525154 184601 525188
rect 184659 525154 184693 525188
rect 184751 525154 184785 525188
rect 184843 525154 184877 525188
rect 184935 525154 184969 525188
rect 185027 525154 185061 525188
rect 185119 525154 185153 525188
rect 185211 525154 185245 525188
rect 185303 525154 185337 525188
rect 185395 525154 185429 525188
rect 185487 525154 185521 525188
rect 185579 525154 185613 525188
rect 185671 525154 185705 525188
rect 185763 525154 185797 525188
rect 185855 525154 185889 525188
rect 185947 525154 185981 525188
rect 186039 525154 186073 525188
rect 186131 525154 186165 525188
rect 186223 525154 186257 525188
rect 186315 525154 186349 525188
rect 186407 525154 186441 525188
rect 186499 525154 186533 525188
rect 186591 525154 186625 525188
rect 186683 525154 186717 525188
rect 186775 525154 186809 525188
rect 186867 525154 186901 525188
rect 186959 525154 186993 525188
rect 187051 525154 187085 525188
rect 187143 525154 187177 525188
rect 187235 525154 187269 525188
rect 187327 525154 187361 525188
rect 187419 525154 187453 525188
rect 172239 524610 172273 524644
rect 172331 524610 172365 524644
rect 172423 524610 172457 524644
rect 172515 524610 172549 524644
rect 172607 524610 172641 524644
rect 172699 524610 172733 524644
rect 172791 524610 172825 524644
rect 172883 524610 172917 524644
rect 172975 524610 173009 524644
rect 173067 524610 173101 524644
rect 173159 524610 173193 524644
rect 173251 524610 173285 524644
rect 173343 524610 173377 524644
rect 173435 524610 173469 524644
rect 173527 524610 173561 524644
rect 173619 524610 173653 524644
rect 173711 524610 173745 524644
rect 173803 524610 173837 524644
rect 173895 524610 173929 524644
rect 173987 524610 174021 524644
rect 174079 524610 174113 524644
rect 174171 524610 174205 524644
rect 174263 524610 174297 524644
rect 174355 524610 174389 524644
rect 174447 524610 174481 524644
rect 174539 524610 174573 524644
rect 174631 524610 174665 524644
rect 174723 524610 174757 524644
rect 174815 524610 174849 524644
rect 174907 524610 174941 524644
rect 174999 524610 175033 524644
rect 175091 524610 175125 524644
rect 175183 524610 175217 524644
rect 175275 524610 175309 524644
rect 175367 524610 175401 524644
rect 175459 524610 175493 524644
rect 175551 524610 175585 524644
rect 175643 524610 175677 524644
rect 175735 524610 175769 524644
rect 175827 524610 175861 524644
rect 175919 524610 175953 524644
rect 176011 524610 176045 524644
rect 176103 524610 176137 524644
rect 176195 524610 176229 524644
rect 176287 524610 176321 524644
rect 176379 524610 176413 524644
rect 176471 524610 176505 524644
rect 176563 524610 176597 524644
rect 176655 524610 176689 524644
rect 176747 524610 176781 524644
rect 176839 524610 176873 524644
rect 176931 524610 176965 524644
rect 177023 524610 177057 524644
rect 177115 524610 177149 524644
rect 177207 524610 177241 524644
rect 177299 524610 177333 524644
rect 177391 524610 177425 524644
rect 177483 524610 177517 524644
rect 177575 524610 177609 524644
rect 177667 524610 177701 524644
rect 177759 524610 177793 524644
rect 177851 524610 177885 524644
rect 177943 524610 177977 524644
rect 178035 524610 178069 524644
rect 178127 524610 178161 524644
rect 178219 524610 178253 524644
rect 178311 524610 178345 524644
rect 178403 524610 178437 524644
rect 178495 524610 178529 524644
rect 178587 524610 178621 524644
rect 178679 524610 178713 524644
rect 178771 524610 178805 524644
rect 178863 524610 178897 524644
rect 178955 524610 178989 524644
rect 179047 524610 179081 524644
rect 179139 524610 179173 524644
rect 179231 524610 179265 524644
rect 179323 524610 179357 524644
rect 179415 524610 179449 524644
rect 179507 524610 179541 524644
rect 179599 524610 179633 524644
rect 179691 524610 179725 524644
rect 179783 524610 179817 524644
rect 179875 524610 179909 524644
rect 179967 524610 180001 524644
rect 180059 524610 180093 524644
rect 180151 524610 180185 524644
rect 180243 524610 180277 524644
rect 180335 524610 180369 524644
rect 180427 524610 180461 524644
rect 180519 524610 180553 524644
rect 180611 524610 180645 524644
rect 180703 524610 180737 524644
rect 180795 524610 180829 524644
rect 180887 524610 180921 524644
rect 180979 524610 181013 524644
rect 181071 524610 181105 524644
rect 181163 524610 181197 524644
rect 181255 524610 181289 524644
rect 181347 524610 181381 524644
rect 181439 524610 181473 524644
rect 181531 524610 181565 524644
rect 181623 524610 181657 524644
rect 181715 524610 181749 524644
rect 181807 524610 181841 524644
rect 181899 524610 181933 524644
rect 181991 524610 182025 524644
rect 182083 524610 182117 524644
rect 182175 524610 182209 524644
rect 182267 524610 182301 524644
rect 182359 524610 182393 524644
rect 182451 524610 182485 524644
rect 182543 524610 182577 524644
rect 182635 524610 182669 524644
rect 182727 524610 182761 524644
rect 182819 524610 182853 524644
rect 182911 524610 182945 524644
rect 183003 524610 183037 524644
rect 183095 524610 183129 524644
rect 183187 524610 183221 524644
rect 183279 524610 183313 524644
rect 183371 524610 183405 524644
rect 183463 524610 183497 524644
rect 183555 524610 183589 524644
rect 183647 524610 183681 524644
rect 183739 524610 183773 524644
rect 183831 524610 183865 524644
rect 183923 524610 183957 524644
rect 184015 524610 184049 524644
rect 184107 524610 184141 524644
rect 184199 524610 184233 524644
rect 184291 524610 184325 524644
rect 184383 524610 184417 524644
rect 184475 524610 184509 524644
rect 184567 524610 184601 524644
rect 184659 524610 184693 524644
rect 184751 524610 184785 524644
rect 184843 524610 184877 524644
rect 184935 524610 184969 524644
rect 185027 524610 185061 524644
rect 185119 524610 185153 524644
rect 185211 524610 185245 524644
rect 185303 524610 185337 524644
rect 185395 524610 185429 524644
rect 185487 524610 185521 524644
rect 185579 524610 185613 524644
rect 185671 524610 185705 524644
rect 185763 524610 185797 524644
rect 185855 524610 185889 524644
rect 185947 524610 185981 524644
rect 186039 524610 186073 524644
rect 186131 524610 186165 524644
rect 186223 524610 186257 524644
rect 186315 524610 186349 524644
rect 186407 524610 186441 524644
rect 186499 524610 186533 524644
rect 186591 524610 186625 524644
rect 186683 524610 186717 524644
rect 186775 524610 186809 524644
rect 186867 524610 186901 524644
rect 186959 524610 186993 524644
rect 187051 524610 187085 524644
rect 187143 524610 187177 524644
rect 187235 524610 187269 524644
rect 187327 524610 187361 524644
rect 187419 524610 187453 524644
rect 172239 524066 172273 524100
rect 172331 524066 172365 524100
rect 172423 524066 172457 524100
rect 172515 524066 172549 524100
rect 172607 524066 172641 524100
rect 172699 524066 172733 524100
rect 172791 524066 172825 524100
rect 172883 524066 172917 524100
rect 172975 524066 173009 524100
rect 173067 524066 173101 524100
rect 173159 524066 173193 524100
rect 173251 524066 173285 524100
rect 173343 524066 173377 524100
rect 173435 524066 173469 524100
rect 173527 524066 173561 524100
rect 173619 524066 173653 524100
rect 173711 524066 173745 524100
rect 173803 524066 173837 524100
rect 173895 524066 173929 524100
rect 173987 524066 174021 524100
rect 174079 524066 174113 524100
rect 174171 524066 174205 524100
rect 174263 524066 174297 524100
rect 174355 524066 174389 524100
rect 174447 524066 174481 524100
rect 174539 524066 174573 524100
rect 174631 524066 174665 524100
rect 174723 524066 174757 524100
rect 174815 524066 174849 524100
rect 174907 524066 174941 524100
rect 174999 524066 175033 524100
rect 175091 524066 175125 524100
rect 175183 524066 175217 524100
rect 175275 524066 175309 524100
rect 175367 524066 175401 524100
rect 175459 524066 175493 524100
rect 175551 524066 175585 524100
rect 175643 524066 175677 524100
rect 175735 524066 175769 524100
rect 175827 524066 175861 524100
rect 175919 524066 175953 524100
rect 176011 524066 176045 524100
rect 176103 524066 176137 524100
rect 176195 524066 176229 524100
rect 176287 524066 176321 524100
rect 176379 524066 176413 524100
rect 176471 524066 176505 524100
rect 176563 524066 176597 524100
rect 176655 524066 176689 524100
rect 176747 524066 176781 524100
rect 176839 524066 176873 524100
rect 176931 524066 176965 524100
rect 177023 524066 177057 524100
rect 177115 524066 177149 524100
rect 177207 524066 177241 524100
rect 177299 524066 177333 524100
rect 177391 524066 177425 524100
rect 177483 524066 177517 524100
rect 177575 524066 177609 524100
rect 177667 524066 177701 524100
rect 177759 524066 177793 524100
rect 177851 524066 177885 524100
rect 177943 524066 177977 524100
rect 178035 524066 178069 524100
rect 178127 524066 178161 524100
rect 178219 524066 178253 524100
rect 178311 524066 178345 524100
rect 178403 524066 178437 524100
rect 178495 524066 178529 524100
rect 178587 524066 178621 524100
rect 178679 524066 178713 524100
rect 178771 524066 178805 524100
rect 178863 524066 178897 524100
rect 178955 524066 178989 524100
rect 179047 524066 179081 524100
rect 179139 524066 179173 524100
rect 179231 524066 179265 524100
rect 179323 524066 179357 524100
rect 179415 524066 179449 524100
rect 179507 524066 179541 524100
rect 179599 524066 179633 524100
rect 179691 524066 179725 524100
rect 179783 524066 179817 524100
rect 179875 524066 179909 524100
rect 179967 524066 180001 524100
rect 180059 524066 180093 524100
rect 180151 524066 180185 524100
rect 180243 524066 180277 524100
rect 180335 524066 180369 524100
rect 180427 524066 180461 524100
rect 180519 524066 180553 524100
rect 180611 524066 180645 524100
rect 180703 524066 180737 524100
rect 180795 524066 180829 524100
rect 180887 524066 180921 524100
rect 180979 524066 181013 524100
rect 181071 524066 181105 524100
rect 181163 524066 181197 524100
rect 181255 524066 181289 524100
rect 181347 524066 181381 524100
rect 181439 524066 181473 524100
rect 181531 524066 181565 524100
rect 181623 524066 181657 524100
rect 181715 524066 181749 524100
rect 181807 524066 181841 524100
rect 181899 524066 181933 524100
rect 181991 524066 182025 524100
rect 182083 524066 182117 524100
rect 182175 524066 182209 524100
rect 182267 524066 182301 524100
rect 182359 524066 182393 524100
rect 182451 524066 182485 524100
rect 182543 524066 182577 524100
rect 182635 524066 182669 524100
rect 182727 524066 182761 524100
rect 182819 524066 182853 524100
rect 182911 524066 182945 524100
rect 183003 524066 183037 524100
rect 183095 524066 183129 524100
rect 183187 524066 183221 524100
rect 183279 524066 183313 524100
rect 183371 524066 183405 524100
rect 183463 524066 183497 524100
rect 183555 524066 183589 524100
rect 183647 524066 183681 524100
rect 183739 524066 183773 524100
rect 183831 524066 183865 524100
rect 183923 524066 183957 524100
rect 184015 524066 184049 524100
rect 184107 524066 184141 524100
rect 184199 524066 184233 524100
rect 184291 524066 184325 524100
rect 184383 524066 184417 524100
rect 184475 524066 184509 524100
rect 184567 524066 184601 524100
rect 184659 524066 184693 524100
rect 184751 524066 184785 524100
rect 184843 524066 184877 524100
rect 184935 524066 184969 524100
rect 185027 524066 185061 524100
rect 185119 524066 185153 524100
rect 185211 524066 185245 524100
rect 185303 524066 185337 524100
rect 185395 524066 185429 524100
rect 185487 524066 185521 524100
rect 185579 524066 185613 524100
rect 185671 524066 185705 524100
rect 185763 524066 185797 524100
rect 185855 524066 185889 524100
rect 185947 524066 185981 524100
rect 186039 524066 186073 524100
rect 186131 524066 186165 524100
rect 186223 524066 186257 524100
rect 186315 524066 186349 524100
rect 186407 524066 186441 524100
rect 186499 524066 186533 524100
rect 186591 524066 186625 524100
rect 186683 524066 186717 524100
rect 186775 524066 186809 524100
rect 186867 524066 186901 524100
rect 186959 524066 186993 524100
rect 187051 524066 187085 524100
rect 187143 524066 187177 524100
rect 187235 524066 187269 524100
rect 187327 524066 187361 524100
rect 187419 524066 187453 524100
rect 172239 523522 172273 523556
rect 172331 523522 172365 523556
rect 172423 523522 172457 523556
rect 172515 523522 172549 523556
rect 172607 523522 172641 523556
rect 172699 523522 172733 523556
rect 172791 523522 172825 523556
rect 172883 523522 172917 523556
rect 172975 523522 173009 523556
rect 173067 523522 173101 523556
rect 173159 523522 173193 523556
rect 173251 523522 173285 523556
rect 173343 523522 173377 523556
rect 173435 523522 173469 523556
rect 173527 523522 173561 523556
rect 173619 523522 173653 523556
rect 173711 523522 173745 523556
rect 173803 523522 173837 523556
rect 173895 523522 173929 523556
rect 173987 523522 174021 523556
rect 174079 523522 174113 523556
rect 174171 523522 174205 523556
rect 174263 523522 174297 523556
rect 174355 523522 174389 523556
rect 174447 523522 174481 523556
rect 174539 523522 174573 523556
rect 174631 523522 174665 523556
rect 174723 523522 174757 523556
rect 174815 523522 174849 523556
rect 174907 523522 174941 523556
rect 174999 523522 175033 523556
rect 175091 523522 175125 523556
rect 175183 523522 175217 523556
rect 175275 523522 175309 523556
rect 175367 523522 175401 523556
rect 175459 523522 175493 523556
rect 175551 523522 175585 523556
rect 175643 523522 175677 523556
rect 175735 523522 175769 523556
rect 175827 523522 175861 523556
rect 175919 523522 175953 523556
rect 176011 523522 176045 523556
rect 176103 523522 176137 523556
rect 176195 523522 176229 523556
rect 176287 523522 176321 523556
rect 176379 523522 176413 523556
rect 176471 523522 176505 523556
rect 176563 523522 176597 523556
rect 176655 523522 176689 523556
rect 176747 523522 176781 523556
rect 176839 523522 176873 523556
rect 176931 523522 176965 523556
rect 177023 523522 177057 523556
rect 177115 523522 177149 523556
rect 177207 523522 177241 523556
rect 177299 523522 177333 523556
rect 177391 523522 177425 523556
rect 177483 523522 177517 523556
rect 177575 523522 177609 523556
rect 177667 523522 177701 523556
rect 177759 523522 177793 523556
rect 177851 523522 177885 523556
rect 177943 523522 177977 523556
rect 178035 523522 178069 523556
rect 178127 523522 178161 523556
rect 178219 523522 178253 523556
rect 178311 523522 178345 523556
rect 178403 523522 178437 523556
rect 178495 523522 178529 523556
rect 178587 523522 178621 523556
rect 178679 523522 178713 523556
rect 178771 523522 178805 523556
rect 178863 523522 178897 523556
rect 178955 523522 178989 523556
rect 179047 523522 179081 523556
rect 179139 523522 179173 523556
rect 179231 523522 179265 523556
rect 179323 523522 179357 523556
rect 179415 523522 179449 523556
rect 179507 523522 179541 523556
rect 179599 523522 179633 523556
rect 179691 523522 179725 523556
rect 179783 523522 179817 523556
rect 179875 523522 179909 523556
rect 179967 523522 180001 523556
rect 180059 523522 180093 523556
rect 180151 523522 180185 523556
rect 180243 523522 180277 523556
rect 180335 523522 180369 523556
rect 180427 523522 180461 523556
rect 180519 523522 180553 523556
rect 180611 523522 180645 523556
rect 180703 523522 180737 523556
rect 180795 523522 180829 523556
rect 180887 523522 180921 523556
rect 180979 523522 181013 523556
rect 181071 523522 181105 523556
rect 181163 523522 181197 523556
rect 181255 523522 181289 523556
rect 181347 523522 181381 523556
rect 181439 523522 181473 523556
rect 181531 523522 181565 523556
rect 181623 523522 181657 523556
rect 181715 523522 181749 523556
rect 181807 523522 181841 523556
rect 181899 523522 181933 523556
rect 181991 523522 182025 523556
rect 182083 523522 182117 523556
rect 182175 523522 182209 523556
rect 182267 523522 182301 523556
rect 182359 523522 182393 523556
rect 182451 523522 182485 523556
rect 182543 523522 182577 523556
rect 182635 523522 182669 523556
rect 182727 523522 182761 523556
rect 182819 523522 182853 523556
rect 182911 523522 182945 523556
rect 183003 523522 183037 523556
rect 183095 523522 183129 523556
rect 183187 523522 183221 523556
rect 183279 523522 183313 523556
rect 183371 523522 183405 523556
rect 183463 523522 183497 523556
rect 183555 523522 183589 523556
rect 183647 523522 183681 523556
rect 183739 523522 183773 523556
rect 183831 523522 183865 523556
rect 183923 523522 183957 523556
rect 184015 523522 184049 523556
rect 184107 523522 184141 523556
rect 184199 523522 184233 523556
rect 184291 523522 184325 523556
rect 184383 523522 184417 523556
rect 184475 523522 184509 523556
rect 184567 523522 184601 523556
rect 184659 523522 184693 523556
rect 184751 523522 184785 523556
rect 184843 523522 184877 523556
rect 184935 523522 184969 523556
rect 185027 523522 185061 523556
rect 185119 523522 185153 523556
rect 185211 523522 185245 523556
rect 185303 523522 185337 523556
rect 185395 523522 185429 523556
rect 185487 523522 185521 523556
rect 185579 523522 185613 523556
rect 185671 523522 185705 523556
rect 185763 523522 185797 523556
rect 185855 523522 185889 523556
rect 185947 523522 185981 523556
rect 186039 523522 186073 523556
rect 186131 523522 186165 523556
rect 186223 523522 186257 523556
rect 186315 523522 186349 523556
rect 186407 523522 186441 523556
rect 186499 523522 186533 523556
rect 186591 523522 186625 523556
rect 186683 523522 186717 523556
rect 186775 523522 186809 523556
rect 186867 523522 186901 523556
rect 186959 523522 186993 523556
rect 187051 523522 187085 523556
rect 187143 523522 187177 523556
rect 187235 523522 187269 523556
rect 187327 523522 187361 523556
rect 187419 523522 187453 523556
rect 172239 522978 172273 523012
rect 172331 522978 172365 523012
rect 172423 522978 172457 523012
rect 172515 522978 172549 523012
rect 172607 522978 172641 523012
rect 172699 522978 172733 523012
rect 172791 522978 172825 523012
rect 172883 522978 172917 523012
rect 172975 522978 173009 523012
rect 173067 522978 173101 523012
rect 173159 522978 173193 523012
rect 173251 522978 173285 523012
rect 173343 522978 173377 523012
rect 173435 522978 173469 523012
rect 173527 522978 173561 523012
rect 173619 522978 173653 523012
rect 173711 522978 173745 523012
rect 173803 522978 173837 523012
rect 173895 522978 173929 523012
rect 173987 522978 174021 523012
rect 174079 522978 174113 523012
rect 174171 522978 174205 523012
rect 174263 522978 174297 523012
rect 174355 522978 174389 523012
rect 174447 522978 174481 523012
rect 174539 522978 174573 523012
rect 174631 522978 174665 523012
rect 174723 522978 174757 523012
rect 174815 522978 174849 523012
rect 174907 522978 174941 523012
rect 174999 522978 175033 523012
rect 175091 522978 175125 523012
rect 175183 522978 175217 523012
rect 175275 522978 175309 523012
rect 175367 522978 175401 523012
rect 175459 522978 175493 523012
rect 175551 522978 175585 523012
rect 175643 522978 175677 523012
rect 175735 522978 175769 523012
rect 175827 522978 175861 523012
rect 175919 522978 175953 523012
rect 176011 522978 176045 523012
rect 176103 522978 176137 523012
rect 176195 522978 176229 523012
rect 176287 522978 176321 523012
rect 176379 522978 176413 523012
rect 176471 522978 176505 523012
rect 176563 522978 176597 523012
rect 176655 522978 176689 523012
rect 176747 522978 176781 523012
rect 176839 522978 176873 523012
rect 176931 522978 176965 523012
rect 177023 522978 177057 523012
rect 177115 522978 177149 523012
rect 177207 522978 177241 523012
rect 177299 522978 177333 523012
rect 177391 522978 177425 523012
rect 177483 522978 177517 523012
rect 177575 522978 177609 523012
rect 177667 522978 177701 523012
rect 177759 522978 177793 523012
rect 177851 522978 177885 523012
rect 177943 522978 177977 523012
rect 178035 522978 178069 523012
rect 178127 522978 178161 523012
rect 178219 522978 178253 523012
rect 178311 522978 178345 523012
rect 178403 522978 178437 523012
rect 178495 522978 178529 523012
rect 178587 522978 178621 523012
rect 178679 522978 178713 523012
rect 178771 522978 178805 523012
rect 178863 522978 178897 523012
rect 178955 522978 178989 523012
rect 179047 522978 179081 523012
rect 179139 522978 179173 523012
rect 179231 522978 179265 523012
rect 179323 522978 179357 523012
rect 179415 522978 179449 523012
rect 179507 522978 179541 523012
rect 179599 522978 179633 523012
rect 179691 522978 179725 523012
rect 179783 522978 179817 523012
rect 179875 522978 179909 523012
rect 179967 522978 180001 523012
rect 180059 522978 180093 523012
rect 180151 522978 180185 523012
rect 180243 522978 180277 523012
rect 180335 522978 180369 523012
rect 180427 522978 180461 523012
rect 180519 522978 180553 523012
rect 180611 522978 180645 523012
rect 180703 522978 180737 523012
rect 180795 522978 180829 523012
rect 180887 522978 180921 523012
rect 180979 522978 181013 523012
rect 181071 522978 181105 523012
rect 181163 522978 181197 523012
rect 181255 522978 181289 523012
rect 181347 522978 181381 523012
rect 181439 522978 181473 523012
rect 181531 522978 181565 523012
rect 181623 522978 181657 523012
rect 181715 522978 181749 523012
rect 181807 522978 181841 523012
rect 181899 522978 181933 523012
rect 181991 522978 182025 523012
rect 182083 522978 182117 523012
rect 182175 522978 182209 523012
rect 182267 522978 182301 523012
rect 182359 522978 182393 523012
rect 182451 522978 182485 523012
rect 182543 522978 182577 523012
rect 182635 522978 182669 523012
rect 182727 522978 182761 523012
rect 182819 522978 182853 523012
rect 182911 522978 182945 523012
rect 183003 522978 183037 523012
rect 183095 522978 183129 523012
rect 183187 522978 183221 523012
rect 183279 522978 183313 523012
rect 183371 522978 183405 523012
rect 183463 522978 183497 523012
rect 183555 522978 183589 523012
rect 183647 522978 183681 523012
rect 183739 522978 183773 523012
rect 183831 522978 183865 523012
rect 183923 522978 183957 523012
rect 184015 522978 184049 523012
rect 184107 522978 184141 523012
rect 184199 522978 184233 523012
rect 184291 522978 184325 523012
rect 184383 522978 184417 523012
rect 184475 522978 184509 523012
rect 184567 522978 184601 523012
rect 184659 522978 184693 523012
rect 184751 522978 184785 523012
rect 184843 522978 184877 523012
rect 184935 522978 184969 523012
rect 185027 522978 185061 523012
rect 185119 522978 185153 523012
rect 185211 522978 185245 523012
rect 185303 522978 185337 523012
rect 185395 522978 185429 523012
rect 185487 522978 185521 523012
rect 185579 522978 185613 523012
rect 185671 522978 185705 523012
rect 185763 522978 185797 523012
rect 185855 522978 185889 523012
rect 185947 522978 185981 523012
rect 186039 522978 186073 523012
rect 186131 522978 186165 523012
rect 186223 522978 186257 523012
rect 186315 522978 186349 523012
rect 186407 522978 186441 523012
rect 186499 522978 186533 523012
rect 186591 522978 186625 523012
rect 186683 522978 186717 523012
rect 186775 522978 186809 523012
rect 186867 522978 186901 523012
rect 186959 522978 186993 523012
rect 187051 522978 187085 523012
rect 187143 522978 187177 523012
rect 187235 522978 187269 523012
rect 187327 522978 187361 523012
rect 187419 522978 187453 523012
rect 172239 522434 172273 522468
rect 172331 522434 172365 522468
rect 172423 522434 172457 522468
rect 172515 522434 172549 522468
rect 172607 522434 172641 522468
rect 172699 522434 172733 522468
rect 172791 522434 172825 522468
rect 172883 522434 172917 522468
rect 172975 522434 173009 522468
rect 173067 522434 173101 522468
rect 173159 522434 173193 522468
rect 173251 522434 173285 522468
rect 173343 522434 173377 522468
rect 173435 522434 173469 522468
rect 173527 522434 173561 522468
rect 173619 522434 173653 522468
rect 173711 522434 173745 522468
rect 173803 522434 173837 522468
rect 173895 522434 173929 522468
rect 173987 522434 174021 522468
rect 174079 522434 174113 522468
rect 174171 522434 174205 522468
rect 174263 522434 174297 522468
rect 174355 522434 174389 522468
rect 174447 522434 174481 522468
rect 174539 522434 174573 522468
rect 174631 522434 174665 522468
rect 174723 522434 174757 522468
rect 174815 522434 174849 522468
rect 174907 522434 174941 522468
rect 174999 522434 175033 522468
rect 175091 522434 175125 522468
rect 175183 522434 175217 522468
rect 175275 522434 175309 522468
rect 175367 522434 175401 522468
rect 175459 522434 175493 522468
rect 175551 522434 175585 522468
rect 175643 522434 175677 522468
rect 175735 522434 175769 522468
rect 175827 522434 175861 522468
rect 175919 522434 175953 522468
rect 176011 522434 176045 522468
rect 176103 522434 176137 522468
rect 176195 522434 176229 522468
rect 176287 522434 176321 522468
rect 176379 522434 176413 522468
rect 176471 522434 176505 522468
rect 176563 522434 176597 522468
rect 176655 522434 176689 522468
rect 176747 522434 176781 522468
rect 176839 522434 176873 522468
rect 176931 522434 176965 522468
rect 177023 522434 177057 522468
rect 177115 522434 177149 522468
rect 177207 522434 177241 522468
rect 177299 522434 177333 522468
rect 177391 522434 177425 522468
rect 177483 522434 177517 522468
rect 177575 522434 177609 522468
rect 177667 522434 177701 522468
rect 177759 522434 177793 522468
rect 177851 522434 177885 522468
rect 177943 522434 177977 522468
rect 178035 522434 178069 522468
rect 178127 522434 178161 522468
rect 178219 522434 178253 522468
rect 178311 522434 178345 522468
rect 178403 522434 178437 522468
rect 178495 522434 178529 522468
rect 178587 522434 178621 522468
rect 178679 522434 178713 522468
rect 178771 522434 178805 522468
rect 178863 522434 178897 522468
rect 178955 522434 178989 522468
rect 179047 522434 179081 522468
rect 179139 522434 179173 522468
rect 179231 522434 179265 522468
rect 179323 522434 179357 522468
rect 179415 522434 179449 522468
rect 179507 522434 179541 522468
rect 179599 522434 179633 522468
rect 179691 522434 179725 522468
rect 179783 522434 179817 522468
rect 179875 522434 179909 522468
rect 179967 522434 180001 522468
rect 180059 522434 180093 522468
rect 180151 522434 180185 522468
rect 180243 522434 180277 522468
rect 180335 522434 180369 522468
rect 180427 522434 180461 522468
rect 180519 522434 180553 522468
rect 180611 522434 180645 522468
rect 180703 522434 180737 522468
rect 180795 522434 180829 522468
rect 180887 522434 180921 522468
rect 180979 522434 181013 522468
rect 181071 522434 181105 522468
rect 181163 522434 181197 522468
rect 181255 522434 181289 522468
rect 181347 522434 181381 522468
rect 181439 522434 181473 522468
rect 181531 522434 181565 522468
rect 181623 522434 181657 522468
rect 181715 522434 181749 522468
rect 181807 522434 181841 522468
rect 181899 522434 181933 522468
rect 181991 522434 182025 522468
rect 182083 522434 182117 522468
rect 182175 522434 182209 522468
rect 182267 522434 182301 522468
rect 182359 522434 182393 522468
rect 182451 522434 182485 522468
rect 182543 522434 182577 522468
rect 182635 522434 182669 522468
rect 182727 522434 182761 522468
rect 182819 522434 182853 522468
rect 182911 522434 182945 522468
rect 183003 522434 183037 522468
rect 183095 522434 183129 522468
rect 183187 522434 183221 522468
rect 183279 522434 183313 522468
rect 183371 522434 183405 522468
rect 183463 522434 183497 522468
rect 183555 522434 183589 522468
rect 183647 522434 183681 522468
rect 183739 522434 183773 522468
rect 183831 522434 183865 522468
rect 183923 522434 183957 522468
rect 184015 522434 184049 522468
rect 184107 522434 184141 522468
rect 184199 522434 184233 522468
rect 184291 522434 184325 522468
rect 184383 522434 184417 522468
rect 184475 522434 184509 522468
rect 184567 522434 184601 522468
rect 184659 522434 184693 522468
rect 184751 522434 184785 522468
rect 184843 522434 184877 522468
rect 184935 522434 184969 522468
rect 185027 522434 185061 522468
rect 185119 522434 185153 522468
rect 185211 522434 185245 522468
rect 185303 522434 185337 522468
rect 185395 522434 185429 522468
rect 185487 522434 185521 522468
rect 185579 522434 185613 522468
rect 185671 522434 185705 522468
rect 185763 522434 185797 522468
rect 185855 522434 185889 522468
rect 185947 522434 185981 522468
rect 186039 522434 186073 522468
rect 186131 522434 186165 522468
rect 186223 522434 186257 522468
rect 186315 522434 186349 522468
rect 186407 522434 186441 522468
rect 186499 522434 186533 522468
rect 186591 522434 186625 522468
rect 186683 522434 186717 522468
rect 186775 522434 186809 522468
rect 186867 522434 186901 522468
rect 186959 522434 186993 522468
rect 187051 522434 187085 522468
rect 187143 522434 187177 522468
rect 187235 522434 187269 522468
rect 187327 522434 187361 522468
rect 187419 522434 187453 522468
rect 172239 521890 172273 521924
rect 172331 521890 172365 521924
rect 172423 521890 172457 521924
rect 172515 521890 172549 521924
rect 172607 521890 172641 521924
rect 172699 521890 172733 521924
rect 172791 521890 172825 521924
rect 172883 521890 172917 521924
rect 172975 521890 173009 521924
rect 173067 521890 173101 521924
rect 173159 521890 173193 521924
rect 173251 521890 173285 521924
rect 173343 521890 173377 521924
rect 173435 521890 173469 521924
rect 173527 521890 173561 521924
rect 173619 521890 173653 521924
rect 173711 521890 173745 521924
rect 173803 521890 173837 521924
rect 173895 521890 173929 521924
rect 173987 521890 174021 521924
rect 174079 521890 174113 521924
rect 174171 521890 174205 521924
rect 174263 521890 174297 521924
rect 174355 521890 174389 521924
rect 174447 521890 174481 521924
rect 174539 521890 174573 521924
rect 174631 521890 174665 521924
rect 174723 521890 174757 521924
rect 174815 521890 174849 521924
rect 174907 521890 174941 521924
rect 174999 521890 175033 521924
rect 175091 521890 175125 521924
rect 175183 521890 175217 521924
rect 175275 521890 175309 521924
rect 175367 521890 175401 521924
rect 175459 521890 175493 521924
rect 175551 521890 175585 521924
rect 175643 521890 175677 521924
rect 175735 521890 175769 521924
rect 175827 521890 175861 521924
rect 175919 521890 175953 521924
rect 176011 521890 176045 521924
rect 176103 521890 176137 521924
rect 176195 521890 176229 521924
rect 176287 521890 176321 521924
rect 176379 521890 176413 521924
rect 176471 521890 176505 521924
rect 176563 521890 176597 521924
rect 176655 521890 176689 521924
rect 176747 521890 176781 521924
rect 176839 521890 176873 521924
rect 176931 521890 176965 521924
rect 177023 521890 177057 521924
rect 177115 521890 177149 521924
rect 177207 521890 177241 521924
rect 177299 521890 177333 521924
rect 177391 521890 177425 521924
rect 177483 521890 177517 521924
rect 177575 521890 177609 521924
rect 177667 521890 177701 521924
rect 177759 521890 177793 521924
rect 177851 521890 177885 521924
rect 177943 521890 177977 521924
rect 178035 521890 178069 521924
rect 178127 521890 178161 521924
rect 178219 521890 178253 521924
rect 178311 521890 178345 521924
rect 178403 521890 178437 521924
rect 178495 521890 178529 521924
rect 178587 521890 178621 521924
rect 178679 521890 178713 521924
rect 178771 521890 178805 521924
rect 178863 521890 178897 521924
rect 178955 521890 178989 521924
rect 179047 521890 179081 521924
rect 179139 521890 179173 521924
rect 179231 521890 179265 521924
rect 179323 521890 179357 521924
rect 179415 521890 179449 521924
rect 179507 521890 179541 521924
rect 179599 521890 179633 521924
rect 179691 521890 179725 521924
rect 179783 521890 179817 521924
rect 179875 521890 179909 521924
rect 179967 521890 180001 521924
rect 180059 521890 180093 521924
rect 180151 521890 180185 521924
rect 180243 521890 180277 521924
rect 180335 521890 180369 521924
rect 180427 521890 180461 521924
rect 180519 521890 180553 521924
rect 180611 521890 180645 521924
rect 180703 521890 180737 521924
rect 180795 521890 180829 521924
rect 180887 521890 180921 521924
rect 180979 521890 181013 521924
rect 181071 521890 181105 521924
rect 181163 521890 181197 521924
rect 181255 521890 181289 521924
rect 181347 521890 181381 521924
rect 181439 521890 181473 521924
rect 181531 521890 181565 521924
rect 181623 521890 181657 521924
rect 181715 521890 181749 521924
rect 181807 521890 181841 521924
rect 181899 521890 181933 521924
rect 181991 521890 182025 521924
rect 182083 521890 182117 521924
rect 182175 521890 182209 521924
rect 182267 521890 182301 521924
rect 182359 521890 182393 521924
rect 182451 521890 182485 521924
rect 182543 521890 182577 521924
rect 182635 521890 182669 521924
rect 182727 521890 182761 521924
rect 182819 521890 182853 521924
rect 182911 521890 182945 521924
rect 183003 521890 183037 521924
rect 183095 521890 183129 521924
rect 183187 521890 183221 521924
rect 183279 521890 183313 521924
rect 183371 521890 183405 521924
rect 183463 521890 183497 521924
rect 183555 521890 183589 521924
rect 183647 521890 183681 521924
rect 183739 521890 183773 521924
rect 183831 521890 183865 521924
rect 183923 521890 183957 521924
rect 184015 521890 184049 521924
rect 184107 521890 184141 521924
rect 184199 521890 184233 521924
rect 184291 521890 184325 521924
rect 184383 521890 184417 521924
rect 184475 521890 184509 521924
rect 184567 521890 184601 521924
rect 184659 521890 184693 521924
rect 184751 521890 184785 521924
rect 184843 521890 184877 521924
rect 184935 521890 184969 521924
rect 185027 521890 185061 521924
rect 185119 521890 185153 521924
rect 185211 521890 185245 521924
rect 185303 521890 185337 521924
rect 185395 521890 185429 521924
rect 185487 521890 185521 521924
rect 185579 521890 185613 521924
rect 185671 521890 185705 521924
rect 185763 521890 185797 521924
rect 185855 521890 185889 521924
rect 185947 521890 185981 521924
rect 186039 521890 186073 521924
rect 186131 521890 186165 521924
rect 186223 521890 186257 521924
rect 186315 521890 186349 521924
rect 186407 521890 186441 521924
rect 186499 521890 186533 521924
rect 186591 521890 186625 521924
rect 186683 521890 186717 521924
rect 186775 521890 186809 521924
rect 186867 521890 186901 521924
rect 186959 521890 186993 521924
rect 187051 521890 187085 521924
rect 187143 521890 187177 521924
rect 187235 521890 187269 521924
rect 187327 521890 187361 521924
rect 187419 521890 187453 521924
rect 172239 521346 172273 521380
rect 172331 521346 172365 521380
rect 172423 521346 172457 521380
rect 172515 521346 172549 521380
rect 172607 521346 172641 521380
rect 172699 521346 172733 521380
rect 172791 521346 172825 521380
rect 172883 521346 172917 521380
rect 172975 521346 173009 521380
rect 173067 521346 173101 521380
rect 173159 521346 173193 521380
rect 173251 521346 173285 521380
rect 173343 521346 173377 521380
rect 173435 521346 173469 521380
rect 173527 521346 173561 521380
rect 173619 521346 173653 521380
rect 173711 521346 173745 521380
rect 173803 521346 173837 521380
rect 173895 521346 173929 521380
rect 173987 521346 174021 521380
rect 174079 521346 174113 521380
rect 174171 521346 174205 521380
rect 174263 521346 174297 521380
rect 174355 521346 174389 521380
rect 174447 521346 174481 521380
rect 174539 521346 174573 521380
rect 174631 521346 174665 521380
rect 174723 521346 174757 521380
rect 174815 521346 174849 521380
rect 174907 521346 174941 521380
rect 174999 521346 175033 521380
rect 175091 521346 175125 521380
rect 175183 521346 175217 521380
rect 175275 521346 175309 521380
rect 175367 521346 175401 521380
rect 175459 521346 175493 521380
rect 175551 521346 175585 521380
rect 175643 521346 175677 521380
rect 175735 521346 175769 521380
rect 175827 521346 175861 521380
rect 175919 521346 175953 521380
rect 176011 521346 176045 521380
rect 176103 521346 176137 521380
rect 176195 521346 176229 521380
rect 176287 521346 176321 521380
rect 176379 521346 176413 521380
rect 176471 521346 176505 521380
rect 176563 521346 176597 521380
rect 176655 521346 176689 521380
rect 176747 521346 176781 521380
rect 176839 521346 176873 521380
rect 176931 521346 176965 521380
rect 177023 521346 177057 521380
rect 177115 521346 177149 521380
rect 177207 521346 177241 521380
rect 177299 521346 177333 521380
rect 177391 521346 177425 521380
rect 177483 521346 177517 521380
rect 177575 521346 177609 521380
rect 177667 521346 177701 521380
rect 177759 521346 177793 521380
rect 177851 521346 177885 521380
rect 177943 521346 177977 521380
rect 178035 521346 178069 521380
rect 178127 521346 178161 521380
rect 178219 521346 178253 521380
rect 178311 521346 178345 521380
rect 178403 521346 178437 521380
rect 178495 521346 178529 521380
rect 178587 521346 178621 521380
rect 178679 521346 178713 521380
rect 178771 521346 178805 521380
rect 178863 521346 178897 521380
rect 178955 521346 178989 521380
rect 179047 521346 179081 521380
rect 179139 521346 179173 521380
rect 179231 521346 179265 521380
rect 179323 521346 179357 521380
rect 179415 521346 179449 521380
rect 179507 521346 179541 521380
rect 179599 521346 179633 521380
rect 179691 521346 179725 521380
rect 179783 521346 179817 521380
rect 179875 521346 179909 521380
rect 179967 521346 180001 521380
rect 180059 521346 180093 521380
rect 180151 521346 180185 521380
rect 180243 521346 180277 521380
rect 180335 521346 180369 521380
rect 180427 521346 180461 521380
rect 180519 521346 180553 521380
rect 180611 521346 180645 521380
rect 180703 521346 180737 521380
rect 180795 521346 180829 521380
rect 180887 521346 180921 521380
rect 180979 521346 181013 521380
rect 181071 521346 181105 521380
rect 181163 521346 181197 521380
rect 181255 521346 181289 521380
rect 181347 521346 181381 521380
rect 181439 521346 181473 521380
rect 181531 521346 181565 521380
rect 181623 521346 181657 521380
rect 181715 521346 181749 521380
rect 181807 521346 181841 521380
rect 181899 521346 181933 521380
rect 181991 521346 182025 521380
rect 182083 521346 182117 521380
rect 182175 521346 182209 521380
rect 182267 521346 182301 521380
rect 182359 521346 182393 521380
rect 182451 521346 182485 521380
rect 182543 521346 182577 521380
rect 182635 521346 182669 521380
rect 182727 521346 182761 521380
rect 182819 521346 182853 521380
rect 182911 521346 182945 521380
rect 183003 521346 183037 521380
rect 183095 521346 183129 521380
rect 183187 521346 183221 521380
rect 183279 521346 183313 521380
rect 183371 521346 183405 521380
rect 183463 521346 183497 521380
rect 183555 521346 183589 521380
rect 183647 521346 183681 521380
rect 183739 521346 183773 521380
rect 183831 521346 183865 521380
rect 183923 521346 183957 521380
rect 184015 521346 184049 521380
rect 184107 521346 184141 521380
rect 184199 521346 184233 521380
rect 184291 521346 184325 521380
rect 184383 521346 184417 521380
rect 184475 521346 184509 521380
rect 184567 521346 184601 521380
rect 184659 521346 184693 521380
rect 184751 521346 184785 521380
rect 184843 521346 184877 521380
rect 184935 521346 184969 521380
rect 185027 521346 185061 521380
rect 185119 521346 185153 521380
rect 185211 521346 185245 521380
rect 185303 521346 185337 521380
rect 185395 521346 185429 521380
rect 185487 521346 185521 521380
rect 185579 521346 185613 521380
rect 185671 521346 185705 521380
rect 185763 521346 185797 521380
rect 185855 521346 185889 521380
rect 185947 521346 185981 521380
rect 186039 521346 186073 521380
rect 186131 521346 186165 521380
rect 186223 521346 186257 521380
rect 186315 521346 186349 521380
rect 186407 521346 186441 521380
rect 186499 521346 186533 521380
rect 186591 521346 186625 521380
rect 186683 521346 186717 521380
rect 186775 521346 186809 521380
rect 186867 521346 186901 521380
rect 186959 521346 186993 521380
rect 187051 521346 187085 521380
rect 187143 521346 187177 521380
rect 187235 521346 187269 521380
rect 187327 521346 187361 521380
rect 187419 521346 187453 521380
rect 172239 520802 172273 520836
rect 172331 520802 172365 520836
rect 172423 520802 172457 520836
rect 172515 520802 172549 520836
rect 172607 520802 172641 520836
rect 172699 520802 172733 520836
rect 172791 520802 172825 520836
rect 172883 520802 172917 520836
rect 172975 520802 173009 520836
rect 173067 520802 173101 520836
rect 173159 520802 173193 520836
rect 173251 520802 173285 520836
rect 173343 520802 173377 520836
rect 173435 520802 173469 520836
rect 173527 520802 173561 520836
rect 173619 520802 173653 520836
rect 173711 520802 173745 520836
rect 173803 520802 173837 520836
rect 173895 520802 173929 520836
rect 173987 520802 174021 520836
rect 174079 520802 174113 520836
rect 174171 520802 174205 520836
rect 174263 520802 174297 520836
rect 174355 520802 174389 520836
rect 174447 520802 174481 520836
rect 174539 520802 174573 520836
rect 174631 520802 174665 520836
rect 174723 520802 174757 520836
rect 174815 520802 174849 520836
rect 174907 520802 174941 520836
rect 174999 520802 175033 520836
rect 175091 520802 175125 520836
rect 175183 520802 175217 520836
rect 175275 520802 175309 520836
rect 175367 520802 175401 520836
rect 175459 520802 175493 520836
rect 175551 520802 175585 520836
rect 175643 520802 175677 520836
rect 175735 520802 175769 520836
rect 175827 520802 175861 520836
rect 175919 520802 175953 520836
rect 176011 520802 176045 520836
rect 176103 520802 176137 520836
rect 176195 520802 176229 520836
rect 176287 520802 176321 520836
rect 176379 520802 176413 520836
rect 176471 520802 176505 520836
rect 176563 520802 176597 520836
rect 176655 520802 176689 520836
rect 176747 520802 176781 520836
rect 176839 520802 176873 520836
rect 176931 520802 176965 520836
rect 177023 520802 177057 520836
rect 177115 520802 177149 520836
rect 177207 520802 177241 520836
rect 177299 520802 177333 520836
rect 177391 520802 177425 520836
rect 177483 520802 177517 520836
rect 177575 520802 177609 520836
rect 177667 520802 177701 520836
rect 177759 520802 177793 520836
rect 177851 520802 177885 520836
rect 177943 520802 177977 520836
rect 178035 520802 178069 520836
rect 178127 520802 178161 520836
rect 178219 520802 178253 520836
rect 178311 520802 178345 520836
rect 178403 520802 178437 520836
rect 178495 520802 178529 520836
rect 178587 520802 178621 520836
rect 178679 520802 178713 520836
rect 178771 520802 178805 520836
rect 178863 520802 178897 520836
rect 178955 520802 178989 520836
rect 179047 520802 179081 520836
rect 179139 520802 179173 520836
rect 179231 520802 179265 520836
rect 179323 520802 179357 520836
rect 179415 520802 179449 520836
rect 179507 520802 179541 520836
rect 179599 520802 179633 520836
rect 179691 520802 179725 520836
rect 179783 520802 179817 520836
rect 179875 520802 179909 520836
rect 179967 520802 180001 520836
rect 180059 520802 180093 520836
rect 180151 520802 180185 520836
rect 180243 520802 180277 520836
rect 180335 520802 180369 520836
rect 180427 520802 180461 520836
rect 180519 520802 180553 520836
rect 180611 520802 180645 520836
rect 180703 520802 180737 520836
rect 180795 520802 180829 520836
rect 180887 520802 180921 520836
rect 180979 520802 181013 520836
rect 181071 520802 181105 520836
rect 181163 520802 181197 520836
rect 181255 520802 181289 520836
rect 181347 520802 181381 520836
rect 181439 520802 181473 520836
rect 181531 520802 181565 520836
rect 181623 520802 181657 520836
rect 181715 520802 181749 520836
rect 181807 520802 181841 520836
rect 181899 520802 181933 520836
rect 181991 520802 182025 520836
rect 182083 520802 182117 520836
rect 182175 520802 182209 520836
rect 182267 520802 182301 520836
rect 182359 520802 182393 520836
rect 182451 520802 182485 520836
rect 182543 520802 182577 520836
rect 182635 520802 182669 520836
rect 182727 520802 182761 520836
rect 182819 520802 182853 520836
rect 182911 520802 182945 520836
rect 183003 520802 183037 520836
rect 183095 520802 183129 520836
rect 183187 520802 183221 520836
rect 183279 520802 183313 520836
rect 183371 520802 183405 520836
rect 183463 520802 183497 520836
rect 183555 520802 183589 520836
rect 183647 520802 183681 520836
rect 183739 520802 183773 520836
rect 183831 520802 183865 520836
rect 183923 520802 183957 520836
rect 184015 520802 184049 520836
rect 184107 520802 184141 520836
rect 184199 520802 184233 520836
rect 184291 520802 184325 520836
rect 184383 520802 184417 520836
rect 184475 520802 184509 520836
rect 184567 520802 184601 520836
rect 184659 520802 184693 520836
rect 184751 520802 184785 520836
rect 184843 520802 184877 520836
rect 184935 520802 184969 520836
rect 185027 520802 185061 520836
rect 185119 520802 185153 520836
rect 185211 520802 185245 520836
rect 185303 520802 185337 520836
rect 185395 520802 185429 520836
rect 185487 520802 185521 520836
rect 185579 520802 185613 520836
rect 185671 520802 185705 520836
rect 185763 520802 185797 520836
rect 185855 520802 185889 520836
rect 185947 520802 185981 520836
rect 186039 520802 186073 520836
rect 186131 520802 186165 520836
rect 186223 520802 186257 520836
rect 186315 520802 186349 520836
rect 186407 520802 186441 520836
rect 186499 520802 186533 520836
rect 186591 520802 186625 520836
rect 186683 520802 186717 520836
rect 186775 520802 186809 520836
rect 186867 520802 186901 520836
rect 186959 520802 186993 520836
rect 187051 520802 187085 520836
rect 187143 520802 187177 520836
rect 187235 520802 187269 520836
rect 187327 520802 187361 520836
rect 187419 520802 187453 520836
rect 172239 520258 172273 520292
rect 172331 520258 172365 520292
rect 172423 520258 172457 520292
rect 172515 520258 172549 520292
rect 172607 520258 172641 520292
rect 172699 520258 172733 520292
rect 172791 520258 172825 520292
rect 172883 520258 172917 520292
rect 172975 520258 173009 520292
rect 173067 520258 173101 520292
rect 173159 520258 173193 520292
rect 173251 520258 173285 520292
rect 173343 520258 173377 520292
rect 173435 520258 173469 520292
rect 173527 520258 173561 520292
rect 173619 520258 173653 520292
rect 173711 520258 173745 520292
rect 173803 520258 173837 520292
rect 173895 520258 173929 520292
rect 173987 520258 174021 520292
rect 174079 520258 174113 520292
rect 174171 520258 174205 520292
rect 174263 520258 174297 520292
rect 174355 520258 174389 520292
rect 174447 520258 174481 520292
rect 174539 520258 174573 520292
rect 174631 520258 174665 520292
rect 174723 520258 174757 520292
rect 174815 520258 174849 520292
rect 174907 520258 174941 520292
rect 174999 520258 175033 520292
rect 175091 520258 175125 520292
rect 175183 520258 175217 520292
rect 175275 520258 175309 520292
rect 175367 520258 175401 520292
rect 175459 520258 175493 520292
rect 175551 520258 175585 520292
rect 175643 520258 175677 520292
rect 175735 520258 175769 520292
rect 175827 520258 175861 520292
rect 175919 520258 175953 520292
rect 176011 520258 176045 520292
rect 176103 520258 176137 520292
rect 176195 520258 176229 520292
rect 176287 520258 176321 520292
rect 176379 520258 176413 520292
rect 176471 520258 176505 520292
rect 176563 520258 176597 520292
rect 176655 520258 176689 520292
rect 176747 520258 176781 520292
rect 176839 520258 176873 520292
rect 176931 520258 176965 520292
rect 177023 520258 177057 520292
rect 177115 520258 177149 520292
rect 177207 520258 177241 520292
rect 177299 520258 177333 520292
rect 177391 520258 177425 520292
rect 177483 520258 177517 520292
rect 177575 520258 177609 520292
rect 177667 520258 177701 520292
rect 177759 520258 177793 520292
rect 177851 520258 177885 520292
rect 177943 520258 177977 520292
rect 178035 520258 178069 520292
rect 178127 520258 178161 520292
rect 178219 520258 178253 520292
rect 178311 520258 178345 520292
rect 178403 520258 178437 520292
rect 178495 520258 178529 520292
rect 178587 520258 178621 520292
rect 178679 520258 178713 520292
rect 178771 520258 178805 520292
rect 178863 520258 178897 520292
rect 178955 520258 178989 520292
rect 179047 520258 179081 520292
rect 179139 520258 179173 520292
rect 179231 520258 179265 520292
rect 179323 520258 179357 520292
rect 179415 520258 179449 520292
rect 179507 520258 179541 520292
rect 179599 520258 179633 520292
rect 179691 520258 179725 520292
rect 179783 520258 179817 520292
rect 179875 520258 179909 520292
rect 179967 520258 180001 520292
rect 180059 520258 180093 520292
rect 180151 520258 180185 520292
rect 180243 520258 180277 520292
rect 180335 520258 180369 520292
rect 180427 520258 180461 520292
rect 180519 520258 180553 520292
rect 180611 520258 180645 520292
rect 180703 520258 180737 520292
rect 180795 520258 180829 520292
rect 180887 520258 180921 520292
rect 180979 520258 181013 520292
rect 181071 520258 181105 520292
rect 181163 520258 181197 520292
rect 181255 520258 181289 520292
rect 181347 520258 181381 520292
rect 181439 520258 181473 520292
rect 181531 520258 181565 520292
rect 181623 520258 181657 520292
rect 181715 520258 181749 520292
rect 181807 520258 181841 520292
rect 181899 520258 181933 520292
rect 181991 520258 182025 520292
rect 182083 520258 182117 520292
rect 182175 520258 182209 520292
rect 182267 520258 182301 520292
rect 182359 520258 182393 520292
rect 182451 520258 182485 520292
rect 182543 520258 182577 520292
rect 182635 520258 182669 520292
rect 182727 520258 182761 520292
rect 182819 520258 182853 520292
rect 182911 520258 182945 520292
rect 183003 520258 183037 520292
rect 183095 520258 183129 520292
rect 183187 520258 183221 520292
rect 183279 520258 183313 520292
rect 183371 520258 183405 520292
rect 183463 520258 183497 520292
rect 183555 520258 183589 520292
rect 183647 520258 183681 520292
rect 183739 520258 183773 520292
rect 183831 520258 183865 520292
rect 183923 520258 183957 520292
rect 184015 520258 184049 520292
rect 184107 520258 184141 520292
rect 184199 520258 184233 520292
rect 184291 520258 184325 520292
rect 184383 520258 184417 520292
rect 184475 520258 184509 520292
rect 184567 520258 184601 520292
rect 184659 520258 184693 520292
rect 184751 520258 184785 520292
rect 184843 520258 184877 520292
rect 184935 520258 184969 520292
rect 185027 520258 185061 520292
rect 185119 520258 185153 520292
rect 185211 520258 185245 520292
rect 185303 520258 185337 520292
rect 185395 520258 185429 520292
rect 185487 520258 185521 520292
rect 185579 520258 185613 520292
rect 185671 520258 185705 520292
rect 185763 520258 185797 520292
rect 185855 520258 185889 520292
rect 185947 520258 185981 520292
rect 186039 520258 186073 520292
rect 186131 520258 186165 520292
rect 186223 520258 186257 520292
rect 186315 520258 186349 520292
rect 186407 520258 186441 520292
rect 186499 520258 186533 520292
rect 186591 520258 186625 520292
rect 186683 520258 186717 520292
rect 186775 520258 186809 520292
rect 186867 520258 186901 520292
rect 186959 520258 186993 520292
rect 187051 520258 187085 520292
rect 187143 520258 187177 520292
rect 187235 520258 187269 520292
rect 187327 520258 187361 520292
rect 187419 520258 187453 520292
rect 172239 519714 172273 519748
rect 172331 519714 172365 519748
rect 172423 519714 172457 519748
rect 172515 519714 172549 519748
rect 172607 519714 172641 519748
rect 172699 519714 172733 519748
rect 172791 519714 172825 519748
rect 172883 519714 172917 519748
rect 172975 519714 173009 519748
rect 173067 519714 173101 519748
rect 173159 519714 173193 519748
rect 173251 519714 173285 519748
rect 173343 519714 173377 519748
rect 173435 519714 173469 519748
rect 173527 519714 173561 519748
rect 173619 519714 173653 519748
rect 173711 519714 173745 519748
rect 173803 519714 173837 519748
rect 173895 519714 173929 519748
rect 173987 519714 174021 519748
rect 174079 519714 174113 519748
rect 174171 519714 174205 519748
rect 174263 519714 174297 519748
rect 174355 519714 174389 519748
rect 174447 519714 174481 519748
rect 174539 519714 174573 519748
rect 174631 519714 174665 519748
rect 174723 519714 174757 519748
rect 174815 519714 174849 519748
rect 174907 519714 174941 519748
rect 174999 519714 175033 519748
rect 175091 519714 175125 519748
rect 175183 519714 175217 519748
rect 175275 519714 175309 519748
rect 175367 519714 175401 519748
rect 175459 519714 175493 519748
rect 175551 519714 175585 519748
rect 175643 519714 175677 519748
rect 175735 519714 175769 519748
rect 175827 519714 175861 519748
rect 175919 519714 175953 519748
rect 176011 519714 176045 519748
rect 176103 519714 176137 519748
rect 176195 519714 176229 519748
rect 176287 519714 176321 519748
rect 176379 519714 176413 519748
rect 176471 519714 176505 519748
rect 176563 519714 176597 519748
rect 176655 519714 176689 519748
rect 176747 519714 176781 519748
rect 176839 519714 176873 519748
rect 176931 519714 176965 519748
rect 177023 519714 177057 519748
rect 177115 519714 177149 519748
rect 177207 519714 177241 519748
rect 177299 519714 177333 519748
rect 177391 519714 177425 519748
rect 177483 519714 177517 519748
rect 177575 519714 177609 519748
rect 177667 519714 177701 519748
rect 177759 519714 177793 519748
rect 177851 519714 177885 519748
rect 177943 519714 177977 519748
rect 178035 519714 178069 519748
rect 178127 519714 178161 519748
rect 178219 519714 178253 519748
rect 178311 519714 178345 519748
rect 178403 519714 178437 519748
rect 178495 519714 178529 519748
rect 178587 519714 178621 519748
rect 178679 519714 178713 519748
rect 178771 519714 178805 519748
rect 178863 519714 178897 519748
rect 178955 519714 178989 519748
rect 179047 519714 179081 519748
rect 179139 519714 179173 519748
rect 179231 519714 179265 519748
rect 179323 519714 179357 519748
rect 179415 519714 179449 519748
rect 179507 519714 179541 519748
rect 179599 519714 179633 519748
rect 179691 519714 179725 519748
rect 179783 519714 179817 519748
rect 179875 519714 179909 519748
rect 179967 519714 180001 519748
rect 180059 519714 180093 519748
rect 180151 519714 180185 519748
rect 180243 519714 180277 519748
rect 180335 519714 180369 519748
rect 180427 519714 180461 519748
rect 180519 519714 180553 519748
rect 180611 519714 180645 519748
rect 180703 519714 180737 519748
rect 180795 519714 180829 519748
rect 180887 519714 180921 519748
rect 180979 519714 181013 519748
rect 181071 519714 181105 519748
rect 181163 519714 181197 519748
rect 181255 519714 181289 519748
rect 181347 519714 181381 519748
rect 181439 519714 181473 519748
rect 181531 519714 181565 519748
rect 181623 519714 181657 519748
rect 181715 519714 181749 519748
rect 181807 519714 181841 519748
rect 181899 519714 181933 519748
rect 181991 519714 182025 519748
rect 182083 519714 182117 519748
rect 182175 519714 182209 519748
rect 182267 519714 182301 519748
rect 182359 519714 182393 519748
rect 182451 519714 182485 519748
rect 182543 519714 182577 519748
rect 182635 519714 182669 519748
rect 182727 519714 182761 519748
rect 182819 519714 182853 519748
rect 182911 519714 182945 519748
rect 183003 519714 183037 519748
rect 183095 519714 183129 519748
rect 183187 519714 183221 519748
rect 183279 519714 183313 519748
rect 183371 519714 183405 519748
rect 183463 519714 183497 519748
rect 183555 519714 183589 519748
rect 183647 519714 183681 519748
rect 183739 519714 183773 519748
rect 183831 519714 183865 519748
rect 183923 519714 183957 519748
rect 184015 519714 184049 519748
rect 184107 519714 184141 519748
rect 184199 519714 184233 519748
rect 184291 519714 184325 519748
rect 184383 519714 184417 519748
rect 184475 519714 184509 519748
rect 184567 519714 184601 519748
rect 184659 519714 184693 519748
rect 184751 519714 184785 519748
rect 184843 519714 184877 519748
rect 184935 519714 184969 519748
rect 185027 519714 185061 519748
rect 185119 519714 185153 519748
rect 185211 519714 185245 519748
rect 185303 519714 185337 519748
rect 185395 519714 185429 519748
rect 185487 519714 185521 519748
rect 185579 519714 185613 519748
rect 185671 519714 185705 519748
rect 185763 519714 185797 519748
rect 185855 519714 185889 519748
rect 185947 519714 185981 519748
rect 186039 519714 186073 519748
rect 186131 519714 186165 519748
rect 186223 519714 186257 519748
rect 186315 519714 186349 519748
rect 186407 519714 186441 519748
rect 186499 519714 186533 519748
rect 186591 519714 186625 519748
rect 186683 519714 186717 519748
rect 186775 519714 186809 519748
rect 186867 519714 186901 519748
rect 186959 519714 186993 519748
rect 187051 519714 187085 519748
rect 187143 519714 187177 519748
rect 187235 519714 187269 519748
rect 187327 519714 187361 519748
rect 187419 519714 187453 519748
rect 172239 519170 172273 519204
rect 172331 519170 172365 519204
rect 172423 519170 172457 519204
rect 172515 519170 172549 519204
rect 172607 519170 172641 519204
rect 172699 519170 172733 519204
rect 172791 519170 172825 519204
rect 172883 519170 172917 519204
rect 172975 519170 173009 519204
rect 173067 519170 173101 519204
rect 173159 519170 173193 519204
rect 173251 519170 173285 519204
rect 173343 519170 173377 519204
rect 173435 519170 173469 519204
rect 173527 519170 173561 519204
rect 173619 519170 173653 519204
rect 173711 519170 173745 519204
rect 173803 519170 173837 519204
rect 173895 519170 173929 519204
rect 173987 519170 174021 519204
rect 174079 519170 174113 519204
rect 174171 519170 174205 519204
rect 174263 519170 174297 519204
rect 174355 519170 174389 519204
rect 174447 519170 174481 519204
rect 174539 519170 174573 519204
rect 174631 519170 174665 519204
rect 174723 519170 174757 519204
rect 174815 519170 174849 519204
rect 174907 519170 174941 519204
rect 174999 519170 175033 519204
rect 175091 519170 175125 519204
rect 175183 519170 175217 519204
rect 175275 519170 175309 519204
rect 175367 519170 175401 519204
rect 175459 519170 175493 519204
rect 175551 519170 175585 519204
rect 175643 519170 175677 519204
rect 175735 519170 175769 519204
rect 175827 519170 175861 519204
rect 175919 519170 175953 519204
rect 176011 519170 176045 519204
rect 176103 519170 176137 519204
rect 176195 519170 176229 519204
rect 176287 519170 176321 519204
rect 176379 519170 176413 519204
rect 176471 519170 176505 519204
rect 176563 519170 176597 519204
rect 176655 519170 176689 519204
rect 176747 519170 176781 519204
rect 176839 519170 176873 519204
rect 176931 519170 176965 519204
rect 177023 519170 177057 519204
rect 177115 519170 177149 519204
rect 177207 519170 177241 519204
rect 177299 519170 177333 519204
rect 177391 519170 177425 519204
rect 177483 519170 177517 519204
rect 177575 519170 177609 519204
rect 177667 519170 177701 519204
rect 177759 519170 177793 519204
rect 177851 519170 177885 519204
rect 177943 519170 177977 519204
rect 178035 519170 178069 519204
rect 178127 519170 178161 519204
rect 178219 519170 178253 519204
rect 178311 519170 178345 519204
rect 178403 519170 178437 519204
rect 178495 519170 178529 519204
rect 178587 519170 178621 519204
rect 178679 519170 178713 519204
rect 178771 519170 178805 519204
rect 178863 519170 178897 519204
rect 178955 519170 178989 519204
rect 179047 519170 179081 519204
rect 179139 519170 179173 519204
rect 179231 519170 179265 519204
rect 179323 519170 179357 519204
rect 179415 519170 179449 519204
rect 179507 519170 179541 519204
rect 179599 519170 179633 519204
rect 179691 519170 179725 519204
rect 179783 519170 179817 519204
rect 179875 519170 179909 519204
rect 179967 519170 180001 519204
rect 180059 519170 180093 519204
rect 180151 519170 180185 519204
rect 180243 519170 180277 519204
rect 180335 519170 180369 519204
rect 180427 519170 180461 519204
rect 180519 519170 180553 519204
rect 180611 519170 180645 519204
rect 180703 519170 180737 519204
rect 180795 519170 180829 519204
rect 180887 519170 180921 519204
rect 180979 519170 181013 519204
rect 181071 519170 181105 519204
rect 181163 519170 181197 519204
rect 181255 519170 181289 519204
rect 181347 519170 181381 519204
rect 181439 519170 181473 519204
rect 181531 519170 181565 519204
rect 181623 519170 181657 519204
rect 181715 519170 181749 519204
rect 181807 519170 181841 519204
rect 181899 519170 181933 519204
rect 181991 519170 182025 519204
rect 182083 519170 182117 519204
rect 182175 519170 182209 519204
rect 182267 519170 182301 519204
rect 182359 519170 182393 519204
rect 182451 519170 182485 519204
rect 182543 519170 182577 519204
rect 182635 519170 182669 519204
rect 182727 519170 182761 519204
rect 182819 519170 182853 519204
rect 182911 519170 182945 519204
rect 183003 519170 183037 519204
rect 183095 519170 183129 519204
rect 183187 519170 183221 519204
rect 183279 519170 183313 519204
rect 183371 519170 183405 519204
rect 183463 519170 183497 519204
rect 183555 519170 183589 519204
rect 183647 519170 183681 519204
rect 183739 519170 183773 519204
rect 183831 519170 183865 519204
rect 183923 519170 183957 519204
rect 184015 519170 184049 519204
rect 184107 519170 184141 519204
rect 184199 519170 184233 519204
rect 184291 519170 184325 519204
rect 184383 519170 184417 519204
rect 184475 519170 184509 519204
rect 184567 519170 184601 519204
rect 184659 519170 184693 519204
rect 184751 519170 184785 519204
rect 184843 519170 184877 519204
rect 184935 519170 184969 519204
rect 185027 519170 185061 519204
rect 185119 519170 185153 519204
rect 185211 519170 185245 519204
rect 185303 519170 185337 519204
rect 185395 519170 185429 519204
rect 185487 519170 185521 519204
rect 185579 519170 185613 519204
rect 185671 519170 185705 519204
rect 185763 519170 185797 519204
rect 185855 519170 185889 519204
rect 185947 519170 185981 519204
rect 186039 519170 186073 519204
rect 186131 519170 186165 519204
rect 186223 519170 186257 519204
rect 186315 519170 186349 519204
rect 186407 519170 186441 519204
rect 186499 519170 186533 519204
rect 186591 519170 186625 519204
rect 186683 519170 186717 519204
rect 186775 519170 186809 519204
rect 186867 519170 186901 519204
rect 186959 519170 186993 519204
rect 187051 519170 187085 519204
rect 187143 519170 187177 519204
rect 187235 519170 187269 519204
rect 187327 519170 187361 519204
rect 187419 519170 187453 519204
rect 172239 518626 172273 518660
rect 172331 518626 172365 518660
rect 172423 518626 172457 518660
rect 172515 518626 172549 518660
rect 172607 518626 172641 518660
rect 172699 518626 172733 518660
rect 172791 518626 172825 518660
rect 172883 518626 172917 518660
rect 172975 518626 173009 518660
rect 173067 518626 173101 518660
rect 173159 518626 173193 518660
rect 173251 518626 173285 518660
rect 173343 518626 173377 518660
rect 173435 518626 173469 518660
rect 173527 518626 173561 518660
rect 173619 518626 173653 518660
rect 173711 518626 173745 518660
rect 173803 518626 173837 518660
rect 173895 518626 173929 518660
rect 173987 518626 174021 518660
rect 174079 518626 174113 518660
rect 174171 518626 174205 518660
rect 174263 518626 174297 518660
rect 174355 518626 174389 518660
rect 174447 518626 174481 518660
rect 174539 518626 174573 518660
rect 174631 518626 174665 518660
rect 174723 518626 174757 518660
rect 174815 518626 174849 518660
rect 174907 518626 174941 518660
rect 174999 518626 175033 518660
rect 175091 518626 175125 518660
rect 175183 518626 175217 518660
rect 175275 518626 175309 518660
rect 175367 518626 175401 518660
rect 175459 518626 175493 518660
rect 175551 518626 175585 518660
rect 175643 518626 175677 518660
rect 175735 518626 175769 518660
rect 175827 518626 175861 518660
rect 175919 518626 175953 518660
rect 176011 518626 176045 518660
rect 176103 518626 176137 518660
rect 176195 518626 176229 518660
rect 176287 518626 176321 518660
rect 176379 518626 176413 518660
rect 176471 518626 176505 518660
rect 176563 518626 176597 518660
rect 176655 518626 176689 518660
rect 176747 518626 176781 518660
rect 176839 518626 176873 518660
rect 176931 518626 176965 518660
rect 177023 518626 177057 518660
rect 177115 518626 177149 518660
rect 177207 518626 177241 518660
rect 177299 518626 177333 518660
rect 177391 518626 177425 518660
rect 177483 518626 177517 518660
rect 177575 518626 177609 518660
rect 177667 518626 177701 518660
rect 177759 518626 177793 518660
rect 177851 518626 177885 518660
rect 177943 518626 177977 518660
rect 178035 518626 178069 518660
rect 178127 518626 178161 518660
rect 178219 518626 178253 518660
rect 178311 518626 178345 518660
rect 178403 518626 178437 518660
rect 178495 518626 178529 518660
rect 178587 518626 178621 518660
rect 178679 518626 178713 518660
rect 178771 518626 178805 518660
rect 178863 518626 178897 518660
rect 178955 518626 178989 518660
rect 179047 518626 179081 518660
rect 179139 518626 179173 518660
rect 179231 518626 179265 518660
rect 179323 518626 179357 518660
rect 179415 518626 179449 518660
rect 179507 518626 179541 518660
rect 179599 518626 179633 518660
rect 179691 518626 179725 518660
rect 179783 518626 179817 518660
rect 179875 518626 179909 518660
rect 179967 518626 180001 518660
rect 180059 518626 180093 518660
rect 180151 518626 180185 518660
rect 180243 518626 180277 518660
rect 180335 518626 180369 518660
rect 180427 518626 180461 518660
rect 180519 518626 180553 518660
rect 180611 518626 180645 518660
rect 180703 518626 180737 518660
rect 180795 518626 180829 518660
rect 180887 518626 180921 518660
rect 180979 518626 181013 518660
rect 181071 518626 181105 518660
rect 181163 518626 181197 518660
rect 181255 518626 181289 518660
rect 181347 518626 181381 518660
rect 181439 518626 181473 518660
rect 181531 518626 181565 518660
rect 181623 518626 181657 518660
rect 181715 518626 181749 518660
rect 181807 518626 181841 518660
rect 181899 518626 181933 518660
rect 181991 518626 182025 518660
rect 182083 518626 182117 518660
rect 182175 518626 182209 518660
rect 182267 518626 182301 518660
rect 182359 518626 182393 518660
rect 182451 518626 182485 518660
rect 182543 518626 182577 518660
rect 182635 518626 182669 518660
rect 182727 518626 182761 518660
rect 182819 518626 182853 518660
rect 182911 518626 182945 518660
rect 183003 518626 183037 518660
rect 183095 518626 183129 518660
rect 183187 518626 183221 518660
rect 183279 518626 183313 518660
rect 183371 518626 183405 518660
rect 183463 518626 183497 518660
rect 183555 518626 183589 518660
rect 183647 518626 183681 518660
rect 183739 518626 183773 518660
rect 183831 518626 183865 518660
rect 183923 518626 183957 518660
rect 184015 518626 184049 518660
rect 184107 518626 184141 518660
rect 184199 518626 184233 518660
rect 184291 518626 184325 518660
rect 184383 518626 184417 518660
rect 184475 518626 184509 518660
rect 184567 518626 184601 518660
rect 184659 518626 184693 518660
rect 184751 518626 184785 518660
rect 184843 518626 184877 518660
rect 184935 518626 184969 518660
rect 185027 518626 185061 518660
rect 185119 518626 185153 518660
rect 185211 518626 185245 518660
rect 185303 518626 185337 518660
rect 185395 518626 185429 518660
rect 185487 518626 185521 518660
rect 185579 518626 185613 518660
rect 185671 518626 185705 518660
rect 185763 518626 185797 518660
rect 185855 518626 185889 518660
rect 185947 518626 185981 518660
rect 186039 518626 186073 518660
rect 186131 518626 186165 518660
rect 186223 518626 186257 518660
rect 186315 518626 186349 518660
rect 186407 518626 186441 518660
rect 186499 518626 186533 518660
rect 186591 518626 186625 518660
rect 186683 518626 186717 518660
rect 186775 518626 186809 518660
rect 186867 518626 186901 518660
rect 186959 518626 186993 518660
rect 187051 518626 187085 518660
rect 187143 518626 187177 518660
rect 187235 518626 187269 518660
rect 187327 518626 187361 518660
rect 187419 518626 187453 518660
rect 172239 518082 172273 518116
rect 172331 518082 172365 518116
rect 172423 518082 172457 518116
rect 172515 518082 172549 518116
rect 172607 518082 172641 518116
rect 172699 518082 172733 518116
rect 172791 518082 172825 518116
rect 172883 518082 172917 518116
rect 172975 518082 173009 518116
rect 173067 518082 173101 518116
rect 173159 518082 173193 518116
rect 173251 518082 173285 518116
rect 173343 518082 173377 518116
rect 173435 518082 173469 518116
rect 173527 518082 173561 518116
rect 173619 518082 173653 518116
rect 173711 518082 173745 518116
rect 173803 518082 173837 518116
rect 173895 518082 173929 518116
rect 173987 518082 174021 518116
rect 174079 518082 174113 518116
rect 174171 518082 174205 518116
rect 174263 518082 174297 518116
rect 174355 518082 174389 518116
rect 174447 518082 174481 518116
rect 174539 518082 174573 518116
rect 174631 518082 174665 518116
rect 174723 518082 174757 518116
rect 174815 518082 174849 518116
rect 174907 518082 174941 518116
rect 174999 518082 175033 518116
rect 175091 518082 175125 518116
rect 175183 518082 175217 518116
rect 175275 518082 175309 518116
rect 175367 518082 175401 518116
rect 175459 518082 175493 518116
rect 175551 518082 175585 518116
rect 175643 518082 175677 518116
rect 175735 518082 175769 518116
rect 175827 518082 175861 518116
rect 175919 518082 175953 518116
rect 176011 518082 176045 518116
rect 176103 518082 176137 518116
rect 176195 518082 176229 518116
rect 176287 518082 176321 518116
rect 176379 518082 176413 518116
rect 176471 518082 176505 518116
rect 176563 518082 176597 518116
rect 176655 518082 176689 518116
rect 176747 518082 176781 518116
rect 176839 518082 176873 518116
rect 176931 518082 176965 518116
rect 177023 518082 177057 518116
rect 177115 518082 177149 518116
rect 177207 518082 177241 518116
rect 177299 518082 177333 518116
rect 177391 518082 177425 518116
rect 177483 518082 177517 518116
rect 177575 518082 177609 518116
rect 177667 518082 177701 518116
rect 177759 518082 177793 518116
rect 177851 518082 177885 518116
rect 177943 518082 177977 518116
rect 178035 518082 178069 518116
rect 178127 518082 178161 518116
rect 178219 518082 178253 518116
rect 178311 518082 178345 518116
rect 178403 518082 178437 518116
rect 178495 518082 178529 518116
rect 178587 518082 178621 518116
rect 178679 518082 178713 518116
rect 178771 518082 178805 518116
rect 178863 518082 178897 518116
rect 178955 518082 178989 518116
rect 179047 518082 179081 518116
rect 179139 518082 179173 518116
rect 179231 518082 179265 518116
rect 179323 518082 179357 518116
rect 179415 518082 179449 518116
rect 179507 518082 179541 518116
rect 179599 518082 179633 518116
rect 179691 518082 179725 518116
rect 179783 518082 179817 518116
rect 179875 518082 179909 518116
rect 179967 518082 180001 518116
rect 180059 518082 180093 518116
rect 180151 518082 180185 518116
rect 180243 518082 180277 518116
rect 180335 518082 180369 518116
rect 180427 518082 180461 518116
rect 180519 518082 180553 518116
rect 180611 518082 180645 518116
rect 180703 518082 180737 518116
rect 180795 518082 180829 518116
rect 180887 518082 180921 518116
rect 180979 518082 181013 518116
rect 181071 518082 181105 518116
rect 181163 518082 181197 518116
rect 181255 518082 181289 518116
rect 181347 518082 181381 518116
rect 181439 518082 181473 518116
rect 181531 518082 181565 518116
rect 181623 518082 181657 518116
rect 181715 518082 181749 518116
rect 181807 518082 181841 518116
rect 181899 518082 181933 518116
rect 181991 518082 182025 518116
rect 182083 518082 182117 518116
rect 182175 518082 182209 518116
rect 182267 518082 182301 518116
rect 182359 518082 182393 518116
rect 182451 518082 182485 518116
rect 182543 518082 182577 518116
rect 182635 518082 182669 518116
rect 182727 518082 182761 518116
rect 182819 518082 182853 518116
rect 182911 518082 182945 518116
rect 183003 518082 183037 518116
rect 183095 518082 183129 518116
rect 183187 518082 183221 518116
rect 183279 518082 183313 518116
rect 183371 518082 183405 518116
rect 183463 518082 183497 518116
rect 183555 518082 183589 518116
rect 183647 518082 183681 518116
rect 183739 518082 183773 518116
rect 183831 518082 183865 518116
rect 183923 518082 183957 518116
rect 184015 518082 184049 518116
rect 184107 518082 184141 518116
rect 184199 518082 184233 518116
rect 184291 518082 184325 518116
rect 184383 518082 184417 518116
rect 184475 518082 184509 518116
rect 184567 518082 184601 518116
rect 184659 518082 184693 518116
rect 184751 518082 184785 518116
rect 184843 518082 184877 518116
rect 184935 518082 184969 518116
rect 185027 518082 185061 518116
rect 185119 518082 185153 518116
rect 185211 518082 185245 518116
rect 185303 518082 185337 518116
rect 185395 518082 185429 518116
rect 185487 518082 185521 518116
rect 185579 518082 185613 518116
rect 185671 518082 185705 518116
rect 185763 518082 185797 518116
rect 185855 518082 185889 518116
rect 185947 518082 185981 518116
rect 186039 518082 186073 518116
rect 186131 518082 186165 518116
rect 186223 518082 186257 518116
rect 186315 518082 186349 518116
rect 186407 518082 186441 518116
rect 186499 518082 186533 518116
rect 186591 518082 186625 518116
rect 186683 518082 186717 518116
rect 186775 518082 186809 518116
rect 186867 518082 186901 518116
rect 186959 518082 186993 518116
rect 187051 518082 187085 518116
rect 187143 518082 187177 518116
rect 187235 518082 187269 518116
rect 187327 518082 187361 518116
rect 187419 518082 187453 518116
rect 172239 517538 172273 517572
rect 172331 517538 172365 517572
rect 172423 517538 172457 517572
rect 172515 517538 172549 517572
rect 172607 517538 172641 517572
rect 172699 517538 172733 517572
rect 172791 517538 172825 517572
rect 172883 517538 172917 517572
rect 172975 517538 173009 517572
rect 173067 517538 173101 517572
rect 173159 517538 173193 517572
rect 173251 517538 173285 517572
rect 173343 517538 173377 517572
rect 173435 517538 173469 517572
rect 173527 517538 173561 517572
rect 173619 517538 173653 517572
rect 173711 517538 173745 517572
rect 173803 517538 173837 517572
rect 173895 517538 173929 517572
rect 173987 517538 174021 517572
rect 174079 517538 174113 517572
rect 174171 517538 174205 517572
rect 174263 517538 174297 517572
rect 174355 517538 174389 517572
rect 174447 517538 174481 517572
rect 174539 517538 174573 517572
rect 174631 517538 174665 517572
rect 174723 517538 174757 517572
rect 174815 517538 174849 517572
rect 174907 517538 174941 517572
rect 174999 517538 175033 517572
rect 175091 517538 175125 517572
rect 175183 517538 175217 517572
rect 175275 517538 175309 517572
rect 175367 517538 175401 517572
rect 175459 517538 175493 517572
rect 175551 517538 175585 517572
rect 175643 517538 175677 517572
rect 175735 517538 175769 517572
rect 175827 517538 175861 517572
rect 175919 517538 175953 517572
rect 176011 517538 176045 517572
rect 176103 517538 176137 517572
rect 176195 517538 176229 517572
rect 176287 517538 176321 517572
rect 176379 517538 176413 517572
rect 176471 517538 176505 517572
rect 176563 517538 176597 517572
rect 176655 517538 176689 517572
rect 176747 517538 176781 517572
rect 176839 517538 176873 517572
rect 176931 517538 176965 517572
rect 177023 517538 177057 517572
rect 177115 517538 177149 517572
rect 177207 517538 177241 517572
rect 177299 517538 177333 517572
rect 177391 517538 177425 517572
rect 177483 517538 177517 517572
rect 177575 517538 177609 517572
rect 177667 517538 177701 517572
rect 177759 517538 177793 517572
rect 177851 517538 177885 517572
rect 177943 517538 177977 517572
rect 178035 517538 178069 517572
rect 178127 517538 178161 517572
rect 178219 517538 178253 517572
rect 178311 517538 178345 517572
rect 178403 517538 178437 517572
rect 178495 517538 178529 517572
rect 178587 517538 178621 517572
rect 178679 517538 178713 517572
rect 178771 517538 178805 517572
rect 178863 517538 178897 517572
rect 178955 517538 178989 517572
rect 179047 517538 179081 517572
rect 179139 517538 179173 517572
rect 179231 517538 179265 517572
rect 179323 517538 179357 517572
rect 179415 517538 179449 517572
rect 179507 517538 179541 517572
rect 179599 517538 179633 517572
rect 179691 517538 179725 517572
rect 179783 517538 179817 517572
rect 179875 517538 179909 517572
rect 179967 517538 180001 517572
rect 180059 517538 180093 517572
rect 180151 517538 180185 517572
rect 180243 517538 180277 517572
rect 180335 517538 180369 517572
rect 180427 517538 180461 517572
rect 180519 517538 180553 517572
rect 180611 517538 180645 517572
rect 180703 517538 180737 517572
rect 180795 517538 180829 517572
rect 180887 517538 180921 517572
rect 180979 517538 181013 517572
rect 181071 517538 181105 517572
rect 181163 517538 181197 517572
rect 181255 517538 181289 517572
rect 181347 517538 181381 517572
rect 181439 517538 181473 517572
rect 181531 517538 181565 517572
rect 181623 517538 181657 517572
rect 181715 517538 181749 517572
rect 181807 517538 181841 517572
rect 181899 517538 181933 517572
rect 181991 517538 182025 517572
rect 182083 517538 182117 517572
rect 182175 517538 182209 517572
rect 182267 517538 182301 517572
rect 182359 517538 182393 517572
rect 182451 517538 182485 517572
rect 182543 517538 182577 517572
rect 182635 517538 182669 517572
rect 182727 517538 182761 517572
rect 182819 517538 182853 517572
rect 182911 517538 182945 517572
rect 183003 517538 183037 517572
rect 183095 517538 183129 517572
rect 183187 517538 183221 517572
rect 183279 517538 183313 517572
rect 183371 517538 183405 517572
rect 183463 517538 183497 517572
rect 183555 517538 183589 517572
rect 183647 517538 183681 517572
rect 183739 517538 183773 517572
rect 183831 517538 183865 517572
rect 183923 517538 183957 517572
rect 184015 517538 184049 517572
rect 184107 517538 184141 517572
rect 184199 517538 184233 517572
rect 184291 517538 184325 517572
rect 184383 517538 184417 517572
rect 184475 517538 184509 517572
rect 184567 517538 184601 517572
rect 184659 517538 184693 517572
rect 184751 517538 184785 517572
rect 184843 517538 184877 517572
rect 184935 517538 184969 517572
rect 185027 517538 185061 517572
rect 185119 517538 185153 517572
rect 185211 517538 185245 517572
rect 185303 517538 185337 517572
rect 185395 517538 185429 517572
rect 185487 517538 185521 517572
rect 185579 517538 185613 517572
rect 185671 517538 185705 517572
rect 185763 517538 185797 517572
rect 185855 517538 185889 517572
rect 185947 517538 185981 517572
rect 186039 517538 186073 517572
rect 186131 517538 186165 517572
rect 186223 517538 186257 517572
rect 186315 517538 186349 517572
rect 186407 517538 186441 517572
rect 186499 517538 186533 517572
rect 186591 517538 186625 517572
rect 186683 517538 186717 517572
rect 186775 517538 186809 517572
rect 186867 517538 186901 517572
rect 186959 517538 186993 517572
rect 187051 517538 187085 517572
rect 187143 517538 187177 517572
rect 187235 517538 187269 517572
rect 187327 517538 187361 517572
rect 187419 517538 187453 517572
rect 172239 516994 172273 517028
rect 172331 516994 172365 517028
rect 172423 516994 172457 517028
rect 172515 516994 172549 517028
rect 172607 516994 172641 517028
rect 172699 516994 172733 517028
rect 172791 516994 172825 517028
rect 172883 516994 172917 517028
rect 172975 516994 173009 517028
rect 173067 516994 173101 517028
rect 173159 516994 173193 517028
rect 173251 516994 173285 517028
rect 173343 516994 173377 517028
rect 173435 516994 173469 517028
rect 173527 516994 173561 517028
rect 173619 516994 173653 517028
rect 173711 516994 173745 517028
rect 173803 516994 173837 517028
rect 173895 516994 173929 517028
rect 173987 516994 174021 517028
rect 174079 516994 174113 517028
rect 174171 516994 174205 517028
rect 174263 516994 174297 517028
rect 174355 516994 174389 517028
rect 174447 516994 174481 517028
rect 174539 516994 174573 517028
rect 174631 516994 174665 517028
rect 174723 516994 174757 517028
rect 174815 516994 174849 517028
rect 174907 516994 174941 517028
rect 174999 516994 175033 517028
rect 175091 516994 175125 517028
rect 175183 516994 175217 517028
rect 175275 516994 175309 517028
rect 175367 516994 175401 517028
rect 175459 516994 175493 517028
rect 175551 516994 175585 517028
rect 175643 516994 175677 517028
rect 175735 516994 175769 517028
rect 175827 516994 175861 517028
rect 175919 516994 175953 517028
rect 176011 516994 176045 517028
rect 176103 516994 176137 517028
rect 176195 516994 176229 517028
rect 176287 516994 176321 517028
rect 176379 516994 176413 517028
rect 176471 516994 176505 517028
rect 176563 516994 176597 517028
rect 176655 516994 176689 517028
rect 176747 516994 176781 517028
rect 176839 516994 176873 517028
rect 176931 516994 176965 517028
rect 177023 516994 177057 517028
rect 177115 516994 177149 517028
rect 177207 516994 177241 517028
rect 177299 516994 177333 517028
rect 177391 516994 177425 517028
rect 177483 516994 177517 517028
rect 177575 516994 177609 517028
rect 177667 516994 177701 517028
rect 177759 516994 177793 517028
rect 177851 516994 177885 517028
rect 177943 516994 177977 517028
rect 178035 516994 178069 517028
rect 178127 516994 178161 517028
rect 178219 516994 178253 517028
rect 178311 516994 178345 517028
rect 178403 516994 178437 517028
rect 178495 516994 178529 517028
rect 178587 516994 178621 517028
rect 178679 516994 178713 517028
rect 178771 516994 178805 517028
rect 178863 516994 178897 517028
rect 178955 516994 178989 517028
rect 179047 516994 179081 517028
rect 179139 516994 179173 517028
rect 179231 516994 179265 517028
rect 179323 516994 179357 517028
rect 179415 516994 179449 517028
rect 179507 516994 179541 517028
rect 179599 516994 179633 517028
rect 179691 516994 179725 517028
rect 179783 516994 179817 517028
rect 179875 516994 179909 517028
rect 179967 516994 180001 517028
rect 180059 516994 180093 517028
rect 180151 516994 180185 517028
rect 180243 516994 180277 517028
rect 180335 516994 180369 517028
rect 180427 516994 180461 517028
rect 180519 516994 180553 517028
rect 180611 516994 180645 517028
rect 180703 516994 180737 517028
rect 180795 516994 180829 517028
rect 180887 516994 180921 517028
rect 180979 516994 181013 517028
rect 181071 516994 181105 517028
rect 181163 516994 181197 517028
rect 181255 516994 181289 517028
rect 181347 516994 181381 517028
rect 181439 516994 181473 517028
rect 181531 516994 181565 517028
rect 181623 516994 181657 517028
rect 181715 516994 181749 517028
rect 181807 516994 181841 517028
rect 181899 516994 181933 517028
rect 181991 516994 182025 517028
rect 182083 516994 182117 517028
rect 182175 516994 182209 517028
rect 182267 516994 182301 517028
rect 182359 516994 182393 517028
rect 182451 516994 182485 517028
rect 182543 516994 182577 517028
rect 182635 516994 182669 517028
rect 182727 516994 182761 517028
rect 182819 516994 182853 517028
rect 182911 516994 182945 517028
rect 183003 516994 183037 517028
rect 183095 516994 183129 517028
rect 183187 516994 183221 517028
rect 183279 516994 183313 517028
rect 183371 516994 183405 517028
rect 183463 516994 183497 517028
rect 183555 516994 183589 517028
rect 183647 516994 183681 517028
rect 183739 516994 183773 517028
rect 183831 516994 183865 517028
rect 183923 516994 183957 517028
rect 184015 516994 184049 517028
rect 184107 516994 184141 517028
rect 184199 516994 184233 517028
rect 184291 516994 184325 517028
rect 184383 516994 184417 517028
rect 184475 516994 184509 517028
rect 184567 516994 184601 517028
rect 184659 516994 184693 517028
rect 184751 516994 184785 517028
rect 184843 516994 184877 517028
rect 184935 516994 184969 517028
rect 185027 516994 185061 517028
rect 185119 516994 185153 517028
rect 185211 516994 185245 517028
rect 185303 516994 185337 517028
rect 185395 516994 185429 517028
rect 185487 516994 185521 517028
rect 185579 516994 185613 517028
rect 185671 516994 185705 517028
rect 185763 516994 185797 517028
rect 185855 516994 185889 517028
rect 185947 516994 185981 517028
rect 186039 516994 186073 517028
rect 186131 516994 186165 517028
rect 186223 516994 186257 517028
rect 186315 516994 186349 517028
rect 186407 516994 186441 517028
rect 186499 516994 186533 517028
rect 186591 516994 186625 517028
rect 186683 516994 186717 517028
rect 186775 516994 186809 517028
rect 186867 516994 186901 517028
rect 186959 516994 186993 517028
rect 187051 516994 187085 517028
rect 187143 516994 187177 517028
rect 187235 516994 187269 517028
rect 187327 516994 187361 517028
rect 187419 516994 187453 517028
rect 172239 516450 172273 516484
rect 172331 516450 172365 516484
rect 172423 516450 172457 516484
rect 172515 516450 172549 516484
rect 172607 516450 172641 516484
rect 172699 516450 172733 516484
rect 172791 516450 172825 516484
rect 172883 516450 172917 516484
rect 172975 516450 173009 516484
rect 173067 516450 173101 516484
rect 173159 516450 173193 516484
rect 173251 516450 173285 516484
rect 173343 516450 173377 516484
rect 173435 516450 173469 516484
rect 173527 516450 173561 516484
rect 173619 516450 173653 516484
rect 173711 516450 173745 516484
rect 173803 516450 173837 516484
rect 173895 516450 173929 516484
rect 173987 516450 174021 516484
rect 174079 516450 174113 516484
rect 174171 516450 174205 516484
rect 174263 516450 174297 516484
rect 174355 516450 174389 516484
rect 174447 516450 174481 516484
rect 174539 516450 174573 516484
rect 174631 516450 174665 516484
rect 174723 516450 174757 516484
rect 174815 516450 174849 516484
rect 174907 516450 174941 516484
rect 174999 516450 175033 516484
rect 175091 516450 175125 516484
rect 175183 516450 175217 516484
rect 175275 516450 175309 516484
rect 175367 516450 175401 516484
rect 175459 516450 175493 516484
rect 175551 516450 175585 516484
rect 175643 516450 175677 516484
rect 175735 516450 175769 516484
rect 175827 516450 175861 516484
rect 175919 516450 175953 516484
rect 176011 516450 176045 516484
rect 176103 516450 176137 516484
rect 176195 516450 176229 516484
rect 176287 516450 176321 516484
rect 176379 516450 176413 516484
rect 176471 516450 176505 516484
rect 176563 516450 176597 516484
rect 176655 516450 176689 516484
rect 176747 516450 176781 516484
rect 176839 516450 176873 516484
rect 176931 516450 176965 516484
rect 177023 516450 177057 516484
rect 177115 516450 177149 516484
rect 177207 516450 177241 516484
rect 177299 516450 177333 516484
rect 177391 516450 177425 516484
rect 177483 516450 177517 516484
rect 177575 516450 177609 516484
rect 177667 516450 177701 516484
rect 177759 516450 177793 516484
rect 177851 516450 177885 516484
rect 177943 516450 177977 516484
rect 178035 516450 178069 516484
rect 178127 516450 178161 516484
rect 178219 516450 178253 516484
rect 178311 516450 178345 516484
rect 178403 516450 178437 516484
rect 178495 516450 178529 516484
rect 178587 516450 178621 516484
rect 178679 516450 178713 516484
rect 178771 516450 178805 516484
rect 178863 516450 178897 516484
rect 178955 516450 178989 516484
rect 179047 516450 179081 516484
rect 179139 516450 179173 516484
rect 179231 516450 179265 516484
rect 179323 516450 179357 516484
rect 179415 516450 179449 516484
rect 179507 516450 179541 516484
rect 179599 516450 179633 516484
rect 179691 516450 179725 516484
rect 179783 516450 179817 516484
rect 179875 516450 179909 516484
rect 179967 516450 180001 516484
rect 180059 516450 180093 516484
rect 180151 516450 180185 516484
rect 180243 516450 180277 516484
rect 180335 516450 180369 516484
rect 180427 516450 180461 516484
rect 180519 516450 180553 516484
rect 180611 516450 180645 516484
rect 180703 516450 180737 516484
rect 180795 516450 180829 516484
rect 180887 516450 180921 516484
rect 180979 516450 181013 516484
rect 181071 516450 181105 516484
rect 181163 516450 181197 516484
rect 181255 516450 181289 516484
rect 181347 516450 181381 516484
rect 181439 516450 181473 516484
rect 181531 516450 181565 516484
rect 181623 516450 181657 516484
rect 181715 516450 181749 516484
rect 181807 516450 181841 516484
rect 181899 516450 181933 516484
rect 181991 516450 182025 516484
rect 182083 516450 182117 516484
rect 182175 516450 182209 516484
rect 182267 516450 182301 516484
rect 182359 516450 182393 516484
rect 182451 516450 182485 516484
rect 182543 516450 182577 516484
rect 182635 516450 182669 516484
rect 182727 516450 182761 516484
rect 182819 516450 182853 516484
rect 182911 516450 182945 516484
rect 183003 516450 183037 516484
rect 183095 516450 183129 516484
rect 183187 516450 183221 516484
rect 183279 516450 183313 516484
rect 183371 516450 183405 516484
rect 183463 516450 183497 516484
rect 183555 516450 183589 516484
rect 183647 516450 183681 516484
rect 183739 516450 183773 516484
rect 183831 516450 183865 516484
rect 183923 516450 183957 516484
rect 184015 516450 184049 516484
rect 184107 516450 184141 516484
rect 184199 516450 184233 516484
rect 184291 516450 184325 516484
rect 184383 516450 184417 516484
rect 184475 516450 184509 516484
rect 184567 516450 184601 516484
rect 184659 516450 184693 516484
rect 184751 516450 184785 516484
rect 184843 516450 184877 516484
rect 184935 516450 184969 516484
rect 185027 516450 185061 516484
rect 185119 516450 185153 516484
rect 185211 516450 185245 516484
rect 185303 516450 185337 516484
rect 185395 516450 185429 516484
rect 185487 516450 185521 516484
rect 185579 516450 185613 516484
rect 185671 516450 185705 516484
rect 185763 516450 185797 516484
rect 185855 516450 185889 516484
rect 185947 516450 185981 516484
rect 186039 516450 186073 516484
rect 186131 516450 186165 516484
rect 186223 516450 186257 516484
rect 186315 516450 186349 516484
rect 186407 516450 186441 516484
rect 186499 516450 186533 516484
rect 186591 516450 186625 516484
rect 186683 516450 186717 516484
rect 186775 516450 186809 516484
rect 186867 516450 186901 516484
rect 186959 516450 186993 516484
rect 187051 516450 187085 516484
rect 187143 516450 187177 516484
rect 187235 516450 187269 516484
rect 187327 516450 187361 516484
rect 187419 516450 187453 516484
rect 172239 515906 172273 515940
rect 172331 515906 172365 515940
rect 172423 515906 172457 515940
rect 172515 515906 172549 515940
rect 172607 515906 172641 515940
rect 172699 515906 172733 515940
rect 172791 515906 172825 515940
rect 172883 515906 172917 515940
rect 172975 515906 173009 515940
rect 173067 515906 173101 515940
rect 173159 515906 173193 515940
rect 173251 515906 173285 515940
rect 173343 515906 173377 515940
rect 173435 515906 173469 515940
rect 173527 515906 173561 515940
rect 173619 515906 173653 515940
rect 173711 515906 173745 515940
rect 173803 515906 173837 515940
rect 173895 515906 173929 515940
rect 173987 515906 174021 515940
rect 174079 515906 174113 515940
rect 174171 515906 174205 515940
rect 174263 515906 174297 515940
rect 174355 515906 174389 515940
rect 174447 515906 174481 515940
rect 174539 515906 174573 515940
rect 174631 515906 174665 515940
rect 174723 515906 174757 515940
rect 174815 515906 174849 515940
rect 174907 515906 174941 515940
rect 174999 515906 175033 515940
rect 175091 515906 175125 515940
rect 175183 515906 175217 515940
rect 175275 515906 175309 515940
rect 175367 515906 175401 515940
rect 175459 515906 175493 515940
rect 175551 515906 175585 515940
rect 175643 515906 175677 515940
rect 175735 515906 175769 515940
rect 175827 515906 175861 515940
rect 175919 515906 175953 515940
rect 176011 515906 176045 515940
rect 176103 515906 176137 515940
rect 176195 515906 176229 515940
rect 176287 515906 176321 515940
rect 176379 515906 176413 515940
rect 176471 515906 176505 515940
rect 176563 515906 176597 515940
rect 176655 515906 176689 515940
rect 176747 515906 176781 515940
rect 176839 515906 176873 515940
rect 176931 515906 176965 515940
rect 177023 515906 177057 515940
rect 177115 515906 177149 515940
rect 177207 515906 177241 515940
rect 177299 515906 177333 515940
rect 177391 515906 177425 515940
rect 177483 515906 177517 515940
rect 177575 515906 177609 515940
rect 177667 515906 177701 515940
rect 177759 515906 177793 515940
rect 177851 515906 177885 515940
rect 177943 515906 177977 515940
rect 178035 515906 178069 515940
rect 178127 515906 178161 515940
rect 178219 515906 178253 515940
rect 178311 515906 178345 515940
rect 178403 515906 178437 515940
rect 178495 515906 178529 515940
rect 178587 515906 178621 515940
rect 178679 515906 178713 515940
rect 178771 515906 178805 515940
rect 178863 515906 178897 515940
rect 178955 515906 178989 515940
rect 179047 515906 179081 515940
rect 179139 515906 179173 515940
rect 179231 515906 179265 515940
rect 179323 515906 179357 515940
rect 179415 515906 179449 515940
rect 179507 515906 179541 515940
rect 179599 515906 179633 515940
rect 179691 515906 179725 515940
rect 179783 515906 179817 515940
rect 179875 515906 179909 515940
rect 179967 515906 180001 515940
rect 180059 515906 180093 515940
rect 180151 515906 180185 515940
rect 180243 515906 180277 515940
rect 180335 515906 180369 515940
rect 180427 515906 180461 515940
rect 180519 515906 180553 515940
rect 180611 515906 180645 515940
rect 180703 515906 180737 515940
rect 180795 515906 180829 515940
rect 180887 515906 180921 515940
rect 180979 515906 181013 515940
rect 181071 515906 181105 515940
rect 181163 515906 181197 515940
rect 181255 515906 181289 515940
rect 181347 515906 181381 515940
rect 181439 515906 181473 515940
rect 181531 515906 181565 515940
rect 181623 515906 181657 515940
rect 181715 515906 181749 515940
rect 181807 515906 181841 515940
rect 181899 515906 181933 515940
rect 181991 515906 182025 515940
rect 182083 515906 182117 515940
rect 182175 515906 182209 515940
rect 182267 515906 182301 515940
rect 182359 515906 182393 515940
rect 182451 515906 182485 515940
rect 182543 515906 182577 515940
rect 182635 515906 182669 515940
rect 182727 515906 182761 515940
rect 182819 515906 182853 515940
rect 182911 515906 182945 515940
rect 183003 515906 183037 515940
rect 183095 515906 183129 515940
rect 183187 515906 183221 515940
rect 183279 515906 183313 515940
rect 183371 515906 183405 515940
rect 183463 515906 183497 515940
rect 183555 515906 183589 515940
rect 183647 515906 183681 515940
rect 183739 515906 183773 515940
rect 183831 515906 183865 515940
rect 183923 515906 183957 515940
rect 184015 515906 184049 515940
rect 184107 515906 184141 515940
rect 184199 515906 184233 515940
rect 184291 515906 184325 515940
rect 184383 515906 184417 515940
rect 184475 515906 184509 515940
rect 184567 515906 184601 515940
rect 184659 515906 184693 515940
rect 184751 515906 184785 515940
rect 184843 515906 184877 515940
rect 184935 515906 184969 515940
rect 185027 515906 185061 515940
rect 185119 515906 185153 515940
rect 185211 515906 185245 515940
rect 185303 515906 185337 515940
rect 185395 515906 185429 515940
rect 185487 515906 185521 515940
rect 185579 515906 185613 515940
rect 185671 515906 185705 515940
rect 185763 515906 185797 515940
rect 185855 515906 185889 515940
rect 185947 515906 185981 515940
rect 186039 515906 186073 515940
rect 186131 515906 186165 515940
rect 186223 515906 186257 515940
rect 186315 515906 186349 515940
rect 186407 515906 186441 515940
rect 186499 515906 186533 515940
rect 186591 515906 186625 515940
rect 186683 515906 186717 515940
rect 186775 515906 186809 515940
rect 186867 515906 186901 515940
rect 186959 515906 186993 515940
rect 187051 515906 187085 515940
rect 187143 515906 187177 515940
rect 187235 515906 187269 515940
rect 187327 515906 187361 515940
rect 187419 515906 187453 515940
rect 173619 515829 173653 515838
rect 173619 515804 173623 515829
rect 173623 515804 173653 515829
rect 173527 515532 173561 515566
rect 182083 515822 182089 515838
rect 182089 515822 182117 515838
rect 182083 515804 182117 515822
rect 182267 515628 182301 515634
rect 182267 515600 182293 515628
rect 182293 515600 182301 515628
rect 186591 515829 186625 515838
rect 186591 515804 186595 515829
rect 186595 515804 186625 515829
rect 186499 515532 186533 515566
rect 172239 515362 172273 515396
rect 172331 515362 172365 515396
rect 172423 515362 172457 515396
rect 172515 515362 172549 515396
rect 172607 515362 172641 515396
rect 172699 515362 172733 515396
rect 172791 515362 172825 515396
rect 172883 515362 172917 515396
rect 172975 515362 173009 515396
rect 173067 515362 173101 515396
rect 173159 515362 173193 515396
rect 173251 515362 173285 515396
rect 173343 515362 173377 515396
rect 173435 515362 173469 515396
rect 173527 515362 173561 515396
rect 173619 515362 173653 515396
rect 173711 515362 173745 515396
rect 173803 515362 173837 515396
rect 173895 515362 173929 515396
rect 173987 515362 174021 515396
rect 174079 515362 174113 515396
rect 174171 515362 174205 515396
rect 174263 515362 174297 515396
rect 174355 515362 174389 515396
rect 174447 515362 174481 515396
rect 174539 515362 174573 515396
rect 174631 515362 174665 515396
rect 174723 515362 174757 515396
rect 174815 515362 174849 515396
rect 174907 515362 174941 515396
rect 174999 515362 175033 515396
rect 175091 515362 175125 515396
rect 175183 515362 175217 515396
rect 175275 515362 175309 515396
rect 175367 515362 175401 515396
rect 175459 515362 175493 515396
rect 175551 515362 175585 515396
rect 175643 515362 175677 515396
rect 175735 515362 175769 515396
rect 175827 515362 175861 515396
rect 175919 515362 175953 515396
rect 176011 515362 176045 515396
rect 176103 515362 176137 515396
rect 176195 515362 176229 515396
rect 176287 515362 176321 515396
rect 176379 515362 176413 515396
rect 176471 515362 176505 515396
rect 176563 515362 176597 515396
rect 176655 515362 176689 515396
rect 176747 515362 176781 515396
rect 176839 515362 176873 515396
rect 176931 515362 176965 515396
rect 177023 515362 177057 515396
rect 177115 515362 177149 515396
rect 177207 515362 177241 515396
rect 177299 515362 177333 515396
rect 177391 515362 177425 515396
rect 177483 515362 177517 515396
rect 177575 515362 177609 515396
rect 177667 515362 177701 515396
rect 177759 515362 177793 515396
rect 177851 515362 177885 515396
rect 177943 515362 177977 515396
rect 178035 515362 178069 515396
rect 178127 515362 178161 515396
rect 178219 515362 178253 515396
rect 178311 515362 178345 515396
rect 178403 515362 178437 515396
rect 178495 515362 178529 515396
rect 178587 515362 178621 515396
rect 178679 515362 178713 515396
rect 178771 515362 178805 515396
rect 178863 515362 178897 515396
rect 178955 515362 178989 515396
rect 179047 515362 179081 515396
rect 179139 515362 179173 515396
rect 179231 515362 179265 515396
rect 179323 515362 179357 515396
rect 179415 515362 179449 515396
rect 179507 515362 179541 515396
rect 179599 515362 179633 515396
rect 179691 515362 179725 515396
rect 179783 515362 179817 515396
rect 179875 515362 179909 515396
rect 179967 515362 180001 515396
rect 180059 515362 180093 515396
rect 180151 515362 180185 515396
rect 180243 515362 180277 515396
rect 180335 515362 180369 515396
rect 180427 515362 180461 515396
rect 180519 515362 180553 515396
rect 180611 515362 180645 515396
rect 180703 515362 180737 515396
rect 180795 515362 180829 515396
rect 180887 515362 180921 515396
rect 180979 515362 181013 515396
rect 181071 515362 181105 515396
rect 181163 515362 181197 515396
rect 181255 515362 181289 515396
rect 181347 515362 181381 515396
rect 181439 515362 181473 515396
rect 181531 515362 181565 515396
rect 181623 515362 181657 515396
rect 181715 515362 181749 515396
rect 181807 515362 181841 515396
rect 181899 515362 181933 515396
rect 181991 515362 182025 515396
rect 182083 515362 182117 515396
rect 182175 515362 182209 515396
rect 182267 515362 182301 515396
rect 182359 515362 182393 515396
rect 182451 515362 182485 515396
rect 182543 515362 182577 515396
rect 182635 515362 182669 515396
rect 182727 515362 182761 515396
rect 182819 515362 182853 515396
rect 182911 515362 182945 515396
rect 183003 515362 183037 515396
rect 183095 515362 183129 515396
rect 183187 515362 183221 515396
rect 183279 515362 183313 515396
rect 183371 515362 183405 515396
rect 183463 515362 183497 515396
rect 183555 515362 183589 515396
rect 183647 515362 183681 515396
rect 183739 515362 183773 515396
rect 183831 515362 183865 515396
rect 183923 515362 183957 515396
rect 184015 515362 184049 515396
rect 184107 515362 184141 515396
rect 184199 515362 184233 515396
rect 184291 515362 184325 515396
rect 184383 515362 184417 515396
rect 184475 515362 184509 515396
rect 184567 515362 184601 515396
rect 184659 515362 184693 515396
rect 184751 515362 184785 515396
rect 184843 515362 184877 515396
rect 184935 515362 184969 515396
rect 185027 515362 185061 515396
rect 185119 515362 185153 515396
rect 185211 515362 185245 515396
rect 185303 515362 185337 515396
rect 185395 515362 185429 515396
rect 185487 515362 185521 515396
rect 185579 515362 185613 515396
rect 185671 515362 185705 515396
rect 185763 515362 185797 515396
rect 185855 515362 185889 515396
rect 185947 515362 185981 515396
rect 186039 515362 186073 515396
rect 186131 515362 186165 515396
rect 186223 515362 186257 515396
rect 186315 515362 186349 515396
rect 186407 515362 186441 515396
rect 186499 515362 186533 515396
rect 186591 515362 186625 515396
rect 186683 515362 186717 515396
rect 186775 515362 186809 515396
rect 186867 515362 186901 515396
rect 186959 515362 186993 515396
rect 187051 515362 187085 515396
rect 187143 515362 187177 515396
rect 187235 515362 187269 515396
rect 187327 515362 187361 515396
rect 187419 515362 187453 515396
<< metal1 >>
rect 17990 699000 18000 701000
rect 20000 699000 20010 701000
rect 69990 699000 70000 701000
rect 72000 699000 72010 701000
rect 121990 699000 122000 701000
rect 124000 699000 124010 701000
rect 18000 687000 20000 699000
rect 70000 691000 72000 699000
rect 122000 695000 124000 699000
rect 122000 693000 156000 695000
rect 70000 689000 152000 691000
rect 18000 685000 148000 687000
rect 2990 682000 3000 684000
rect 5000 682000 11000 684000
rect 9000 533000 11000 682000
rect 146000 628000 148000 685000
rect 145990 626000 146000 628000
rect 148000 626000 148010 628000
rect 150000 549000 152000 689000
rect 154000 553000 156000 693000
rect 153990 551000 154000 553000
rect 156000 551000 156010 553000
rect 150000 547000 179000 549000
rect 145990 544000 146000 546000
rect 148000 544000 163800 546000
rect 177000 544000 179000 547000
rect 163500 543230 163800 544000
rect 153990 538000 154000 540000
rect 156000 538000 156010 540000
rect 163030 538897 163230 538907
rect 163020 538867 163030 538897
rect 158680 538747 163030 538867
rect 158680 538617 158980 538747
rect 158670 538537 158980 538617
rect 158670 538501 158960 538537
rect 158670 538467 158728 538501
rect 158896 538467 158960 538501
rect 158670 538429 158960 538467
rect 158660 538417 158964 538429
rect 158660 538241 158666 538417
rect 158700 538387 158924 538417
rect 158700 538241 158706 538387
rect 158660 538229 158706 538241
rect 158918 538241 158924 538387
rect 158958 538241 158964 538417
rect 159030 538427 159060 538747
rect 161380 538697 161530 538707
rect 161380 538577 161390 538697
rect 161510 538577 161530 538697
rect 161380 538567 161530 538577
rect 159092 538501 159284 538507
rect 159092 538467 159104 538501
rect 159272 538467 159284 538501
rect 159092 538461 159284 538467
rect 159350 538501 159542 538507
rect 159350 538467 159362 538501
rect 159530 538467 159542 538501
rect 159350 538461 159542 538467
rect 159608 538501 159800 538507
rect 159608 538467 159620 538501
rect 159788 538467 159800 538501
rect 159608 538461 159800 538467
rect 159866 538501 160058 538507
rect 159866 538467 159878 538501
rect 160046 538467 160058 538501
rect 159866 538461 160058 538467
rect 160124 538501 160316 538507
rect 160124 538467 160136 538501
rect 160304 538467 160316 538501
rect 160124 538461 160316 538467
rect 160382 538501 160574 538507
rect 160382 538467 160394 538501
rect 160562 538467 160574 538501
rect 160382 538461 160574 538467
rect 160640 538501 160832 538507
rect 160640 538467 160652 538501
rect 160820 538467 160832 538501
rect 160640 538461 160832 538467
rect 160898 538501 161090 538507
rect 160898 538467 160910 538501
rect 161078 538467 161090 538501
rect 160898 538461 161090 538467
rect 161156 538501 161348 538507
rect 161156 538467 161168 538501
rect 161336 538467 161348 538501
rect 161156 538461 161348 538467
rect 161440 538429 161500 538567
rect 161536 538501 161728 538507
rect 161536 538467 161548 538501
rect 161716 538467 161728 538501
rect 161536 538461 161728 538467
rect 161810 538437 161850 538747
rect 162260 538737 162560 538747
rect 162260 538697 162270 538737
rect 162530 538697 162560 538737
rect 163020 538697 163030 538747
rect 163330 538697 163340 538897
rect 161936 538501 162128 538507
rect 161936 538467 161948 538501
rect 162116 538467 162128 538501
rect 161936 538461 162128 538467
rect 162260 538501 162560 538697
rect 162260 538467 162328 538501
rect 162496 538467 162560 538501
rect 161750 538429 161910 538437
rect 162260 538429 162560 538467
rect 159030 538400 161150 538427
rect 159030 538387 159042 538400
rect 159036 538312 159042 538387
rect 159076 538387 159558 538400
rect 159076 538312 159082 538387
rect 159036 538300 159082 538312
rect 159294 538346 159340 538358
rect 159294 538267 159300 538346
rect 158918 538229 158964 538241
rect 159290 538258 159300 538267
rect 159334 538267 159340 538346
rect 159390 538327 159490 538337
rect 159390 538267 159400 538327
rect 159334 538258 159400 538267
rect 159290 538247 159400 538258
rect 159480 538267 159490 538327
rect 159552 538312 159558 538387
rect 159592 538387 160074 538400
rect 159592 538312 159598 538387
rect 159552 538300 159598 538312
rect 159810 538346 159856 538358
rect 159810 538267 159816 538346
rect 159480 538258 159816 538267
rect 159850 538267 159856 538346
rect 160068 538312 160074 538387
rect 160108 538387 160590 538400
rect 160108 538312 160114 538387
rect 160068 538300 160114 538312
rect 160326 538346 160372 538358
rect 160326 538267 160332 538346
rect 159850 538258 160332 538267
rect 160366 538267 160372 538346
rect 160584 538312 160590 538387
rect 160624 538387 161106 538400
rect 160624 538312 160630 538387
rect 160584 538300 160630 538312
rect 160842 538346 160888 538358
rect 160842 538267 160848 538346
rect 160366 538258 160848 538267
rect 160882 538267 160888 538346
rect 161100 538312 161106 538387
rect 161140 538387 161150 538400
rect 161440 538417 161526 538429
rect 161140 538312 161146 538387
rect 161100 538300 161146 538312
rect 161358 538346 161404 538358
rect 161358 538267 161364 538346
rect 160882 538258 161364 538267
rect 161398 538258 161404 538346
rect 159480 538247 161404 538258
rect 159290 538246 161404 538247
rect 159290 538227 161390 538246
rect 161440 538241 161486 538417
rect 161520 538241 161526 538417
rect 161440 538229 161526 538241
rect 161738 538417 161926 538429
rect 161738 538241 161744 538417
rect 161778 538241 161886 538417
rect 161920 538377 161926 538417
rect 162138 538417 162184 538429
rect 161920 538337 161930 538377
rect 161920 538241 161926 538337
rect 161738 538237 161926 538241
rect 161738 538229 161784 538237
rect 161880 538229 161926 538237
rect 162138 538241 162144 538417
rect 162178 538397 162184 538417
rect 162260 538417 162564 538429
rect 162178 538257 162190 538397
rect 162178 538241 162210 538257
rect 162138 538229 162210 538241
rect 162260 538241 162266 538417
rect 162300 538337 162524 538417
rect 162300 538241 162306 538337
rect 162260 538229 162306 538241
rect 162518 538241 162524 538337
rect 162558 538241 162564 538417
rect 162518 538229 162564 538241
rect 161440 538227 161500 538229
rect 158716 538191 158908 538197
rect 158716 538157 158728 538191
rect 158896 538157 158908 538191
rect 159092 538191 159284 538197
rect 159092 538187 159104 538191
rect 158716 538151 158908 538157
rect 159090 538157 159104 538187
rect 159272 538187 159284 538191
rect 159350 538191 159542 538197
rect 159350 538187 159362 538191
rect 159272 538157 159362 538187
rect 159530 538187 159542 538191
rect 159608 538191 159800 538197
rect 159608 538187 159620 538191
rect 159530 538157 159620 538187
rect 159788 538187 159800 538191
rect 159866 538191 160058 538197
rect 159866 538187 159878 538191
rect 159788 538157 159878 538187
rect 160046 538187 160058 538191
rect 160124 538191 160316 538197
rect 160124 538187 160136 538191
rect 160046 538157 160136 538187
rect 160304 538187 160316 538191
rect 160382 538191 160574 538197
rect 160382 538187 160394 538191
rect 160304 538157 160394 538187
rect 160562 538187 160574 538191
rect 160640 538191 160832 538197
rect 160640 538187 160652 538191
rect 160562 538157 160652 538187
rect 160820 538187 160832 538191
rect 160898 538191 161090 538197
rect 160898 538187 160910 538191
rect 160820 538157 160910 538187
rect 161078 538187 161090 538191
rect 161156 538191 161348 538197
rect 161156 538187 161168 538191
rect 161078 538157 161168 538187
rect 161336 538187 161348 538191
rect 161450 538187 161490 538227
rect 162170 538197 162210 538229
rect 161336 538157 161490 538187
rect 161530 538191 162210 538197
rect 161530 538157 161548 538191
rect 161716 538157 161948 538191
rect 162116 538157 162210 538191
rect 159090 538147 161490 538157
rect 161536 538151 161728 538157
rect 161936 538151 162128 538157
rect 154000 537000 156000 538000
rect 161450 537997 161490 538147
rect 162170 537997 162210 538157
rect 162316 538191 162508 538197
rect 162316 538157 162328 538191
rect 162496 538157 162508 538191
rect 162316 538151 162508 538157
rect 163530 538067 163730 543230
rect 178100 543004 178400 544000
rect 178180 541737 178380 543004
rect 164280 541537 188980 541737
rect 164280 540997 164480 541537
rect 164720 541157 164780 541167
rect 165020 541162 166040 541187
rect 165020 541158 166255 541162
rect 164680 541151 164820 541157
rect 164680 541117 164730 541151
rect 164764 541117 164820 541151
rect 165020 541127 165033 541158
rect 165021 541124 165033 541127
rect 165067 541127 165225 541158
rect 165067 541124 165079 541127
rect 165021 541118 165079 541124
rect 165213 541124 165225 541127
rect 165259 541127 165417 541158
rect 165259 541124 165271 541127
rect 165213 541118 165271 541124
rect 165405 541124 165417 541127
rect 165451 541127 165609 541158
rect 165451 541124 165463 541127
rect 165405 541118 165463 541124
rect 165597 541124 165609 541127
rect 165643 541127 165801 541158
rect 165643 541124 165655 541127
rect 165597 541118 165655 541124
rect 165789 541124 165801 541127
rect 165835 541127 165993 541158
rect 165835 541124 165847 541127
rect 165789 541118 165847 541124
rect 165981 541124 165993 541127
rect 166027 541124 166255 541158
rect 165981 541118 166255 541124
rect 164680 541050 164820 541117
rect 166025 541112 166255 541118
rect 164680 540997 164686 541050
rect 164280 540917 164686 540997
rect 164280 540867 164480 540917
rect 164680 540562 164686 540917
rect 164720 540917 164774 541050
rect 164720 540562 164726 540917
rect 164680 540550 164726 540562
rect 164768 540562 164774 540917
rect 164808 540997 164820 541050
rect 164979 541057 165025 541069
rect 165171 541057 165217 541069
rect 165363 541057 165409 541069
rect 165555 541057 165601 541069
rect 165747 541057 165793 541069
rect 165939 541057 165985 541069
rect 164979 540997 164985 541057
rect 164808 540917 164985 540997
rect 164808 540562 164814 540917
rect 164768 540550 164814 540562
rect 164883 540603 164929 540615
rect 164883 540317 164889 540603
rect 164850 540115 164889 540317
rect 164923 540317 164929 540603
rect 164979 540569 164985 540917
rect 165019 540667 165177 541057
rect 165019 540569 165025 540667
rect 164979 540557 165025 540569
rect 165075 540603 165121 540615
rect 165075 540317 165081 540603
rect 164923 540115 165081 540317
rect 165115 540317 165121 540603
rect 165171 540569 165177 540667
rect 165211 540667 165369 541057
rect 165211 540569 165217 540667
rect 165171 540557 165217 540569
rect 165267 540603 165313 540615
rect 165267 540317 165273 540603
rect 165115 540115 165273 540317
rect 165307 540317 165313 540603
rect 165363 540569 165369 540667
rect 165403 540667 165561 541057
rect 165403 540569 165409 540667
rect 165363 540557 165409 540569
rect 165459 540603 165505 540615
rect 165459 540317 165465 540603
rect 165307 540115 165465 540317
rect 165499 540317 165505 540603
rect 165555 540569 165561 540667
rect 165595 540667 165753 541057
rect 165595 540569 165601 540667
rect 165555 540557 165601 540569
rect 165651 540603 165697 540615
rect 165651 540317 165657 540603
rect 165499 540115 165657 540317
rect 165691 540317 165697 540603
rect 165747 540569 165753 540667
rect 165787 541027 165945 541057
rect 165979 541027 166010 541057
rect 165787 540927 165890 541027
rect 166000 540927 166010 541027
rect 165787 540907 165945 540927
rect 165979 540907 166010 540927
rect 165787 540807 165890 540907
rect 166000 540807 166010 540907
rect 166205 540862 166255 541112
rect 166398 541151 166460 541157
rect 166398 541117 166410 541151
rect 166444 541117 166460 541151
rect 166398 541111 166460 541117
rect 166400 541097 166460 541111
rect 168080 540997 168280 541537
rect 168520 541157 168580 541167
rect 168820 541162 169840 541187
rect 168820 541158 170055 541162
rect 168480 541151 168620 541157
rect 168480 541117 168530 541151
rect 168564 541117 168620 541151
rect 168820 541127 168833 541158
rect 168821 541124 168833 541127
rect 168867 541127 169025 541158
rect 168867 541124 168879 541127
rect 168821 541118 168879 541124
rect 169013 541124 169025 541127
rect 169059 541127 169217 541158
rect 169059 541124 169071 541127
rect 169013 541118 169071 541124
rect 169205 541124 169217 541127
rect 169251 541127 169409 541158
rect 169251 541124 169263 541127
rect 169205 541118 169263 541124
rect 169397 541124 169409 541127
rect 169443 541127 169601 541158
rect 169443 541124 169455 541127
rect 169397 541118 169455 541124
rect 169589 541124 169601 541127
rect 169635 541127 169793 541158
rect 169635 541124 169647 541127
rect 169589 541118 169647 541124
rect 169781 541124 169793 541127
rect 169827 541124 170055 541158
rect 169781 541118 170055 541124
rect 168480 541050 168620 541117
rect 169825 541112 170055 541118
rect 168480 540997 168486 541050
rect 166680 540862 167720 540927
rect 168080 540917 168486 540997
rect 168080 540867 168280 540917
rect 165787 540787 165945 540807
rect 165979 540787 166010 540807
rect 165787 540687 165890 540787
rect 166000 540687 166010 540787
rect 165787 540667 165945 540687
rect 165787 540569 165793 540667
rect 165747 540557 165793 540569
rect 165843 540603 165889 540615
rect 165843 540317 165849 540603
rect 165691 540115 165849 540317
rect 165883 540317 165889 540603
rect 165939 540569 165945 540667
rect 165979 540667 166010 540687
rect 166200 540812 167720 540862
rect 165979 540569 165985 540667
rect 165939 540557 165985 540569
rect 166035 540603 166081 540615
rect 166035 540317 166041 540603
rect 165883 540115 166041 540317
rect 166075 540115 166081 540603
rect 166200 540367 166250 540812
rect 166680 540727 167720 540812
rect 166360 540596 166406 540608
rect 166200 540357 166260 540367
rect 166198 540351 166260 540357
rect 166198 540317 166210 540351
rect 166244 540317 166260 540351
rect 166198 540311 166260 540317
rect 166200 540307 166260 540311
rect 166160 540267 166206 540279
rect 166160 540187 166166 540267
rect 164850 540107 166081 540115
rect 164850 540103 164929 540107
rect 165075 540103 165121 540107
rect 165267 540103 165313 540107
rect 165459 540103 165505 540107
rect 165651 540103 165697 540107
rect 165843 540103 165889 540107
rect 166035 540103 166081 540107
rect 164850 540097 164920 540103
rect 164710 540041 164780 540057
rect 164710 540007 164730 540041
rect 164764 540007 164780 540041
rect 164710 539987 164780 540007
rect 164850 539787 164880 540097
rect 166140 540091 166166 540187
rect 166200 540091 166206 540267
rect 166140 540079 166206 540091
rect 166248 540267 166294 540279
rect 166248 540091 166254 540267
rect 166288 540257 166294 540267
rect 166360 540257 166366 540596
rect 166288 540108 166366 540257
rect 166400 540267 166406 540596
rect 166448 540596 166494 540608
rect 166448 540267 166454 540596
rect 166400 540108 166454 540267
rect 166488 540267 166494 540596
rect 166670 540277 166890 540287
rect 166488 540257 166510 540267
rect 166670 540257 166690 540277
rect 166488 540247 166690 540257
rect 166488 540117 166570 540247
rect 166630 540117 166690 540247
rect 166488 540108 166690 540117
rect 166288 540107 166690 540108
rect 166288 540091 166294 540107
rect 166360 540096 166494 540107
rect 166670 540097 166690 540107
rect 166870 540097 166890 540277
rect 166248 540079 166294 540091
rect 164925 540048 164983 540054
rect 164925 540047 164937 540048
rect 164920 540014 164937 540047
rect 164971 540047 164983 540048
rect 165117 540048 165175 540054
rect 165117 540047 165129 540048
rect 164971 540014 165129 540047
rect 165163 540047 165175 540048
rect 165309 540048 165367 540054
rect 165309 540047 165321 540048
rect 165163 540014 165321 540047
rect 165355 540047 165367 540048
rect 165501 540048 165559 540054
rect 165501 540047 165513 540048
rect 165355 540014 165513 540047
rect 165547 540047 165559 540048
rect 165693 540048 165751 540054
rect 165693 540047 165705 540048
rect 165547 540014 165705 540047
rect 165739 540047 165751 540048
rect 165885 540048 165943 540054
rect 165885 540047 165897 540048
rect 165739 540014 165897 540047
rect 165931 540014 165943 540048
rect 164920 540008 165943 540014
rect 164920 539987 165940 540008
rect 161450 537957 161650 537997
rect 161290 537738 161350 537757
rect 161290 537704 161304 537738
rect 161338 537704 161350 537738
rect 161290 537697 161350 537704
rect 161490 537744 161550 537757
rect 161490 537738 161554 537744
rect 161490 537704 161508 537738
rect 161542 537704 161554 537738
rect 161490 537698 161554 537704
rect 161490 537697 161550 537698
rect 161610 537657 161650 537957
rect 162010 537957 162210 537997
rect 162870 537977 162950 537987
rect 161680 537767 161760 537777
rect 161680 537707 161690 537767
rect 161750 537707 161760 537767
rect 161680 537704 161700 537707
rect 161734 537704 161760 537707
rect 161680 537697 161760 537704
rect 161890 537744 161950 537757
rect 161890 537738 161954 537744
rect 161890 537704 161908 537738
rect 161942 537704 161954 537738
rect 161890 537698 161954 537704
rect 161890 537697 161950 537698
rect 161550 537640 161770 537657
rect 162010 537640 162050 537957
rect 162870 537917 162880 537977
rect 162940 537967 162950 537977
rect 163020 537967 163730 538067
rect 162940 537917 163730 537967
rect 162870 537907 162950 537917
rect 163020 537867 163730 537917
rect 164280 539687 164880 539787
rect 164280 537963 164480 539687
rect 164640 539638 164880 539687
rect 164640 539604 164714 539638
rect 164748 539604 164880 539638
rect 164640 539545 164880 539604
rect 165020 539651 166030 539657
rect 165020 539645 166043 539651
rect 165020 539611 165037 539645
rect 165071 539611 165229 539645
rect 165263 539611 165421 539645
rect 165455 539611 165613 539645
rect 165647 539611 165805 539645
rect 165839 539611 165997 539645
rect 166031 539611 166043 539645
rect 165020 539605 166043 539611
rect 165020 539597 166030 539605
rect 166140 539557 166170 540079
rect 166198 540041 166260 540047
rect 166198 540007 166210 540041
rect 166244 540007 166260 540041
rect 166198 540001 166260 540007
rect 166200 539638 166260 540001
rect 166370 540041 166490 540096
rect 166670 540087 166890 540097
rect 166370 540007 166410 540041
rect 166444 540007 166490 540041
rect 166370 539987 166490 540007
rect 166200 539604 166214 539638
rect 166248 539604 166260 539638
rect 166200 539597 166260 539604
rect 166400 539638 166480 539657
rect 166400 539604 166414 539638
rect 166448 539604 166480 539638
rect 166400 539597 166480 539604
rect 164640 539447 164670 539545
rect 164664 538569 164670 539447
rect 164704 539447 164758 539545
rect 164704 538569 164710 539447
rect 164664 538557 164710 538569
rect 164752 538569 164758 539447
rect 164792 539527 164880 539545
rect 164983 539535 165029 539547
rect 164792 539517 164950 539527
rect 164983 539517 164989 539535
rect 164792 539447 164989 539517
rect 164792 538569 164798 539447
rect 164850 539237 164989 539447
rect 164887 539081 164933 539093
rect 164887 538593 164893 539081
rect 164927 538967 164933 539081
rect 164983 539047 164989 539237
rect 165023 539517 165029 539535
rect 165175 539535 165221 539547
rect 165175 539517 165181 539535
rect 165023 539237 165181 539517
rect 165023 539047 165029 539237
rect 164983 539035 165029 539047
rect 165079 539081 165125 539093
rect 165079 538967 165085 539081
rect 164927 538593 165085 538967
rect 165119 538967 165125 539081
rect 165175 539047 165181 539237
rect 165215 539517 165221 539535
rect 165367 539535 165413 539547
rect 165367 539517 165373 539535
rect 165215 539237 165373 539517
rect 165215 539047 165221 539237
rect 165175 539035 165221 539047
rect 165271 539081 165317 539093
rect 165271 538967 165277 539081
rect 165119 538593 165277 538967
rect 165311 538967 165317 539081
rect 165367 539047 165373 539237
rect 165407 539517 165413 539535
rect 165559 539535 165605 539547
rect 165559 539517 165565 539535
rect 165407 539237 165565 539517
rect 165407 539047 165413 539237
rect 165367 539035 165413 539047
rect 165463 539081 165509 539093
rect 165463 538967 165469 539081
rect 165311 538593 165469 538967
rect 165503 538967 165509 539081
rect 165559 539047 165565 539237
rect 165599 539517 165605 539535
rect 165751 539535 165797 539547
rect 165751 539517 165757 539535
rect 165599 539237 165757 539517
rect 165599 539047 165605 539237
rect 165559 539035 165605 539047
rect 165655 539081 165701 539093
rect 165655 538967 165661 539081
rect 165503 538593 165661 538967
rect 165695 538967 165701 539081
rect 165751 539047 165757 539237
rect 165791 539517 165797 539535
rect 165943 539535 165989 539547
rect 165943 539517 165949 539535
rect 165791 539237 165949 539517
rect 165791 539047 165797 539237
rect 165751 539035 165797 539047
rect 165847 539081 165893 539093
rect 165847 538967 165853 539081
rect 165695 538593 165853 538967
rect 165887 538967 165893 539081
rect 165943 539047 165949 539237
rect 165983 539517 165989 539535
rect 166140 539545 166210 539557
rect 165983 539237 166000 539517
rect 166140 539407 166170 539545
rect 165983 539047 165989 539237
rect 165943 539035 165989 539047
rect 166039 539081 166085 539093
rect 166039 538967 166045 539081
rect 165887 538837 166045 538967
rect 165887 538737 165900 538837
rect 166040 538737 166045 538837
rect 165887 538593 166045 538737
rect 166079 538593 166085 539081
rect 166164 539067 166170 539407
rect 164887 538587 166085 538593
rect 164887 538581 164933 538587
rect 165079 538581 165125 538587
rect 165271 538581 165317 538587
rect 165463 538581 165509 538587
rect 165655 538581 165701 538587
rect 165847 538581 165893 538587
rect 166039 538581 166085 538587
rect 166130 538969 166170 539067
rect 166204 538969 166210 539545
rect 166130 538957 166210 538969
rect 166252 539545 166298 539557
rect 166252 538969 166258 539545
rect 166292 539537 166298 539545
rect 166292 539307 166410 539537
rect 166670 539337 166890 539347
rect 166670 539307 166690 539337
rect 166292 539297 166690 539307
rect 166292 539207 166570 539297
rect 166620 539207 166690 539297
rect 166292 539197 166690 539207
rect 166292 539074 166410 539197
rect 166670 539157 166690 539197
rect 166870 539157 166890 539337
rect 166670 539147 166890 539157
rect 166292 538969 166370 539074
rect 166252 538967 166370 538969
rect 166252 538957 166298 538967
rect 164752 538557 164798 538569
rect 164929 538517 164987 538523
rect 165121 538517 165179 538523
rect 165313 538517 165371 538523
rect 165505 538517 165563 538523
rect 165697 538517 165755 538523
rect 165889 538517 165947 538523
rect 166130 538517 166170 538957
rect 166200 538910 166260 538917
rect 166200 538876 166214 538910
rect 166248 538876 166260 538910
rect 166200 538857 166260 538876
rect 166364 538607 166370 538967
rect 164700 538510 164760 538517
rect 164700 538476 164714 538510
rect 164748 538476 164760 538510
rect 164700 538457 164760 538476
rect 164920 538483 164941 538517
rect 164975 538483 165133 538517
rect 165167 538483 165325 538517
rect 165359 538483 165517 538517
rect 165551 538483 165709 538517
rect 165743 538483 165901 538517
rect 165935 538483 166170 538517
rect 164920 538457 166170 538483
rect 166360 538586 166370 538607
rect 166404 538607 166410 539074
rect 166452 539074 166498 539086
rect 166452 538607 166458 539074
rect 166404 538586 166458 538607
rect 166492 538586 166498 539074
rect 166360 538574 166498 538586
rect 166360 538510 166480 538574
rect 166360 538477 166414 538510
rect 166400 538476 166414 538477
rect 166448 538477 166480 538510
rect 166448 538476 166460 538477
rect 166400 538457 166460 538476
rect 166560 537975 167305 537977
rect 164280 537847 164334 537963
rect 162090 537744 162150 537757
rect 162088 537738 162150 537744
rect 162088 537704 162100 537738
rect 162134 537704 162150 537738
rect 162088 537698 162150 537704
rect 162090 537697 162150 537698
rect 162310 537738 162370 537757
rect 162310 537704 162324 537738
rect 162358 537704 162370 537738
rect 162310 537697 162370 537704
rect 161550 537628 161788 537640
rect 161254 537374 161300 537386
rect 161254 537257 161260 537374
rect 161250 537107 161260 537257
rect 161254 537086 161260 537107
rect 161294 537257 161300 537374
rect 161342 537374 161388 537386
rect 161342 537257 161348 537374
rect 161294 537086 161348 537257
rect 161382 537257 161388 537374
rect 161454 537374 161500 537386
rect 161454 537257 161460 537374
rect 161382 537107 161460 537257
rect 161382 537086 161388 537107
rect 161254 537074 161388 537086
rect 161454 537086 161460 537107
rect 161494 537257 161500 537374
rect 161550 537340 161556 537628
rect 161590 537497 161748 537628
rect 161590 537340 161596 537497
rect 161550 537328 161596 537340
rect 161646 537374 161692 537386
rect 161646 537257 161652 537374
rect 161494 537097 161652 537257
rect 161494 537086 161500 537097
rect 161454 537074 161500 537086
rect 161646 537086 161652 537097
rect 161686 537257 161692 537374
rect 161742 537340 161748 537497
rect 161782 537340 161788 537628
rect 161742 537328 161788 537340
rect 161854 537637 161900 537640
rect 162010 537637 162092 537640
rect 161854 537628 162092 537637
rect 161854 537340 161860 537628
rect 161894 537497 162052 537628
rect 161894 537340 161900 537497
rect 161854 537328 161900 537340
rect 161950 537374 161996 537386
rect 161950 537257 161956 537374
rect 161686 537097 161956 537257
rect 161686 537086 161692 537097
rect 161646 537074 161692 537086
rect 161280 537010 161360 537074
rect 154000 536997 156802 537000
rect 154000 536987 157000 536997
rect 154000 536967 157400 536987
rect 161280 536977 161304 537010
rect 161290 536976 161304 536977
rect 161338 536977 161360 537010
rect 161590 537010 161650 537017
rect 161338 536976 161350 536977
rect 154000 536957 157525 536967
rect 161290 536957 161350 536976
rect 161590 536976 161604 537010
rect 161638 536976 161650 537010
rect 161590 536957 161650 536976
rect 154000 536877 157420 536957
rect 157510 536877 157525 536957
rect 154000 536857 157525 536877
rect 161770 536937 161870 537097
rect 161950 537086 161956 537097
rect 161990 537257 161996 537374
rect 162046 537340 162052 537497
rect 162086 537340 162092 537628
rect 164328 537566 164334 537847
rect 164372 537847 164480 537963
rect 164646 537967 164696 537975
rect 164964 537967 165014 537975
rect 164646 537963 165014 537967
rect 164372 537566 164378 537847
rect 164328 537554 164378 537566
rect 164646 537566 164652 537963
rect 164690 537567 164970 537963
rect 164690 537566 164696 537567
rect 164646 537554 164696 537566
rect 164964 537566 164970 537567
rect 165008 537566 165014 537963
rect 164964 537554 165014 537566
rect 165282 537963 165332 537975
rect 165282 537566 165288 537963
rect 165326 537957 165332 537963
rect 165600 537963 165650 537975
rect 165600 537957 165606 537963
rect 165326 537597 165606 537957
rect 165326 537566 165332 537597
rect 165282 537554 165332 537566
rect 165600 537566 165606 537597
rect 165644 537566 165650 537963
rect 165600 537554 165650 537566
rect 165918 537963 165968 537975
rect 165918 537566 165924 537963
rect 165962 537957 165968 537963
rect 166236 537963 166286 537975
rect 166236 537957 166242 537963
rect 165962 537597 166242 537957
rect 165962 537566 165968 537597
rect 165918 537554 165968 537566
rect 166236 537566 166242 537597
rect 166280 537566 166286 537963
rect 166236 537554 166286 537566
rect 166554 537963 167305 537975
rect 166554 537566 166560 537963
rect 166598 537566 167305 537963
rect 166554 537554 167305 537566
rect 166560 537547 167305 537554
rect 162046 537328 162092 537340
rect 162142 537374 162188 537386
rect 162142 537257 162148 537374
rect 161990 537097 162148 537257
rect 161990 537086 161996 537097
rect 161950 537074 161996 537086
rect 162142 537086 162148 537097
rect 162182 537237 162188 537374
rect 162274 537374 162320 537386
rect 162274 537237 162280 537374
rect 162182 537117 162280 537237
rect 162182 537086 162188 537117
rect 162142 537074 162188 537086
rect 162274 537086 162280 537117
rect 162314 537127 162320 537374
rect 162362 537374 162408 537386
rect 162362 537127 162368 537374
rect 162314 537086 162368 537127
rect 162402 537127 162408 537374
rect 163020 537167 163730 537227
rect 162402 537086 162410 537127
rect 162274 537074 162410 537086
rect 161770 536857 161790 536937
rect 161850 536857 161870 536937
rect 154000 536800 157400 536857
rect 161770 536837 161870 536857
rect 161990 537010 162050 537017
rect 161990 536976 162004 537010
rect 162038 537007 162050 537010
rect 162280 537010 162410 537074
rect 162038 536976 162060 537007
rect 161990 536917 162060 536976
rect 162280 536976 162324 537010
rect 162358 536976 162410 537010
rect 162280 536967 162410 536976
rect 162910 537097 163730 537167
rect 162310 536957 162370 536967
rect 162910 536917 162960 537097
rect 163020 537027 163730 537097
rect 161990 536847 162960 536917
rect 156614 536798 157400 536800
rect 156800 536797 157400 536798
rect 157200 536787 157400 536797
rect 162300 536757 162720 536817
rect 162300 536737 162360 536757
rect 157800 536718 157992 536724
rect 157800 536684 157812 536718
rect 157980 536684 157992 536718
rect 157800 536678 157992 536684
rect 158150 536718 162360 536737
rect 162660 536737 162720 536757
rect 163030 536737 163230 536797
rect 158150 536684 158190 536718
rect 158358 536684 158448 536718
rect 158616 536684 158706 536718
rect 158874 536684 158964 536718
rect 159132 536684 159222 536718
rect 159390 536684 159480 536718
rect 159648 536684 159738 536718
rect 159906 536684 159996 536718
rect 160164 536684 160254 536718
rect 160422 536684 160512 536718
rect 160680 536684 160896 536718
rect 161064 536684 161154 536718
rect 161322 536684 161412 536718
rect 161580 536684 161794 536718
rect 161962 536684 162052 536718
rect 162220 536684 162360 536718
rect 158150 536677 162360 536684
rect 162420 536718 162612 536724
rect 162420 536684 162432 536718
rect 162600 536684 162612 536718
rect 162420 536678 162612 536684
rect 162660 536677 163230 536737
rect 157744 536625 157790 536637
rect 157744 536157 157750 536625
rect 157740 536049 157750 536157
rect 157784 536157 157790 536625
rect 158002 536625 158048 536637
rect 158002 536157 158008 536625
rect 157784 536049 158008 536157
rect 158042 536157 158048 536625
rect 161990 536620 162030 536677
rect 158380 536608 158426 536620
rect 158122 536354 158168 536366
rect 158042 536049 158050 536157
rect 158122 536066 158128 536354
rect 158162 536177 158168 536354
rect 158380 536320 158386 536608
rect 158420 536597 158426 536608
rect 158896 536608 158942 536620
rect 158896 536597 158902 536608
rect 158420 536587 158902 536597
rect 158420 536487 158480 536587
rect 158420 536320 158426 536487
rect 158470 536427 158480 536487
rect 158580 536487 158902 536587
rect 158580 536427 158600 536487
rect 158470 536407 158600 536427
rect 158380 536308 158426 536320
rect 158638 536354 158684 536366
rect 158638 536177 158644 536354
rect 158162 536077 158644 536177
rect 158162 536066 158168 536077
rect 158122 536054 158168 536066
rect 158638 536066 158644 536077
rect 158678 536177 158684 536354
rect 158896 536320 158902 536487
rect 158936 536597 158942 536608
rect 159412 536608 159458 536620
rect 159412 536597 159418 536608
rect 158936 536487 159418 536597
rect 158936 536320 158942 536487
rect 158896 536308 158942 536320
rect 159154 536354 159200 536366
rect 159154 536177 159160 536354
rect 158678 536077 159160 536177
rect 158678 536066 158684 536077
rect 158638 536054 158684 536066
rect 159154 536066 159160 536077
rect 159194 536177 159200 536354
rect 159412 536320 159418 536487
rect 159452 536597 159458 536608
rect 159928 536608 159974 536620
rect 159928 536597 159934 536608
rect 159452 536487 159934 536597
rect 159452 536320 159458 536487
rect 159412 536308 159458 536320
rect 159670 536354 159716 536366
rect 159670 536177 159676 536354
rect 159194 536077 159676 536177
rect 159194 536066 159200 536077
rect 159154 536054 159200 536066
rect 159670 536066 159676 536077
rect 159710 536177 159716 536354
rect 159928 536320 159934 536487
rect 159968 536597 159974 536608
rect 160444 536608 160490 536620
rect 160444 536597 160450 536608
rect 159968 536487 160450 536597
rect 159968 536320 159974 536487
rect 159928 536308 159974 536320
rect 160186 536354 160232 536366
rect 160186 536177 160192 536354
rect 159710 536077 160192 536177
rect 159710 536066 159716 536077
rect 159670 536054 159716 536066
rect 160186 536066 160192 536077
rect 160226 536177 160232 536354
rect 160444 536320 160450 536487
rect 160484 536597 160490 536608
rect 160828 536617 160874 536620
rect 161344 536617 161390 536620
rect 160828 536608 161390 536617
rect 160484 536487 160510 536597
rect 160484 536320 160490 536487
rect 160444 536308 160490 536320
rect 160702 536354 160748 536366
rect 160702 536177 160708 536354
rect 160226 536077 160708 536177
rect 160226 536066 160232 536077
rect 160186 536054 160232 536066
rect 160702 536066 160708 536077
rect 160742 536177 160748 536354
rect 160828 536320 160834 536608
rect 160868 536577 161350 536608
rect 160868 536497 161090 536577
rect 161170 536497 161350 536577
rect 160868 536457 161350 536497
rect 160868 536320 160874 536457
rect 160828 536308 160874 536320
rect 161086 536354 161132 536366
rect 161086 536197 161092 536354
rect 160742 536066 160770 536177
rect 161070 536077 161092 536197
rect 160702 536054 160770 536066
rect 161086 536066 161092 536077
rect 161126 536197 161132 536354
rect 161344 536320 161350 536457
rect 161384 536320 161390 536608
rect 161984 536608 162030 536620
rect 161344 536308 161390 536320
rect 161602 536354 161648 536366
rect 161602 536197 161608 536354
rect 161126 536077 161608 536197
rect 161126 536066 161132 536077
rect 161086 536054 161132 536066
rect 161602 536066 161608 536077
rect 161642 536197 161648 536354
rect 161726 536354 161772 536366
rect 161642 536066 161670 536197
rect 161602 536054 161670 536066
rect 161726 536066 161732 536354
rect 161766 536217 161772 536354
rect 161984 536320 161990 536608
rect 162024 536320 162030 536608
rect 162364 536625 162410 536637
rect 161984 536308 162030 536320
rect 162242 536354 162288 536366
rect 162242 536217 162248 536354
rect 161766 536097 162248 536217
rect 161766 536066 161772 536097
rect 161726 536054 161772 536066
rect 162242 536066 162248 536097
rect 162282 536217 162288 536354
rect 162282 536066 162310 536217
rect 162242 536054 162310 536066
rect 157740 535990 158050 536049
rect 157740 535956 157812 535990
rect 157980 535956 158050 535990
rect 157740 535837 158050 535956
rect 158178 535990 158370 535996
rect 158178 535956 158190 535990
rect 158358 535956 158370 535990
rect 158178 535950 158370 535956
rect 158436 535990 158628 535996
rect 158436 535956 158448 535990
rect 158616 535956 158628 535990
rect 158436 535950 158628 535956
rect 158694 535990 158886 535996
rect 158694 535956 158706 535990
rect 158874 535956 158886 535990
rect 158694 535950 158886 535956
rect 158952 535990 159144 535996
rect 158952 535956 158964 535990
rect 159132 535956 159144 535990
rect 158952 535950 159144 535956
rect 159210 535990 159402 535996
rect 159210 535956 159222 535990
rect 159390 535956 159402 535990
rect 159210 535950 159402 535956
rect 159468 535990 159660 535996
rect 159468 535956 159480 535990
rect 159648 535956 159660 535990
rect 159468 535950 159660 535956
rect 159726 535990 159918 535996
rect 159726 535956 159738 535990
rect 159906 535956 159918 535990
rect 159726 535950 159918 535956
rect 159984 535990 160176 535996
rect 159984 535956 159996 535990
rect 160164 535956 160176 535990
rect 159984 535950 160176 535956
rect 160242 535990 160434 535996
rect 160242 535956 160254 535990
rect 160422 535956 160434 535990
rect 160242 535950 160434 535956
rect 160500 535990 160692 535996
rect 160500 535956 160512 535990
rect 160680 535956 160692 535990
rect 160500 535950 160692 535956
rect 160730 535837 160770 536054
rect 160884 535990 161076 535996
rect 160884 535956 160896 535990
rect 161064 535956 161076 535990
rect 160884 535950 161076 535956
rect 161142 535990 161334 535996
rect 161142 535956 161154 535990
rect 161322 535956 161334 535990
rect 161142 535950 161334 535956
rect 161400 535990 161592 535996
rect 161400 535956 161412 535990
rect 161580 535956 161592 535990
rect 161400 535950 161592 535956
rect 161630 535837 161670 536054
rect 161782 535990 161974 535996
rect 161782 535956 161794 535990
rect 161962 535956 161974 535990
rect 161782 535950 161974 535956
rect 162040 535990 162232 535996
rect 162040 535956 162052 535990
rect 162220 535956 162232 535990
rect 162040 535950 162232 535956
rect 162270 535837 162310 536054
rect 162364 536049 162370 536625
rect 162404 536117 162410 536625
rect 162622 536625 162668 536637
rect 162622 536117 162628 536625
rect 162404 536049 162628 536117
rect 162662 536117 162668 536625
rect 162662 536049 162670 536117
rect 162364 536037 162670 536049
rect 162380 535990 162670 536037
rect 162380 535956 162432 535990
rect 162600 535956 162670 535990
rect 162380 535837 162670 535956
rect 157740 535797 162710 535837
rect 157750 535777 162710 535797
rect 157750 535737 162050 535777
rect 162650 535737 162710 535777
rect 157750 535717 162710 535737
rect 160210 535617 160330 535717
rect 160180 535607 160380 535617
rect 160180 535467 160200 535607
rect 160350 535467 160380 535607
rect 160180 535247 160380 535467
rect 163030 533000 163230 536677
rect 163530 536307 163730 537027
rect 164328 536448 164378 536460
rect 163530 536267 164100 536307
rect 163530 535937 163840 536267
rect 164050 535937 164100 536267
rect 164328 536051 164334 536448
rect 164372 536447 164378 536448
rect 164646 536448 164696 536460
rect 164646 536447 164652 536448
rect 164372 536051 164652 536447
rect 164690 536051 164696 536448
rect 164328 536047 164696 536051
rect 164328 536039 164378 536047
rect 164646 536039 164696 536047
rect 164964 536448 165014 536460
rect 164964 536051 164970 536448
rect 165008 536447 165014 536448
rect 165282 536448 165332 536460
rect 165282 536447 165288 536448
rect 165008 536051 165288 536447
rect 165326 536051 165332 536448
rect 164964 536047 165332 536051
rect 164964 536039 165014 536047
rect 165282 536039 165332 536047
rect 165600 536448 165650 536460
rect 165600 536051 165606 536448
rect 165644 536447 165650 536448
rect 165918 536448 165968 536460
rect 165918 536447 165924 536448
rect 165644 536087 165924 536447
rect 165644 536051 165650 536087
rect 165600 536039 165650 536051
rect 165918 536051 165924 536087
rect 165962 536051 165968 536448
rect 165918 536039 165968 536051
rect 166236 536448 166286 536460
rect 166236 536051 166242 536448
rect 166280 536427 166286 536448
rect 166554 536448 166604 536460
rect 166554 536427 166560 536448
rect 166280 536067 166560 536427
rect 166280 536051 166286 536067
rect 166236 536039 166286 536051
rect 166554 536051 166560 536067
rect 166598 536051 166604 536448
rect 166554 536039 166604 536051
rect 166875 536297 167305 537547
rect 166875 536077 166930 536297
rect 167260 536077 167305 536297
rect 166875 536012 167305 536077
rect 163530 535917 164100 535937
rect 163530 535667 163800 535917
rect 163530 535623 164380 535667
rect 163530 535267 164304 535623
rect 163530 535257 163800 535267
rect 164298 535226 164304 535267
rect 164342 535267 164380 535623
rect 164616 535627 164666 535635
rect 164934 535627 164984 535635
rect 164616 535623 164984 535627
rect 164342 535226 164348 535267
rect 164298 535214 164348 535226
rect 164616 535226 164622 535623
rect 164660 535257 164940 535623
rect 164660 535226 164666 535257
rect 164616 535214 164666 535226
rect 164934 535226 164940 535257
rect 164978 535226 164984 535623
rect 164934 535214 164984 535226
rect 165252 535627 165302 535635
rect 165570 535627 165620 535635
rect 165252 535623 165620 535627
rect 165252 535226 165258 535623
rect 165296 535257 165576 535623
rect 165296 535226 165302 535257
rect 165252 535214 165302 535226
rect 165570 535226 165576 535257
rect 165614 535226 165620 535623
rect 165570 535214 165620 535226
rect 165888 535623 165938 535635
rect 165888 535226 165894 535623
rect 165932 535607 165938 535623
rect 166206 535623 166256 535635
rect 166206 535607 166212 535623
rect 165932 535237 166212 535607
rect 165932 535226 165938 535237
rect 165888 535214 165938 535226
rect 166206 535226 166212 535237
rect 166250 535226 166256 535623
rect 166500 535623 167265 535647
rect 166500 535237 166530 535623
rect 166206 535214 166256 535226
rect 166524 535226 166530 535237
rect 166568 535587 167265 535623
rect 166568 535457 166720 535587
rect 166850 535577 167265 535587
rect 166850 535457 166900 535577
rect 166568 535447 166900 535457
rect 167030 535557 167265 535577
rect 167030 535447 167080 535557
rect 166568 535427 167080 535447
rect 167210 535427 167265 535557
rect 166568 535397 167265 535427
rect 166568 535267 166700 535397
rect 166830 535387 167265 535397
rect 166830 535267 166890 535387
rect 166568 535257 166890 535267
rect 167020 535377 167265 535387
rect 167020 535257 167090 535377
rect 166568 535247 167090 535257
rect 167220 535247 167265 535377
rect 166568 535237 167265 535247
rect 166568 535226 166574 535237
rect 166524 535214 166574 535226
rect 164298 534108 164348 534120
rect 164298 533711 164304 534108
rect 164342 534097 164348 534108
rect 164616 534108 164666 534120
rect 164616 534097 164622 534108
rect 164342 533727 164622 534097
rect 164342 533711 164348 533727
rect 164298 533699 164348 533711
rect 164616 533711 164622 533727
rect 164660 534097 164666 534108
rect 164934 534108 164984 534120
rect 164660 533727 164670 534097
rect 164660 533711 164666 533727
rect 164616 533699 164666 533711
rect 164934 533711 164940 534108
rect 164978 534097 164984 534108
rect 165252 534108 165302 534120
rect 165252 534097 165258 534108
rect 164978 533727 165258 534097
rect 164978 533711 164984 533727
rect 164934 533699 164984 533711
rect 165252 533711 165258 533727
rect 165296 533711 165302 534108
rect 165252 533699 165302 533711
rect 165570 534108 165620 534120
rect 165570 533711 165576 534108
rect 165614 534097 165620 534108
rect 165888 534108 165938 534120
rect 165888 534097 165894 534108
rect 165614 533727 165894 534097
rect 165614 533711 165620 533727
rect 165570 533699 165620 533711
rect 165888 533711 165894 533727
rect 165932 533711 165938 534108
rect 165888 533699 165938 533711
rect 166206 534108 166256 534120
rect 166206 533711 166212 534108
rect 166250 534087 166256 534108
rect 166524 534108 166574 534120
rect 166524 534087 166530 534108
rect 166250 533717 166530 534087
rect 166250 533711 166256 533717
rect 166206 533699 166256 533711
rect 166524 533711 166530 533717
rect 166568 533711 166574 534108
rect 166524 533699 166574 533711
rect 9000 531000 163230 533000
rect 167520 532787 167720 540727
rect 168480 540562 168486 540917
rect 168520 540917 168574 541050
rect 168520 540562 168526 540917
rect 168480 540550 168526 540562
rect 168568 540562 168574 540917
rect 168608 540997 168620 541050
rect 168779 541057 168825 541069
rect 168971 541057 169017 541069
rect 169163 541057 169209 541069
rect 169355 541057 169401 541069
rect 169547 541057 169593 541069
rect 169739 541057 169785 541069
rect 168779 540997 168785 541057
rect 168608 540917 168785 540997
rect 168608 540562 168614 540917
rect 168568 540550 168614 540562
rect 168683 540603 168729 540615
rect 168683 540317 168689 540603
rect 168650 540115 168689 540317
rect 168723 540317 168729 540603
rect 168779 540569 168785 540917
rect 168819 540667 168977 541057
rect 168819 540569 168825 540667
rect 168779 540557 168825 540569
rect 168875 540603 168921 540615
rect 168875 540317 168881 540603
rect 168723 540115 168881 540317
rect 168915 540317 168921 540603
rect 168971 540569 168977 540667
rect 169011 540667 169169 541057
rect 169011 540569 169017 540667
rect 168971 540557 169017 540569
rect 169067 540603 169113 540615
rect 169067 540317 169073 540603
rect 168915 540115 169073 540317
rect 169107 540317 169113 540603
rect 169163 540569 169169 540667
rect 169203 540667 169361 541057
rect 169203 540569 169209 540667
rect 169163 540557 169209 540569
rect 169259 540603 169305 540615
rect 169259 540317 169265 540603
rect 169107 540115 169265 540317
rect 169299 540317 169305 540603
rect 169355 540569 169361 540667
rect 169395 540667 169553 541057
rect 169395 540569 169401 540667
rect 169355 540557 169401 540569
rect 169451 540603 169497 540615
rect 169451 540317 169457 540603
rect 169299 540115 169457 540317
rect 169491 540317 169497 540603
rect 169547 540569 169553 540667
rect 169587 541027 169745 541057
rect 169779 541027 169810 541057
rect 169587 540927 169690 541027
rect 169800 540927 169810 541027
rect 169587 540907 169745 540927
rect 169779 540907 169810 540927
rect 169587 540807 169690 540907
rect 169800 540807 169810 540907
rect 170005 540862 170055 541112
rect 170198 541151 170260 541157
rect 170198 541117 170210 541151
rect 170244 541117 170260 541151
rect 170198 541111 170260 541117
rect 170200 541097 170260 541111
rect 171780 540997 171980 541537
rect 172220 541157 172280 541167
rect 172520 541162 173540 541187
rect 172520 541158 173755 541162
rect 172180 541151 172320 541157
rect 172180 541117 172230 541151
rect 172264 541117 172320 541151
rect 172520 541127 172533 541158
rect 172521 541124 172533 541127
rect 172567 541127 172725 541158
rect 172567 541124 172579 541127
rect 172521 541118 172579 541124
rect 172713 541124 172725 541127
rect 172759 541127 172917 541158
rect 172759 541124 172771 541127
rect 172713 541118 172771 541124
rect 172905 541124 172917 541127
rect 172951 541127 173109 541158
rect 172951 541124 172963 541127
rect 172905 541118 172963 541124
rect 173097 541124 173109 541127
rect 173143 541127 173301 541158
rect 173143 541124 173155 541127
rect 173097 541118 173155 541124
rect 173289 541124 173301 541127
rect 173335 541127 173493 541158
rect 173335 541124 173347 541127
rect 173289 541118 173347 541124
rect 173481 541124 173493 541127
rect 173527 541124 173755 541158
rect 173481 541118 173755 541124
rect 172180 541050 172320 541117
rect 173525 541112 173755 541118
rect 172180 540997 172186 541050
rect 170480 540862 171250 540927
rect 171780 540917 172186 540997
rect 171780 540867 171980 540917
rect 169587 540787 169745 540807
rect 169779 540787 169810 540807
rect 169587 540687 169690 540787
rect 169800 540687 169810 540787
rect 169587 540667 169745 540687
rect 169587 540569 169593 540667
rect 169547 540557 169593 540569
rect 169643 540603 169689 540615
rect 169643 540317 169649 540603
rect 169491 540115 169649 540317
rect 169683 540317 169689 540603
rect 169739 540569 169745 540667
rect 169779 540667 169810 540687
rect 170000 540812 171250 540862
rect 169779 540569 169785 540667
rect 169739 540557 169785 540569
rect 169835 540603 169881 540615
rect 169835 540317 169841 540603
rect 169683 540115 169841 540317
rect 169875 540115 169881 540603
rect 170000 540367 170050 540812
rect 170480 540727 171250 540812
rect 170160 540596 170206 540608
rect 170000 540357 170060 540367
rect 169998 540351 170060 540357
rect 169998 540317 170010 540351
rect 170044 540317 170060 540351
rect 169998 540311 170060 540317
rect 170000 540307 170060 540311
rect 169960 540267 170006 540279
rect 169960 540187 169966 540267
rect 168650 540107 169881 540115
rect 168650 540103 168729 540107
rect 168875 540103 168921 540107
rect 169067 540103 169113 540107
rect 169259 540103 169305 540107
rect 169451 540103 169497 540107
rect 169643 540103 169689 540107
rect 169835 540103 169881 540107
rect 168650 540097 168720 540103
rect 168510 540041 168580 540057
rect 168510 540007 168530 540041
rect 168564 540007 168580 540041
rect 168510 539987 168580 540007
rect 168650 539787 168680 540097
rect 169940 540091 169966 540187
rect 170000 540091 170006 540267
rect 169940 540079 170006 540091
rect 170048 540267 170094 540279
rect 170048 540091 170054 540267
rect 170088 540257 170094 540267
rect 170160 540257 170166 540596
rect 170088 540108 170166 540257
rect 170200 540267 170206 540596
rect 170248 540596 170294 540608
rect 170248 540267 170254 540596
rect 170200 540108 170254 540267
rect 170288 540267 170294 540596
rect 170470 540277 170690 540287
rect 170288 540257 170310 540267
rect 170470 540257 170490 540277
rect 170288 540247 170490 540257
rect 170288 540117 170370 540247
rect 170430 540117 170490 540247
rect 170288 540108 170490 540117
rect 170088 540107 170490 540108
rect 170088 540091 170094 540107
rect 170160 540096 170294 540107
rect 170470 540097 170490 540107
rect 170670 540097 170690 540277
rect 170048 540079 170094 540091
rect 168725 540048 168783 540054
rect 168725 540047 168737 540048
rect 168720 540014 168737 540047
rect 168771 540047 168783 540048
rect 168917 540048 168975 540054
rect 168917 540047 168929 540048
rect 168771 540014 168929 540047
rect 168963 540047 168975 540048
rect 169109 540048 169167 540054
rect 169109 540047 169121 540048
rect 168963 540014 169121 540047
rect 169155 540047 169167 540048
rect 169301 540048 169359 540054
rect 169301 540047 169313 540048
rect 169155 540014 169313 540047
rect 169347 540047 169359 540048
rect 169493 540048 169551 540054
rect 169493 540047 169505 540048
rect 169347 540014 169505 540047
rect 169539 540047 169551 540048
rect 169685 540048 169743 540054
rect 169685 540047 169697 540048
rect 169539 540014 169697 540047
rect 169731 540014 169743 540048
rect 168720 540008 169743 540014
rect 168720 539987 169740 540008
rect 168080 539687 168680 539787
rect 168080 537963 168280 539687
rect 168440 539638 168680 539687
rect 168440 539604 168514 539638
rect 168548 539604 168680 539638
rect 168440 539545 168680 539604
rect 168820 539651 169830 539657
rect 168820 539645 169843 539651
rect 168820 539611 168837 539645
rect 168871 539611 169029 539645
rect 169063 539611 169221 539645
rect 169255 539611 169413 539645
rect 169447 539611 169605 539645
rect 169639 539611 169797 539645
rect 169831 539611 169843 539645
rect 168820 539605 169843 539611
rect 168820 539597 169830 539605
rect 169940 539557 169970 540079
rect 169998 540041 170060 540047
rect 169998 540007 170010 540041
rect 170044 540007 170060 540041
rect 169998 540001 170060 540007
rect 170000 539638 170060 540001
rect 170170 540041 170290 540096
rect 170470 540087 170690 540097
rect 170170 540007 170210 540041
rect 170244 540007 170290 540041
rect 170170 539987 170290 540007
rect 170000 539604 170014 539638
rect 170048 539604 170060 539638
rect 170000 539597 170060 539604
rect 170200 539638 170280 539657
rect 170200 539604 170214 539638
rect 170248 539604 170280 539638
rect 170200 539597 170280 539604
rect 168440 539447 168470 539545
rect 168464 538569 168470 539447
rect 168504 539447 168558 539545
rect 168504 538569 168510 539447
rect 168464 538557 168510 538569
rect 168552 538569 168558 539447
rect 168592 539527 168680 539545
rect 168783 539535 168829 539547
rect 168592 539517 168750 539527
rect 168783 539517 168789 539535
rect 168592 539447 168789 539517
rect 168592 538569 168598 539447
rect 168650 539237 168789 539447
rect 168687 539081 168733 539093
rect 168687 538593 168693 539081
rect 168727 538967 168733 539081
rect 168783 539047 168789 539237
rect 168823 539517 168829 539535
rect 168975 539535 169021 539547
rect 168975 539517 168981 539535
rect 168823 539237 168981 539517
rect 168823 539047 168829 539237
rect 168783 539035 168829 539047
rect 168879 539081 168925 539093
rect 168879 538967 168885 539081
rect 168727 538593 168885 538967
rect 168919 538967 168925 539081
rect 168975 539047 168981 539237
rect 169015 539517 169021 539535
rect 169167 539535 169213 539547
rect 169167 539517 169173 539535
rect 169015 539237 169173 539517
rect 169015 539047 169021 539237
rect 168975 539035 169021 539047
rect 169071 539081 169117 539093
rect 169071 538967 169077 539081
rect 168919 538593 169077 538967
rect 169111 538967 169117 539081
rect 169167 539047 169173 539237
rect 169207 539517 169213 539535
rect 169359 539535 169405 539547
rect 169359 539517 169365 539535
rect 169207 539237 169365 539517
rect 169207 539047 169213 539237
rect 169167 539035 169213 539047
rect 169263 539081 169309 539093
rect 169263 538967 169269 539081
rect 169111 538593 169269 538967
rect 169303 538967 169309 539081
rect 169359 539047 169365 539237
rect 169399 539517 169405 539535
rect 169551 539535 169597 539547
rect 169551 539517 169557 539535
rect 169399 539237 169557 539517
rect 169399 539047 169405 539237
rect 169359 539035 169405 539047
rect 169455 539081 169501 539093
rect 169455 538967 169461 539081
rect 169303 538593 169461 538967
rect 169495 538967 169501 539081
rect 169551 539047 169557 539237
rect 169591 539517 169597 539535
rect 169743 539535 169789 539547
rect 169743 539517 169749 539535
rect 169591 539237 169749 539517
rect 169591 539047 169597 539237
rect 169551 539035 169597 539047
rect 169647 539081 169693 539093
rect 169647 538967 169653 539081
rect 169495 538593 169653 538967
rect 169687 538967 169693 539081
rect 169743 539047 169749 539237
rect 169783 539517 169789 539535
rect 169940 539545 170010 539557
rect 169783 539237 169800 539517
rect 169940 539407 169970 539545
rect 169783 539047 169789 539237
rect 169743 539035 169789 539047
rect 169839 539081 169885 539093
rect 169839 538967 169845 539081
rect 169687 538837 169845 538967
rect 169687 538737 169700 538837
rect 169840 538737 169845 538837
rect 169687 538593 169845 538737
rect 169879 538593 169885 539081
rect 169964 539067 169970 539407
rect 168687 538587 169885 538593
rect 168687 538581 168733 538587
rect 168879 538581 168925 538587
rect 169071 538581 169117 538587
rect 169263 538581 169309 538587
rect 169455 538581 169501 538587
rect 169647 538581 169693 538587
rect 169839 538581 169885 538587
rect 169930 538969 169970 539067
rect 170004 538969 170010 539545
rect 169930 538957 170010 538969
rect 170052 539545 170098 539557
rect 170052 538969 170058 539545
rect 170092 539537 170098 539545
rect 170092 539307 170210 539537
rect 170470 539337 170690 539347
rect 170470 539307 170490 539337
rect 170092 539297 170490 539307
rect 170092 539207 170370 539297
rect 170420 539207 170490 539297
rect 170092 539197 170490 539207
rect 170092 539074 170210 539197
rect 170470 539157 170490 539197
rect 170670 539157 170690 539337
rect 170470 539147 170690 539157
rect 170092 538969 170170 539074
rect 170052 538967 170170 538969
rect 170052 538957 170098 538967
rect 168552 538557 168598 538569
rect 168729 538517 168787 538523
rect 168921 538517 168979 538523
rect 169113 538517 169171 538523
rect 169305 538517 169363 538523
rect 169497 538517 169555 538523
rect 169689 538517 169747 538523
rect 169930 538517 169970 538957
rect 170000 538910 170060 538917
rect 170000 538876 170014 538910
rect 170048 538876 170060 538910
rect 170000 538857 170060 538876
rect 170164 538607 170170 538967
rect 168500 538510 168560 538517
rect 168500 538476 168514 538510
rect 168548 538476 168560 538510
rect 168500 538457 168560 538476
rect 168720 538483 168741 538517
rect 168775 538483 168933 538517
rect 168967 538483 169125 538517
rect 169159 538483 169317 538517
rect 169351 538483 169509 538517
rect 169543 538483 169701 538517
rect 169735 538483 169970 538517
rect 168720 538457 169970 538483
rect 170160 538586 170170 538607
rect 170204 538607 170210 539074
rect 170252 539074 170298 539086
rect 170252 538607 170258 539074
rect 170204 538586 170258 538607
rect 170292 538586 170298 539074
rect 170160 538574 170298 538586
rect 170160 538510 170280 538574
rect 170160 538477 170214 538510
rect 170200 538476 170214 538477
rect 170248 538477 170280 538510
rect 170248 538476 170260 538477
rect 170200 538457 170260 538476
rect 168440 537975 168770 537977
rect 169070 537975 169915 537977
rect 168080 537847 168106 537963
rect 168100 537566 168106 537847
rect 168144 537847 168280 537963
rect 168418 537963 168786 537975
rect 168144 537566 168150 537847
rect 168100 537554 168150 537566
rect 168418 537566 168424 537963
rect 168462 537617 168742 537963
rect 168462 537566 168468 537617
rect 168418 537554 168468 537566
rect 168736 537566 168742 537617
rect 168780 537566 168786 537963
rect 168736 537554 168786 537566
rect 169054 537963 169915 537975
rect 169054 537566 169060 537963
rect 169098 537567 169915 537963
rect 169098 537566 169104 537567
rect 169054 537554 169104 537566
rect 168100 536448 168150 536460
rect 168100 536051 168106 536448
rect 168144 536437 168150 536448
rect 168418 536448 168468 536460
rect 168418 536437 168424 536448
rect 168144 536077 168424 536437
rect 168144 536051 168150 536077
rect 168100 536039 168150 536051
rect 168418 536051 168424 536077
rect 168462 536051 168468 536448
rect 168418 536039 168468 536051
rect 168736 536457 168786 536460
rect 169054 536457 169104 536460
rect 168736 536448 169104 536457
rect 168736 536051 168742 536448
rect 168780 536097 169060 536448
rect 168780 536051 168786 536097
rect 168736 536039 168786 536051
rect 169054 536051 169060 536097
rect 169098 536051 169104 536448
rect 169054 536039 169104 536051
rect 169505 536287 169915 537567
rect 169505 536007 169570 536287
rect 169870 536007 169915 536287
rect 169505 535942 169915 536007
rect 171050 533537 171250 540727
rect 172180 540562 172186 540917
rect 172220 540917 172274 541050
rect 172220 540562 172226 540917
rect 172180 540550 172226 540562
rect 172268 540562 172274 540917
rect 172308 540997 172320 541050
rect 172479 541057 172525 541069
rect 172671 541057 172717 541069
rect 172863 541057 172909 541069
rect 173055 541057 173101 541069
rect 173247 541057 173293 541069
rect 173439 541057 173485 541069
rect 172479 540997 172485 541057
rect 172308 540917 172485 540997
rect 172308 540562 172314 540917
rect 172268 540550 172314 540562
rect 172383 540603 172429 540615
rect 172383 540317 172389 540603
rect 172350 540115 172389 540317
rect 172423 540317 172429 540603
rect 172479 540569 172485 540917
rect 172519 540667 172677 541057
rect 172519 540569 172525 540667
rect 172479 540557 172525 540569
rect 172575 540603 172621 540615
rect 172575 540317 172581 540603
rect 172423 540115 172581 540317
rect 172615 540317 172621 540603
rect 172671 540569 172677 540667
rect 172711 540667 172869 541057
rect 172711 540569 172717 540667
rect 172671 540557 172717 540569
rect 172767 540603 172813 540615
rect 172767 540317 172773 540603
rect 172615 540115 172773 540317
rect 172807 540317 172813 540603
rect 172863 540569 172869 540667
rect 172903 540667 173061 541057
rect 172903 540569 172909 540667
rect 172863 540557 172909 540569
rect 172959 540603 173005 540615
rect 172959 540317 172965 540603
rect 172807 540115 172965 540317
rect 172999 540317 173005 540603
rect 173055 540569 173061 540667
rect 173095 540667 173253 541057
rect 173095 540569 173101 540667
rect 173055 540557 173101 540569
rect 173151 540603 173197 540615
rect 173151 540317 173157 540603
rect 172999 540115 173157 540317
rect 173191 540317 173197 540603
rect 173247 540569 173253 540667
rect 173287 541027 173445 541057
rect 173479 541027 173510 541057
rect 173287 540927 173390 541027
rect 173500 540927 173510 541027
rect 173287 540907 173445 540927
rect 173479 540907 173510 540927
rect 173287 540807 173390 540907
rect 173500 540807 173510 540907
rect 173705 540862 173755 541112
rect 173898 541151 173960 541157
rect 173898 541117 173910 541151
rect 173944 541117 173960 541151
rect 173898 541111 173960 541117
rect 173900 541097 173960 541111
rect 175280 540997 175480 541537
rect 175720 541157 175780 541167
rect 176020 541162 177040 541187
rect 176020 541158 177255 541162
rect 175680 541151 175820 541157
rect 175680 541117 175730 541151
rect 175764 541117 175820 541151
rect 176020 541127 176033 541158
rect 176021 541124 176033 541127
rect 176067 541127 176225 541158
rect 176067 541124 176079 541127
rect 176021 541118 176079 541124
rect 176213 541124 176225 541127
rect 176259 541127 176417 541158
rect 176259 541124 176271 541127
rect 176213 541118 176271 541124
rect 176405 541124 176417 541127
rect 176451 541127 176609 541158
rect 176451 541124 176463 541127
rect 176405 541118 176463 541124
rect 176597 541124 176609 541127
rect 176643 541127 176801 541158
rect 176643 541124 176655 541127
rect 176597 541118 176655 541124
rect 176789 541124 176801 541127
rect 176835 541127 176993 541158
rect 176835 541124 176847 541127
rect 176789 541118 176847 541124
rect 176981 541124 176993 541127
rect 177027 541124 177255 541158
rect 176981 541118 177255 541124
rect 175680 541050 175820 541117
rect 177025 541112 177255 541118
rect 175680 540997 175686 541050
rect 174180 540862 174880 540927
rect 175280 540917 175686 540997
rect 175280 540867 175480 540917
rect 173287 540787 173445 540807
rect 173479 540787 173510 540807
rect 173287 540687 173390 540787
rect 173500 540687 173510 540787
rect 173287 540667 173445 540687
rect 173287 540569 173293 540667
rect 173247 540557 173293 540569
rect 173343 540603 173389 540615
rect 173343 540317 173349 540603
rect 173191 540115 173349 540317
rect 173383 540317 173389 540603
rect 173439 540569 173445 540667
rect 173479 540667 173510 540687
rect 173700 540812 174880 540862
rect 173479 540569 173485 540667
rect 173439 540557 173485 540569
rect 173535 540603 173581 540615
rect 173535 540317 173541 540603
rect 173383 540115 173541 540317
rect 173575 540115 173581 540603
rect 173700 540367 173750 540812
rect 174180 540727 174880 540812
rect 173860 540596 173906 540608
rect 173700 540357 173760 540367
rect 173698 540351 173760 540357
rect 173698 540317 173710 540351
rect 173744 540317 173760 540351
rect 173698 540311 173760 540317
rect 173700 540307 173760 540311
rect 173660 540267 173706 540279
rect 173660 540187 173666 540267
rect 172350 540107 173581 540115
rect 172350 540103 172429 540107
rect 172575 540103 172621 540107
rect 172767 540103 172813 540107
rect 172959 540103 173005 540107
rect 173151 540103 173197 540107
rect 173343 540103 173389 540107
rect 173535 540103 173581 540107
rect 172350 540097 172420 540103
rect 172210 540041 172280 540057
rect 172210 540007 172230 540041
rect 172264 540007 172280 540041
rect 172210 539987 172280 540007
rect 172350 539787 172380 540097
rect 173640 540091 173666 540187
rect 173700 540091 173706 540267
rect 173640 540079 173706 540091
rect 173748 540267 173794 540279
rect 173748 540091 173754 540267
rect 173788 540257 173794 540267
rect 173860 540257 173866 540596
rect 173788 540108 173866 540257
rect 173900 540267 173906 540596
rect 173948 540596 173994 540608
rect 173948 540267 173954 540596
rect 173900 540108 173954 540267
rect 173988 540267 173994 540596
rect 174180 540287 174380 540297
rect 173988 540257 174010 540267
rect 174170 540257 174190 540287
rect 173988 540247 174190 540257
rect 173988 540117 174070 540247
rect 174130 540117 174190 540247
rect 173988 540108 174190 540117
rect 173788 540107 174190 540108
rect 174370 540107 174390 540287
rect 173788 540091 173794 540107
rect 173860 540096 173994 540107
rect 173748 540079 173794 540091
rect 172425 540048 172483 540054
rect 172425 540047 172437 540048
rect 172420 540014 172437 540047
rect 172471 540047 172483 540048
rect 172617 540048 172675 540054
rect 172617 540047 172629 540048
rect 172471 540014 172629 540047
rect 172663 540047 172675 540048
rect 172809 540048 172867 540054
rect 172809 540047 172821 540048
rect 172663 540014 172821 540047
rect 172855 540047 172867 540048
rect 173001 540048 173059 540054
rect 173001 540047 173013 540048
rect 172855 540014 173013 540047
rect 173047 540047 173059 540048
rect 173193 540048 173251 540054
rect 173193 540047 173205 540048
rect 173047 540014 173205 540047
rect 173239 540047 173251 540048
rect 173385 540048 173443 540054
rect 173385 540047 173397 540048
rect 173239 540014 173397 540047
rect 173431 540014 173443 540048
rect 172420 540008 173443 540014
rect 172420 539987 173440 540008
rect 171780 539687 172380 539787
rect 171780 537963 171980 539687
rect 172140 539638 172380 539687
rect 172140 539604 172214 539638
rect 172248 539604 172380 539638
rect 172140 539545 172380 539604
rect 172520 539651 173530 539657
rect 172520 539645 173543 539651
rect 172520 539611 172537 539645
rect 172571 539611 172729 539645
rect 172763 539611 172921 539645
rect 172955 539611 173113 539645
rect 173147 539611 173305 539645
rect 173339 539611 173497 539645
rect 173531 539611 173543 539645
rect 172520 539605 173543 539611
rect 172520 539597 173530 539605
rect 173640 539557 173670 540079
rect 173698 540041 173760 540047
rect 173698 540007 173710 540041
rect 173744 540007 173760 540041
rect 173698 540001 173760 540007
rect 173700 539638 173760 540001
rect 173870 540041 173990 540096
rect 174170 540087 174390 540107
rect 173870 540007 173910 540041
rect 173944 540007 173990 540041
rect 173870 539987 173990 540007
rect 173700 539604 173714 539638
rect 173748 539604 173760 539638
rect 173700 539597 173760 539604
rect 173900 539638 173980 539657
rect 173900 539604 173914 539638
rect 173948 539604 173980 539638
rect 173900 539597 173980 539604
rect 172140 539447 172170 539545
rect 172164 538569 172170 539447
rect 172204 539447 172258 539545
rect 172204 538569 172210 539447
rect 172164 538557 172210 538569
rect 172252 538569 172258 539447
rect 172292 539527 172380 539545
rect 172483 539535 172529 539547
rect 172292 539517 172450 539527
rect 172483 539517 172489 539535
rect 172292 539447 172489 539517
rect 172292 538569 172298 539447
rect 172350 539237 172489 539447
rect 172387 539081 172433 539093
rect 172387 538593 172393 539081
rect 172427 538967 172433 539081
rect 172483 539047 172489 539237
rect 172523 539517 172529 539535
rect 172675 539535 172721 539547
rect 172675 539517 172681 539535
rect 172523 539237 172681 539517
rect 172523 539047 172529 539237
rect 172483 539035 172529 539047
rect 172579 539081 172625 539093
rect 172579 538967 172585 539081
rect 172427 538593 172585 538967
rect 172619 538967 172625 539081
rect 172675 539047 172681 539237
rect 172715 539517 172721 539535
rect 172867 539535 172913 539547
rect 172867 539517 172873 539535
rect 172715 539237 172873 539517
rect 172715 539047 172721 539237
rect 172675 539035 172721 539047
rect 172771 539081 172817 539093
rect 172771 538967 172777 539081
rect 172619 538593 172777 538967
rect 172811 538967 172817 539081
rect 172867 539047 172873 539237
rect 172907 539517 172913 539535
rect 173059 539535 173105 539547
rect 173059 539517 173065 539535
rect 172907 539237 173065 539517
rect 172907 539047 172913 539237
rect 172867 539035 172913 539047
rect 172963 539081 173009 539093
rect 172963 538967 172969 539081
rect 172811 538593 172969 538967
rect 173003 538967 173009 539081
rect 173059 539047 173065 539237
rect 173099 539517 173105 539535
rect 173251 539535 173297 539547
rect 173251 539517 173257 539535
rect 173099 539237 173257 539517
rect 173099 539047 173105 539237
rect 173059 539035 173105 539047
rect 173155 539081 173201 539093
rect 173155 538967 173161 539081
rect 173003 538593 173161 538967
rect 173195 538967 173201 539081
rect 173251 539047 173257 539237
rect 173291 539517 173297 539535
rect 173443 539535 173489 539547
rect 173443 539517 173449 539535
rect 173291 539237 173449 539517
rect 173291 539047 173297 539237
rect 173251 539035 173297 539047
rect 173347 539081 173393 539093
rect 173347 538967 173353 539081
rect 173195 538593 173353 538967
rect 173387 538967 173393 539081
rect 173443 539047 173449 539237
rect 173483 539517 173489 539535
rect 173640 539545 173710 539557
rect 173483 539237 173500 539517
rect 173640 539407 173670 539545
rect 173483 539047 173489 539237
rect 173443 539035 173489 539047
rect 173539 539081 173585 539093
rect 173539 538967 173545 539081
rect 173387 538837 173545 538967
rect 173387 538737 173400 538837
rect 173540 538737 173545 538837
rect 173387 538593 173545 538737
rect 173579 538593 173585 539081
rect 173664 539067 173670 539407
rect 172387 538587 173585 538593
rect 172387 538581 172433 538587
rect 172579 538581 172625 538587
rect 172771 538581 172817 538587
rect 172963 538581 173009 538587
rect 173155 538581 173201 538587
rect 173347 538581 173393 538587
rect 173539 538581 173585 538587
rect 173630 538969 173670 539067
rect 173704 538969 173710 539545
rect 173630 538957 173710 538969
rect 173752 539545 173798 539557
rect 173752 538969 173758 539545
rect 173792 539537 173798 539545
rect 173792 539307 173910 539537
rect 174170 539337 174390 539347
rect 174170 539307 174190 539337
rect 173792 539297 174190 539307
rect 173792 539207 174070 539297
rect 174120 539207 174190 539297
rect 173792 539197 174190 539207
rect 173792 539074 173910 539197
rect 174170 539157 174190 539197
rect 174370 539157 174390 539337
rect 174170 539147 174390 539157
rect 173792 538969 173870 539074
rect 173752 538967 173870 538969
rect 173752 538957 173798 538967
rect 172252 538557 172298 538569
rect 172429 538517 172487 538523
rect 172621 538517 172679 538523
rect 172813 538517 172871 538523
rect 173005 538517 173063 538523
rect 173197 538517 173255 538523
rect 173389 538517 173447 538523
rect 173630 538517 173670 538957
rect 173700 538910 173760 538917
rect 173700 538876 173714 538910
rect 173748 538876 173760 538910
rect 173700 538857 173760 538876
rect 173864 538607 173870 538967
rect 172200 538510 172260 538517
rect 172200 538476 172214 538510
rect 172248 538476 172260 538510
rect 172200 538457 172260 538476
rect 172420 538483 172441 538517
rect 172475 538483 172633 538517
rect 172667 538483 172825 538517
rect 172859 538483 173017 538517
rect 173051 538483 173209 538517
rect 173243 538483 173401 538517
rect 173435 538483 173670 538517
rect 172420 538457 173670 538483
rect 173860 538586 173870 538607
rect 173904 538607 173910 539074
rect 173952 539074 173998 539086
rect 173952 538607 173958 539074
rect 173904 538586 173958 538607
rect 173992 538586 173998 539074
rect 173860 538574 173998 538586
rect 173860 538510 173980 538574
rect 173860 538477 173914 538510
rect 173900 538476 173914 538477
rect 173948 538477 173980 538510
rect 173948 538476 173960 538477
rect 173900 538457 173960 538476
rect 171780 537847 171842 537963
rect 171836 537566 171842 537847
rect 171880 537847 171980 537963
rect 172154 537967 172204 537975
rect 172154 537963 172980 537967
rect 171880 537566 171886 537847
rect 171836 537554 171886 537566
rect 172154 537566 172160 537963
rect 172198 537566 172980 537963
rect 172154 537554 172980 537566
rect 172170 537547 172980 537554
rect 171836 536448 171886 536460
rect 171836 536051 171842 536448
rect 171880 536437 171886 536448
rect 172154 536448 172204 536460
rect 172154 536437 172160 536448
rect 171880 536077 172160 536437
rect 171880 536051 171886 536077
rect 171836 536039 171886 536051
rect 172154 536051 172160 536077
rect 172198 536051 172204 536448
rect 172154 536039 172204 536051
rect 172560 536297 172980 537547
rect 172560 536007 172610 536297
rect 172940 536007 172980 536297
rect 172560 535947 172980 536007
rect 174680 533537 174880 540727
rect 175680 540562 175686 540917
rect 175720 540917 175774 541050
rect 175720 540562 175726 540917
rect 175680 540550 175726 540562
rect 175768 540562 175774 540917
rect 175808 540997 175820 541050
rect 175979 541057 176025 541069
rect 176171 541057 176217 541069
rect 176363 541057 176409 541069
rect 176555 541057 176601 541069
rect 176747 541057 176793 541069
rect 176939 541057 176985 541069
rect 175979 540997 175985 541057
rect 175808 540917 175985 540997
rect 175808 540562 175814 540917
rect 175768 540550 175814 540562
rect 175883 540603 175929 540615
rect 175883 540317 175889 540603
rect 175850 540115 175889 540317
rect 175923 540317 175929 540603
rect 175979 540569 175985 540917
rect 176019 540667 176177 541057
rect 176019 540569 176025 540667
rect 175979 540557 176025 540569
rect 176075 540603 176121 540615
rect 176075 540317 176081 540603
rect 175923 540115 176081 540317
rect 176115 540317 176121 540603
rect 176171 540569 176177 540667
rect 176211 540667 176369 541057
rect 176211 540569 176217 540667
rect 176171 540557 176217 540569
rect 176267 540603 176313 540615
rect 176267 540317 176273 540603
rect 176115 540115 176273 540317
rect 176307 540317 176313 540603
rect 176363 540569 176369 540667
rect 176403 540667 176561 541057
rect 176403 540569 176409 540667
rect 176363 540557 176409 540569
rect 176459 540603 176505 540615
rect 176459 540317 176465 540603
rect 176307 540115 176465 540317
rect 176499 540317 176505 540603
rect 176555 540569 176561 540667
rect 176595 540667 176753 541057
rect 176595 540569 176601 540667
rect 176555 540557 176601 540569
rect 176651 540603 176697 540615
rect 176651 540317 176657 540603
rect 176499 540115 176657 540317
rect 176691 540317 176697 540603
rect 176747 540569 176753 540667
rect 176787 541027 176945 541057
rect 176979 541027 177010 541057
rect 176787 540927 176890 541027
rect 177000 540927 177010 541027
rect 176787 540907 176945 540927
rect 176979 540907 177010 540927
rect 176787 540807 176890 540907
rect 177000 540807 177010 540907
rect 177205 540862 177255 541112
rect 177398 541151 177460 541157
rect 177398 541117 177410 541151
rect 177444 541117 177460 541151
rect 177398 541111 177460 541117
rect 177400 541097 177460 541111
rect 178880 540997 179080 541537
rect 179320 541157 179380 541167
rect 179620 541162 180640 541187
rect 179620 541158 180855 541162
rect 179280 541151 179420 541157
rect 179280 541117 179330 541151
rect 179364 541117 179420 541151
rect 179620 541127 179633 541158
rect 179621 541124 179633 541127
rect 179667 541127 179825 541158
rect 179667 541124 179679 541127
rect 179621 541118 179679 541124
rect 179813 541124 179825 541127
rect 179859 541127 180017 541158
rect 179859 541124 179871 541127
rect 179813 541118 179871 541124
rect 180005 541124 180017 541127
rect 180051 541127 180209 541158
rect 180051 541124 180063 541127
rect 180005 541118 180063 541124
rect 180197 541124 180209 541127
rect 180243 541127 180401 541158
rect 180243 541124 180255 541127
rect 180197 541118 180255 541124
rect 180389 541124 180401 541127
rect 180435 541127 180593 541158
rect 180435 541124 180447 541127
rect 180389 541118 180447 541124
rect 180581 541124 180593 541127
rect 180627 541124 180855 541158
rect 180581 541118 180855 541124
rect 179280 541050 179420 541117
rect 180625 541112 180855 541118
rect 179280 540997 179286 541050
rect 177680 540862 178420 540927
rect 178880 540917 179286 540997
rect 178880 540867 179080 540917
rect 176787 540787 176945 540807
rect 176979 540787 177010 540807
rect 176787 540687 176890 540787
rect 177000 540687 177010 540787
rect 176787 540667 176945 540687
rect 176787 540569 176793 540667
rect 176747 540557 176793 540569
rect 176843 540603 176889 540615
rect 176843 540317 176849 540603
rect 176691 540115 176849 540317
rect 176883 540317 176889 540603
rect 176939 540569 176945 540667
rect 176979 540667 177010 540687
rect 177200 540812 178420 540862
rect 176979 540569 176985 540667
rect 176939 540557 176985 540569
rect 177035 540603 177081 540615
rect 177035 540317 177041 540603
rect 176883 540115 177041 540317
rect 177075 540115 177081 540603
rect 177200 540367 177250 540812
rect 177680 540727 178420 540812
rect 177360 540596 177406 540608
rect 177200 540357 177260 540367
rect 177198 540351 177260 540357
rect 177198 540317 177210 540351
rect 177244 540317 177260 540351
rect 177198 540311 177260 540317
rect 177200 540307 177260 540311
rect 177160 540267 177206 540279
rect 177160 540187 177166 540267
rect 175850 540107 177081 540115
rect 175850 540103 175929 540107
rect 176075 540103 176121 540107
rect 176267 540103 176313 540107
rect 176459 540103 176505 540107
rect 176651 540103 176697 540107
rect 176843 540103 176889 540107
rect 177035 540103 177081 540107
rect 175850 540097 175920 540103
rect 175710 540041 175780 540057
rect 175710 540007 175730 540041
rect 175764 540007 175780 540041
rect 175710 539987 175780 540007
rect 175850 539787 175880 540097
rect 177140 540091 177166 540187
rect 177200 540091 177206 540267
rect 177140 540079 177206 540091
rect 177248 540267 177294 540279
rect 177248 540091 177254 540267
rect 177288 540257 177294 540267
rect 177360 540257 177366 540596
rect 177288 540108 177366 540257
rect 177400 540267 177406 540596
rect 177448 540596 177494 540608
rect 177448 540267 177454 540596
rect 177400 540108 177454 540267
rect 177488 540267 177494 540596
rect 177670 540277 177890 540287
rect 177488 540257 177510 540267
rect 177670 540257 177700 540277
rect 177488 540247 177700 540257
rect 177488 540117 177570 540247
rect 177630 540117 177700 540247
rect 177488 540108 177700 540117
rect 177288 540107 177700 540108
rect 177288 540091 177294 540107
rect 177360 540096 177494 540107
rect 177670 540097 177700 540107
rect 177880 540097 177890 540277
rect 177248 540079 177294 540091
rect 175925 540048 175983 540054
rect 175925 540047 175937 540048
rect 175920 540014 175937 540047
rect 175971 540047 175983 540048
rect 176117 540048 176175 540054
rect 176117 540047 176129 540048
rect 175971 540014 176129 540047
rect 176163 540047 176175 540048
rect 176309 540048 176367 540054
rect 176309 540047 176321 540048
rect 176163 540014 176321 540047
rect 176355 540047 176367 540048
rect 176501 540048 176559 540054
rect 176501 540047 176513 540048
rect 176355 540014 176513 540047
rect 176547 540047 176559 540048
rect 176693 540048 176751 540054
rect 176693 540047 176705 540048
rect 176547 540014 176705 540047
rect 176739 540047 176751 540048
rect 176885 540048 176943 540054
rect 176885 540047 176897 540048
rect 176739 540014 176897 540047
rect 176931 540014 176943 540048
rect 175920 540008 176943 540014
rect 175920 539987 176940 540008
rect 175280 539687 175880 539787
rect 175280 537963 175480 539687
rect 175640 539638 175880 539687
rect 175640 539604 175714 539638
rect 175748 539604 175880 539638
rect 175640 539545 175880 539604
rect 176020 539651 177030 539657
rect 176020 539645 177043 539651
rect 176020 539611 176037 539645
rect 176071 539611 176229 539645
rect 176263 539611 176421 539645
rect 176455 539611 176613 539645
rect 176647 539611 176805 539645
rect 176839 539611 176997 539645
rect 177031 539611 177043 539645
rect 176020 539605 177043 539611
rect 176020 539597 177030 539605
rect 177140 539557 177170 540079
rect 177198 540041 177260 540047
rect 177198 540007 177210 540041
rect 177244 540007 177260 540041
rect 177198 540001 177260 540007
rect 177200 539638 177260 540001
rect 177370 540041 177490 540096
rect 177670 540087 177890 540097
rect 177370 540007 177410 540041
rect 177444 540007 177490 540041
rect 177370 539987 177490 540007
rect 177200 539604 177214 539638
rect 177248 539604 177260 539638
rect 177200 539597 177260 539604
rect 177400 539638 177480 539657
rect 177400 539604 177414 539638
rect 177448 539604 177480 539638
rect 177400 539597 177480 539604
rect 175640 539447 175670 539545
rect 175664 538569 175670 539447
rect 175704 539447 175758 539545
rect 175704 538569 175710 539447
rect 175664 538557 175710 538569
rect 175752 538569 175758 539447
rect 175792 539527 175880 539545
rect 175983 539535 176029 539547
rect 175792 539517 175950 539527
rect 175983 539517 175989 539535
rect 175792 539447 175989 539517
rect 175792 538569 175798 539447
rect 175850 539237 175989 539447
rect 175887 539081 175933 539093
rect 175887 538593 175893 539081
rect 175927 538967 175933 539081
rect 175983 539047 175989 539237
rect 176023 539517 176029 539535
rect 176175 539535 176221 539547
rect 176175 539517 176181 539535
rect 176023 539237 176181 539517
rect 176023 539047 176029 539237
rect 175983 539035 176029 539047
rect 176079 539081 176125 539093
rect 176079 538967 176085 539081
rect 175927 538593 176085 538967
rect 176119 538967 176125 539081
rect 176175 539047 176181 539237
rect 176215 539517 176221 539535
rect 176367 539535 176413 539547
rect 176367 539517 176373 539535
rect 176215 539237 176373 539517
rect 176215 539047 176221 539237
rect 176175 539035 176221 539047
rect 176271 539081 176317 539093
rect 176271 538967 176277 539081
rect 176119 538593 176277 538967
rect 176311 538967 176317 539081
rect 176367 539047 176373 539237
rect 176407 539517 176413 539535
rect 176559 539535 176605 539547
rect 176559 539517 176565 539535
rect 176407 539237 176565 539517
rect 176407 539047 176413 539237
rect 176367 539035 176413 539047
rect 176463 539081 176509 539093
rect 176463 538967 176469 539081
rect 176311 538593 176469 538967
rect 176503 538967 176509 539081
rect 176559 539047 176565 539237
rect 176599 539517 176605 539535
rect 176751 539535 176797 539547
rect 176751 539517 176757 539535
rect 176599 539237 176757 539517
rect 176599 539047 176605 539237
rect 176559 539035 176605 539047
rect 176655 539081 176701 539093
rect 176655 538967 176661 539081
rect 176503 538593 176661 538967
rect 176695 538967 176701 539081
rect 176751 539047 176757 539237
rect 176791 539517 176797 539535
rect 176943 539535 176989 539547
rect 176943 539517 176949 539535
rect 176791 539237 176949 539517
rect 176791 539047 176797 539237
rect 176751 539035 176797 539047
rect 176847 539081 176893 539093
rect 176847 538967 176853 539081
rect 176695 538593 176853 538967
rect 176887 538967 176893 539081
rect 176943 539047 176949 539237
rect 176983 539517 176989 539535
rect 177140 539545 177210 539557
rect 176983 539237 177000 539517
rect 177140 539407 177170 539545
rect 176983 539047 176989 539237
rect 176943 539035 176989 539047
rect 177039 539081 177085 539093
rect 177039 538967 177045 539081
rect 176887 538837 177045 538967
rect 176887 538737 176900 538837
rect 177040 538737 177045 538837
rect 176887 538593 177045 538737
rect 177079 538593 177085 539081
rect 177164 539067 177170 539407
rect 175887 538587 177085 538593
rect 175887 538581 175933 538587
rect 176079 538581 176125 538587
rect 176271 538581 176317 538587
rect 176463 538581 176509 538587
rect 176655 538581 176701 538587
rect 176847 538581 176893 538587
rect 177039 538581 177085 538587
rect 177130 538969 177170 539067
rect 177204 538969 177210 539545
rect 177130 538957 177210 538969
rect 177252 539545 177298 539557
rect 177252 538969 177258 539545
rect 177292 539537 177298 539545
rect 177292 539307 177410 539537
rect 177670 539337 177890 539347
rect 177670 539307 177690 539337
rect 177292 539297 177690 539307
rect 177292 539207 177570 539297
rect 177620 539207 177690 539297
rect 177292 539197 177690 539207
rect 177292 539074 177410 539197
rect 177670 539157 177690 539197
rect 177870 539157 177890 539337
rect 177670 539147 177890 539157
rect 177292 538969 177370 539074
rect 177252 538967 177370 538969
rect 177252 538957 177298 538967
rect 175752 538557 175798 538569
rect 175929 538517 175987 538523
rect 176121 538517 176179 538523
rect 176313 538517 176371 538523
rect 176505 538517 176563 538523
rect 176697 538517 176755 538523
rect 176889 538517 176947 538523
rect 177130 538517 177170 538957
rect 177200 538910 177260 538917
rect 177200 538876 177214 538910
rect 177248 538876 177260 538910
rect 177200 538857 177260 538876
rect 177364 538607 177370 538967
rect 175700 538510 175760 538517
rect 175700 538476 175714 538510
rect 175748 538476 175760 538510
rect 175700 538457 175760 538476
rect 175920 538483 175941 538517
rect 175975 538483 176133 538517
rect 176167 538483 176325 538517
rect 176359 538483 176517 538517
rect 176551 538483 176709 538517
rect 176743 538483 176901 538517
rect 176935 538483 177170 538517
rect 175920 538457 177170 538483
rect 177360 538586 177370 538607
rect 177404 538607 177410 539074
rect 177452 539074 177498 539086
rect 177452 538607 177458 539074
rect 177404 538586 177458 538607
rect 177492 538586 177498 539074
rect 177360 538574 177498 538586
rect 177360 538510 177480 538574
rect 177360 538477 177414 538510
rect 177400 538476 177414 538477
rect 177448 538477 177480 538510
rect 177448 538476 177460 538477
rect 177400 538457 177460 538476
rect 175280 537847 175360 537963
rect 175354 537566 175360 537847
rect 175398 537847 175480 537963
rect 175398 537566 175404 537847
rect 175354 537554 175404 537566
rect 175354 536448 175404 536460
rect 175354 536327 175360 536448
rect 175230 536287 175360 536327
rect 175398 536327 175404 536448
rect 175398 536287 175580 536327
rect 175230 535977 175280 536287
rect 175500 535977 175580 536287
rect 175230 535927 175580 535977
rect 171050 533337 173930 533537
rect 174680 533337 176730 533537
rect 173730 532787 173930 533337
rect 167520 532767 172530 532787
rect 167520 532597 172360 532767
rect 172490 532597 172530 532767
rect 167520 532587 172530 532597
rect 173730 532777 174730 532787
rect 173730 532607 174490 532777
rect 174620 532607 174730 532777
rect 173730 532587 174730 532607
rect 176530 532767 176730 533337
rect 176530 532597 176580 532767
rect 176710 532597 176730 532767
rect 176530 532487 176730 532597
rect 178220 532787 178420 540727
rect 179280 540562 179286 540917
rect 179320 540917 179374 541050
rect 179320 540562 179326 540917
rect 179280 540550 179326 540562
rect 179368 540562 179374 540917
rect 179408 540997 179420 541050
rect 179579 541057 179625 541069
rect 179771 541057 179817 541069
rect 179963 541057 180009 541069
rect 180155 541057 180201 541069
rect 180347 541057 180393 541069
rect 180539 541057 180585 541069
rect 179579 540997 179585 541057
rect 179408 540917 179585 540997
rect 179408 540562 179414 540917
rect 179368 540550 179414 540562
rect 179483 540603 179529 540615
rect 179483 540317 179489 540603
rect 179450 540115 179489 540317
rect 179523 540317 179529 540603
rect 179579 540569 179585 540917
rect 179619 540667 179777 541057
rect 179619 540569 179625 540667
rect 179579 540557 179625 540569
rect 179675 540603 179721 540615
rect 179675 540317 179681 540603
rect 179523 540115 179681 540317
rect 179715 540317 179721 540603
rect 179771 540569 179777 540667
rect 179811 540667 179969 541057
rect 179811 540569 179817 540667
rect 179771 540557 179817 540569
rect 179867 540603 179913 540615
rect 179867 540317 179873 540603
rect 179715 540115 179873 540317
rect 179907 540317 179913 540603
rect 179963 540569 179969 540667
rect 180003 540667 180161 541057
rect 180003 540569 180009 540667
rect 179963 540557 180009 540569
rect 180059 540603 180105 540615
rect 180059 540317 180065 540603
rect 179907 540115 180065 540317
rect 180099 540317 180105 540603
rect 180155 540569 180161 540667
rect 180195 540667 180353 541057
rect 180195 540569 180201 540667
rect 180155 540557 180201 540569
rect 180251 540603 180297 540615
rect 180251 540317 180257 540603
rect 180099 540115 180257 540317
rect 180291 540317 180297 540603
rect 180347 540569 180353 540667
rect 180387 541027 180545 541057
rect 180579 541027 180610 541057
rect 180387 540927 180490 541027
rect 180600 540927 180610 541027
rect 180387 540907 180545 540927
rect 180579 540907 180610 540927
rect 180387 540807 180490 540907
rect 180600 540807 180610 540907
rect 180805 540862 180855 541112
rect 180998 541151 181060 541157
rect 180998 541117 181010 541151
rect 181044 541117 181060 541151
rect 180998 541111 181060 541117
rect 181000 541097 181060 541111
rect 182180 540997 182380 541537
rect 182620 541157 182680 541167
rect 182920 541162 183940 541187
rect 182920 541158 184155 541162
rect 182580 541151 182720 541157
rect 182580 541117 182630 541151
rect 182664 541117 182720 541151
rect 182920 541127 182933 541158
rect 182921 541124 182933 541127
rect 182967 541127 183125 541158
rect 182967 541124 182979 541127
rect 182921 541118 182979 541124
rect 183113 541124 183125 541127
rect 183159 541127 183317 541158
rect 183159 541124 183171 541127
rect 183113 541118 183171 541124
rect 183305 541124 183317 541127
rect 183351 541127 183509 541158
rect 183351 541124 183363 541127
rect 183305 541118 183363 541124
rect 183497 541124 183509 541127
rect 183543 541127 183701 541158
rect 183543 541124 183555 541127
rect 183497 541118 183555 541124
rect 183689 541124 183701 541127
rect 183735 541127 183893 541158
rect 183735 541124 183747 541127
rect 183689 541118 183747 541124
rect 183881 541124 183893 541127
rect 183927 541124 184155 541158
rect 183881 541118 184155 541124
rect 182580 541050 182720 541117
rect 183925 541112 184155 541118
rect 182580 540997 182586 541050
rect 181280 540862 181930 540927
rect 182180 540917 182586 540997
rect 182180 540867 182380 540917
rect 180387 540787 180545 540807
rect 180579 540787 180610 540807
rect 180387 540687 180490 540787
rect 180600 540687 180610 540787
rect 180387 540667 180545 540687
rect 180387 540569 180393 540667
rect 180347 540557 180393 540569
rect 180443 540603 180489 540615
rect 180443 540317 180449 540603
rect 180291 540115 180449 540317
rect 180483 540317 180489 540603
rect 180539 540569 180545 540667
rect 180579 540667 180610 540687
rect 180800 540812 181930 540862
rect 180579 540569 180585 540667
rect 180539 540557 180585 540569
rect 180635 540603 180681 540615
rect 180635 540317 180641 540603
rect 180483 540115 180641 540317
rect 180675 540115 180681 540603
rect 180800 540367 180850 540812
rect 181280 540727 181930 540812
rect 180960 540596 181006 540608
rect 180800 540357 180860 540367
rect 180798 540351 180860 540357
rect 180798 540317 180810 540351
rect 180844 540317 180860 540351
rect 180798 540311 180860 540317
rect 180800 540307 180860 540311
rect 180760 540267 180806 540279
rect 180760 540187 180766 540267
rect 179450 540107 180681 540115
rect 179450 540103 179529 540107
rect 179675 540103 179721 540107
rect 179867 540103 179913 540107
rect 180059 540103 180105 540107
rect 180251 540103 180297 540107
rect 180443 540103 180489 540107
rect 180635 540103 180681 540107
rect 179450 540097 179520 540103
rect 179310 540041 179380 540057
rect 179310 540007 179330 540041
rect 179364 540007 179380 540041
rect 179310 539987 179380 540007
rect 179450 539787 179480 540097
rect 180740 540091 180766 540187
rect 180800 540091 180806 540267
rect 180740 540079 180806 540091
rect 180848 540267 180894 540279
rect 180848 540091 180854 540267
rect 180888 540257 180894 540267
rect 180960 540257 180966 540596
rect 180888 540108 180966 540257
rect 181000 540267 181006 540596
rect 181048 540596 181094 540608
rect 181048 540267 181054 540596
rect 181000 540108 181054 540267
rect 181088 540267 181094 540596
rect 181270 540277 181490 540287
rect 181088 540257 181110 540267
rect 181270 540257 181290 540277
rect 181088 540247 181290 540257
rect 181088 540117 181170 540247
rect 181230 540117 181290 540247
rect 181088 540108 181290 540117
rect 180888 540107 181290 540108
rect 180888 540091 180894 540107
rect 180960 540096 181094 540107
rect 181270 540097 181290 540107
rect 181470 540097 181490 540277
rect 180848 540079 180894 540091
rect 179525 540048 179583 540054
rect 179525 540047 179537 540048
rect 179520 540014 179537 540047
rect 179571 540047 179583 540048
rect 179717 540048 179775 540054
rect 179717 540047 179729 540048
rect 179571 540014 179729 540047
rect 179763 540047 179775 540048
rect 179909 540048 179967 540054
rect 179909 540047 179921 540048
rect 179763 540014 179921 540047
rect 179955 540047 179967 540048
rect 180101 540048 180159 540054
rect 180101 540047 180113 540048
rect 179955 540014 180113 540047
rect 180147 540047 180159 540048
rect 180293 540048 180351 540054
rect 180293 540047 180305 540048
rect 180147 540014 180305 540047
rect 180339 540047 180351 540048
rect 180485 540048 180543 540054
rect 180485 540047 180497 540048
rect 180339 540014 180497 540047
rect 180531 540014 180543 540048
rect 179520 540008 180543 540014
rect 179520 539987 180540 540008
rect 178880 539687 179480 539787
rect 178880 537963 179080 539687
rect 179240 539638 179480 539687
rect 179240 539604 179314 539638
rect 179348 539604 179480 539638
rect 179240 539545 179480 539604
rect 179620 539651 180630 539657
rect 179620 539645 180643 539651
rect 179620 539611 179637 539645
rect 179671 539611 179829 539645
rect 179863 539611 180021 539645
rect 180055 539611 180213 539645
rect 180247 539611 180405 539645
rect 180439 539611 180597 539645
rect 180631 539611 180643 539645
rect 179620 539605 180643 539611
rect 179620 539597 180630 539605
rect 180740 539557 180770 540079
rect 180798 540041 180860 540047
rect 180798 540007 180810 540041
rect 180844 540007 180860 540041
rect 180798 540001 180860 540007
rect 180800 539638 180860 540001
rect 180970 540041 181090 540096
rect 181270 540087 181490 540097
rect 180970 540007 181010 540041
rect 181044 540007 181090 540041
rect 180970 539987 181090 540007
rect 180800 539604 180814 539638
rect 180848 539604 180860 539638
rect 180800 539597 180860 539604
rect 181000 539638 181080 539657
rect 181000 539604 181014 539638
rect 181048 539604 181080 539638
rect 181000 539597 181080 539604
rect 179240 539447 179270 539545
rect 179264 538569 179270 539447
rect 179304 539447 179358 539545
rect 179304 538569 179310 539447
rect 179264 538557 179310 538569
rect 179352 538569 179358 539447
rect 179392 539527 179480 539545
rect 179583 539535 179629 539547
rect 179392 539517 179550 539527
rect 179583 539517 179589 539535
rect 179392 539447 179589 539517
rect 179392 538569 179398 539447
rect 179450 539237 179589 539447
rect 179487 539081 179533 539093
rect 179487 538593 179493 539081
rect 179527 538967 179533 539081
rect 179583 539047 179589 539237
rect 179623 539517 179629 539535
rect 179775 539535 179821 539547
rect 179775 539517 179781 539535
rect 179623 539237 179781 539517
rect 179623 539047 179629 539237
rect 179583 539035 179629 539047
rect 179679 539081 179725 539093
rect 179679 538967 179685 539081
rect 179527 538593 179685 538967
rect 179719 538967 179725 539081
rect 179775 539047 179781 539237
rect 179815 539517 179821 539535
rect 179967 539535 180013 539547
rect 179967 539517 179973 539535
rect 179815 539237 179973 539517
rect 179815 539047 179821 539237
rect 179775 539035 179821 539047
rect 179871 539081 179917 539093
rect 179871 538967 179877 539081
rect 179719 538593 179877 538967
rect 179911 538967 179917 539081
rect 179967 539047 179973 539237
rect 180007 539517 180013 539535
rect 180159 539535 180205 539547
rect 180159 539517 180165 539535
rect 180007 539237 180165 539517
rect 180007 539047 180013 539237
rect 179967 539035 180013 539047
rect 180063 539081 180109 539093
rect 180063 538967 180069 539081
rect 179911 538593 180069 538967
rect 180103 538967 180109 539081
rect 180159 539047 180165 539237
rect 180199 539517 180205 539535
rect 180351 539535 180397 539547
rect 180351 539517 180357 539535
rect 180199 539237 180357 539517
rect 180199 539047 180205 539237
rect 180159 539035 180205 539047
rect 180255 539081 180301 539093
rect 180255 538967 180261 539081
rect 180103 538593 180261 538967
rect 180295 538967 180301 539081
rect 180351 539047 180357 539237
rect 180391 539517 180397 539535
rect 180543 539535 180589 539547
rect 180543 539517 180549 539535
rect 180391 539237 180549 539517
rect 180391 539047 180397 539237
rect 180351 539035 180397 539047
rect 180447 539081 180493 539093
rect 180447 538967 180453 539081
rect 180295 538593 180453 538967
rect 180487 538967 180493 539081
rect 180543 539047 180549 539237
rect 180583 539517 180589 539535
rect 180740 539545 180810 539557
rect 180583 539237 180600 539517
rect 180740 539407 180770 539545
rect 180583 539047 180589 539237
rect 180543 539035 180589 539047
rect 180639 539081 180685 539093
rect 180639 538967 180645 539081
rect 180487 538837 180645 538967
rect 180487 538737 180500 538837
rect 180640 538737 180645 538837
rect 180487 538593 180645 538737
rect 180679 538593 180685 539081
rect 180764 539067 180770 539407
rect 179487 538587 180685 538593
rect 179487 538581 179533 538587
rect 179679 538581 179725 538587
rect 179871 538581 179917 538587
rect 180063 538581 180109 538587
rect 180255 538581 180301 538587
rect 180447 538581 180493 538587
rect 180639 538581 180685 538587
rect 180730 538969 180770 539067
rect 180804 538969 180810 539545
rect 180730 538957 180810 538969
rect 180852 539545 180898 539557
rect 180852 538969 180858 539545
rect 180892 539537 180898 539545
rect 180892 539307 181010 539537
rect 181270 539337 181490 539347
rect 181270 539307 181290 539337
rect 180892 539297 181290 539307
rect 180892 539207 181170 539297
rect 181220 539207 181290 539297
rect 180892 539197 181290 539207
rect 180892 539074 181010 539197
rect 181270 539157 181290 539197
rect 181470 539157 181490 539337
rect 181270 539147 181490 539157
rect 180892 538969 180970 539074
rect 180852 538967 180970 538969
rect 180852 538957 180898 538967
rect 179352 538557 179398 538569
rect 179529 538517 179587 538523
rect 179721 538517 179779 538523
rect 179913 538517 179971 538523
rect 180105 538517 180163 538523
rect 180297 538517 180355 538523
rect 180489 538517 180547 538523
rect 180730 538517 180770 538957
rect 180800 538910 180860 538917
rect 180800 538876 180814 538910
rect 180848 538876 180860 538910
rect 180800 538857 180860 538876
rect 180964 538607 180970 538967
rect 179300 538510 179360 538517
rect 179300 538476 179314 538510
rect 179348 538476 179360 538510
rect 179300 538457 179360 538476
rect 179520 538483 179541 538517
rect 179575 538483 179733 538517
rect 179767 538483 179925 538517
rect 179959 538483 180117 538517
rect 180151 538483 180309 538517
rect 180343 538483 180501 538517
rect 180535 538483 180770 538517
rect 179520 538457 180770 538483
rect 180960 538586 180970 538607
rect 181004 538607 181010 539074
rect 181052 539074 181098 539086
rect 181052 538607 181058 539074
rect 181004 538586 181058 538607
rect 181092 538586 181098 539074
rect 180960 538574 181098 538586
rect 180960 538510 181080 538574
rect 180960 538477 181014 538510
rect 181000 538476 181014 538477
rect 181048 538477 181080 538510
rect 181048 538476 181060 538477
rect 181000 538457 181060 538476
rect 178880 537847 178960 537963
rect 178954 537566 178960 537847
rect 178998 537847 179080 537963
rect 178998 537566 179004 537847
rect 178954 537554 179004 537566
rect 178954 537008 179004 537020
rect 178954 536997 178960 537008
rect 178820 536611 178960 536997
rect 178998 536997 179004 537008
rect 178998 536611 179120 536997
rect 178820 536307 179120 536611
rect 178820 535997 178870 536307
rect 179070 535997 179120 536307
rect 178820 535897 179120 535997
rect 181730 533537 181930 540727
rect 182580 540562 182586 540917
rect 182620 540917 182674 541050
rect 182620 540562 182626 540917
rect 182580 540550 182626 540562
rect 182668 540562 182674 540917
rect 182708 540997 182720 541050
rect 182879 541057 182925 541069
rect 183071 541057 183117 541069
rect 183263 541057 183309 541069
rect 183455 541057 183501 541069
rect 183647 541057 183693 541069
rect 183839 541057 183885 541069
rect 182879 540997 182885 541057
rect 182708 540917 182885 540997
rect 182708 540562 182714 540917
rect 182668 540550 182714 540562
rect 182783 540603 182829 540615
rect 182783 540317 182789 540603
rect 182750 540115 182789 540317
rect 182823 540317 182829 540603
rect 182879 540569 182885 540917
rect 182919 540667 183077 541057
rect 182919 540569 182925 540667
rect 182879 540557 182925 540569
rect 182975 540603 183021 540615
rect 182975 540317 182981 540603
rect 182823 540115 182981 540317
rect 183015 540317 183021 540603
rect 183071 540569 183077 540667
rect 183111 540667 183269 541057
rect 183111 540569 183117 540667
rect 183071 540557 183117 540569
rect 183167 540603 183213 540615
rect 183167 540317 183173 540603
rect 183015 540115 183173 540317
rect 183207 540317 183213 540603
rect 183263 540569 183269 540667
rect 183303 540667 183461 541057
rect 183303 540569 183309 540667
rect 183263 540557 183309 540569
rect 183359 540603 183405 540615
rect 183359 540317 183365 540603
rect 183207 540115 183365 540317
rect 183399 540317 183405 540603
rect 183455 540569 183461 540667
rect 183495 540667 183653 541057
rect 183495 540569 183501 540667
rect 183455 540557 183501 540569
rect 183551 540603 183597 540615
rect 183551 540317 183557 540603
rect 183399 540115 183557 540317
rect 183591 540317 183597 540603
rect 183647 540569 183653 540667
rect 183687 541027 183845 541057
rect 183879 541027 183910 541057
rect 183687 540927 183790 541027
rect 183900 540927 183910 541027
rect 183687 540907 183845 540927
rect 183879 540907 183910 540927
rect 183687 540807 183790 540907
rect 183900 540807 183910 540907
rect 184105 540862 184155 541112
rect 184298 541151 184360 541157
rect 184298 541117 184310 541151
rect 184344 541117 184360 541151
rect 184298 541111 184360 541117
rect 184300 541097 184360 541111
rect 185480 540997 185680 541537
rect 185920 541157 185980 541167
rect 186220 541162 187240 541187
rect 186220 541158 187455 541162
rect 185880 541151 186020 541157
rect 185880 541117 185930 541151
rect 185964 541117 186020 541151
rect 186220 541127 186233 541158
rect 186221 541124 186233 541127
rect 186267 541127 186425 541158
rect 186267 541124 186279 541127
rect 186221 541118 186279 541124
rect 186413 541124 186425 541127
rect 186459 541127 186617 541158
rect 186459 541124 186471 541127
rect 186413 541118 186471 541124
rect 186605 541124 186617 541127
rect 186651 541127 186809 541158
rect 186651 541124 186663 541127
rect 186605 541118 186663 541124
rect 186797 541124 186809 541127
rect 186843 541127 187001 541158
rect 186843 541124 186855 541127
rect 186797 541118 186855 541124
rect 186989 541124 187001 541127
rect 187035 541127 187193 541158
rect 187035 541124 187047 541127
rect 186989 541118 187047 541124
rect 187181 541124 187193 541127
rect 187227 541124 187455 541158
rect 187181 541118 187455 541124
rect 185880 541050 186020 541117
rect 187225 541112 187455 541118
rect 185880 540997 185886 541050
rect 184580 540862 185170 540927
rect 185480 540917 185886 540997
rect 185480 540867 185680 540917
rect 183687 540787 183845 540807
rect 183879 540787 183910 540807
rect 183687 540687 183790 540787
rect 183900 540687 183910 540787
rect 183687 540667 183845 540687
rect 183687 540569 183693 540667
rect 183647 540557 183693 540569
rect 183743 540603 183789 540615
rect 183743 540317 183749 540603
rect 183591 540115 183749 540317
rect 183783 540317 183789 540603
rect 183839 540569 183845 540667
rect 183879 540667 183910 540687
rect 184100 540812 185170 540862
rect 183879 540569 183885 540667
rect 183839 540557 183885 540569
rect 183935 540603 183981 540615
rect 183935 540317 183941 540603
rect 183783 540115 183941 540317
rect 183975 540115 183981 540603
rect 184100 540367 184150 540812
rect 184580 540727 185170 540812
rect 184260 540596 184306 540608
rect 184100 540357 184160 540367
rect 184098 540351 184160 540357
rect 184098 540317 184110 540351
rect 184144 540317 184160 540351
rect 184098 540311 184160 540317
rect 184100 540307 184160 540311
rect 184060 540267 184106 540279
rect 184060 540187 184066 540267
rect 182750 540107 183981 540115
rect 182750 540103 182829 540107
rect 182975 540103 183021 540107
rect 183167 540103 183213 540107
rect 183359 540103 183405 540107
rect 183551 540103 183597 540107
rect 183743 540103 183789 540107
rect 183935 540103 183981 540107
rect 182750 540097 182820 540103
rect 182610 540041 182680 540057
rect 182610 540007 182630 540041
rect 182664 540007 182680 540041
rect 182610 539987 182680 540007
rect 182750 539787 182780 540097
rect 184040 540091 184066 540187
rect 184100 540091 184106 540267
rect 184040 540079 184106 540091
rect 184148 540267 184194 540279
rect 184148 540091 184154 540267
rect 184188 540257 184194 540267
rect 184260 540257 184266 540596
rect 184188 540108 184266 540257
rect 184300 540267 184306 540596
rect 184348 540596 184394 540608
rect 184348 540267 184354 540596
rect 184300 540108 184354 540267
rect 184388 540267 184394 540596
rect 184570 540277 184790 540287
rect 184388 540257 184410 540267
rect 184570 540257 184590 540277
rect 184388 540247 184590 540257
rect 184388 540117 184470 540247
rect 184530 540117 184590 540247
rect 184388 540108 184590 540117
rect 184188 540107 184590 540108
rect 184188 540091 184194 540107
rect 184260 540096 184394 540107
rect 184570 540097 184590 540107
rect 184770 540097 184790 540277
rect 184148 540079 184194 540091
rect 182825 540048 182883 540054
rect 182825 540047 182837 540048
rect 182820 540014 182837 540047
rect 182871 540047 182883 540048
rect 183017 540048 183075 540054
rect 183017 540047 183029 540048
rect 182871 540014 183029 540047
rect 183063 540047 183075 540048
rect 183209 540048 183267 540054
rect 183209 540047 183221 540048
rect 183063 540014 183221 540047
rect 183255 540047 183267 540048
rect 183401 540048 183459 540054
rect 183401 540047 183413 540048
rect 183255 540014 183413 540047
rect 183447 540047 183459 540048
rect 183593 540048 183651 540054
rect 183593 540047 183605 540048
rect 183447 540014 183605 540047
rect 183639 540047 183651 540048
rect 183785 540048 183843 540054
rect 183785 540047 183797 540048
rect 183639 540014 183797 540047
rect 183831 540014 183843 540048
rect 182820 540008 183843 540014
rect 182820 539987 183840 540008
rect 182180 539687 182780 539787
rect 182180 537963 182380 539687
rect 182540 539638 182780 539687
rect 182540 539604 182614 539638
rect 182648 539604 182780 539638
rect 182540 539545 182780 539604
rect 182920 539651 183930 539657
rect 182920 539645 183943 539651
rect 182920 539611 182937 539645
rect 182971 539611 183129 539645
rect 183163 539611 183321 539645
rect 183355 539611 183513 539645
rect 183547 539611 183705 539645
rect 183739 539611 183897 539645
rect 183931 539611 183943 539645
rect 182920 539605 183943 539611
rect 182920 539597 183930 539605
rect 184040 539557 184070 540079
rect 184098 540041 184160 540047
rect 184098 540007 184110 540041
rect 184144 540007 184160 540041
rect 184098 540001 184160 540007
rect 184100 539638 184160 540001
rect 184270 540041 184390 540096
rect 184570 540087 184790 540097
rect 184270 540007 184310 540041
rect 184344 540007 184390 540041
rect 184270 539987 184390 540007
rect 184100 539604 184114 539638
rect 184148 539604 184160 539638
rect 184100 539597 184160 539604
rect 184300 539638 184380 539657
rect 184300 539604 184314 539638
rect 184348 539604 184380 539638
rect 184300 539597 184380 539604
rect 182540 539447 182570 539545
rect 182564 538569 182570 539447
rect 182604 539447 182658 539545
rect 182604 538569 182610 539447
rect 182564 538557 182610 538569
rect 182652 538569 182658 539447
rect 182692 539527 182780 539545
rect 182883 539535 182929 539547
rect 182692 539517 182850 539527
rect 182883 539517 182889 539535
rect 182692 539447 182889 539517
rect 182692 538569 182698 539447
rect 182750 539237 182889 539447
rect 182787 539081 182833 539093
rect 182787 538593 182793 539081
rect 182827 538967 182833 539081
rect 182883 539047 182889 539237
rect 182923 539517 182929 539535
rect 183075 539535 183121 539547
rect 183075 539517 183081 539535
rect 182923 539237 183081 539517
rect 182923 539047 182929 539237
rect 182883 539035 182929 539047
rect 182979 539081 183025 539093
rect 182979 538967 182985 539081
rect 182827 538593 182985 538967
rect 183019 538967 183025 539081
rect 183075 539047 183081 539237
rect 183115 539517 183121 539535
rect 183267 539535 183313 539547
rect 183267 539517 183273 539535
rect 183115 539237 183273 539517
rect 183115 539047 183121 539237
rect 183075 539035 183121 539047
rect 183171 539081 183217 539093
rect 183171 538967 183177 539081
rect 183019 538593 183177 538967
rect 183211 538967 183217 539081
rect 183267 539047 183273 539237
rect 183307 539517 183313 539535
rect 183459 539535 183505 539547
rect 183459 539517 183465 539535
rect 183307 539237 183465 539517
rect 183307 539047 183313 539237
rect 183267 539035 183313 539047
rect 183363 539081 183409 539093
rect 183363 538967 183369 539081
rect 183211 538593 183369 538967
rect 183403 538967 183409 539081
rect 183459 539047 183465 539237
rect 183499 539517 183505 539535
rect 183651 539535 183697 539547
rect 183651 539517 183657 539535
rect 183499 539237 183657 539517
rect 183499 539047 183505 539237
rect 183459 539035 183505 539047
rect 183555 539081 183601 539093
rect 183555 538967 183561 539081
rect 183403 538593 183561 538967
rect 183595 538967 183601 539081
rect 183651 539047 183657 539237
rect 183691 539517 183697 539535
rect 183843 539535 183889 539547
rect 183843 539517 183849 539535
rect 183691 539237 183849 539517
rect 183691 539047 183697 539237
rect 183651 539035 183697 539047
rect 183747 539081 183793 539093
rect 183747 538967 183753 539081
rect 183595 538593 183753 538967
rect 183787 538967 183793 539081
rect 183843 539047 183849 539237
rect 183883 539517 183889 539535
rect 184040 539545 184110 539557
rect 183883 539237 183900 539517
rect 184040 539407 184070 539545
rect 183883 539047 183889 539237
rect 183843 539035 183889 539047
rect 183939 539081 183985 539093
rect 183939 538967 183945 539081
rect 183787 538837 183945 538967
rect 183787 538737 183800 538837
rect 183940 538737 183945 538837
rect 183787 538593 183945 538737
rect 183979 538593 183985 539081
rect 184064 539067 184070 539407
rect 182787 538587 183985 538593
rect 182787 538581 182833 538587
rect 182979 538581 183025 538587
rect 183171 538581 183217 538587
rect 183363 538581 183409 538587
rect 183555 538581 183601 538587
rect 183747 538581 183793 538587
rect 183939 538581 183985 538587
rect 184030 538969 184070 539067
rect 184104 538969 184110 539545
rect 184030 538957 184110 538969
rect 184152 539545 184198 539557
rect 184152 538969 184158 539545
rect 184192 539537 184198 539545
rect 184192 539307 184310 539537
rect 184570 539337 184790 539347
rect 184570 539307 184590 539337
rect 184192 539297 184590 539307
rect 184192 539207 184470 539297
rect 184520 539207 184590 539297
rect 184192 539197 184590 539207
rect 184192 539074 184310 539197
rect 184570 539157 184590 539197
rect 184770 539157 184790 539337
rect 184570 539147 184790 539157
rect 184192 538969 184270 539074
rect 184152 538967 184270 538969
rect 184152 538957 184198 538967
rect 182652 538557 182698 538569
rect 182829 538517 182887 538523
rect 183021 538517 183079 538523
rect 183213 538517 183271 538523
rect 183405 538517 183463 538523
rect 183597 538517 183655 538523
rect 183789 538517 183847 538523
rect 184030 538517 184070 538957
rect 184100 538910 184160 538917
rect 184100 538876 184114 538910
rect 184148 538876 184160 538910
rect 184100 538857 184160 538876
rect 184264 538607 184270 538967
rect 182600 538510 182660 538517
rect 182600 538476 182614 538510
rect 182648 538476 182660 538510
rect 182600 538457 182660 538476
rect 182820 538483 182841 538517
rect 182875 538483 183033 538517
rect 183067 538483 183225 538517
rect 183259 538483 183417 538517
rect 183451 538483 183609 538517
rect 183643 538483 183801 538517
rect 183835 538483 184070 538517
rect 182820 538457 184070 538483
rect 184260 538586 184270 538607
rect 184304 538607 184310 539074
rect 184352 539074 184398 539086
rect 184352 538607 184358 539074
rect 184304 538586 184358 538607
rect 184392 538586 184398 539074
rect 184260 538574 184398 538586
rect 184260 538510 184380 538574
rect 184260 538477 184314 538510
rect 184300 538476 184314 538477
rect 184348 538477 184380 538510
rect 184348 538476 184360 538477
rect 184300 538457 184360 538476
rect 182180 537847 182260 537963
rect 182254 537566 182260 537847
rect 182298 537847 182380 537963
rect 182298 537566 182304 537847
rect 182254 537554 182304 537566
rect 182254 537288 182304 537300
rect 182254 537117 182260 537288
rect 182130 536891 182260 537117
rect 182298 537117 182304 537288
rect 182298 536891 182430 537117
rect 182130 536317 182430 536891
rect 182130 536057 182190 536317
rect 182390 536057 182430 536317
rect 182130 536017 182430 536057
rect 184970 533587 185170 540727
rect 185880 540562 185886 540917
rect 185920 540917 185974 541050
rect 185920 540562 185926 540917
rect 185880 540550 185926 540562
rect 185968 540562 185974 540917
rect 186008 540997 186020 541050
rect 186179 541057 186225 541069
rect 186371 541057 186417 541069
rect 186563 541057 186609 541069
rect 186755 541057 186801 541069
rect 186947 541057 186993 541069
rect 187139 541057 187185 541069
rect 186179 540997 186185 541057
rect 186008 540917 186185 540997
rect 186008 540562 186014 540917
rect 185968 540550 186014 540562
rect 186083 540603 186129 540615
rect 186083 540317 186089 540603
rect 186050 540115 186089 540317
rect 186123 540317 186129 540603
rect 186179 540569 186185 540917
rect 186219 540667 186377 541057
rect 186219 540569 186225 540667
rect 186179 540557 186225 540569
rect 186275 540603 186321 540615
rect 186275 540317 186281 540603
rect 186123 540115 186281 540317
rect 186315 540317 186321 540603
rect 186371 540569 186377 540667
rect 186411 540667 186569 541057
rect 186411 540569 186417 540667
rect 186371 540557 186417 540569
rect 186467 540603 186513 540615
rect 186467 540317 186473 540603
rect 186315 540115 186473 540317
rect 186507 540317 186513 540603
rect 186563 540569 186569 540667
rect 186603 540667 186761 541057
rect 186603 540569 186609 540667
rect 186563 540557 186609 540569
rect 186659 540603 186705 540615
rect 186659 540317 186665 540603
rect 186507 540115 186665 540317
rect 186699 540317 186705 540603
rect 186755 540569 186761 540667
rect 186795 540667 186953 541057
rect 186795 540569 186801 540667
rect 186755 540557 186801 540569
rect 186851 540603 186897 540615
rect 186851 540317 186857 540603
rect 186699 540115 186857 540317
rect 186891 540317 186897 540603
rect 186947 540569 186953 540667
rect 186987 541027 187145 541057
rect 187179 541027 187210 541057
rect 186987 540927 187090 541027
rect 187200 540927 187210 541027
rect 186987 540907 187145 540927
rect 187179 540907 187210 540927
rect 186987 540807 187090 540907
rect 187200 540807 187210 540907
rect 187405 540862 187455 541112
rect 187598 541151 187660 541157
rect 187598 541117 187610 541151
rect 187644 541117 187660 541151
rect 187598 541111 187660 541117
rect 187600 541097 187660 541111
rect 188780 540997 188980 541537
rect 189220 541157 189280 541167
rect 189520 541162 190540 541187
rect 189520 541158 190755 541162
rect 189180 541151 189320 541157
rect 189180 541117 189230 541151
rect 189264 541117 189320 541151
rect 189520 541127 189533 541158
rect 189521 541124 189533 541127
rect 189567 541127 189725 541158
rect 189567 541124 189579 541127
rect 189521 541118 189579 541124
rect 189713 541124 189725 541127
rect 189759 541127 189917 541158
rect 189759 541124 189771 541127
rect 189713 541118 189771 541124
rect 189905 541124 189917 541127
rect 189951 541127 190109 541158
rect 189951 541124 189963 541127
rect 189905 541118 189963 541124
rect 190097 541124 190109 541127
rect 190143 541127 190301 541158
rect 190143 541124 190155 541127
rect 190097 541118 190155 541124
rect 190289 541124 190301 541127
rect 190335 541127 190493 541158
rect 190335 541124 190347 541127
rect 190289 541118 190347 541124
rect 190481 541124 190493 541127
rect 190527 541124 190755 541158
rect 190481 541118 190755 541124
rect 189180 541050 189320 541117
rect 190525 541112 190755 541118
rect 189180 540997 189186 541050
rect 187880 540862 188400 540927
rect 188780 540917 189186 540997
rect 188780 540867 188980 540917
rect 186987 540787 187145 540807
rect 187179 540787 187210 540807
rect 186987 540687 187090 540787
rect 187200 540687 187210 540787
rect 186987 540667 187145 540687
rect 186987 540569 186993 540667
rect 186947 540557 186993 540569
rect 187043 540603 187089 540615
rect 187043 540317 187049 540603
rect 186891 540115 187049 540317
rect 187083 540317 187089 540603
rect 187139 540569 187145 540667
rect 187179 540667 187210 540687
rect 187400 540812 188400 540862
rect 187179 540569 187185 540667
rect 187139 540557 187185 540569
rect 187235 540603 187281 540615
rect 187235 540317 187241 540603
rect 187083 540115 187241 540317
rect 187275 540115 187281 540603
rect 187400 540367 187450 540812
rect 187880 540727 188400 540812
rect 187560 540596 187606 540608
rect 187400 540357 187460 540367
rect 187398 540351 187460 540357
rect 187398 540317 187410 540351
rect 187444 540317 187460 540351
rect 187398 540311 187460 540317
rect 187400 540307 187460 540311
rect 187360 540267 187406 540279
rect 187360 540187 187366 540267
rect 186050 540107 187281 540115
rect 186050 540103 186129 540107
rect 186275 540103 186321 540107
rect 186467 540103 186513 540107
rect 186659 540103 186705 540107
rect 186851 540103 186897 540107
rect 187043 540103 187089 540107
rect 187235 540103 187281 540107
rect 186050 540097 186120 540103
rect 185910 540041 185980 540057
rect 185910 540007 185930 540041
rect 185964 540007 185980 540041
rect 185910 539987 185980 540007
rect 186050 539787 186080 540097
rect 187340 540091 187366 540187
rect 187400 540091 187406 540267
rect 187340 540079 187406 540091
rect 187448 540267 187494 540279
rect 187448 540091 187454 540267
rect 187488 540257 187494 540267
rect 187560 540257 187566 540596
rect 187488 540108 187566 540257
rect 187600 540267 187606 540596
rect 187648 540596 187694 540608
rect 187648 540267 187654 540596
rect 187600 540108 187654 540267
rect 187688 540267 187694 540596
rect 187870 540277 188090 540287
rect 187688 540257 187710 540267
rect 187870 540257 187900 540277
rect 187688 540247 187900 540257
rect 187688 540117 187770 540247
rect 187830 540117 187900 540247
rect 187688 540108 187900 540117
rect 187488 540107 187900 540108
rect 187488 540091 187494 540107
rect 187560 540096 187694 540107
rect 187870 540097 187900 540107
rect 188080 540097 188090 540277
rect 187448 540079 187494 540091
rect 186125 540048 186183 540054
rect 186125 540047 186137 540048
rect 186120 540014 186137 540047
rect 186171 540047 186183 540048
rect 186317 540048 186375 540054
rect 186317 540047 186329 540048
rect 186171 540014 186329 540047
rect 186363 540047 186375 540048
rect 186509 540048 186567 540054
rect 186509 540047 186521 540048
rect 186363 540014 186521 540047
rect 186555 540047 186567 540048
rect 186701 540048 186759 540054
rect 186701 540047 186713 540048
rect 186555 540014 186713 540047
rect 186747 540047 186759 540048
rect 186893 540048 186951 540054
rect 186893 540047 186905 540048
rect 186747 540014 186905 540047
rect 186939 540047 186951 540048
rect 187085 540048 187143 540054
rect 187085 540047 187097 540048
rect 186939 540014 187097 540047
rect 187131 540014 187143 540048
rect 186120 540008 187143 540014
rect 186120 539987 187140 540008
rect 185480 539687 186080 539787
rect 185480 537963 185680 539687
rect 185840 539638 186080 539687
rect 185840 539604 185914 539638
rect 185948 539604 186080 539638
rect 185840 539545 186080 539604
rect 186220 539651 187230 539657
rect 186220 539645 187243 539651
rect 186220 539611 186237 539645
rect 186271 539611 186429 539645
rect 186463 539611 186621 539645
rect 186655 539611 186813 539645
rect 186847 539611 187005 539645
rect 187039 539611 187197 539645
rect 187231 539611 187243 539645
rect 186220 539605 187243 539611
rect 186220 539597 187230 539605
rect 187340 539557 187370 540079
rect 187398 540041 187460 540047
rect 187398 540007 187410 540041
rect 187444 540007 187460 540041
rect 187398 540001 187460 540007
rect 187400 539638 187460 540001
rect 187570 540041 187690 540096
rect 187870 540087 188090 540097
rect 187570 540007 187610 540041
rect 187644 540007 187690 540041
rect 187570 539987 187690 540007
rect 187400 539604 187414 539638
rect 187448 539604 187460 539638
rect 187400 539597 187460 539604
rect 187600 539638 187680 539657
rect 187600 539604 187614 539638
rect 187648 539604 187680 539638
rect 187600 539597 187680 539604
rect 185840 539447 185870 539545
rect 185864 538569 185870 539447
rect 185904 539447 185958 539545
rect 185904 538569 185910 539447
rect 185864 538557 185910 538569
rect 185952 538569 185958 539447
rect 185992 539527 186080 539545
rect 186183 539535 186229 539547
rect 185992 539517 186150 539527
rect 186183 539517 186189 539535
rect 185992 539447 186189 539517
rect 185992 538569 185998 539447
rect 186050 539237 186189 539447
rect 186087 539081 186133 539093
rect 186087 538593 186093 539081
rect 186127 538967 186133 539081
rect 186183 539047 186189 539237
rect 186223 539517 186229 539535
rect 186375 539535 186421 539547
rect 186375 539517 186381 539535
rect 186223 539237 186381 539517
rect 186223 539047 186229 539237
rect 186183 539035 186229 539047
rect 186279 539081 186325 539093
rect 186279 538967 186285 539081
rect 186127 538593 186285 538967
rect 186319 538967 186325 539081
rect 186375 539047 186381 539237
rect 186415 539517 186421 539535
rect 186567 539535 186613 539547
rect 186567 539517 186573 539535
rect 186415 539237 186573 539517
rect 186415 539047 186421 539237
rect 186375 539035 186421 539047
rect 186471 539081 186517 539093
rect 186471 538967 186477 539081
rect 186319 538593 186477 538967
rect 186511 538967 186517 539081
rect 186567 539047 186573 539237
rect 186607 539517 186613 539535
rect 186759 539535 186805 539547
rect 186759 539517 186765 539535
rect 186607 539237 186765 539517
rect 186607 539047 186613 539237
rect 186567 539035 186613 539047
rect 186663 539081 186709 539093
rect 186663 538967 186669 539081
rect 186511 538593 186669 538967
rect 186703 538967 186709 539081
rect 186759 539047 186765 539237
rect 186799 539517 186805 539535
rect 186951 539535 186997 539547
rect 186951 539517 186957 539535
rect 186799 539237 186957 539517
rect 186799 539047 186805 539237
rect 186759 539035 186805 539047
rect 186855 539081 186901 539093
rect 186855 538967 186861 539081
rect 186703 538593 186861 538967
rect 186895 538967 186901 539081
rect 186951 539047 186957 539237
rect 186991 539517 186997 539535
rect 187143 539535 187189 539547
rect 187143 539517 187149 539535
rect 186991 539237 187149 539517
rect 186991 539047 186997 539237
rect 186951 539035 186997 539047
rect 187047 539081 187093 539093
rect 187047 538967 187053 539081
rect 186895 538593 187053 538967
rect 187087 538967 187093 539081
rect 187143 539047 187149 539237
rect 187183 539517 187189 539535
rect 187340 539545 187410 539557
rect 187183 539237 187200 539517
rect 187340 539407 187370 539545
rect 187183 539047 187189 539237
rect 187143 539035 187189 539047
rect 187239 539081 187285 539093
rect 187239 538967 187245 539081
rect 187087 538837 187245 538967
rect 187087 538737 187100 538837
rect 187240 538737 187245 538837
rect 187087 538593 187245 538737
rect 187279 538593 187285 539081
rect 187364 539067 187370 539407
rect 186087 538587 187285 538593
rect 186087 538581 186133 538587
rect 186279 538581 186325 538587
rect 186471 538581 186517 538587
rect 186663 538581 186709 538587
rect 186855 538581 186901 538587
rect 187047 538581 187093 538587
rect 187239 538581 187285 538587
rect 187330 538969 187370 539067
rect 187404 538969 187410 539545
rect 187330 538957 187410 538969
rect 187452 539545 187498 539557
rect 187452 538969 187458 539545
rect 187492 539537 187498 539545
rect 187492 539307 187610 539537
rect 187870 539337 188090 539347
rect 187870 539307 187890 539337
rect 187492 539297 187890 539307
rect 187492 539207 187770 539297
rect 187820 539207 187890 539297
rect 187492 539197 187890 539207
rect 187492 539074 187610 539197
rect 187870 539157 187890 539197
rect 188070 539157 188090 539337
rect 187870 539147 188090 539157
rect 187492 538969 187570 539074
rect 187452 538967 187570 538969
rect 187452 538957 187498 538967
rect 185952 538557 185998 538569
rect 186129 538517 186187 538523
rect 186321 538517 186379 538523
rect 186513 538517 186571 538523
rect 186705 538517 186763 538523
rect 186897 538517 186955 538523
rect 187089 538517 187147 538523
rect 187330 538517 187370 538957
rect 187400 538910 187460 538917
rect 187400 538876 187414 538910
rect 187448 538876 187460 538910
rect 187400 538857 187460 538876
rect 187564 538607 187570 538967
rect 185900 538510 185960 538517
rect 185900 538476 185914 538510
rect 185948 538476 185960 538510
rect 185900 538457 185960 538476
rect 186120 538483 186141 538517
rect 186175 538483 186333 538517
rect 186367 538483 186525 538517
rect 186559 538483 186717 538517
rect 186751 538483 186909 538517
rect 186943 538483 187101 538517
rect 187135 538483 187370 538517
rect 186120 538457 187370 538483
rect 187560 538586 187570 538607
rect 187604 538607 187610 539074
rect 187652 539074 187698 539086
rect 187652 538607 187658 539074
rect 187604 538586 187658 538607
rect 187692 538586 187698 539074
rect 187560 538574 187698 538586
rect 187560 538510 187680 538574
rect 187560 538477 187614 538510
rect 187600 538476 187614 538477
rect 187648 538477 187680 538510
rect 187648 538476 187660 538477
rect 187600 538457 187660 538476
rect 185480 537847 185560 537963
rect 185554 537566 185560 537847
rect 185598 537847 185680 537963
rect 185598 537566 185604 537847
rect 185554 537554 185604 537566
rect 185554 537428 185604 537440
rect 185554 537237 185560 537428
rect 185430 537031 185560 537237
rect 185598 537237 185604 537428
rect 185598 537031 185730 537237
rect 185430 536297 185730 537031
rect 185430 536177 185490 536297
rect 185700 536177 185730 536297
rect 185430 536137 185730 536177
rect 180830 533337 181930 533537
rect 182930 533387 185170 533587
rect 178220 532767 178930 532787
rect 178220 532597 178700 532767
rect 178830 532597 178930 532767
rect 178220 532587 178930 532597
rect 180830 532767 181030 533337
rect 180830 532597 180870 532767
rect 181000 532597 181030 532767
rect 180830 532487 181030 532597
rect 182930 532767 183130 533387
rect 184970 533337 185170 533387
rect 188200 533287 188400 540727
rect 189180 540562 189186 540917
rect 189220 540917 189274 541050
rect 189220 540562 189226 540917
rect 189180 540550 189226 540562
rect 189268 540562 189274 540917
rect 189308 540997 189320 541050
rect 189479 541057 189525 541069
rect 189671 541057 189717 541069
rect 189863 541057 189909 541069
rect 190055 541057 190101 541069
rect 190247 541057 190293 541069
rect 190439 541057 190485 541069
rect 189479 540997 189485 541057
rect 189308 540917 189485 540997
rect 189308 540562 189314 540917
rect 189268 540550 189314 540562
rect 189383 540603 189429 540615
rect 189383 540317 189389 540603
rect 189350 540115 189389 540317
rect 189423 540317 189429 540603
rect 189479 540569 189485 540917
rect 189519 540667 189677 541057
rect 189519 540569 189525 540667
rect 189479 540557 189525 540569
rect 189575 540603 189621 540615
rect 189575 540317 189581 540603
rect 189423 540115 189581 540317
rect 189615 540317 189621 540603
rect 189671 540569 189677 540667
rect 189711 540667 189869 541057
rect 189711 540569 189717 540667
rect 189671 540557 189717 540569
rect 189767 540603 189813 540615
rect 189767 540317 189773 540603
rect 189615 540115 189773 540317
rect 189807 540317 189813 540603
rect 189863 540569 189869 540667
rect 189903 540667 190061 541057
rect 189903 540569 189909 540667
rect 189863 540557 189909 540569
rect 189959 540603 190005 540615
rect 189959 540317 189965 540603
rect 189807 540115 189965 540317
rect 189999 540317 190005 540603
rect 190055 540569 190061 540667
rect 190095 540667 190253 541057
rect 190095 540569 190101 540667
rect 190055 540557 190101 540569
rect 190151 540603 190197 540615
rect 190151 540317 190157 540603
rect 189999 540115 190157 540317
rect 190191 540317 190197 540603
rect 190247 540569 190253 540667
rect 190287 541027 190445 541057
rect 190479 541027 190510 541057
rect 190287 540927 190390 541027
rect 190500 540927 190510 541027
rect 190287 540907 190445 540927
rect 190479 540907 190510 540927
rect 190287 540807 190390 540907
rect 190500 540807 190510 540907
rect 190705 540862 190755 541112
rect 190898 541151 190960 541157
rect 190898 541117 190910 541151
rect 190944 541117 190960 541151
rect 190898 541111 190960 541117
rect 190900 541097 190960 541111
rect 191180 540862 191680 540927
rect 190287 540787 190445 540807
rect 190479 540787 190510 540807
rect 190287 540687 190390 540787
rect 190500 540687 190510 540787
rect 190287 540667 190445 540687
rect 190287 540569 190293 540667
rect 190247 540557 190293 540569
rect 190343 540603 190389 540615
rect 190343 540317 190349 540603
rect 190191 540115 190349 540317
rect 190383 540317 190389 540603
rect 190439 540569 190445 540667
rect 190479 540667 190510 540687
rect 190700 540812 191680 540862
rect 190479 540569 190485 540667
rect 190439 540557 190485 540569
rect 190535 540603 190581 540615
rect 190535 540317 190541 540603
rect 190383 540115 190541 540317
rect 190575 540115 190581 540603
rect 190700 540367 190750 540812
rect 191180 540727 191680 540812
rect 190860 540596 190906 540608
rect 190700 540357 190760 540367
rect 190698 540351 190760 540357
rect 190698 540317 190710 540351
rect 190744 540317 190760 540351
rect 190698 540311 190760 540317
rect 190700 540307 190760 540311
rect 190660 540267 190706 540279
rect 190660 540187 190666 540267
rect 189350 540107 190581 540115
rect 189350 540103 189429 540107
rect 189575 540103 189621 540107
rect 189767 540103 189813 540107
rect 189959 540103 190005 540107
rect 190151 540103 190197 540107
rect 190343 540103 190389 540107
rect 190535 540103 190581 540107
rect 189350 540097 189420 540103
rect 189210 540041 189280 540057
rect 189210 540007 189230 540041
rect 189264 540007 189280 540041
rect 189210 539987 189280 540007
rect 189350 539787 189380 540097
rect 190640 540091 190666 540187
rect 190700 540091 190706 540267
rect 190640 540079 190706 540091
rect 190748 540267 190794 540279
rect 190748 540091 190754 540267
rect 190788 540257 190794 540267
rect 190860 540257 190866 540596
rect 190788 540108 190866 540257
rect 190900 540267 190906 540596
rect 190948 540596 190994 540608
rect 190948 540267 190954 540596
rect 190900 540108 190954 540267
rect 190988 540267 190994 540596
rect 191170 540277 191390 540287
rect 190988 540257 191010 540267
rect 191170 540257 191190 540277
rect 190988 540247 191190 540257
rect 190988 540117 191070 540247
rect 191130 540117 191190 540247
rect 190988 540108 191190 540117
rect 190788 540107 191190 540108
rect 190788 540091 190794 540107
rect 190860 540096 190994 540107
rect 191170 540097 191190 540107
rect 191370 540097 191390 540277
rect 190748 540079 190794 540091
rect 189425 540048 189483 540054
rect 189425 540047 189437 540048
rect 189420 540014 189437 540047
rect 189471 540047 189483 540048
rect 189617 540048 189675 540054
rect 189617 540047 189629 540048
rect 189471 540014 189629 540047
rect 189663 540047 189675 540048
rect 189809 540048 189867 540054
rect 189809 540047 189821 540048
rect 189663 540014 189821 540047
rect 189855 540047 189867 540048
rect 190001 540048 190059 540054
rect 190001 540047 190013 540048
rect 189855 540014 190013 540047
rect 190047 540047 190059 540048
rect 190193 540048 190251 540054
rect 190193 540047 190205 540048
rect 190047 540014 190205 540047
rect 190239 540047 190251 540048
rect 190385 540048 190443 540054
rect 190385 540047 190397 540048
rect 190239 540014 190397 540047
rect 190431 540014 190443 540048
rect 189420 540008 190443 540014
rect 189420 539987 190440 540008
rect 188780 539687 189380 539787
rect 188780 537963 188980 539687
rect 189140 539638 189380 539687
rect 189140 539604 189214 539638
rect 189248 539604 189380 539638
rect 189140 539545 189380 539604
rect 189520 539651 190530 539657
rect 189520 539645 190543 539651
rect 189520 539611 189537 539645
rect 189571 539611 189729 539645
rect 189763 539611 189921 539645
rect 189955 539611 190113 539645
rect 190147 539611 190305 539645
rect 190339 539611 190497 539645
rect 190531 539611 190543 539645
rect 189520 539605 190543 539611
rect 189520 539597 190530 539605
rect 190640 539557 190670 540079
rect 190698 540041 190760 540047
rect 190698 540007 190710 540041
rect 190744 540007 190760 540041
rect 190698 540001 190760 540007
rect 190700 539638 190760 540001
rect 190870 540041 190990 540096
rect 191170 540087 191390 540097
rect 190870 540007 190910 540041
rect 190944 540007 190990 540041
rect 190870 539987 190990 540007
rect 190700 539604 190714 539638
rect 190748 539604 190760 539638
rect 190700 539597 190760 539604
rect 190900 539638 190980 539657
rect 190900 539604 190914 539638
rect 190948 539604 190980 539638
rect 190900 539597 190980 539604
rect 189140 539447 189170 539545
rect 189164 538569 189170 539447
rect 189204 539447 189258 539545
rect 189204 538569 189210 539447
rect 189164 538557 189210 538569
rect 189252 538569 189258 539447
rect 189292 539527 189380 539545
rect 189483 539535 189529 539547
rect 189292 539517 189450 539527
rect 189483 539517 189489 539535
rect 189292 539447 189489 539517
rect 189292 538569 189298 539447
rect 189350 539237 189489 539447
rect 189387 539081 189433 539093
rect 189387 538593 189393 539081
rect 189427 538967 189433 539081
rect 189483 539047 189489 539237
rect 189523 539517 189529 539535
rect 189675 539535 189721 539547
rect 189675 539517 189681 539535
rect 189523 539237 189681 539517
rect 189523 539047 189529 539237
rect 189483 539035 189529 539047
rect 189579 539081 189625 539093
rect 189579 538967 189585 539081
rect 189427 538593 189585 538967
rect 189619 538967 189625 539081
rect 189675 539047 189681 539237
rect 189715 539517 189721 539535
rect 189867 539535 189913 539547
rect 189867 539517 189873 539535
rect 189715 539237 189873 539517
rect 189715 539047 189721 539237
rect 189675 539035 189721 539047
rect 189771 539081 189817 539093
rect 189771 538967 189777 539081
rect 189619 538593 189777 538967
rect 189811 538967 189817 539081
rect 189867 539047 189873 539237
rect 189907 539517 189913 539535
rect 190059 539535 190105 539547
rect 190059 539517 190065 539535
rect 189907 539237 190065 539517
rect 189907 539047 189913 539237
rect 189867 539035 189913 539047
rect 189963 539081 190009 539093
rect 189963 538967 189969 539081
rect 189811 538593 189969 538967
rect 190003 538967 190009 539081
rect 190059 539047 190065 539237
rect 190099 539517 190105 539535
rect 190251 539535 190297 539547
rect 190251 539517 190257 539535
rect 190099 539237 190257 539517
rect 190099 539047 190105 539237
rect 190059 539035 190105 539047
rect 190155 539081 190201 539093
rect 190155 538967 190161 539081
rect 190003 538593 190161 538967
rect 190195 538967 190201 539081
rect 190251 539047 190257 539237
rect 190291 539517 190297 539535
rect 190443 539535 190489 539547
rect 190443 539517 190449 539535
rect 190291 539237 190449 539517
rect 190291 539047 190297 539237
rect 190251 539035 190297 539047
rect 190347 539081 190393 539093
rect 190347 538967 190353 539081
rect 190195 538593 190353 538967
rect 190387 538967 190393 539081
rect 190443 539047 190449 539237
rect 190483 539517 190489 539535
rect 190640 539545 190710 539557
rect 190483 539237 190500 539517
rect 190640 539407 190670 539545
rect 190483 539047 190489 539237
rect 190443 539035 190489 539047
rect 190539 539081 190585 539093
rect 190539 538967 190545 539081
rect 190387 538837 190545 538967
rect 190387 538737 190400 538837
rect 190540 538737 190545 538837
rect 190387 538593 190545 538737
rect 190579 538593 190585 539081
rect 190664 539067 190670 539407
rect 189387 538587 190585 538593
rect 189387 538581 189433 538587
rect 189579 538581 189625 538587
rect 189771 538581 189817 538587
rect 189963 538581 190009 538587
rect 190155 538581 190201 538587
rect 190347 538581 190393 538587
rect 190539 538581 190585 538587
rect 190630 538969 190670 539067
rect 190704 538969 190710 539545
rect 190630 538957 190710 538969
rect 190752 539545 190798 539557
rect 190752 538969 190758 539545
rect 190792 539537 190798 539545
rect 190792 539307 190910 539537
rect 191190 539347 191390 539357
rect 191170 539307 191200 539347
rect 190792 539297 191200 539307
rect 190792 539207 191070 539297
rect 191120 539207 191200 539297
rect 190792 539197 191200 539207
rect 190792 539074 190910 539197
rect 191170 539167 191200 539197
rect 191380 539167 191390 539347
rect 191170 539147 191390 539167
rect 190792 538969 190870 539074
rect 190752 538967 190870 538969
rect 190752 538957 190798 538967
rect 189252 538557 189298 538569
rect 189429 538517 189487 538523
rect 189621 538517 189679 538523
rect 189813 538517 189871 538523
rect 190005 538517 190063 538523
rect 190197 538517 190255 538523
rect 190389 538517 190447 538523
rect 190630 538517 190670 538957
rect 190700 538910 190760 538917
rect 190700 538876 190714 538910
rect 190748 538876 190760 538910
rect 190700 538857 190760 538876
rect 190864 538607 190870 538967
rect 189200 538510 189260 538517
rect 189200 538476 189214 538510
rect 189248 538476 189260 538510
rect 189200 538457 189260 538476
rect 189420 538483 189441 538517
rect 189475 538483 189633 538517
rect 189667 538483 189825 538517
rect 189859 538483 190017 538517
rect 190051 538483 190209 538517
rect 190243 538483 190401 538517
rect 190435 538483 190670 538517
rect 189420 538457 190670 538483
rect 190860 538586 190870 538607
rect 190904 538607 190910 539074
rect 190952 539074 190998 539086
rect 190952 538607 190958 539074
rect 190904 538586 190958 538607
rect 190992 538586 190998 539074
rect 190860 538574 190998 538586
rect 190860 538510 190980 538574
rect 190860 538477 190914 538510
rect 190900 538476 190914 538477
rect 190948 538477 190980 538510
rect 190948 538476 190960 538477
rect 190900 538457 190960 538476
rect 188780 537847 188860 537963
rect 188854 537566 188860 537847
rect 188898 537847 188980 537963
rect 188898 537566 188904 537847
rect 188854 537554 188904 537566
rect 188854 537332 188904 537344
rect 188854 537137 188860 537332
rect 188730 536935 188860 537137
rect 188898 537137 188904 537332
rect 188898 536935 189030 537137
rect 188730 536307 189030 536935
rect 188730 536067 188780 536307
rect 189000 536067 189030 536307
rect 188730 536037 189030 536067
rect 182930 532597 182960 532767
rect 183090 532597 183130 532767
rect 182930 532487 183130 532597
rect 185030 533087 188400 533287
rect 185030 532807 185230 533087
rect 185030 532637 185060 532807
rect 185190 532637 185230 532807
rect 191480 532787 191680 540727
rect 193000 540296 195000 542036
rect 192630 540287 195000 540296
rect 191750 540277 195000 540287
rect 191750 540097 191810 540277
rect 191990 540097 195000 540277
rect 191750 540087 192230 540097
rect 192430 540087 195000 540097
rect 192630 540086 195000 540087
rect 193000 540036 195000 540086
rect 192630 539347 195000 539356
rect 191810 539337 195000 539347
rect 191810 539157 191820 539337
rect 192000 539157 195000 539337
rect 191810 539147 195000 539157
rect 192630 539146 195000 539147
rect 193000 537356 195000 539146
rect 185030 532587 185230 532637
rect 187130 532767 191680 532787
rect 187130 532627 187170 532767
rect 187270 532627 191680 532767
rect 187130 532587 191680 532627
rect 172210 530637 187482 530659
rect 172210 530628 174625 530637
rect 172210 530594 172239 530628
rect 172273 530594 172331 530628
rect 172365 530594 172423 530628
rect 172457 530594 172515 530628
rect 172549 530594 172607 530628
rect 172641 530594 172699 530628
rect 172733 530594 172791 530628
rect 172825 530594 172883 530628
rect 172917 530594 172975 530628
rect 173009 530594 173067 530628
rect 173101 530594 173159 530628
rect 173193 530594 173251 530628
rect 173285 530594 173343 530628
rect 173377 530594 173435 530628
rect 173469 530594 173527 530628
rect 173561 530594 173619 530628
rect 173653 530594 173711 530628
rect 173745 530594 173803 530628
rect 173837 530594 173895 530628
rect 173929 530594 173987 530628
rect 174021 530594 174079 530628
rect 174113 530594 174171 530628
rect 174205 530594 174263 530628
rect 174297 530594 174355 530628
rect 174389 530594 174447 530628
rect 174481 530594 174539 530628
rect 174573 530594 174625 530628
rect 172210 530585 174625 530594
rect 174677 530585 174689 530637
rect 174741 530628 174753 530637
rect 174805 530628 174817 530637
rect 174805 530594 174815 530628
rect 174741 530585 174753 530594
rect 174805 530585 174817 530594
rect 174869 530585 174881 530637
rect 174933 530628 178443 530637
rect 174941 530594 174999 530628
rect 175033 530594 175091 530628
rect 175125 530594 175183 530628
rect 175217 530594 175275 530628
rect 175309 530594 175367 530628
rect 175401 530594 175459 530628
rect 175493 530594 175551 530628
rect 175585 530594 175643 530628
rect 175677 530594 175735 530628
rect 175769 530594 175827 530628
rect 175861 530594 175919 530628
rect 175953 530594 176011 530628
rect 176045 530594 176103 530628
rect 176137 530594 176195 530628
rect 176229 530594 176287 530628
rect 176321 530594 176379 530628
rect 176413 530594 176471 530628
rect 176505 530594 176563 530628
rect 176597 530594 176655 530628
rect 176689 530594 176747 530628
rect 176781 530594 176839 530628
rect 176873 530594 176931 530628
rect 176965 530594 177023 530628
rect 177057 530594 177115 530628
rect 177149 530594 177207 530628
rect 177241 530594 177299 530628
rect 177333 530594 177391 530628
rect 177425 530594 177483 530628
rect 177517 530594 177575 530628
rect 177609 530594 177667 530628
rect 177701 530594 177759 530628
rect 177793 530594 177851 530628
rect 177885 530594 177943 530628
rect 177977 530594 178035 530628
rect 178069 530594 178127 530628
rect 178161 530594 178219 530628
rect 178253 530594 178311 530628
rect 178345 530594 178403 530628
rect 178437 530594 178443 530628
rect 174933 530585 178443 530594
rect 178495 530628 178507 530637
rect 178495 530585 178507 530594
rect 178559 530585 178571 530637
rect 178623 530585 178635 530637
rect 178687 530628 178699 530637
rect 178751 530628 182261 530637
rect 178751 530594 178771 530628
rect 178805 530594 178863 530628
rect 178897 530594 178955 530628
rect 178989 530594 179047 530628
rect 179081 530594 179139 530628
rect 179173 530594 179231 530628
rect 179265 530594 179323 530628
rect 179357 530594 179415 530628
rect 179449 530594 179507 530628
rect 179541 530594 179599 530628
rect 179633 530594 179691 530628
rect 179725 530594 179783 530628
rect 179817 530594 179875 530628
rect 179909 530594 179967 530628
rect 180001 530594 180059 530628
rect 180093 530594 180151 530628
rect 180185 530594 180243 530628
rect 180277 530594 180335 530628
rect 180369 530594 180427 530628
rect 180461 530594 180519 530628
rect 180553 530594 180611 530628
rect 180645 530594 180703 530628
rect 180737 530594 180795 530628
rect 180829 530594 180887 530628
rect 180921 530594 180979 530628
rect 181013 530594 181071 530628
rect 181105 530594 181163 530628
rect 181197 530594 181255 530628
rect 181289 530594 181347 530628
rect 181381 530594 181439 530628
rect 181473 530594 181531 530628
rect 181565 530594 181623 530628
rect 181657 530594 181715 530628
rect 181749 530594 181807 530628
rect 181841 530594 181899 530628
rect 181933 530594 181991 530628
rect 182025 530594 182083 530628
rect 182117 530594 182175 530628
rect 182209 530594 182261 530628
rect 178687 530585 178699 530594
rect 178751 530585 182261 530594
rect 182313 530585 182325 530637
rect 182377 530628 182389 530637
rect 182441 530628 182453 530637
rect 182441 530594 182451 530628
rect 182377 530585 182389 530594
rect 182441 530585 182453 530594
rect 182505 530585 182517 530637
rect 182569 530628 186079 530637
rect 182577 530594 182635 530628
rect 182669 530594 182727 530628
rect 182761 530594 182819 530628
rect 182853 530594 182911 530628
rect 182945 530594 183003 530628
rect 183037 530594 183095 530628
rect 183129 530594 183187 530628
rect 183221 530594 183279 530628
rect 183313 530594 183371 530628
rect 183405 530594 183463 530628
rect 183497 530594 183555 530628
rect 183589 530594 183647 530628
rect 183681 530594 183739 530628
rect 183773 530594 183831 530628
rect 183865 530594 183923 530628
rect 183957 530594 184015 530628
rect 184049 530594 184107 530628
rect 184141 530594 184199 530628
rect 184233 530594 184291 530628
rect 184325 530594 184383 530628
rect 184417 530594 184475 530628
rect 184509 530594 184567 530628
rect 184601 530594 184659 530628
rect 184693 530594 184751 530628
rect 184785 530594 184843 530628
rect 184877 530594 184935 530628
rect 184969 530594 185027 530628
rect 185061 530594 185119 530628
rect 185153 530594 185211 530628
rect 185245 530594 185303 530628
rect 185337 530594 185395 530628
rect 185429 530594 185487 530628
rect 185521 530594 185579 530628
rect 185613 530594 185671 530628
rect 185705 530594 185763 530628
rect 185797 530594 185855 530628
rect 185889 530594 185947 530628
rect 185981 530594 186039 530628
rect 186073 530594 186079 530628
rect 182569 530585 186079 530594
rect 186131 530628 186143 530637
rect 186131 530585 186143 530594
rect 186195 530585 186207 530637
rect 186259 530585 186271 530637
rect 186323 530628 186335 530637
rect 186387 530628 187482 530637
rect 186387 530594 186407 530628
rect 186441 530594 186499 530628
rect 186533 530594 186591 530628
rect 186625 530594 186683 530628
rect 186717 530594 186775 530628
rect 186809 530594 186867 530628
rect 186901 530594 186959 530628
rect 186993 530594 187051 530628
rect 187085 530594 187143 530628
rect 187177 530594 187235 530628
rect 187269 530594 187327 530628
rect 187361 530594 187419 530628
rect 187453 530594 187482 530628
rect 186323 530585 186335 530594
rect 186387 530585 187482 530594
rect 172210 530563 187482 530585
rect 176824 530523 176830 530535
rect 176658 530495 176830 530523
rect 172408 530415 172414 530467
rect 172466 530455 172472 530467
rect 172503 530458 172561 530464
rect 172503 530455 172515 530458
rect 172466 530427 172515 530455
rect 172466 530415 172472 530427
rect 172503 530424 172515 530427
rect 172549 530424 172561 530458
rect 172503 530418 172561 530424
rect 174524 530415 174530 530467
rect 174582 530455 174588 530467
rect 174895 530458 174953 530464
rect 174895 530455 174907 530458
rect 174582 530427 174907 530455
rect 174582 530415 174588 530427
rect 174895 530424 174907 530427
rect 174941 530424 174953 530458
rect 174895 530418 174953 530424
rect 175835 530458 175893 530464
rect 175835 530424 175847 530458
rect 175881 530455 175893 530458
rect 176483 530458 176613 530464
rect 176483 530455 176495 530458
rect 175881 530427 176495 530455
rect 175881 530424 175953 530427
rect 175835 530418 175953 530424
rect 176483 530424 176495 530427
rect 176529 530424 176567 530458
rect 176601 530455 176613 530458
rect 176658 530455 176686 530495
rect 176824 530483 176830 530495
rect 176882 530483 176888 530535
rect 178756 530483 178762 530535
rect 178814 530483 178820 530535
rect 179403 530526 179461 530532
rect 179403 530523 179415 530526
rect 178866 530495 179415 530523
rect 176601 530427 176686 530455
rect 176601 530424 176613 530427
rect 176483 530418 176613 530424
rect 172871 530390 172929 530396
rect 172871 530356 172883 530390
rect 172917 530387 172929 530390
rect 174800 530387 174806 530399
rect 172917 530359 174806 530387
rect 172917 530356 172929 530359
rect 172871 530350 172929 530356
rect 174800 530347 174806 530359
rect 174858 530347 174864 530399
rect 175263 530390 175321 530396
rect 175263 530356 175275 530390
rect 175309 530387 175321 530390
rect 175444 530387 175450 530399
rect 175309 530359 175450 530387
rect 175309 530356 175321 530359
rect 175263 530350 175321 530356
rect 175444 530347 175450 530359
rect 175502 530347 175508 530399
rect 175895 530395 175953 530418
rect 176732 530415 176738 530467
rect 176790 530455 176796 530467
rect 178866 530455 178894 530495
rect 179403 530492 179415 530495
rect 179449 530492 179461 530526
rect 179403 530486 179461 530492
rect 179492 530483 179498 530535
rect 179550 530523 179556 530535
rect 180691 530526 180749 530532
rect 180691 530523 180703 530526
rect 179550 530495 180703 530523
rect 179550 530483 179556 530495
rect 180691 530492 180703 530495
rect 180737 530492 180749 530526
rect 180691 530486 180749 530492
rect 176790 530427 178894 530455
rect 180706 530455 180734 530486
rect 182988 530483 182994 530535
rect 183046 530523 183052 530535
rect 183267 530526 183325 530532
rect 183267 530523 183279 530526
rect 183046 530495 183279 530523
rect 183046 530483 183052 530495
rect 183267 530492 183279 530495
rect 183313 530492 183325 530526
rect 183267 530486 183325 530492
rect 185104 530483 185110 530535
rect 185162 530523 185168 530535
rect 185383 530526 185441 530532
rect 185383 530523 185395 530526
rect 185162 530495 185395 530523
rect 185162 530483 185168 530495
rect 185383 530492 185395 530495
rect 185429 530492 185441 530526
rect 185383 530486 185441 530492
rect 182071 530458 182129 530464
rect 182071 530455 182083 530458
rect 180706 530427 182083 530455
rect 176790 530415 176796 530427
rect 182071 530424 182083 530427
rect 182117 530424 182129 530458
rect 185291 530458 185349 530464
rect 185291 530455 185303 530458
rect 182071 530418 182129 530424
rect 182638 530427 185303 530455
rect 175895 530361 175907 530395
rect 175941 530361 175953 530395
rect 175895 530355 175953 530361
rect 176111 530390 176169 530396
rect 176111 530356 176123 530390
rect 176157 530387 176169 530390
rect 176827 530390 176885 530396
rect 176827 530387 176839 530390
rect 176157 530359 176839 530387
rect 176157 530356 176169 530359
rect 176111 530350 176169 530356
rect 176827 530356 176839 530359
rect 176873 530387 176885 530390
rect 177194 530390 177252 530396
rect 177194 530387 177206 530390
rect 176873 530359 177206 530387
rect 176873 530356 176885 530359
rect 176827 530350 176885 530356
rect 177194 530356 177206 530359
rect 177240 530356 177252 530390
rect 177194 530350 177252 530356
rect 178575 530390 178633 530396
rect 178575 530356 178587 530390
rect 178621 530387 178633 530390
rect 178940 530387 178946 530399
rect 178621 530359 178946 530387
rect 178621 530356 178633 530359
rect 178575 530350 178633 530356
rect 178940 530347 178946 530359
rect 178998 530347 179004 530399
rect 179035 530390 179093 530396
rect 179035 530356 179047 530390
rect 179081 530387 179093 530390
rect 179216 530387 179222 530399
rect 179081 530359 179222 530387
rect 179081 530356 179093 530359
rect 179035 530350 179093 530356
rect 179216 530347 179222 530359
rect 179274 530347 179280 530399
rect 179311 530390 179369 530396
rect 179311 530356 179323 530390
rect 179357 530356 179369 530390
rect 179311 530350 179369 530356
rect 180599 530390 180657 530396
rect 180599 530356 180611 530390
rect 180645 530387 180657 530390
rect 181519 530390 181577 530396
rect 180645 530359 181470 530387
rect 180645 530356 180657 530359
rect 180599 530350 180657 530356
rect 174818 530319 174846 530347
rect 175539 530322 175597 530328
rect 175539 530319 175551 530322
rect 174818 530291 175551 530319
rect 175539 530288 175551 530291
rect 175585 530288 175597 530322
rect 175539 530282 175597 530288
rect 176640 530279 176646 530331
rect 176698 530319 176704 530331
rect 177011 530322 177069 530328
rect 177011 530319 177023 530322
rect 176698 530291 177023 530319
rect 176698 530279 176704 530291
rect 177011 530288 177023 530291
rect 177057 530288 177069 530322
rect 177011 530282 177069 530288
rect 177284 530279 177290 530331
rect 177342 530279 177348 530331
rect 178204 530279 178210 530331
rect 178262 530319 178268 530331
rect 179326 530319 179354 530350
rect 178262 530291 179354 530319
rect 178262 530279 178268 530291
rect 180688 530279 180694 530331
rect 180746 530319 180752 530331
rect 181442 530328 181470 530359
rect 181519 530356 181531 530390
rect 181565 530387 181577 530390
rect 182252 530387 182258 530399
rect 181565 530359 182258 530387
rect 181565 530356 181577 530359
rect 181519 530350 181577 530356
rect 182252 530347 182258 530359
rect 182310 530387 182316 530399
rect 182638 530387 182666 530427
rect 185291 530424 185303 530427
rect 185337 530424 185349 530458
rect 185291 530418 185349 530424
rect 182310 530359 182666 530387
rect 182310 530347 182316 530359
rect 183172 530347 183178 530399
rect 183230 530347 183236 530399
rect 187128 530347 187134 530399
rect 187186 530347 187192 530399
rect 180783 530322 180841 530328
rect 180783 530319 180795 530322
rect 180746 530291 180795 530319
rect 180746 530279 180752 530291
rect 180783 530288 180795 530291
rect 180829 530319 180841 530322
rect 181243 530322 181301 530328
rect 181243 530319 181255 530322
rect 180829 530291 181255 530319
rect 180829 530288 180841 530291
rect 180783 530282 180841 530288
rect 181243 530288 181255 530291
rect 181289 530288 181301 530322
rect 181243 530282 181301 530288
rect 181427 530322 181485 530328
rect 181427 530288 181439 530322
rect 181473 530319 181485 530322
rect 182620 530319 182626 530331
rect 181473 530291 182626 530319
rect 181473 530288 181485 530291
rect 181427 530282 181485 530288
rect 182620 530279 182626 530291
rect 182678 530279 182684 530331
rect 176111 530254 176169 530260
rect 176111 530220 176123 530254
rect 176157 530251 176169 530254
rect 176735 530254 176793 530260
rect 176735 530251 176747 530254
rect 176157 530223 176747 530251
rect 176157 530220 176169 530223
rect 176111 530214 176169 530220
rect 176735 530220 176747 530223
rect 176781 530251 176793 530254
rect 177113 530254 177171 530260
rect 177113 530251 177125 530254
rect 176781 530223 177125 530251
rect 176781 530220 176793 530223
rect 176735 530214 176793 530220
rect 177113 530220 177125 530223
rect 177159 530220 177171 530254
rect 177113 530214 177171 530220
rect 181887 530254 181945 530260
rect 181887 530220 181899 530254
rect 181933 530251 181945 530254
rect 181933 530223 182758 530251
rect 181933 530220 181945 530223
rect 181887 530214 181945 530220
rect 182730 530195 182758 530223
rect 177652 530143 177658 530195
rect 177710 530143 177716 530195
rect 178296 530143 178302 530195
rect 178354 530183 178360 530195
rect 178391 530186 178449 530192
rect 178391 530183 178403 530186
rect 178354 530155 178403 530183
rect 178354 530143 178360 530155
rect 178391 530152 178403 530155
rect 178437 530152 178449 530186
rect 178391 530146 178449 530152
rect 179676 530143 179682 530195
rect 179734 530183 179740 530195
rect 180231 530186 180289 530192
rect 180231 530183 180243 530186
rect 179734 530155 180243 530183
rect 179734 530143 179740 530155
rect 180231 530152 180243 530155
rect 180277 530152 180289 530186
rect 180231 530146 180289 530152
rect 182160 530143 182166 530195
rect 182218 530143 182224 530195
rect 182712 530143 182718 530195
rect 182770 530143 182776 530195
rect 172210 530093 187482 530115
rect 172210 530084 173965 530093
rect 174017 530084 174029 530093
rect 174081 530084 174093 530093
rect 172210 530050 172239 530084
rect 172273 530050 172331 530084
rect 172365 530050 172423 530084
rect 172457 530050 172515 530084
rect 172549 530050 172607 530084
rect 172641 530050 172699 530084
rect 172733 530050 172791 530084
rect 172825 530050 172883 530084
rect 172917 530050 172975 530084
rect 173009 530050 173067 530084
rect 173101 530050 173159 530084
rect 173193 530050 173251 530084
rect 173285 530050 173343 530084
rect 173377 530050 173435 530084
rect 173469 530050 173527 530084
rect 173561 530050 173619 530084
rect 173653 530050 173711 530084
rect 173745 530050 173803 530084
rect 173837 530050 173895 530084
rect 173929 530050 173965 530084
rect 174021 530050 174029 530084
rect 172210 530041 173965 530050
rect 174017 530041 174029 530050
rect 174081 530041 174093 530050
rect 174145 530041 174157 530093
rect 174209 530041 174221 530093
rect 174273 530084 177783 530093
rect 174297 530050 174355 530084
rect 174389 530050 174447 530084
rect 174481 530050 174539 530084
rect 174573 530050 174631 530084
rect 174665 530050 174723 530084
rect 174757 530050 174815 530084
rect 174849 530050 174907 530084
rect 174941 530050 174999 530084
rect 175033 530050 175091 530084
rect 175125 530050 175183 530084
rect 175217 530050 175275 530084
rect 175309 530050 175367 530084
rect 175401 530050 175459 530084
rect 175493 530050 175551 530084
rect 175585 530050 175643 530084
rect 175677 530050 175735 530084
rect 175769 530050 175827 530084
rect 175861 530050 175919 530084
rect 175953 530050 176011 530084
rect 176045 530050 176103 530084
rect 176137 530050 176195 530084
rect 176229 530050 176287 530084
rect 176321 530050 176379 530084
rect 176413 530050 176471 530084
rect 176505 530050 176563 530084
rect 176597 530050 176655 530084
rect 176689 530050 176747 530084
rect 176781 530050 176839 530084
rect 176873 530050 176931 530084
rect 176965 530050 177023 530084
rect 177057 530050 177115 530084
rect 177149 530050 177207 530084
rect 177241 530050 177299 530084
rect 177333 530050 177391 530084
rect 177425 530050 177483 530084
rect 177517 530050 177575 530084
rect 177609 530050 177667 530084
rect 177701 530050 177759 530084
rect 174273 530041 177783 530050
rect 177835 530041 177847 530093
rect 177899 530041 177911 530093
rect 177963 530084 177975 530093
rect 178027 530084 178039 530093
rect 178091 530084 181601 530093
rect 181653 530084 181665 530093
rect 181717 530084 181729 530093
rect 178027 530050 178035 530084
rect 178091 530050 178127 530084
rect 178161 530050 178219 530084
rect 178253 530050 178311 530084
rect 178345 530050 178403 530084
rect 178437 530050 178495 530084
rect 178529 530050 178587 530084
rect 178621 530050 178679 530084
rect 178713 530050 178771 530084
rect 178805 530050 178863 530084
rect 178897 530050 178955 530084
rect 178989 530050 179047 530084
rect 179081 530050 179139 530084
rect 179173 530050 179231 530084
rect 179265 530050 179323 530084
rect 179357 530050 179415 530084
rect 179449 530050 179507 530084
rect 179541 530050 179599 530084
rect 179633 530050 179691 530084
rect 179725 530050 179783 530084
rect 179817 530050 179875 530084
rect 179909 530050 179967 530084
rect 180001 530050 180059 530084
rect 180093 530050 180151 530084
rect 180185 530050 180243 530084
rect 180277 530050 180335 530084
rect 180369 530050 180427 530084
rect 180461 530050 180519 530084
rect 180553 530050 180611 530084
rect 180645 530050 180703 530084
rect 180737 530050 180795 530084
rect 180829 530050 180887 530084
rect 180921 530050 180979 530084
rect 181013 530050 181071 530084
rect 181105 530050 181163 530084
rect 181197 530050 181255 530084
rect 181289 530050 181347 530084
rect 181381 530050 181439 530084
rect 181473 530050 181531 530084
rect 181565 530050 181601 530084
rect 181657 530050 181665 530084
rect 177963 530041 177975 530050
rect 178027 530041 178039 530050
rect 178091 530041 181601 530050
rect 181653 530041 181665 530050
rect 181717 530041 181729 530050
rect 181781 530041 181793 530093
rect 181845 530041 181857 530093
rect 181909 530084 185419 530093
rect 181933 530050 181991 530084
rect 182025 530050 182083 530084
rect 182117 530050 182175 530084
rect 182209 530050 182267 530084
rect 182301 530050 182359 530084
rect 182393 530050 182451 530084
rect 182485 530050 182543 530084
rect 182577 530050 182635 530084
rect 182669 530050 182727 530084
rect 182761 530050 182819 530084
rect 182853 530050 182911 530084
rect 182945 530050 183003 530084
rect 183037 530050 183095 530084
rect 183129 530050 183187 530084
rect 183221 530050 183279 530084
rect 183313 530050 183371 530084
rect 183405 530050 183463 530084
rect 183497 530050 183555 530084
rect 183589 530050 183647 530084
rect 183681 530050 183739 530084
rect 183773 530050 183831 530084
rect 183865 530050 183923 530084
rect 183957 530050 184015 530084
rect 184049 530050 184107 530084
rect 184141 530050 184199 530084
rect 184233 530050 184291 530084
rect 184325 530050 184383 530084
rect 184417 530050 184475 530084
rect 184509 530050 184567 530084
rect 184601 530050 184659 530084
rect 184693 530050 184751 530084
rect 184785 530050 184843 530084
rect 184877 530050 184935 530084
rect 184969 530050 185027 530084
rect 185061 530050 185119 530084
rect 185153 530050 185211 530084
rect 185245 530050 185303 530084
rect 185337 530050 185395 530084
rect 181909 530041 185419 530050
rect 185471 530041 185483 530093
rect 185535 530041 185547 530093
rect 185599 530084 185611 530093
rect 185663 530084 185675 530093
rect 185727 530084 187482 530093
rect 185663 530050 185671 530084
rect 185727 530050 185763 530084
rect 185797 530050 185855 530084
rect 185889 530050 185947 530084
rect 185981 530050 186039 530084
rect 186073 530050 186131 530084
rect 186165 530050 186223 530084
rect 186257 530050 186315 530084
rect 186349 530050 186407 530084
rect 186441 530050 186499 530084
rect 186533 530050 186591 530084
rect 186625 530050 186683 530084
rect 186717 530050 186775 530084
rect 186809 530050 186867 530084
rect 186901 530050 186959 530084
rect 186993 530050 187051 530084
rect 187085 530050 187143 530084
rect 187177 530050 187235 530084
rect 187269 530050 187327 530084
rect 187361 530050 187419 530084
rect 187453 530050 187482 530084
rect 185599 530041 185611 530050
rect 185663 530041 185675 530050
rect 185727 530041 187482 530050
rect 172210 530019 187482 530041
rect 177287 529982 177345 529988
rect 177287 529948 177299 529982
rect 177333 529979 177345 529982
rect 178204 529979 178210 529991
rect 177333 529951 178210 529979
rect 177333 529948 177345 529951
rect 177287 529942 177345 529948
rect 178204 529939 178210 529951
rect 178262 529939 178268 529991
rect 178391 529982 178449 529988
rect 178391 529948 178403 529982
rect 178437 529979 178449 529982
rect 179492 529979 179498 529991
rect 178437 529951 179498 529979
rect 178437 529948 178449 529951
rect 178391 529942 178449 529948
rect 179492 529939 179498 529951
rect 179550 529939 179556 529991
rect 180872 529939 180878 529991
rect 180930 529979 180936 529991
rect 182160 529979 182166 529991
rect 180930 529951 182166 529979
rect 180930 529939 180936 529951
rect 182160 529939 182166 529951
rect 182218 529939 182224 529991
rect 182620 529939 182626 529991
rect 182678 529939 182684 529991
rect 175713 529914 175771 529920
rect 175713 529880 175725 529914
rect 175759 529911 175771 529914
rect 176091 529914 176149 529920
rect 176091 529911 176103 529914
rect 175759 529883 176103 529911
rect 175759 529880 175771 529883
rect 175713 529874 175771 529880
rect 176091 529880 176103 529883
rect 176137 529911 176149 529914
rect 176715 529914 176773 529920
rect 176715 529911 176727 529914
rect 176137 529883 176727 529911
rect 176137 529880 176149 529883
rect 176091 529874 176149 529880
rect 176715 529880 176727 529883
rect 176761 529880 176773 529914
rect 176715 529874 176773 529880
rect 178112 529871 178118 529923
rect 178170 529911 178176 529923
rect 178299 529914 178357 529920
rect 178299 529911 178311 529914
rect 178170 529883 178311 529911
rect 178170 529871 178176 529883
rect 178299 529880 178311 529883
rect 178345 529880 178357 529914
rect 178299 529874 178357 529880
rect 178963 529914 179021 529920
rect 178963 529880 178975 529914
rect 179009 529911 179021 529914
rect 179587 529914 179645 529920
rect 179587 529911 179599 529914
rect 179009 529883 179599 529911
rect 179009 529880 179021 529883
rect 178963 529874 179021 529880
rect 179587 529880 179599 529883
rect 179633 529911 179645 529914
rect 179965 529914 180023 529920
rect 179965 529911 179977 529914
rect 179633 529883 179977 529911
rect 179633 529880 179645 529883
rect 179587 529874 179645 529880
rect 179965 529880 179977 529883
rect 180011 529880 180023 529914
rect 179965 529874 180023 529880
rect 180405 529914 180463 529920
rect 180405 529880 180417 529914
rect 180451 529911 180463 529914
rect 180783 529914 180841 529920
rect 180783 529911 180795 529914
rect 180451 529883 180795 529911
rect 180451 529880 180463 529883
rect 180405 529874 180463 529880
rect 180783 529880 180795 529883
rect 180829 529911 180841 529914
rect 181407 529914 181465 529920
rect 181407 529911 181419 529914
rect 180829 529883 181419 529911
rect 180829 529880 180841 529883
rect 180783 529874 180841 529880
rect 181407 529880 181419 529883
rect 181453 529880 181465 529914
rect 181407 529874 181465 529880
rect 174800 529803 174806 529855
rect 174858 529803 174864 529855
rect 175815 529846 175873 529852
rect 175815 529812 175827 529846
rect 175861 529843 175873 529846
rect 177655 529846 177713 529852
rect 177655 529843 177667 529846
rect 175861 529815 177422 529843
rect 175861 529812 175873 529815
rect 175815 529806 175873 529812
rect 175539 529778 175597 529784
rect 175539 529744 175551 529778
rect 175585 529744 175597 529778
rect 175539 529738 175597 529744
rect 175632 529778 175690 529784
rect 175632 529744 175644 529778
rect 175678 529775 175690 529778
rect 175999 529778 176057 529784
rect 175999 529775 176011 529778
rect 175678 529747 176011 529775
rect 175678 529744 175690 529747
rect 175632 529738 175690 529744
rect 175999 529744 176011 529747
rect 176045 529775 176057 529778
rect 176715 529778 176773 529784
rect 176715 529775 176727 529778
rect 176045 529747 176727 529775
rect 176045 529744 176057 529747
rect 175999 529738 176057 529744
rect 176715 529744 176727 529747
rect 176761 529744 176773 529778
rect 176715 529738 176773 529744
rect 175554 529707 175582 529738
rect 176824 529735 176830 529787
rect 176882 529775 176888 529787
rect 176931 529775 176989 529779
rect 176882 529773 176989 529775
rect 176882 529747 176943 529773
rect 176882 529735 176888 529747
rect 176931 529739 176943 529747
rect 176977 529739 176989 529773
rect 176931 529716 176989 529739
rect 177394 529719 177422 529815
rect 177578 529815 177667 529843
rect 177578 529719 177606 529815
rect 177655 529812 177667 529815
rect 177701 529812 177713 529846
rect 179308 529843 179314 529855
rect 177655 529806 177713 529812
rect 177946 529815 179314 529843
rect 177946 529784 177974 529815
rect 179308 529803 179314 529815
rect 179366 529803 179372 529855
rect 179860 529803 179866 529855
rect 179918 529803 179924 529855
rect 180507 529846 180565 529852
rect 180507 529812 180519 529846
rect 180553 529843 180565 529846
rect 181979 529846 182037 529852
rect 180553 529815 181838 529843
rect 180553 529812 180565 529815
rect 180507 529806 180565 529812
rect 177931 529778 177989 529784
rect 177931 529744 177943 529778
rect 177977 529744 177989 529778
rect 177931 529738 177989 529744
rect 178747 529773 178805 529779
rect 178747 529739 178759 529773
rect 178793 529739 178805 529773
rect 176271 529710 176401 529716
rect 175554 529679 176134 529707
rect 176106 529651 176134 529679
rect 176271 529676 176283 529710
rect 176317 529676 176355 529710
rect 176389 529707 176401 529710
rect 176931 529710 177049 529716
rect 176931 529707 177003 529710
rect 176389 529679 177003 529707
rect 176389 529676 176401 529679
rect 176271 529670 176401 529676
rect 175352 529599 175358 529651
rect 175410 529639 175416 529651
rect 175447 529642 175505 529648
rect 175447 529639 175459 529642
rect 175410 529611 175459 529639
rect 175410 529599 175416 529611
rect 175447 529608 175459 529611
rect 175493 529608 175505 529642
rect 175447 529602 175505 529608
rect 176088 529599 176094 529651
rect 176146 529599 176152 529651
rect 176934 529639 176962 529679
rect 176991 529676 177003 529679
rect 177037 529676 177049 529710
rect 176991 529670 177049 529676
rect 177376 529667 177382 529719
rect 177434 529667 177440 529719
rect 177560 529667 177566 529719
rect 177618 529667 177624 529719
rect 177652 529667 177658 529719
rect 177710 529707 177716 529719
rect 178747 529716 178805 529739
rect 178963 529778 179021 529784
rect 178963 529744 178975 529778
rect 179009 529775 179021 529778
rect 179679 529778 179737 529784
rect 179679 529775 179691 529778
rect 179009 529747 179691 529775
rect 179009 529744 179021 529747
rect 178963 529738 179021 529744
rect 179679 529744 179691 529747
rect 179725 529775 179737 529778
rect 180046 529778 180104 529784
rect 180046 529775 180058 529778
rect 179725 529747 180058 529775
rect 179725 529744 179737 529747
rect 179679 529738 179737 529744
rect 180046 529744 180058 529747
rect 180092 529744 180104 529778
rect 180046 529738 180104 529744
rect 180139 529778 180197 529784
rect 180139 529744 180151 529778
rect 180185 529775 180197 529778
rect 180231 529778 180289 529784
rect 180231 529775 180243 529778
rect 180185 529747 180243 529775
rect 180185 529744 180197 529747
rect 180139 529738 180197 529744
rect 180231 529744 180243 529747
rect 180277 529744 180289 529778
rect 180231 529738 180289 529744
rect 180324 529778 180382 529784
rect 180324 529744 180336 529778
rect 180370 529775 180382 529778
rect 180691 529778 180749 529784
rect 180691 529775 180703 529778
rect 180370 529747 180703 529775
rect 180370 529744 180382 529747
rect 180324 529738 180382 529744
rect 180691 529744 180703 529747
rect 180737 529775 180749 529778
rect 181407 529778 181465 529784
rect 181407 529775 181419 529778
rect 180737 529747 181419 529775
rect 180737 529744 180749 529747
rect 180691 529738 180749 529744
rect 181407 529744 181419 529747
rect 181453 529744 181465 529778
rect 181407 529738 181465 529744
rect 181623 529773 181681 529779
rect 181623 529739 181635 529773
rect 181669 529739 181681 529773
rect 177839 529710 177897 529716
rect 177839 529707 177851 529710
rect 177710 529679 177851 529707
rect 177710 529667 177716 529679
rect 177839 529676 177851 529679
rect 177885 529676 177897 529710
rect 178687 529710 178805 529716
rect 178687 529707 178699 529710
rect 177839 529670 177897 529676
rect 178406 529679 178699 529707
rect 177928 529639 177934 529651
rect 176934 529611 177934 529639
rect 177928 529599 177934 529611
rect 177986 529639 177992 529651
rect 178406 529639 178434 529679
rect 178687 529676 178699 529679
rect 178733 529707 178805 529710
rect 179335 529710 179465 529716
rect 179335 529707 179347 529710
rect 178733 529679 179347 529707
rect 178733 529676 178745 529679
rect 178687 529670 178745 529676
rect 179335 529676 179347 529679
rect 179381 529676 179419 529710
rect 179453 529676 179465 529710
rect 180246 529707 180274 529738
rect 180963 529710 181093 529716
rect 180246 529679 180550 529707
rect 179335 529670 179465 529676
rect 180522 529651 180550 529679
rect 180963 529676 180975 529710
rect 181009 529676 181047 529710
rect 181081 529707 181093 529710
rect 181516 529707 181522 529719
rect 181081 529679 181522 529707
rect 181081 529676 181093 529679
rect 180963 529670 181093 529676
rect 181516 529667 181522 529679
rect 181574 529707 181580 529719
rect 181623 529716 181681 529739
rect 181623 529710 181741 529716
rect 181623 529707 181695 529710
rect 181574 529679 181695 529707
rect 181574 529667 181580 529679
rect 181683 529676 181695 529679
rect 181729 529676 181741 529710
rect 181683 529670 181741 529676
rect 181810 529651 181838 529815
rect 181979 529812 181991 529846
rect 182025 529843 182037 529846
rect 183172 529843 183178 529855
rect 182025 529815 183178 529843
rect 182025 529812 182037 529815
rect 181979 529806 182037 529812
rect 183172 529803 183178 529815
rect 183230 529803 183236 529855
rect 177986 529611 178434 529639
rect 177986 529599 177992 529611
rect 180504 529599 180510 529651
rect 180562 529599 180568 529651
rect 181792 529599 181798 529651
rect 181850 529599 181856 529651
rect 172210 529549 187482 529571
rect 172210 529540 174625 529549
rect 172210 529506 172239 529540
rect 172273 529506 172331 529540
rect 172365 529506 172423 529540
rect 172457 529506 172515 529540
rect 172549 529506 172607 529540
rect 172641 529506 172699 529540
rect 172733 529506 172791 529540
rect 172825 529506 172883 529540
rect 172917 529506 172975 529540
rect 173009 529506 173067 529540
rect 173101 529506 173159 529540
rect 173193 529506 173251 529540
rect 173285 529506 173343 529540
rect 173377 529506 173435 529540
rect 173469 529506 173527 529540
rect 173561 529506 173619 529540
rect 173653 529506 173711 529540
rect 173745 529506 173803 529540
rect 173837 529506 173895 529540
rect 173929 529506 173987 529540
rect 174021 529506 174079 529540
rect 174113 529506 174171 529540
rect 174205 529506 174263 529540
rect 174297 529506 174355 529540
rect 174389 529506 174447 529540
rect 174481 529506 174539 529540
rect 174573 529506 174625 529540
rect 172210 529497 174625 529506
rect 174677 529497 174689 529549
rect 174741 529540 174753 529549
rect 174805 529540 174817 529549
rect 174805 529506 174815 529540
rect 174741 529497 174753 529506
rect 174805 529497 174817 529506
rect 174869 529497 174881 529549
rect 174933 529540 178443 529549
rect 174941 529506 174999 529540
rect 175033 529506 175091 529540
rect 175125 529506 175183 529540
rect 175217 529506 175275 529540
rect 175309 529506 175367 529540
rect 175401 529506 175459 529540
rect 175493 529506 175551 529540
rect 175585 529506 175643 529540
rect 175677 529506 175735 529540
rect 175769 529506 175827 529540
rect 175861 529506 175919 529540
rect 175953 529506 176011 529540
rect 176045 529506 176103 529540
rect 176137 529506 176195 529540
rect 176229 529506 176287 529540
rect 176321 529506 176379 529540
rect 176413 529506 176471 529540
rect 176505 529506 176563 529540
rect 176597 529506 176655 529540
rect 176689 529506 176747 529540
rect 176781 529506 176839 529540
rect 176873 529506 176931 529540
rect 176965 529506 177023 529540
rect 177057 529506 177115 529540
rect 177149 529506 177207 529540
rect 177241 529506 177299 529540
rect 177333 529506 177391 529540
rect 177425 529506 177483 529540
rect 177517 529506 177575 529540
rect 177609 529506 177667 529540
rect 177701 529506 177759 529540
rect 177793 529506 177851 529540
rect 177885 529506 177943 529540
rect 177977 529506 178035 529540
rect 178069 529506 178127 529540
rect 178161 529506 178219 529540
rect 178253 529506 178311 529540
rect 178345 529506 178403 529540
rect 178437 529506 178443 529540
rect 174933 529497 178443 529506
rect 178495 529540 178507 529549
rect 178495 529497 178507 529506
rect 178559 529497 178571 529549
rect 178623 529497 178635 529549
rect 178687 529540 178699 529549
rect 178751 529540 182261 529549
rect 178751 529506 178771 529540
rect 178805 529506 178863 529540
rect 178897 529506 178955 529540
rect 178989 529506 179047 529540
rect 179081 529506 179139 529540
rect 179173 529506 179231 529540
rect 179265 529506 179323 529540
rect 179357 529506 179415 529540
rect 179449 529506 179507 529540
rect 179541 529506 179599 529540
rect 179633 529506 179691 529540
rect 179725 529506 179783 529540
rect 179817 529506 179875 529540
rect 179909 529506 179967 529540
rect 180001 529506 180059 529540
rect 180093 529506 180151 529540
rect 180185 529506 180243 529540
rect 180277 529506 180335 529540
rect 180369 529506 180427 529540
rect 180461 529506 180519 529540
rect 180553 529506 180611 529540
rect 180645 529506 180703 529540
rect 180737 529506 180795 529540
rect 180829 529506 180887 529540
rect 180921 529506 180979 529540
rect 181013 529506 181071 529540
rect 181105 529506 181163 529540
rect 181197 529506 181255 529540
rect 181289 529506 181347 529540
rect 181381 529506 181439 529540
rect 181473 529506 181531 529540
rect 181565 529506 181623 529540
rect 181657 529506 181715 529540
rect 181749 529506 181807 529540
rect 181841 529506 181899 529540
rect 181933 529506 181991 529540
rect 182025 529506 182083 529540
rect 182117 529506 182175 529540
rect 182209 529506 182261 529540
rect 178687 529497 178699 529506
rect 178751 529497 182261 529506
rect 182313 529497 182325 529549
rect 182377 529540 182389 529549
rect 182441 529540 182453 529549
rect 182441 529506 182451 529540
rect 182377 529497 182389 529506
rect 182441 529497 182453 529506
rect 182505 529497 182517 529549
rect 182569 529540 186079 529549
rect 182577 529506 182635 529540
rect 182669 529506 182727 529540
rect 182761 529506 182819 529540
rect 182853 529506 182911 529540
rect 182945 529506 183003 529540
rect 183037 529506 183095 529540
rect 183129 529506 183187 529540
rect 183221 529506 183279 529540
rect 183313 529506 183371 529540
rect 183405 529506 183463 529540
rect 183497 529506 183555 529540
rect 183589 529506 183647 529540
rect 183681 529506 183739 529540
rect 183773 529506 183831 529540
rect 183865 529506 183923 529540
rect 183957 529506 184015 529540
rect 184049 529506 184107 529540
rect 184141 529506 184199 529540
rect 184233 529506 184291 529540
rect 184325 529506 184383 529540
rect 184417 529506 184475 529540
rect 184509 529506 184567 529540
rect 184601 529506 184659 529540
rect 184693 529506 184751 529540
rect 184785 529506 184843 529540
rect 184877 529506 184935 529540
rect 184969 529506 185027 529540
rect 185061 529506 185119 529540
rect 185153 529506 185211 529540
rect 185245 529506 185303 529540
rect 185337 529506 185395 529540
rect 185429 529506 185487 529540
rect 185521 529506 185579 529540
rect 185613 529506 185671 529540
rect 185705 529506 185763 529540
rect 185797 529506 185855 529540
rect 185889 529506 185947 529540
rect 185981 529506 186039 529540
rect 186073 529506 186079 529540
rect 182569 529497 186079 529506
rect 186131 529540 186143 529549
rect 186131 529497 186143 529506
rect 186195 529497 186207 529549
rect 186259 529497 186271 529549
rect 186323 529540 186335 529549
rect 186387 529540 187482 529549
rect 186387 529506 186407 529540
rect 186441 529506 186499 529540
rect 186533 529506 186591 529540
rect 186625 529506 186683 529540
rect 186717 529506 186775 529540
rect 186809 529506 186867 529540
rect 186901 529506 186959 529540
rect 186993 529506 187051 529540
rect 187085 529506 187143 529540
rect 187177 529506 187235 529540
rect 187269 529506 187327 529540
rect 187361 529506 187419 529540
rect 187453 529506 187482 529540
rect 186323 529497 186335 529506
rect 186387 529497 187482 529506
rect 172210 529475 187482 529497
rect 175352 529395 175358 529447
rect 175410 529395 175416 529447
rect 177928 529395 177934 529447
rect 177986 529435 177992 529447
rect 177986 529407 179354 529435
rect 177986 529395 177992 529407
rect 178023 529370 178081 529376
rect 178023 529336 178035 529370
rect 178069 529367 178081 529370
rect 178296 529367 178302 529379
rect 178069 529339 178302 529367
rect 178069 529336 178081 529339
rect 178023 529330 178081 529336
rect 178296 529327 178302 529339
rect 178354 529327 178360 529379
rect 178479 529370 178609 529376
rect 178479 529336 178491 529370
rect 178525 529336 178563 529370
rect 178597 529367 178609 529370
rect 179199 529370 179257 529376
rect 179199 529367 179211 529370
rect 178597 529339 179211 529367
rect 178597 529336 178609 529339
rect 178479 529330 178609 529336
rect 179139 529336 179211 529339
rect 179245 529367 179257 529370
rect 179326 529367 179354 529407
rect 179860 529395 179866 529447
rect 179918 529395 179924 529447
rect 181792 529395 181798 529447
rect 181850 529435 181856 529447
rect 182531 529438 182589 529444
rect 182531 529435 182543 529438
rect 181850 529407 182543 529435
rect 181850 529395 181856 529407
rect 182531 529404 182543 529407
rect 182577 529404 182589 529438
rect 182531 529398 182589 529404
rect 179245 529339 181562 529367
rect 179245 529336 179257 529339
rect 179139 529330 179257 529336
rect 175444 529259 175450 529311
rect 175502 529299 175508 529311
rect 176732 529299 176738 529311
rect 175502 529271 176738 529299
rect 175502 529259 175508 529271
rect 176732 529259 176738 529271
rect 176790 529259 176796 529311
rect 177652 529259 177658 529311
rect 177710 529259 177716 529311
rect 177840 529302 177898 529308
rect 177840 529268 177852 529302
rect 177886 529299 177898 529302
rect 178207 529302 178265 529308
rect 178207 529299 178219 529302
rect 177886 529271 178219 529299
rect 177886 529268 177898 529271
rect 177840 529262 177898 529268
rect 178207 529268 178219 529271
rect 178253 529299 178265 529302
rect 178923 529302 178981 529308
rect 178923 529299 178935 529302
rect 178253 529271 178935 529299
rect 178253 529268 178265 529271
rect 178207 529262 178265 529268
rect 178923 529268 178935 529271
rect 178969 529268 178981 529302
rect 178923 529262 178981 529268
rect 179139 529307 179197 529330
rect 181534 529311 181562 529339
rect 179139 529273 179151 529307
rect 179185 529273 179197 529307
rect 179139 529267 179197 529273
rect 179676 529259 179682 529311
rect 179734 529259 179740 529311
rect 180691 529302 180749 529308
rect 180691 529268 180703 529302
rect 180737 529268 180749 529302
rect 180691 529262 180749 529268
rect 173604 529191 173610 529243
rect 173662 529231 173668 529243
rect 175260 529231 175266 529243
rect 173662 529203 175266 529231
rect 173662 529191 173668 529203
rect 175260 529191 175266 529203
rect 175318 529191 175324 529243
rect 177284 529231 177290 529243
rect 176198 529203 177290 529231
rect 175815 529098 175873 529104
rect 175815 529064 175827 529098
rect 175861 529095 175873 529098
rect 175904 529095 175910 529107
rect 175861 529067 175910 529095
rect 175861 529064 175873 529067
rect 175815 529058 175873 529064
rect 175904 529055 175910 529067
rect 175962 529055 175968 529107
rect 176088 529055 176094 529107
rect 176146 529095 176152 529107
rect 176198 529104 176226 529203
rect 177284 529191 177290 529203
rect 177342 529231 177348 529243
rect 177747 529234 177805 529240
rect 177747 529231 177759 529234
rect 177342 529203 177759 529231
rect 177342 529191 177348 529203
rect 177747 529200 177759 529203
rect 177793 529200 177805 529234
rect 180706 529231 180734 529262
rect 181516 529259 181522 529311
rect 181574 529259 181580 529311
rect 182712 529259 182718 529311
rect 182770 529259 182776 529311
rect 177747 529194 177805 529200
rect 179694 529203 180734 529231
rect 177921 529166 177979 529172
rect 177921 529132 177933 529166
rect 177967 529163 177979 529166
rect 178299 529166 178357 529172
rect 178299 529163 178311 529166
rect 177967 529135 178311 529163
rect 177967 529132 177979 529135
rect 177921 529126 177979 529132
rect 178299 529132 178311 529135
rect 178345 529163 178357 529166
rect 178923 529166 178981 529172
rect 178923 529163 178935 529166
rect 178345 529135 178935 529163
rect 178345 529132 178357 529135
rect 178299 529126 178357 529132
rect 178923 529132 178935 529135
rect 178969 529132 178981 529166
rect 178923 529126 178981 529132
rect 179694 529107 179722 529203
rect 176183 529098 176241 529104
rect 176183 529095 176195 529098
rect 176146 529067 176195 529095
rect 176146 529055 176152 529067
rect 176183 529064 176195 529067
rect 176229 529064 176241 529098
rect 176183 529058 176241 529064
rect 179308 529055 179314 529107
rect 179366 529095 179372 529107
rect 179495 529098 179553 529104
rect 179495 529095 179507 529098
rect 179366 529067 179507 529095
rect 179366 529055 179372 529067
rect 179495 529064 179507 529067
rect 179541 529064 179553 529098
rect 179495 529058 179553 529064
rect 179676 529055 179682 529107
rect 179734 529055 179740 529107
rect 180504 529055 180510 529107
rect 180562 529095 180568 529107
rect 181979 529098 182037 529104
rect 181979 529095 181991 529098
rect 180562 529067 181991 529095
rect 180562 529055 180568 529067
rect 181979 529064 181991 529067
rect 182025 529064 182037 529098
rect 181979 529058 182037 529064
rect 172210 529005 187482 529027
rect 172210 528996 173965 529005
rect 174017 528996 174029 529005
rect 174081 528996 174093 529005
rect 172210 528962 172239 528996
rect 172273 528962 172331 528996
rect 172365 528962 172423 528996
rect 172457 528962 172515 528996
rect 172549 528962 172607 528996
rect 172641 528962 172699 528996
rect 172733 528962 172791 528996
rect 172825 528962 172883 528996
rect 172917 528962 172975 528996
rect 173009 528962 173067 528996
rect 173101 528962 173159 528996
rect 173193 528962 173251 528996
rect 173285 528962 173343 528996
rect 173377 528962 173435 528996
rect 173469 528962 173527 528996
rect 173561 528962 173619 528996
rect 173653 528962 173711 528996
rect 173745 528962 173803 528996
rect 173837 528962 173895 528996
rect 173929 528962 173965 528996
rect 174021 528962 174029 528996
rect 172210 528953 173965 528962
rect 174017 528953 174029 528962
rect 174081 528953 174093 528962
rect 174145 528953 174157 529005
rect 174209 528953 174221 529005
rect 174273 528996 177783 529005
rect 174297 528962 174355 528996
rect 174389 528962 174447 528996
rect 174481 528962 174539 528996
rect 174573 528962 174631 528996
rect 174665 528962 174723 528996
rect 174757 528962 174815 528996
rect 174849 528962 174907 528996
rect 174941 528962 174999 528996
rect 175033 528962 175091 528996
rect 175125 528962 175183 528996
rect 175217 528962 175275 528996
rect 175309 528962 175367 528996
rect 175401 528962 175459 528996
rect 175493 528962 175551 528996
rect 175585 528962 175643 528996
rect 175677 528962 175735 528996
rect 175769 528962 175827 528996
rect 175861 528962 175919 528996
rect 175953 528962 176011 528996
rect 176045 528962 176103 528996
rect 176137 528962 176195 528996
rect 176229 528962 176287 528996
rect 176321 528962 176379 528996
rect 176413 528962 176471 528996
rect 176505 528962 176563 528996
rect 176597 528962 176655 528996
rect 176689 528962 176747 528996
rect 176781 528962 176839 528996
rect 176873 528962 176931 528996
rect 176965 528962 177023 528996
rect 177057 528962 177115 528996
rect 177149 528962 177207 528996
rect 177241 528962 177299 528996
rect 177333 528962 177391 528996
rect 177425 528962 177483 528996
rect 177517 528962 177575 528996
rect 177609 528962 177667 528996
rect 177701 528962 177759 528996
rect 174273 528953 177783 528962
rect 177835 528953 177847 529005
rect 177899 528953 177911 529005
rect 177963 528996 177975 529005
rect 178027 528996 178039 529005
rect 178091 528996 181601 529005
rect 181653 528996 181665 529005
rect 181717 528996 181729 529005
rect 178027 528962 178035 528996
rect 178091 528962 178127 528996
rect 178161 528962 178219 528996
rect 178253 528962 178311 528996
rect 178345 528962 178403 528996
rect 178437 528962 178495 528996
rect 178529 528962 178587 528996
rect 178621 528962 178679 528996
rect 178713 528962 178771 528996
rect 178805 528962 178863 528996
rect 178897 528962 178955 528996
rect 178989 528962 179047 528996
rect 179081 528962 179139 528996
rect 179173 528962 179231 528996
rect 179265 528962 179323 528996
rect 179357 528962 179415 528996
rect 179449 528962 179507 528996
rect 179541 528962 179599 528996
rect 179633 528962 179691 528996
rect 179725 528962 179783 528996
rect 179817 528962 179875 528996
rect 179909 528962 179967 528996
rect 180001 528962 180059 528996
rect 180093 528962 180151 528996
rect 180185 528962 180243 528996
rect 180277 528962 180335 528996
rect 180369 528962 180427 528996
rect 180461 528962 180519 528996
rect 180553 528962 180611 528996
rect 180645 528962 180703 528996
rect 180737 528962 180795 528996
rect 180829 528962 180887 528996
rect 180921 528962 180979 528996
rect 181013 528962 181071 528996
rect 181105 528962 181163 528996
rect 181197 528962 181255 528996
rect 181289 528962 181347 528996
rect 181381 528962 181439 528996
rect 181473 528962 181531 528996
rect 181565 528962 181601 528996
rect 181657 528962 181665 528996
rect 177963 528953 177975 528962
rect 178027 528953 178039 528962
rect 178091 528953 181601 528962
rect 181653 528953 181665 528962
rect 181717 528953 181729 528962
rect 181781 528953 181793 529005
rect 181845 528953 181857 529005
rect 181909 528996 185419 529005
rect 181933 528962 181991 528996
rect 182025 528962 182083 528996
rect 182117 528962 182175 528996
rect 182209 528962 182267 528996
rect 182301 528962 182359 528996
rect 182393 528962 182451 528996
rect 182485 528962 182543 528996
rect 182577 528962 182635 528996
rect 182669 528962 182727 528996
rect 182761 528962 182819 528996
rect 182853 528962 182911 528996
rect 182945 528962 183003 528996
rect 183037 528962 183095 528996
rect 183129 528962 183187 528996
rect 183221 528962 183279 528996
rect 183313 528962 183371 528996
rect 183405 528962 183463 528996
rect 183497 528962 183555 528996
rect 183589 528962 183647 528996
rect 183681 528962 183739 528996
rect 183773 528962 183831 528996
rect 183865 528962 183923 528996
rect 183957 528962 184015 528996
rect 184049 528962 184107 528996
rect 184141 528962 184199 528996
rect 184233 528962 184291 528996
rect 184325 528962 184383 528996
rect 184417 528962 184475 528996
rect 184509 528962 184567 528996
rect 184601 528962 184659 528996
rect 184693 528962 184751 528996
rect 184785 528962 184843 528996
rect 184877 528962 184935 528996
rect 184969 528962 185027 528996
rect 185061 528962 185119 528996
rect 185153 528962 185211 528996
rect 185245 528962 185303 528996
rect 185337 528962 185395 528996
rect 181909 528953 185419 528962
rect 185471 528953 185483 529005
rect 185535 528953 185547 529005
rect 185599 528996 185611 529005
rect 185663 528996 185675 529005
rect 185727 528996 187482 529005
rect 185663 528962 185671 528996
rect 185727 528962 185763 528996
rect 185797 528962 185855 528996
rect 185889 528962 185947 528996
rect 185981 528962 186039 528996
rect 186073 528962 186131 528996
rect 186165 528962 186223 528996
rect 186257 528962 186315 528996
rect 186349 528962 186407 528996
rect 186441 528962 186499 528996
rect 186533 528962 186591 528996
rect 186625 528962 186683 528996
rect 186717 528962 186775 528996
rect 186809 528962 186867 528996
rect 186901 528962 186959 528996
rect 186993 528962 187051 528996
rect 187085 528962 187143 528996
rect 187177 528962 187235 528996
rect 187269 528962 187327 528996
rect 187361 528962 187419 528996
rect 187453 528962 187482 528996
rect 185599 528953 185611 528962
rect 185663 528953 185675 528962
rect 185727 528953 187482 528962
rect 172210 528931 187482 528953
rect 175260 528851 175266 528903
rect 175318 528851 175324 528903
rect 176091 528894 176149 528900
rect 176091 528860 176103 528894
rect 176137 528891 176149 528894
rect 176640 528891 176646 528903
rect 176137 528863 176646 528891
rect 176137 528860 176149 528863
rect 176091 528854 176149 528860
rect 176640 528851 176646 528863
rect 176698 528851 176704 528903
rect 177652 528851 177658 528903
rect 177710 528891 177716 528903
rect 179676 528891 179682 528903
rect 177710 528863 179682 528891
rect 177710 528851 177716 528863
rect 179676 528851 179682 528863
rect 179734 528851 179740 528903
rect 180430 528863 180642 528891
rect 175278 528755 175306 528851
rect 180430 528832 180458 528863
rect 180415 528826 180473 528832
rect 180415 528792 180427 528826
rect 180461 528792 180473 528826
rect 180415 528786 180473 528792
rect 176551 528758 176609 528764
rect 176551 528755 176563 528758
rect 175278 528727 176563 528755
rect 176551 528724 176563 528727
rect 176597 528755 176609 528758
rect 177560 528755 177566 528767
rect 176597 528727 177566 528755
rect 176597 528724 176609 528727
rect 176551 528718 176609 528724
rect 177560 528715 177566 528727
rect 177618 528755 177624 528767
rect 178020 528755 178026 528767
rect 177618 528727 178026 528755
rect 177618 528715 177624 528727
rect 178020 528715 178026 528727
rect 178078 528715 178084 528767
rect 178115 528758 178173 528764
rect 178115 528724 178127 528758
rect 178161 528755 178173 528758
rect 178204 528755 178210 528767
rect 178161 528727 178210 528755
rect 178161 528724 178173 528727
rect 178115 528718 178173 528724
rect 178204 528715 178210 528727
rect 178262 528715 178268 528767
rect 180504 528715 180510 528767
rect 180562 528715 180568 528767
rect 180614 528755 180642 528863
rect 182160 528851 182166 528903
rect 182218 528891 182224 528903
rect 182255 528894 182313 528900
rect 182255 528891 182267 528894
rect 182218 528863 182267 528891
rect 182218 528851 182224 528863
rect 182255 528860 182267 528863
rect 182301 528860 182313 528894
rect 182255 528854 182313 528860
rect 180681 528826 180739 528832
rect 180681 528792 180693 528826
rect 180727 528823 180739 528826
rect 181059 528826 181117 528832
rect 181059 528823 181071 528826
rect 180727 528795 181071 528823
rect 180727 528792 180739 528795
rect 180681 528786 180739 528792
rect 181059 528792 181071 528795
rect 181105 528823 181117 528826
rect 181683 528826 181741 528832
rect 181683 528823 181695 528826
rect 181105 528795 181695 528823
rect 181105 528792 181117 528795
rect 181059 528786 181117 528792
rect 181683 528792 181695 528795
rect 181729 528792 181741 528826
rect 181683 528786 181741 528792
rect 180783 528758 180841 528764
rect 180783 528755 180795 528758
rect 180614 528727 180795 528755
rect 180783 528724 180795 528727
rect 180829 528724 180841 528758
rect 180783 528718 180841 528724
rect 181516 528715 181522 528767
rect 181574 528755 181580 528767
rect 181574 528727 182022 528755
rect 181574 528715 181580 528727
rect 175904 528647 175910 528699
rect 175962 528647 175968 528699
rect 176183 528690 176241 528696
rect 176183 528656 176195 528690
rect 176229 528687 176241 528690
rect 176827 528690 176885 528696
rect 176229 528659 176318 528687
rect 176229 528656 176241 528659
rect 176183 528650 176241 528656
rect 176290 528563 176318 528659
rect 176827 528656 176839 528690
rect 176873 528687 176885 528690
rect 177471 528690 177529 528696
rect 177471 528687 177483 528690
rect 176873 528659 177483 528687
rect 176873 528656 176885 528659
rect 176827 528650 176885 528656
rect 177471 528656 177483 528659
rect 177517 528656 177529 528690
rect 177471 528650 177529 528656
rect 180231 528690 180289 528696
rect 180231 528656 180243 528690
rect 180277 528687 180289 528690
rect 180600 528690 180658 528696
rect 180277 528659 180550 528687
rect 180277 528656 180289 528659
rect 180231 528650 180289 528656
rect 178388 528579 178394 528631
rect 178446 528579 178452 528631
rect 180522 528619 180550 528659
rect 180600 528656 180612 528690
rect 180646 528687 180658 528690
rect 180967 528690 181025 528696
rect 180967 528687 180979 528690
rect 180646 528659 180979 528687
rect 180646 528656 180658 528659
rect 180600 528650 180658 528656
rect 180967 528656 180979 528659
rect 181013 528687 181025 528690
rect 181683 528690 181741 528696
rect 181683 528687 181695 528690
rect 181013 528659 181695 528687
rect 181013 528656 181025 528659
rect 180967 528650 181025 528656
rect 181683 528656 181695 528659
rect 181729 528656 181741 528690
rect 181683 528650 181741 528656
rect 181899 528685 181957 528691
rect 181899 528651 181911 528685
rect 181945 528651 181957 528685
rect 181899 528628 181957 528651
rect 181994 528628 182022 528727
rect 181239 528622 181369 528628
rect 180522 528591 181010 528619
rect 180982 528563 181010 528591
rect 181239 528588 181251 528622
rect 181285 528588 181323 528622
rect 181357 528619 181369 528622
rect 181899 528622 182022 528628
rect 181899 528619 181971 528622
rect 181357 528591 181971 528619
rect 181357 528588 181369 528591
rect 181239 528582 181369 528588
rect 181959 528588 181971 528591
rect 182005 528619 182022 528622
rect 186576 528619 186582 528631
rect 182005 528591 186582 528619
rect 182005 528588 182017 528591
rect 181959 528582 182017 528588
rect 186576 528579 186582 528591
rect 186634 528579 186640 528631
rect 176272 528511 176278 528563
rect 176330 528511 176336 528563
rect 176364 528511 176370 528563
rect 176422 528511 176428 528563
rect 176732 528511 176738 528563
rect 176790 528511 176796 528563
rect 177008 528511 177014 528563
rect 177066 528551 177072 528563
rect 177195 528554 177253 528560
rect 177195 528551 177207 528554
rect 177066 528523 177207 528551
rect 177066 528511 177072 528523
rect 177195 528520 177207 528523
rect 177241 528520 177253 528554
rect 177195 528514 177253 528520
rect 180964 528511 180970 528563
rect 181022 528511 181028 528563
rect 172210 528461 187482 528483
rect 172210 528452 174625 528461
rect 172210 528418 172239 528452
rect 172273 528418 172331 528452
rect 172365 528418 172423 528452
rect 172457 528418 172515 528452
rect 172549 528418 172607 528452
rect 172641 528418 172699 528452
rect 172733 528418 172791 528452
rect 172825 528418 172883 528452
rect 172917 528418 172975 528452
rect 173009 528418 173067 528452
rect 173101 528418 173159 528452
rect 173193 528418 173251 528452
rect 173285 528418 173343 528452
rect 173377 528418 173435 528452
rect 173469 528418 173527 528452
rect 173561 528418 173619 528452
rect 173653 528418 173711 528452
rect 173745 528418 173803 528452
rect 173837 528418 173895 528452
rect 173929 528418 173987 528452
rect 174021 528418 174079 528452
rect 174113 528418 174171 528452
rect 174205 528418 174263 528452
rect 174297 528418 174355 528452
rect 174389 528418 174447 528452
rect 174481 528418 174539 528452
rect 174573 528418 174625 528452
rect 172210 528409 174625 528418
rect 174677 528409 174689 528461
rect 174741 528452 174753 528461
rect 174805 528452 174817 528461
rect 174805 528418 174815 528452
rect 174741 528409 174753 528418
rect 174805 528409 174817 528418
rect 174869 528409 174881 528461
rect 174933 528452 178443 528461
rect 174941 528418 174999 528452
rect 175033 528418 175091 528452
rect 175125 528418 175183 528452
rect 175217 528418 175275 528452
rect 175309 528418 175367 528452
rect 175401 528418 175459 528452
rect 175493 528418 175551 528452
rect 175585 528418 175643 528452
rect 175677 528418 175735 528452
rect 175769 528418 175827 528452
rect 175861 528418 175919 528452
rect 175953 528418 176011 528452
rect 176045 528418 176103 528452
rect 176137 528418 176195 528452
rect 176229 528418 176287 528452
rect 176321 528418 176379 528452
rect 176413 528418 176471 528452
rect 176505 528418 176563 528452
rect 176597 528418 176655 528452
rect 176689 528418 176747 528452
rect 176781 528418 176839 528452
rect 176873 528418 176931 528452
rect 176965 528418 177023 528452
rect 177057 528418 177115 528452
rect 177149 528418 177207 528452
rect 177241 528418 177299 528452
rect 177333 528418 177391 528452
rect 177425 528418 177483 528452
rect 177517 528418 177575 528452
rect 177609 528418 177667 528452
rect 177701 528418 177759 528452
rect 177793 528418 177851 528452
rect 177885 528418 177943 528452
rect 177977 528418 178035 528452
rect 178069 528418 178127 528452
rect 178161 528418 178219 528452
rect 178253 528418 178311 528452
rect 178345 528418 178403 528452
rect 178437 528418 178443 528452
rect 174933 528409 178443 528418
rect 178495 528452 178507 528461
rect 178495 528409 178507 528418
rect 178559 528409 178571 528461
rect 178623 528409 178635 528461
rect 178687 528452 178699 528461
rect 178751 528452 182261 528461
rect 178751 528418 178771 528452
rect 178805 528418 178863 528452
rect 178897 528418 178955 528452
rect 178989 528418 179047 528452
rect 179081 528418 179139 528452
rect 179173 528418 179231 528452
rect 179265 528418 179323 528452
rect 179357 528418 179415 528452
rect 179449 528418 179507 528452
rect 179541 528418 179599 528452
rect 179633 528418 179691 528452
rect 179725 528418 179783 528452
rect 179817 528418 179875 528452
rect 179909 528418 179967 528452
rect 180001 528418 180059 528452
rect 180093 528418 180151 528452
rect 180185 528418 180243 528452
rect 180277 528418 180335 528452
rect 180369 528418 180427 528452
rect 180461 528418 180519 528452
rect 180553 528418 180611 528452
rect 180645 528418 180703 528452
rect 180737 528418 180795 528452
rect 180829 528418 180887 528452
rect 180921 528418 180979 528452
rect 181013 528418 181071 528452
rect 181105 528418 181163 528452
rect 181197 528418 181255 528452
rect 181289 528418 181347 528452
rect 181381 528418 181439 528452
rect 181473 528418 181531 528452
rect 181565 528418 181623 528452
rect 181657 528418 181715 528452
rect 181749 528418 181807 528452
rect 181841 528418 181899 528452
rect 181933 528418 181991 528452
rect 182025 528418 182083 528452
rect 182117 528418 182175 528452
rect 182209 528418 182261 528452
rect 178687 528409 178699 528418
rect 178751 528409 182261 528418
rect 182313 528409 182325 528461
rect 182377 528452 182389 528461
rect 182441 528452 182453 528461
rect 182441 528418 182451 528452
rect 182377 528409 182389 528418
rect 182441 528409 182453 528418
rect 182505 528409 182517 528461
rect 182569 528452 186079 528461
rect 182577 528418 182635 528452
rect 182669 528418 182727 528452
rect 182761 528418 182819 528452
rect 182853 528418 182911 528452
rect 182945 528418 183003 528452
rect 183037 528418 183095 528452
rect 183129 528418 183187 528452
rect 183221 528418 183279 528452
rect 183313 528418 183371 528452
rect 183405 528418 183463 528452
rect 183497 528418 183555 528452
rect 183589 528418 183647 528452
rect 183681 528418 183739 528452
rect 183773 528418 183831 528452
rect 183865 528418 183923 528452
rect 183957 528418 184015 528452
rect 184049 528418 184107 528452
rect 184141 528418 184199 528452
rect 184233 528418 184291 528452
rect 184325 528418 184383 528452
rect 184417 528418 184475 528452
rect 184509 528418 184567 528452
rect 184601 528418 184659 528452
rect 184693 528418 184751 528452
rect 184785 528418 184843 528452
rect 184877 528418 184935 528452
rect 184969 528418 185027 528452
rect 185061 528418 185119 528452
rect 185153 528418 185211 528452
rect 185245 528418 185303 528452
rect 185337 528418 185395 528452
rect 185429 528418 185487 528452
rect 185521 528418 185579 528452
rect 185613 528418 185671 528452
rect 185705 528418 185763 528452
rect 185797 528418 185855 528452
rect 185889 528418 185947 528452
rect 185981 528418 186039 528452
rect 186073 528418 186079 528452
rect 182569 528409 186079 528418
rect 186131 528452 186143 528461
rect 186131 528409 186143 528418
rect 186195 528409 186207 528461
rect 186259 528409 186271 528461
rect 186323 528452 186335 528461
rect 186387 528452 187482 528461
rect 186387 528418 186407 528452
rect 186441 528418 186499 528452
rect 186533 528418 186591 528452
rect 186625 528418 186683 528452
rect 186717 528418 186775 528452
rect 186809 528418 186867 528452
rect 186901 528418 186959 528452
rect 186993 528418 187051 528452
rect 187085 528418 187143 528452
rect 187177 528418 187235 528452
rect 187269 528418 187327 528452
rect 187361 528418 187419 528452
rect 187453 528418 187482 528452
rect 186323 528409 186335 528418
rect 186387 528409 187482 528418
rect 172210 528387 187482 528409
rect 176732 528307 176738 528359
rect 176790 528347 176796 528359
rect 177839 528350 177897 528356
rect 177839 528347 177851 528350
rect 176790 528319 177851 528347
rect 176790 528307 176796 528319
rect 177839 528316 177851 528319
rect 177885 528316 177897 528350
rect 177839 528310 177897 528316
rect 178020 528307 178026 528359
rect 178078 528307 178084 528359
rect 178940 528307 178946 528359
rect 178998 528307 179004 528359
rect 179308 528307 179314 528359
rect 179366 528347 179372 528359
rect 179403 528350 179461 528356
rect 179403 528347 179415 528350
rect 179366 528319 179415 528347
rect 179366 528307 179372 528319
rect 179403 528316 179415 528319
rect 179449 528316 179461 528350
rect 179403 528310 179461 528316
rect 180964 528307 180970 528359
rect 181022 528307 181028 528359
rect 181427 528350 181485 528356
rect 181427 528316 181439 528350
rect 181473 528347 181485 528350
rect 182160 528347 182166 528359
rect 181473 528319 182166 528347
rect 181473 528316 181485 528319
rect 181427 528310 181485 528316
rect 182160 528307 182166 528319
rect 182218 528307 182224 528359
rect 176364 528239 176370 528291
rect 176422 528239 176428 528291
rect 176824 528288 176830 528291
rect 176823 528242 176830 528288
rect 176882 528288 176888 528291
rect 176882 528282 176953 528288
rect 176882 528248 176907 528282
rect 176941 528279 176953 528282
rect 177543 528282 177601 528288
rect 177543 528279 177555 528282
rect 176941 528251 177555 528279
rect 176941 528248 176953 528251
rect 176824 528239 176830 528242
rect 176882 528242 176953 528248
rect 177483 528248 177555 528251
rect 177589 528248 177601 528282
rect 178038 528279 178066 528307
rect 178038 528251 179538 528279
rect 177483 528242 177601 528248
rect 176882 528239 176888 528242
rect 176088 528171 176094 528223
rect 176146 528171 176152 528223
rect 176184 528214 176242 528220
rect 176184 528180 176196 528214
rect 176230 528211 176242 528214
rect 176551 528214 176609 528220
rect 176551 528211 176563 528214
rect 176230 528183 176563 528211
rect 176230 528180 176242 528183
rect 176184 528174 176242 528180
rect 176551 528180 176563 528183
rect 176597 528211 176609 528214
rect 177267 528214 177325 528220
rect 177267 528211 177279 528214
rect 176597 528183 177279 528211
rect 176597 528180 176609 528183
rect 176551 528174 176609 528180
rect 177267 528180 177279 528183
rect 177313 528180 177325 528214
rect 177267 528174 177325 528180
rect 177483 528219 177541 528242
rect 177483 528185 177495 528219
rect 177529 528185 177541 528219
rect 177483 528179 177541 528185
rect 178112 528171 178118 528223
rect 178170 528171 178176 528223
rect 179311 528214 179369 528220
rect 179311 528180 179323 528214
rect 179357 528180 179369 528214
rect 179311 528174 179369 528180
rect 176265 528078 176323 528084
rect 176265 528044 176277 528078
rect 176311 528075 176323 528078
rect 176643 528078 176701 528084
rect 176643 528075 176655 528078
rect 176311 528047 176655 528075
rect 176311 528044 176323 528047
rect 176265 528038 176323 528044
rect 176643 528044 176655 528047
rect 176689 528075 176701 528078
rect 177267 528078 177325 528084
rect 177267 528075 177279 528078
rect 176689 528047 177279 528075
rect 176689 528044 176701 528047
rect 176643 528038 176701 528044
rect 177267 528044 177279 528047
rect 177313 528044 177325 528078
rect 177267 528038 177325 528044
rect 177376 528035 177382 528087
rect 177434 528075 177440 528087
rect 177931 528078 177989 528084
rect 177931 528075 177943 528078
rect 177434 528047 177943 528075
rect 177434 528035 177440 528047
rect 177931 528044 177943 528047
rect 177977 528044 177989 528078
rect 177931 528038 177989 528044
rect 178940 527967 178946 528019
rect 178998 528007 179004 528019
rect 179326 528007 179354 528174
rect 179510 528152 179538 528251
rect 181332 528171 181338 528223
rect 181390 528171 181396 528223
rect 179495 528146 179553 528152
rect 179495 528112 179507 528146
rect 179541 528143 179553 528146
rect 180688 528143 180694 528155
rect 179541 528115 180694 528143
rect 179541 528112 179553 528115
rect 179495 528106 179553 528112
rect 180688 528103 180694 528115
rect 180746 528143 180752 528155
rect 181519 528146 181577 528152
rect 181519 528143 181531 528146
rect 180746 528115 181531 528143
rect 180746 528103 180752 528115
rect 181519 528112 181531 528115
rect 181565 528112 181577 528146
rect 181519 528106 181577 528112
rect 178998 527979 179354 528007
rect 178998 527967 179004 527979
rect 172210 527917 187482 527939
rect 172210 527908 173965 527917
rect 174017 527908 174029 527917
rect 174081 527908 174093 527917
rect 172210 527874 172239 527908
rect 172273 527874 172331 527908
rect 172365 527874 172423 527908
rect 172457 527874 172515 527908
rect 172549 527874 172607 527908
rect 172641 527874 172699 527908
rect 172733 527874 172791 527908
rect 172825 527874 172883 527908
rect 172917 527874 172975 527908
rect 173009 527874 173067 527908
rect 173101 527874 173159 527908
rect 173193 527874 173251 527908
rect 173285 527874 173343 527908
rect 173377 527874 173435 527908
rect 173469 527874 173527 527908
rect 173561 527874 173619 527908
rect 173653 527874 173711 527908
rect 173745 527874 173803 527908
rect 173837 527874 173895 527908
rect 173929 527874 173965 527908
rect 174021 527874 174029 527908
rect 172210 527865 173965 527874
rect 174017 527865 174029 527874
rect 174081 527865 174093 527874
rect 174145 527865 174157 527917
rect 174209 527865 174221 527917
rect 174273 527908 177783 527917
rect 174297 527874 174355 527908
rect 174389 527874 174447 527908
rect 174481 527874 174539 527908
rect 174573 527874 174631 527908
rect 174665 527874 174723 527908
rect 174757 527874 174815 527908
rect 174849 527874 174907 527908
rect 174941 527874 174999 527908
rect 175033 527874 175091 527908
rect 175125 527874 175183 527908
rect 175217 527874 175275 527908
rect 175309 527874 175367 527908
rect 175401 527874 175459 527908
rect 175493 527874 175551 527908
rect 175585 527874 175643 527908
rect 175677 527874 175735 527908
rect 175769 527874 175827 527908
rect 175861 527874 175919 527908
rect 175953 527874 176011 527908
rect 176045 527874 176103 527908
rect 176137 527874 176195 527908
rect 176229 527874 176287 527908
rect 176321 527874 176379 527908
rect 176413 527874 176471 527908
rect 176505 527874 176563 527908
rect 176597 527874 176655 527908
rect 176689 527874 176747 527908
rect 176781 527874 176839 527908
rect 176873 527874 176931 527908
rect 176965 527874 177023 527908
rect 177057 527874 177115 527908
rect 177149 527874 177207 527908
rect 177241 527874 177299 527908
rect 177333 527874 177391 527908
rect 177425 527874 177483 527908
rect 177517 527874 177575 527908
rect 177609 527874 177667 527908
rect 177701 527874 177759 527908
rect 174273 527865 177783 527874
rect 177835 527865 177847 527917
rect 177899 527865 177911 527917
rect 177963 527908 177975 527917
rect 178027 527908 178039 527917
rect 178091 527908 181601 527917
rect 181653 527908 181665 527917
rect 181717 527908 181729 527917
rect 178027 527874 178035 527908
rect 178091 527874 178127 527908
rect 178161 527874 178219 527908
rect 178253 527874 178311 527908
rect 178345 527874 178403 527908
rect 178437 527874 178495 527908
rect 178529 527874 178587 527908
rect 178621 527874 178679 527908
rect 178713 527874 178771 527908
rect 178805 527874 178863 527908
rect 178897 527874 178955 527908
rect 178989 527874 179047 527908
rect 179081 527874 179139 527908
rect 179173 527874 179231 527908
rect 179265 527874 179323 527908
rect 179357 527874 179415 527908
rect 179449 527874 179507 527908
rect 179541 527874 179599 527908
rect 179633 527874 179691 527908
rect 179725 527874 179783 527908
rect 179817 527874 179875 527908
rect 179909 527874 179967 527908
rect 180001 527874 180059 527908
rect 180093 527874 180151 527908
rect 180185 527874 180243 527908
rect 180277 527874 180335 527908
rect 180369 527874 180427 527908
rect 180461 527874 180519 527908
rect 180553 527874 180611 527908
rect 180645 527874 180703 527908
rect 180737 527874 180795 527908
rect 180829 527874 180887 527908
rect 180921 527874 180979 527908
rect 181013 527874 181071 527908
rect 181105 527874 181163 527908
rect 181197 527874 181255 527908
rect 181289 527874 181347 527908
rect 181381 527874 181439 527908
rect 181473 527874 181531 527908
rect 181565 527874 181601 527908
rect 181657 527874 181665 527908
rect 177963 527865 177975 527874
rect 178027 527865 178039 527874
rect 178091 527865 181601 527874
rect 181653 527865 181665 527874
rect 181717 527865 181729 527874
rect 181781 527865 181793 527917
rect 181845 527865 181857 527917
rect 181909 527908 185419 527917
rect 181933 527874 181991 527908
rect 182025 527874 182083 527908
rect 182117 527874 182175 527908
rect 182209 527874 182267 527908
rect 182301 527874 182359 527908
rect 182393 527874 182451 527908
rect 182485 527874 182543 527908
rect 182577 527874 182635 527908
rect 182669 527874 182727 527908
rect 182761 527874 182819 527908
rect 182853 527874 182911 527908
rect 182945 527874 183003 527908
rect 183037 527874 183095 527908
rect 183129 527874 183187 527908
rect 183221 527874 183279 527908
rect 183313 527874 183371 527908
rect 183405 527874 183463 527908
rect 183497 527874 183555 527908
rect 183589 527874 183647 527908
rect 183681 527874 183739 527908
rect 183773 527874 183831 527908
rect 183865 527874 183923 527908
rect 183957 527874 184015 527908
rect 184049 527874 184107 527908
rect 184141 527874 184199 527908
rect 184233 527874 184291 527908
rect 184325 527874 184383 527908
rect 184417 527874 184475 527908
rect 184509 527874 184567 527908
rect 184601 527874 184659 527908
rect 184693 527874 184751 527908
rect 184785 527874 184843 527908
rect 184877 527874 184935 527908
rect 184969 527874 185027 527908
rect 185061 527874 185119 527908
rect 185153 527874 185211 527908
rect 185245 527874 185303 527908
rect 185337 527874 185395 527908
rect 181909 527865 185419 527874
rect 185471 527865 185483 527917
rect 185535 527865 185547 527917
rect 185599 527908 185611 527917
rect 185663 527908 185675 527917
rect 185727 527908 187482 527917
rect 185663 527874 185671 527908
rect 185727 527874 185763 527908
rect 185797 527874 185855 527908
rect 185889 527874 185947 527908
rect 185981 527874 186039 527908
rect 186073 527874 186131 527908
rect 186165 527874 186223 527908
rect 186257 527874 186315 527908
rect 186349 527874 186407 527908
rect 186441 527874 186499 527908
rect 186533 527874 186591 527908
rect 186625 527874 186683 527908
rect 186717 527874 186775 527908
rect 186809 527874 186867 527908
rect 186901 527874 186959 527908
rect 186993 527874 187051 527908
rect 187085 527874 187143 527908
rect 187177 527874 187235 527908
rect 187269 527874 187327 527908
rect 187361 527874 187419 527908
rect 187453 527874 187482 527908
rect 185599 527865 185611 527874
rect 185663 527865 185675 527874
rect 185727 527865 187482 527874
rect 172210 527843 187482 527865
rect 176272 527763 176278 527815
rect 176330 527803 176336 527815
rect 176367 527806 176425 527812
rect 176367 527803 176379 527806
rect 176330 527775 176379 527803
rect 176330 527763 176336 527775
rect 176367 527772 176379 527775
rect 176413 527772 176425 527806
rect 176367 527766 176425 527772
rect 178940 527763 178946 527815
rect 178998 527763 179004 527815
rect 177008 527627 177014 527679
rect 177066 527627 177072 527679
rect 179492 527627 179498 527679
rect 179550 527627 179556 527679
rect 172210 527373 187482 527395
rect 172210 527364 174625 527373
rect 172210 527330 172239 527364
rect 172273 527330 172331 527364
rect 172365 527330 172423 527364
rect 172457 527330 172515 527364
rect 172549 527330 172607 527364
rect 172641 527330 172699 527364
rect 172733 527330 172791 527364
rect 172825 527330 172883 527364
rect 172917 527330 172975 527364
rect 173009 527330 173067 527364
rect 173101 527330 173159 527364
rect 173193 527330 173251 527364
rect 173285 527330 173343 527364
rect 173377 527330 173435 527364
rect 173469 527330 173527 527364
rect 173561 527330 173619 527364
rect 173653 527330 173711 527364
rect 173745 527330 173803 527364
rect 173837 527330 173895 527364
rect 173929 527330 173987 527364
rect 174021 527330 174079 527364
rect 174113 527330 174171 527364
rect 174205 527330 174263 527364
rect 174297 527330 174355 527364
rect 174389 527330 174447 527364
rect 174481 527330 174539 527364
rect 174573 527330 174625 527364
rect 172210 527321 174625 527330
rect 174677 527321 174689 527373
rect 174741 527364 174753 527373
rect 174805 527364 174817 527373
rect 174805 527330 174815 527364
rect 174741 527321 174753 527330
rect 174805 527321 174817 527330
rect 174869 527321 174881 527373
rect 174933 527364 178443 527373
rect 174941 527330 174999 527364
rect 175033 527330 175091 527364
rect 175125 527330 175183 527364
rect 175217 527330 175275 527364
rect 175309 527330 175367 527364
rect 175401 527330 175459 527364
rect 175493 527330 175551 527364
rect 175585 527330 175643 527364
rect 175677 527330 175735 527364
rect 175769 527330 175827 527364
rect 175861 527330 175919 527364
rect 175953 527330 176011 527364
rect 176045 527330 176103 527364
rect 176137 527330 176195 527364
rect 176229 527330 176287 527364
rect 176321 527330 176379 527364
rect 176413 527330 176471 527364
rect 176505 527330 176563 527364
rect 176597 527330 176655 527364
rect 176689 527330 176747 527364
rect 176781 527330 176839 527364
rect 176873 527330 176931 527364
rect 176965 527330 177023 527364
rect 177057 527330 177115 527364
rect 177149 527330 177207 527364
rect 177241 527330 177299 527364
rect 177333 527330 177391 527364
rect 177425 527330 177483 527364
rect 177517 527330 177575 527364
rect 177609 527330 177667 527364
rect 177701 527330 177759 527364
rect 177793 527330 177851 527364
rect 177885 527330 177943 527364
rect 177977 527330 178035 527364
rect 178069 527330 178127 527364
rect 178161 527330 178219 527364
rect 178253 527330 178311 527364
rect 178345 527330 178403 527364
rect 178437 527330 178443 527364
rect 174933 527321 178443 527330
rect 178495 527364 178507 527373
rect 178495 527321 178507 527330
rect 178559 527321 178571 527373
rect 178623 527321 178635 527373
rect 178687 527364 178699 527373
rect 178751 527364 182261 527373
rect 178751 527330 178771 527364
rect 178805 527330 178863 527364
rect 178897 527330 178955 527364
rect 178989 527330 179047 527364
rect 179081 527330 179139 527364
rect 179173 527330 179231 527364
rect 179265 527330 179323 527364
rect 179357 527330 179415 527364
rect 179449 527330 179507 527364
rect 179541 527330 179599 527364
rect 179633 527330 179691 527364
rect 179725 527330 179783 527364
rect 179817 527330 179875 527364
rect 179909 527330 179967 527364
rect 180001 527330 180059 527364
rect 180093 527330 180151 527364
rect 180185 527330 180243 527364
rect 180277 527330 180335 527364
rect 180369 527330 180427 527364
rect 180461 527330 180519 527364
rect 180553 527330 180611 527364
rect 180645 527330 180703 527364
rect 180737 527330 180795 527364
rect 180829 527330 180887 527364
rect 180921 527330 180979 527364
rect 181013 527330 181071 527364
rect 181105 527330 181163 527364
rect 181197 527330 181255 527364
rect 181289 527330 181347 527364
rect 181381 527330 181439 527364
rect 181473 527330 181531 527364
rect 181565 527330 181623 527364
rect 181657 527330 181715 527364
rect 181749 527330 181807 527364
rect 181841 527330 181899 527364
rect 181933 527330 181991 527364
rect 182025 527330 182083 527364
rect 182117 527330 182175 527364
rect 182209 527330 182261 527364
rect 178687 527321 178699 527330
rect 178751 527321 182261 527330
rect 182313 527321 182325 527373
rect 182377 527364 182389 527373
rect 182441 527364 182453 527373
rect 182441 527330 182451 527364
rect 182377 527321 182389 527330
rect 182441 527321 182453 527330
rect 182505 527321 182517 527373
rect 182569 527364 186079 527373
rect 182577 527330 182635 527364
rect 182669 527330 182727 527364
rect 182761 527330 182819 527364
rect 182853 527330 182911 527364
rect 182945 527330 183003 527364
rect 183037 527330 183095 527364
rect 183129 527330 183187 527364
rect 183221 527330 183279 527364
rect 183313 527330 183371 527364
rect 183405 527330 183463 527364
rect 183497 527330 183555 527364
rect 183589 527330 183647 527364
rect 183681 527330 183739 527364
rect 183773 527330 183831 527364
rect 183865 527330 183923 527364
rect 183957 527330 184015 527364
rect 184049 527330 184107 527364
rect 184141 527330 184199 527364
rect 184233 527330 184291 527364
rect 184325 527330 184383 527364
rect 184417 527330 184475 527364
rect 184509 527330 184567 527364
rect 184601 527330 184659 527364
rect 184693 527330 184751 527364
rect 184785 527330 184843 527364
rect 184877 527330 184935 527364
rect 184969 527330 185027 527364
rect 185061 527330 185119 527364
rect 185153 527330 185211 527364
rect 185245 527330 185303 527364
rect 185337 527330 185395 527364
rect 185429 527330 185487 527364
rect 185521 527330 185579 527364
rect 185613 527330 185671 527364
rect 185705 527330 185763 527364
rect 185797 527330 185855 527364
rect 185889 527330 185947 527364
rect 185981 527330 186039 527364
rect 186073 527330 186079 527364
rect 182569 527321 186079 527330
rect 186131 527364 186143 527373
rect 186131 527321 186143 527330
rect 186195 527321 186207 527373
rect 186259 527321 186271 527373
rect 186323 527364 186335 527373
rect 186387 527364 187482 527373
rect 186387 527330 186407 527364
rect 186441 527330 186499 527364
rect 186533 527330 186591 527364
rect 186625 527330 186683 527364
rect 186717 527330 186775 527364
rect 186809 527330 186867 527364
rect 186901 527330 186959 527364
rect 186993 527330 187051 527364
rect 187085 527330 187143 527364
rect 187177 527330 187235 527364
rect 187269 527330 187327 527364
rect 187361 527330 187419 527364
rect 187453 527330 187482 527364
rect 186323 527321 186335 527330
rect 186387 527321 187482 527330
rect 172210 527299 187482 527321
rect 172210 526829 187482 526851
rect 172210 526820 173965 526829
rect 174017 526820 174029 526829
rect 174081 526820 174093 526829
rect 172210 526786 172239 526820
rect 172273 526786 172331 526820
rect 172365 526786 172423 526820
rect 172457 526786 172515 526820
rect 172549 526786 172607 526820
rect 172641 526786 172699 526820
rect 172733 526786 172791 526820
rect 172825 526786 172883 526820
rect 172917 526786 172975 526820
rect 173009 526786 173067 526820
rect 173101 526786 173159 526820
rect 173193 526786 173251 526820
rect 173285 526786 173343 526820
rect 173377 526786 173435 526820
rect 173469 526786 173527 526820
rect 173561 526786 173619 526820
rect 173653 526786 173711 526820
rect 173745 526786 173803 526820
rect 173837 526786 173895 526820
rect 173929 526786 173965 526820
rect 174021 526786 174029 526820
rect 172210 526777 173965 526786
rect 174017 526777 174029 526786
rect 174081 526777 174093 526786
rect 174145 526777 174157 526829
rect 174209 526777 174221 526829
rect 174273 526820 177783 526829
rect 174297 526786 174355 526820
rect 174389 526786 174447 526820
rect 174481 526786 174539 526820
rect 174573 526786 174631 526820
rect 174665 526786 174723 526820
rect 174757 526786 174815 526820
rect 174849 526786 174907 526820
rect 174941 526786 174999 526820
rect 175033 526786 175091 526820
rect 175125 526786 175183 526820
rect 175217 526786 175275 526820
rect 175309 526786 175367 526820
rect 175401 526786 175459 526820
rect 175493 526786 175551 526820
rect 175585 526786 175643 526820
rect 175677 526786 175735 526820
rect 175769 526786 175827 526820
rect 175861 526786 175919 526820
rect 175953 526786 176011 526820
rect 176045 526786 176103 526820
rect 176137 526786 176195 526820
rect 176229 526786 176287 526820
rect 176321 526786 176379 526820
rect 176413 526786 176471 526820
rect 176505 526786 176563 526820
rect 176597 526786 176655 526820
rect 176689 526786 176747 526820
rect 176781 526786 176839 526820
rect 176873 526786 176931 526820
rect 176965 526786 177023 526820
rect 177057 526786 177115 526820
rect 177149 526786 177207 526820
rect 177241 526786 177299 526820
rect 177333 526786 177391 526820
rect 177425 526786 177483 526820
rect 177517 526786 177575 526820
rect 177609 526786 177667 526820
rect 177701 526786 177759 526820
rect 174273 526777 177783 526786
rect 177835 526777 177847 526829
rect 177899 526777 177911 526829
rect 177963 526820 177975 526829
rect 178027 526820 178039 526829
rect 178091 526820 181601 526829
rect 181653 526820 181665 526829
rect 181717 526820 181729 526829
rect 178027 526786 178035 526820
rect 178091 526786 178127 526820
rect 178161 526786 178219 526820
rect 178253 526786 178311 526820
rect 178345 526786 178403 526820
rect 178437 526786 178495 526820
rect 178529 526786 178587 526820
rect 178621 526786 178679 526820
rect 178713 526786 178771 526820
rect 178805 526786 178863 526820
rect 178897 526786 178955 526820
rect 178989 526786 179047 526820
rect 179081 526786 179139 526820
rect 179173 526786 179231 526820
rect 179265 526786 179323 526820
rect 179357 526786 179415 526820
rect 179449 526786 179507 526820
rect 179541 526786 179599 526820
rect 179633 526786 179691 526820
rect 179725 526786 179783 526820
rect 179817 526786 179875 526820
rect 179909 526786 179967 526820
rect 180001 526786 180059 526820
rect 180093 526786 180151 526820
rect 180185 526786 180243 526820
rect 180277 526786 180335 526820
rect 180369 526786 180427 526820
rect 180461 526786 180519 526820
rect 180553 526786 180611 526820
rect 180645 526786 180703 526820
rect 180737 526786 180795 526820
rect 180829 526786 180887 526820
rect 180921 526786 180979 526820
rect 181013 526786 181071 526820
rect 181105 526786 181163 526820
rect 181197 526786 181255 526820
rect 181289 526786 181347 526820
rect 181381 526786 181439 526820
rect 181473 526786 181531 526820
rect 181565 526786 181601 526820
rect 181657 526786 181665 526820
rect 177963 526777 177975 526786
rect 178027 526777 178039 526786
rect 178091 526777 181601 526786
rect 181653 526777 181665 526786
rect 181717 526777 181729 526786
rect 181781 526777 181793 526829
rect 181845 526777 181857 526829
rect 181909 526820 185419 526829
rect 181933 526786 181991 526820
rect 182025 526786 182083 526820
rect 182117 526786 182175 526820
rect 182209 526786 182267 526820
rect 182301 526786 182359 526820
rect 182393 526786 182451 526820
rect 182485 526786 182543 526820
rect 182577 526786 182635 526820
rect 182669 526786 182727 526820
rect 182761 526786 182819 526820
rect 182853 526786 182911 526820
rect 182945 526786 183003 526820
rect 183037 526786 183095 526820
rect 183129 526786 183187 526820
rect 183221 526786 183279 526820
rect 183313 526786 183371 526820
rect 183405 526786 183463 526820
rect 183497 526786 183555 526820
rect 183589 526786 183647 526820
rect 183681 526786 183739 526820
rect 183773 526786 183831 526820
rect 183865 526786 183923 526820
rect 183957 526786 184015 526820
rect 184049 526786 184107 526820
rect 184141 526786 184199 526820
rect 184233 526786 184291 526820
rect 184325 526786 184383 526820
rect 184417 526786 184475 526820
rect 184509 526786 184567 526820
rect 184601 526786 184659 526820
rect 184693 526786 184751 526820
rect 184785 526786 184843 526820
rect 184877 526786 184935 526820
rect 184969 526786 185027 526820
rect 185061 526786 185119 526820
rect 185153 526786 185211 526820
rect 185245 526786 185303 526820
rect 185337 526786 185395 526820
rect 181909 526777 185419 526786
rect 185471 526777 185483 526829
rect 185535 526777 185547 526829
rect 185599 526820 185611 526829
rect 185663 526820 185675 526829
rect 185727 526820 187482 526829
rect 185663 526786 185671 526820
rect 185727 526786 185763 526820
rect 185797 526786 185855 526820
rect 185889 526786 185947 526820
rect 185981 526786 186039 526820
rect 186073 526786 186131 526820
rect 186165 526786 186223 526820
rect 186257 526786 186315 526820
rect 186349 526786 186407 526820
rect 186441 526786 186499 526820
rect 186533 526786 186591 526820
rect 186625 526786 186683 526820
rect 186717 526786 186775 526820
rect 186809 526786 186867 526820
rect 186901 526786 186959 526820
rect 186993 526786 187051 526820
rect 187085 526786 187143 526820
rect 187177 526786 187235 526820
rect 187269 526786 187327 526820
rect 187361 526786 187419 526820
rect 187453 526786 187482 526820
rect 185599 526777 185611 526786
rect 185663 526777 185675 526786
rect 185727 526777 187482 526786
rect 172210 526755 187482 526777
rect 172210 526285 187482 526307
rect 172210 526276 174625 526285
rect 172210 526242 172239 526276
rect 172273 526242 172331 526276
rect 172365 526242 172423 526276
rect 172457 526242 172515 526276
rect 172549 526242 172607 526276
rect 172641 526242 172699 526276
rect 172733 526242 172791 526276
rect 172825 526242 172883 526276
rect 172917 526242 172975 526276
rect 173009 526242 173067 526276
rect 173101 526242 173159 526276
rect 173193 526242 173251 526276
rect 173285 526242 173343 526276
rect 173377 526242 173435 526276
rect 173469 526242 173527 526276
rect 173561 526242 173619 526276
rect 173653 526242 173711 526276
rect 173745 526242 173803 526276
rect 173837 526242 173895 526276
rect 173929 526242 173987 526276
rect 174021 526242 174079 526276
rect 174113 526242 174171 526276
rect 174205 526242 174263 526276
rect 174297 526242 174355 526276
rect 174389 526242 174447 526276
rect 174481 526242 174539 526276
rect 174573 526242 174625 526276
rect 172210 526233 174625 526242
rect 174677 526233 174689 526285
rect 174741 526276 174753 526285
rect 174805 526276 174817 526285
rect 174805 526242 174815 526276
rect 174741 526233 174753 526242
rect 174805 526233 174817 526242
rect 174869 526233 174881 526285
rect 174933 526276 178443 526285
rect 174941 526242 174999 526276
rect 175033 526242 175091 526276
rect 175125 526242 175183 526276
rect 175217 526242 175275 526276
rect 175309 526242 175367 526276
rect 175401 526242 175459 526276
rect 175493 526242 175551 526276
rect 175585 526242 175643 526276
rect 175677 526242 175735 526276
rect 175769 526242 175827 526276
rect 175861 526242 175919 526276
rect 175953 526242 176011 526276
rect 176045 526242 176103 526276
rect 176137 526242 176195 526276
rect 176229 526242 176287 526276
rect 176321 526242 176379 526276
rect 176413 526242 176471 526276
rect 176505 526242 176563 526276
rect 176597 526242 176655 526276
rect 176689 526242 176747 526276
rect 176781 526242 176839 526276
rect 176873 526242 176931 526276
rect 176965 526242 177023 526276
rect 177057 526242 177115 526276
rect 177149 526242 177207 526276
rect 177241 526242 177299 526276
rect 177333 526242 177391 526276
rect 177425 526242 177483 526276
rect 177517 526242 177575 526276
rect 177609 526242 177667 526276
rect 177701 526242 177759 526276
rect 177793 526242 177851 526276
rect 177885 526242 177943 526276
rect 177977 526242 178035 526276
rect 178069 526242 178127 526276
rect 178161 526242 178219 526276
rect 178253 526242 178311 526276
rect 178345 526242 178403 526276
rect 178437 526242 178443 526276
rect 174933 526233 178443 526242
rect 178495 526276 178507 526285
rect 178495 526233 178507 526242
rect 178559 526233 178571 526285
rect 178623 526233 178635 526285
rect 178687 526276 178699 526285
rect 178751 526276 182261 526285
rect 178751 526242 178771 526276
rect 178805 526242 178863 526276
rect 178897 526242 178955 526276
rect 178989 526242 179047 526276
rect 179081 526242 179139 526276
rect 179173 526242 179231 526276
rect 179265 526242 179323 526276
rect 179357 526242 179415 526276
rect 179449 526242 179507 526276
rect 179541 526242 179599 526276
rect 179633 526242 179691 526276
rect 179725 526242 179783 526276
rect 179817 526242 179875 526276
rect 179909 526242 179967 526276
rect 180001 526242 180059 526276
rect 180093 526242 180151 526276
rect 180185 526242 180243 526276
rect 180277 526242 180335 526276
rect 180369 526242 180427 526276
rect 180461 526242 180519 526276
rect 180553 526242 180611 526276
rect 180645 526242 180703 526276
rect 180737 526242 180795 526276
rect 180829 526242 180887 526276
rect 180921 526242 180979 526276
rect 181013 526242 181071 526276
rect 181105 526242 181163 526276
rect 181197 526242 181255 526276
rect 181289 526242 181347 526276
rect 181381 526242 181439 526276
rect 181473 526242 181531 526276
rect 181565 526242 181623 526276
rect 181657 526242 181715 526276
rect 181749 526242 181807 526276
rect 181841 526242 181899 526276
rect 181933 526242 181991 526276
rect 182025 526242 182083 526276
rect 182117 526242 182175 526276
rect 182209 526242 182261 526276
rect 178687 526233 178699 526242
rect 178751 526233 182261 526242
rect 182313 526233 182325 526285
rect 182377 526276 182389 526285
rect 182441 526276 182453 526285
rect 182441 526242 182451 526276
rect 182377 526233 182389 526242
rect 182441 526233 182453 526242
rect 182505 526233 182517 526285
rect 182569 526276 186079 526285
rect 182577 526242 182635 526276
rect 182669 526242 182727 526276
rect 182761 526242 182819 526276
rect 182853 526242 182911 526276
rect 182945 526242 183003 526276
rect 183037 526242 183095 526276
rect 183129 526242 183187 526276
rect 183221 526242 183279 526276
rect 183313 526242 183371 526276
rect 183405 526242 183463 526276
rect 183497 526242 183555 526276
rect 183589 526242 183647 526276
rect 183681 526242 183739 526276
rect 183773 526242 183831 526276
rect 183865 526242 183923 526276
rect 183957 526242 184015 526276
rect 184049 526242 184107 526276
rect 184141 526242 184199 526276
rect 184233 526242 184291 526276
rect 184325 526242 184383 526276
rect 184417 526242 184475 526276
rect 184509 526242 184567 526276
rect 184601 526242 184659 526276
rect 184693 526242 184751 526276
rect 184785 526242 184843 526276
rect 184877 526242 184935 526276
rect 184969 526242 185027 526276
rect 185061 526242 185119 526276
rect 185153 526242 185211 526276
rect 185245 526242 185303 526276
rect 185337 526242 185395 526276
rect 185429 526242 185487 526276
rect 185521 526242 185579 526276
rect 185613 526242 185671 526276
rect 185705 526242 185763 526276
rect 185797 526242 185855 526276
rect 185889 526242 185947 526276
rect 185981 526242 186039 526276
rect 186073 526242 186079 526276
rect 182569 526233 186079 526242
rect 186131 526276 186143 526285
rect 186131 526233 186143 526242
rect 186195 526233 186207 526285
rect 186259 526233 186271 526285
rect 186323 526276 186335 526285
rect 186387 526276 187482 526285
rect 186387 526242 186407 526276
rect 186441 526242 186499 526276
rect 186533 526242 186591 526276
rect 186625 526242 186683 526276
rect 186717 526242 186775 526276
rect 186809 526242 186867 526276
rect 186901 526242 186959 526276
rect 186993 526242 187051 526276
rect 187085 526242 187143 526276
rect 187177 526242 187235 526276
rect 187269 526242 187327 526276
rect 187361 526242 187419 526276
rect 187453 526242 187482 526276
rect 186323 526233 186335 526242
rect 186387 526233 187482 526242
rect 172210 526211 187482 526233
rect 172210 525741 187482 525763
rect 172210 525732 173965 525741
rect 174017 525732 174029 525741
rect 174081 525732 174093 525741
rect 172210 525698 172239 525732
rect 172273 525698 172331 525732
rect 172365 525698 172423 525732
rect 172457 525698 172515 525732
rect 172549 525698 172607 525732
rect 172641 525698 172699 525732
rect 172733 525698 172791 525732
rect 172825 525698 172883 525732
rect 172917 525698 172975 525732
rect 173009 525698 173067 525732
rect 173101 525698 173159 525732
rect 173193 525698 173251 525732
rect 173285 525698 173343 525732
rect 173377 525698 173435 525732
rect 173469 525698 173527 525732
rect 173561 525698 173619 525732
rect 173653 525698 173711 525732
rect 173745 525698 173803 525732
rect 173837 525698 173895 525732
rect 173929 525698 173965 525732
rect 174021 525698 174029 525732
rect 172210 525689 173965 525698
rect 174017 525689 174029 525698
rect 174081 525689 174093 525698
rect 174145 525689 174157 525741
rect 174209 525689 174221 525741
rect 174273 525732 177783 525741
rect 174297 525698 174355 525732
rect 174389 525698 174447 525732
rect 174481 525698 174539 525732
rect 174573 525698 174631 525732
rect 174665 525698 174723 525732
rect 174757 525698 174815 525732
rect 174849 525698 174907 525732
rect 174941 525698 174999 525732
rect 175033 525698 175091 525732
rect 175125 525698 175183 525732
rect 175217 525698 175275 525732
rect 175309 525698 175367 525732
rect 175401 525698 175459 525732
rect 175493 525698 175551 525732
rect 175585 525698 175643 525732
rect 175677 525698 175735 525732
rect 175769 525698 175827 525732
rect 175861 525698 175919 525732
rect 175953 525698 176011 525732
rect 176045 525698 176103 525732
rect 176137 525698 176195 525732
rect 176229 525698 176287 525732
rect 176321 525698 176379 525732
rect 176413 525698 176471 525732
rect 176505 525698 176563 525732
rect 176597 525698 176655 525732
rect 176689 525698 176747 525732
rect 176781 525698 176839 525732
rect 176873 525698 176931 525732
rect 176965 525698 177023 525732
rect 177057 525698 177115 525732
rect 177149 525698 177207 525732
rect 177241 525698 177299 525732
rect 177333 525698 177391 525732
rect 177425 525698 177483 525732
rect 177517 525698 177575 525732
rect 177609 525698 177667 525732
rect 177701 525698 177759 525732
rect 174273 525689 177783 525698
rect 177835 525689 177847 525741
rect 177899 525689 177911 525741
rect 177963 525732 177975 525741
rect 178027 525732 178039 525741
rect 178091 525732 181601 525741
rect 181653 525732 181665 525741
rect 181717 525732 181729 525741
rect 178027 525698 178035 525732
rect 178091 525698 178127 525732
rect 178161 525698 178219 525732
rect 178253 525698 178311 525732
rect 178345 525698 178403 525732
rect 178437 525698 178495 525732
rect 178529 525698 178587 525732
rect 178621 525698 178679 525732
rect 178713 525698 178771 525732
rect 178805 525698 178863 525732
rect 178897 525698 178955 525732
rect 178989 525698 179047 525732
rect 179081 525698 179139 525732
rect 179173 525698 179231 525732
rect 179265 525698 179323 525732
rect 179357 525698 179415 525732
rect 179449 525698 179507 525732
rect 179541 525698 179599 525732
rect 179633 525698 179691 525732
rect 179725 525698 179783 525732
rect 179817 525698 179875 525732
rect 179909 525698 179967 525732
rect 180001 525698 180059 525732
rect 180093 525698 180151 525732
rect 180185 525698 180243 525732
rect 180277 525698 180335 525732
rect 180369 525698 180427 525732
rect 180461 525698 180519 525732
rect 180553 525698 180611 525732
rect 180645 525698 180703 525732
rect 180737 525698 180795 525732
rect 180829 525698 180887 525732
rect 180921 525698 180979 525732
rect 181013 525698 181071 525732
rect 181105 525698 181163 525732
rect 181197 525698 181255 525732
rect 181289 525698 181347 525732
rect 181381 525698 181439 525732
rect 181473 525698 181531 525732
rect 181565 525698 181601 525732
rect 181657 525698 181665 525732
rect 177963 525689 177975 525698
rect 178027 525689 178039 525698
rect 178091 525689 181601 525698
rect 181653 525689 181665 525698
rect 181717 525689 181729 525698
rect 181781 525689 181793 525741
rect 181845 525689 181857 525741
rect 181909 525732 185419 525741
rect 181933 525698 181991 525732
rect 182025 525698 182083 525732
rect 182117 525698 182175 525732
rect 182209 525698 182267 525732
rect 182301 525698 182359 525732
rect 182393 525698 182451 525732
rect 182485 525698 182543 525732
rect 182577 525698 182635 525732
rect 182669 525698 182727 525732
rect 182761 525698 182819 525732
rect 182853 525698 182911 525732
rect 182945 525698 183003 525732
rect 183037 525698 183095 525732
rect 183129 525698 183187 525732
rect 183221 525698 183279 525732
rect 183313 525698 183371 525732
rect 183405 525698 183463 525732
rect 183497 525698 183555 525732
rect 183589 525698 183647 525732
rect 183681 525698 183739 525732
rect 183773 525698 183831 525732
rect 183865 525698 183923 525732
rect 183957 525698 184015 525732
rect 184049 525698 184107 525732
rect 184141 525698 184199 525732
rect 184233 525698 184291 525732
rect 184325 525698 184383 525732
rect 184417 525698 184475 525732
rect 184509 525698 184567 525732
rect 184601 525698 184659 525732
rect 184693 525698 184751 525732
rect 184785 525698 184843 525732
rect 184877 525698 184935 525732
rect 184969 525698 185027 525732
rect 185061 525698 185119 525732
rect 185153 525698 185211 525732
rect 185245 525698 185303 525732
rect 185337 525698 185395 525732
rect 181909 525689 185419 525698
rect 185471 525689 185483 525741
rect 185535 525689 185547 525741
rect 185599 525732 185611 525741
rect 185663 525732 185675 525741
rect 185727 525732 187482 525741
rect 185663 525698 185671 525732
rect 185727 525698 185763 525732
rect 185797 525698 185855 525732
rect 185889 525698 185947 525732
rect 185981 525698 186039 525732
rect 186073 525698 186131 525732
rect 186165 525698 186223 525732
rect 186257 525698 186315 525732
rect 186349 525698 186407 525732
rect 186441 525698 186499 525732
rect 186533 525698 186591 525732
rect 186625 525698 186683 525732
rect 186717 525698 186775 525732
rect 186809 525698 186867 525732
rect 186901 525698 186959 525732
rect 186993 525698 187051 525732
rect 187085 525698 187143 525732
rect 187177 525698 187235 525732
rect 187269 525698 187327 525732
rect 187361 525698 187419 525732
rect 187453 525698 187482 525732
rect 185599 525689 185611 525698
rect 185663 525689 185675 525698
rect 185727 525689 187482 525698
rect 172210 525667 187482 525689
rect 172210 525197 187482 525219
rect 172210 525188 174625 525197
rect 172210 525154 172239 525188
rect 172273 525154 172331 525188
rect 172365 525154 172423 525188
rect 172457 525154 172515 525188
rect 172549 525154 172607 525188
rect 172641 525154 172699 525188
rect 172733 525154 172791 525188
rect 172825 525154 172883 525188
rect 172917 525154 172975 525188
rect 173009 525154 173067 525188
rect 173101 525154 173159 525188
rect 173193 525154 173251 525188
rect 173285 525154 173343 525188
rect 173377 525154 173435 525188
rect 173469 525154 173527 525188
rect 173561 525154 173619 525188
rect 173653 525154 173711 525188
rect 173745 525154 173803 525188
rect 173837 525154 173895 525188
rect 173929 525154 173987 525188
rect 174021 525154 174079 525188
rect 174113 525154 174171 525188
rect 174205 525154 174263 525188
rect 174297 525154 174355 525188
rect 174389 525154 174447 525188
rect 174481 525154 174539 525188
rect 174573 525154 174625 525188
rect 172210 525145 174625 525154
rect 174677 525145 174689 525197
rect 174741 525188 174753 525197
rect 174805 525188 174817 525197
rect 174805 525154 174815 525188
rect 174741 525145 174753 525154
rect 174805 525145 174817 525154
rect 174869 525145 174881 525197
rect 174933 525188 178443 525197
rect 174941 525154 174999 525188
rect 175033 525154 175091 525188
rect 175125 525154 175183 525188
rect 175217 525154 175275 525188
rect 175309 525154 175367 525188
rect 175401 525154 175459 525188
rect 175493 525154 175551 525188
rect 175585 525154 175643 525188
rect 175677 525154 175735 525188
rect 175769 525154 175827 525188
rect 175861 525154 175919 525188
rect 175953 525154 176011 525188
rect 176045 525154 176103 525188
rect 176137 525154 176195 525188
rect 176229 525154 176287 525188
rect 176321 525154 176379 525188
rect 176413 525154 176471 525188
rect 176505 525154 176563 525188
rect 176597 525154 176655 525188
rect 176689 525154 176747 525188
rect 176781 525154 176839 525188
rect 176873 525154 176931 525188
rect 176965 525154 177023 525188
rect 177057 525154 177115 525188
rect 177149 525154 177207 525188
rect 177241 525154 177299 525188
rect 177333 525154 177391 525188
rect 177425 525154 177483 525188
rect 177517 525154 177575 525188
rect 177609 525154 177667 525188
rect 177701 525154 177759 525188
rect 177793 525154 177851 525188
rect 177885 525154 177943 525188
rect 177977 525154 178035 525188
rect 178069 525154 178127 525188
rect 178161 525154 178219 525188
rect 178253 525154 178311 525188
rect 178345 525154 178403 525188
rect 178437 525154 178443 525188
rect 174933 525145 178443 525154
rect 178495 525188 178507 525197
rect 178495 525145 178507 525154
rect 178559 525145 178571 525197
rect 178623 525145 178635 525197
rect 178687 525188 178699 525197
rect 178751 525188 182261 525197
rect 178751 525154 178771 525188
rect 178805 525154 178863 525188
rect 178897 525154 178955 525188
rect 178989 525154 179047 525188
rect 179081 525154 179139 525188
rect 179173 525154 179231 525188
rect 179265 525154 179323 525188
rect 179357 525154 179415 525188
rect 179449 525154 179507 525188
rect 179541 525154 179599 525188
rect 179633 525154 179691 525188
rect 179725 525154 179783 525188
rect 179817 525154 179875 525188
rect 179909 525154 179967 525188
rect 180001 525154 180059 525188
rect 180093 525154 180151 525188
rect 180185 525154 180243 525188
rect 180277 525154 180335 525188
rect 180369 525154 180427 525188
rect 180461 525154 180519 525188
rect 180553 525154 180611 525188
rect 180645 525154 180703 525188
rect 180737 525154 180795 525188
rect 180829 525154 180887 525188
rect 180921 525154 180979 525188
rect 181013 525154 181071 525188
rect 181105 525154 181163 525188
rect 181197 525154 181255 525188
rect 181289 525154 181347 525188
rect 181381 525154 181439 525188
rect 181473 525154 181531 525188
rect 181565 525154 181623 525188
rect 181657 525154 181715 525188
rect 181749 525154 181807 525188
rect 181841 525154 181899 525188
rect 181933 525154 181991 525188
rect 182025 525154 182083 525188
rect 182117 525154 182175 525188
rect 182209 525154 182261 525188
rect 178687 525145 178699 525154
rect 178751 525145 182261 525154
rect 182313 525145 182325 525197
rect 182377 525188 182389 525197
rect 182441 525188 182453 525197
rect 182441 525154 182451 525188
rect 182377 525145 182389 525154
rect 182441 525145 182453 525154
rect 182505 525145 182517 525197
rect 182569 525188 186079 525197
rect 182577 525154 182635 525188
rect 182669 525154 182727 525188
rect 182761 525154 182819 525188
rect 182853 525154 182911 525188
rect 182945 525154 183003 525188
rect 183037 525154 183095 525188
rect 183129 525154 183187 525188
rect 183221 525154 183279 525188
rect 183313 525154 183371 525188
rect 183405 525154 183463 525188
rect 183497 525154 183555 525188
rect 183589 525154 183647 525188
rect 183681 525154 183739 525188
rect 183773 525154 183831 525188
rect 183865 525154 183923 525188
rect 183957 525154 184015 525188
rect 184049 525154 184107 525188
rect 184141 525154 184199 525188
rect 184233 525154 184291 525188
rect 184325 525154 184383 525188
rect 184417 525154 184475 525188
rect 184509 525154 184567 525188
rect 184601 525154 184659 525188
rect 184693 525154 184751 525188
rect 184785 525154 184843 525188
rect 184877 525154 184935 525188
rect 184969 525154 185027 525188
rect 185061 525154 185119 525188
rect 185153 525154 185211 525188
rect 185245 525154 185303 525188
rect 185337 525154 185395 525188
rect 185429 525154 185487 525188
rect 185521 525154 185579 525188
rect 185613 525154 185671 525188
rect 185705 525154 185763 525188
rect 185797 525154 185855 525188
rect 185889 525154 185947 525188
rect 185981 525154 186039 525188
rect 186073 525154 186079 525188
rect 182569 525145 186079 525154
rect 186131 525188 186143 525197
rect 186131 525145 186143 525154
rect 186195 525145 186207 525197
rect 186259 525145 186271 525197
rect 186323 525188 186335 525197
rect 186387 525188 187482 525197
rect 186387 525154 186407 525188
rect 186441 525154 186499 525188
rect 186533 525154 186591 525188
rect 186625 525154 186683 525188
rect 186717 525154 186775 525188
rect 186809 525154 186867 525188
rect 186901 525154 186959 525188
rect 186993 525154 187051 525188
rect 187085 525154 187143 525188
rect 187177 525154 187235 525188
rect 187269 525154 187327 525188
rect 187361 525154 187419 525188
rect 187453 525154 187482 525188
rect 186323 525145 186335 525154
rect 186387 525145 187482 525154
rect 172210 525123 187482 525145
rect 172210 524653 187482 524675
rect 172210 524644 173965 524653
rect 174017 524644 174029 524653
rect 174081 524644 174093 524653
rect 172210 524610 172239 524644
rect 172273 524610 172331 524644
rect 172365 524610 172423 524644
rect 172457 524610 172515 524644
rect 172549 524610 172607 524644
rect 172641 524610 172699 524644
rect 172733 524610 172791 524644
rect 172825 524610 172883 524644
rect 172917 524610 172975 524644
rect 173009 524610 173067 524644
rect 173101 524610 173159 524644
rect 173193 524610 173251 524644
rect 173285 524610 173343 524644
rect 173377 524610 173435 524644
rect 173469 524610 173527 524644
rect 173561 524610 173619 524644
rect 173653 524610 173711 524644
rect 173745 524610 173803 524644
rect 173837 524610 173895 524644
rect 173929 524610 173965 524644
rect 174021 524610 174029 524644
rect 172210 524601 173965 524610
rect 174017 524601 174029 524610
rect 174081 524601 174093 524610
rect 174145 524601 174157 524653
rect 174209 524601 174221 524653
rect 174273 524644 177783 524653
rect 174297 524610 174355 524644
rect 174389 524610 174447 524644
rect 174481 524610 174539 524644
rect 174573 524610 174631 524644
rect 174665 524610 174723 524644
rect 174757 524610 174815 524644
rect 174849 524610 174907 524644
rect 174941 524610 174999 524644
rect 175033 524610 175091 524644
rect 175125 524610 175183 524644
rect 175217 524610 175275 524644
rect 175309 524610 175367 524644
rect 175401 524610 175459 524644
rect 175493 524610 175551 524644
rect 175585 524610 175643 524644
rect 175677 524610 175735 524644
rect 175769 524610 175827 524644
rect 175861 524610 175919 524644
rect 175953 524610 176011 524644
rect 176045 524610 176103 524644
rect 176137 524610 176195 524644
rect 176229 524610 176287 524644
rect 176321 524610 176379 524644
rect 176413 524610 176471 524644
rect 176505 524610 176563 524644
rect 176597 524610 176655 524644
rect 176689 524610 176747 524644
rect 176781 524610 176839 524644
rect 176873 524610 176931 524644
rect 176965 524610 177023 524644
rect 177057 524610 177115 524644
rect 177149 524610 177207 524644
rect 177241 524610 177299 524644
rect 177333 524610 177391 524644
rect 177425 524610 177483 524644
rect 177517 524610 177575 524644
rect 177609 524610 177667 524644
rect 177701 524610 177759 524644
rect 174273 524601 177783 524610
rect 177835 524601 177847 524653
rect 177899 524601 177911 524653
rect 177963 524644 177975 524653
rect 178027 524644 178039 524653
rect 178091 524644 181601 524653
rect 181653 524644 181665 524653
rect 181717 524644 181729 524653
rect 178027 524610 178035 524644
rect 178091 524610 178127 524644
rect 178161 524610 178219 524644
rect 178253 524610 178311 524644
rect 178345 524610 178403 524644
rect 178437 524610 178495 524644
rect 178529 524610 178587 524644
rect 178621 524610 178679 524644
rect 178713 524610 178771 524644
rect 178805 524610 178863 524644
rect 178897 524610 178955 524644
rect 178989 524610 179047 524644
rect 179081 524610 179139 524644
rect 179173 524610 179231 524644
rect 179265 524610 179323 524644
rect 179357 524610 179415 524644
rect 179449 524610 179507 524644
rect 179541 524610 179599 524644
rect 179633 524610 179691 524644
rect 179725 524610 179783 524644
rect 179817 524610 179875 524644
rect 179909 524610 179967 524644
rect 180001 524610 180059 524644
rect 180093 524610 180151 524644
rect 180185 524610 180243 524644
rect 180277 524610 180335 524644
rect 180369 524610 180427 524644
rect 180461 524610 180519 524644
rect 180553 524610 180611 524644
rect 180645 524610 180703 524644
rect 180737 524610 180795 524644
rect 180829 524610 180887 524644
rect 180921 524610 180979 524644
rect 181013 524610 181071 524644
rect 181105 524610 181163 524644
rect 181197 524610 181255 524644
rect 181289 524610 181347 524644
rect 181381 524610 181439 524644
rect 181473 524610 181531 524644
rect 181565 524610 181601 524644
rect 181657 524610 181665 524644
rect 177963 524601 177975 524610
rect 178027 524601 178039 524610
rect 178091 524601 181601 524610
rect 181653 524601 181665 524610
rect 181717 524601 181729 524610
rect 181781 524601 181793 524653
rect 181845 524601 181857 524653
rect 181909 524644 185419 524653
rect 181933 524610 181991 524644
rect 182025 524610 182083 524644
rect 182117 524610 182175 524644
rect 182209 524610 182267 524644
rect 182301 524610 182359 524644
rect 182393 524610 182451 524644
rect 182485 524610 182543 524644
rect 182577 524610 182635 524644
rect 182669 524610 182727 524644
rect 182761 524610 182819 524644
rect 182853 524610 182911 524644
rect 182945 524610 183003 524644
rect 183037 524610 183095 524644
rect 183129 524610 183187 524644
rect 183221 524610 183279 524644
rect 183313 524610 183371 524644
rect 183405 524610 183463 524644
rect 183497 524610 183555 524644
rect 183589 524610 183647 524644
rect 183681 524610 183739 524644
rect 183773 524610 183831 524644
rect 183865 524610 183923 524644
rect 183957 524610 184015 524644
rect 184049 524610 184107 524644
rect 184141 524610 184199 524644
rect 184233 524610 184291 524644
rect 184325 524610 184383 524644
rect 184417 524610 184475 524644
rect 184509 524610 184567 524644
rect 184601 524610 184659 524644
rect 184693 524610 184751 524644
rect 184785 524610 184843 524644
rect 184877 524610 184935 524644
rect 184969 524610 185027 524644
rect 185061 524610 185119 524644
rect 185153 524610 185211 524644
rect 185245 524610 185303 524644
rect 185337 524610 185395 524644
rect 181909 524601 185419 524610
rect 185471 524601 185483 524653
rect 185535 524601 185547 524653
rect 185599 524644 185611 524653
rect 185663 524644 185675 524653
rect 185727 524644 187482 524653
rect 185663 524610 185671 524644
rect 185727 524610 185763 524644
rect 185797 524610 185855 524644
rect 185889 524610 185947 524644
rect 185981 524610 186039 524644
rect 186073 524610 186131 524644
rect 186165 524610 186223 524644
rect 186257 524610 186315 524644
rect 186349 524610 186407 524644
rect 186441 524610 186499 524644
rect 186533 524610 186591 524644
rect 186625 524610 186683 524644
rect 186717 524610 186775 524644
rect 186809 524610 186867 524644
rect 186901 524610 186959 524644
rect 186993 524610 187051 524644
rect 187085 524610 187143 524644
rect 187177 524610 187235 524644
rect 187269 524610 187327 524644
rect 187361 524610 187419 524644
rect 187453 524610 187482 524644
rect 185599 524601 185611 524610
rect 185663 524601 185675 524610
rect 185727 524601 187482 524610
rect 172210 524579 187482 524601
rect 172210 524109 187482 524131
rect 172210 524100 174625 524109
rect 172210 524066 172239 524100
rect 172273 524066 172331 524100
rect 172365 524066 172423 524100
rect 172457 524066 172515 524100
rect 172549 524066 172607 524100
rect 172641 524066 172699 524100
rect 172733 524066 172791 524100
rect 172825 524066 172883 524100
rect 172917 524066 172975 524100
rect 173009 524066 173067 524100
rect 173101 524066 173159 524100
rect 173193 524066 173251 524100
rect 173285 524066 173343 524100
rect 173377 524066 173435 524100
rect 173469 524066 173527 524100
rect 173561 524066 173619 524100
rect 173653 524066 173711 524100
rect 173745 524066 173803 524100
rect 173837 524066 173895 524100
rect 173929 524066 173987 524100
rect 174021 524066 174079 524100
rect 174113 524066 174171 524100
rect 174205 524066 174263 524100
rect 174297 524066 174355 524100
rect 174389 524066 174447 524100
rect 174481 524066 174539 524100
rect 174573 524066 174625 524100
rect 172210 524057 174625 524066
rect 174677 524057 174689 524109
rect 174741 524100 174753 524109
rect 174805 524100 174817 524109
rect 174805 524066 174815 524100
rect 174741 524057 174753 524066
rect 174805 524057 174817 524066
rect 174869 524057 174881 524109
rect 174933 524100 178443 524109
rect 174941 524066 174999 524100
rect 175033 524066 175091 524100
rect 175125 524066 175183 524100
rect 175217 524066 175275 524100
rect 175309 524066 175367 524100
rect 175401 524066 175459 524100
rect 175493 524066 175551 524100
rect 175585 524066 175643 524100
rect 175677 524066 175735 524100
rect 175769 524066 175827 524100
rect 175861 524066 175919 524100
rect 175953 524066 176011 524100
rect 176045 524066 176103 524100
rect 176137 524066 176195 524100
rect 176229 524066 176287 524100
rect 176321 524066 176379 524100
rect 176413 524066 176471 524100
rect 176505 524066 176563 524100
rect 176597 524066 176655 524100
rect 176689 524066 176747 524100
rect 176781 524066 176839 524100
rect 176873 524066 176931 524100
rect 176965 524066 177023 524100
rect 177057 524066 177115 524100
rect 177149 524066 177207 524100
rect 177241 524066 177299 524100
rect 177333 524066 177391 524100
rect 177425 524066 177483 524100
rect 177517 524066 177575 524100
rect 177609 524066 177667 524100
rect 177701 524066 177759 524100
rect 177793 524066 177851 524100
rect 177885 524066 177943 524100
rect 177977 524066 178035 524100
rect 178069 524066 178127 524100
rect 178161 524066 178219 524100
rect 178253 524066 178311 524100
rect 178345 524066 178403 524100
rect 178437 524066 178443 524100
rect 174933 524057 178443 524066
rect 178495 524100 178507 524109
rect 178495 524057 178507 524066
rect 178559 524057 178571 524109
rect 178623 524057 178635 524109
rect 178687 524100 178699 524109
rect 178751 524100 182261 524109
rect 178751 524066 178771 524100
rect 178805 524066 178863 524100
rect 178897 524066 178955 524100
rect 178989 524066 179047 524100
rect 179081 524066 179139 524100
rect 179173 524066 179231 524100
rect 179265 524066 179323 524100
rect 179357 524066 179415 524100
rect 179449 524066 179507 524100
rect 179541 524066 179599 524100
rect 179633 524066 179691 524100
rect 179725 524066 179783 524100
rect 179817 524066 179875 524100
rect 179909 524066 179967 524100
rect 180001 524066 180059 524100
rect 180093 524066 180151 524100
rect 180185 524066 180243 524100
rect 180277 524066 180335 524100
rect 180369 524066 180427 524100
rect 180461 524066 180519 524100
rect 180553 524066 180611 524100
rect 180645 524066 180703 524100
rect 180737 524066 180795 524100
rect 180829 524066 180887 524100
rect 180921 524066 180979 524100
rect 181013 524066 181071 524100
rect 181105 524066 181163 524100
rect 181197 524066 181255 524100
rect 181289 524066 181347 524100
rect 181381 524066 181439 524100
rect 181473 524066 181531 524100
rect 181565 524066 181623 524100
rect 181657 524066 181715 524100
rect 181749 524066 181807 524100
rect 181841 524066 181899 524100
rect 181933 524066 181991 524100
rect 182025 524066 182083 524100
rect 182117 524066 182175 524100
rect 182209 524066 182261 524100
rect 178687 524057 178699 524066
rect 178751 524057 182261 524066
rect 182313 524057 182325 524109
rect 182377 524100 182389 524109
rect 182441 524100 182453 524109
rect 182441 524066 182451 524100
rect 182377 524057 182389 524066
rect 182441 524057 182453 524066
rect 182505 524057 182517 524109
rect 182569 524100 186079 524109
rect 182577 524066 182635 524100
rect 182669 524066 182727 524100
rect 182761 524066 182819 524100
rect 182853 524066 182911 524100
rect 182945 524066 183003 524100
rect 183037 524066 183095 524100
rect 183129 524066 183187 524100
rect 183221 524066 183279 524100
rect 183313 524066 183371 524100
rect 183405 524066 183463 524100
rect 183497 524066 183555 524100
rect 183589 524066 183647 524100
rect 183681 524066 183739 524100
rect 183773 524066 183831 524100
rect 183865 524066 183923 524100
rect 183957 524066 184015 524100
rect 184049 524066 184107 524100
rect 184141 524066 184199 524100
rect 184233 524066 184291 524100
rect 184325 524066 184383 524100
rect 184417 524066 184475 524100
rect 184509 524066 184567 524100
rect 184601 524066 184659 524100
rect 184693 524066 184751 524100
rect 184785 524066 184843 524100
rect 184877 524066 184935 524100
rect 184969 524066 185027 524100
rect 185061 524066 185119 524100
rect 185153 524066 185211 524100
rect 185245 524066 185303 524100
rect 185337 524066 185395 524100
rect 185429 524066 185487 524100
rect 185521 524066 185579 524100
rect 185613 524066 185671 524100
rect 185705 524066 185763 524100
rect 185797 524066 185855 524100
rect 185889 524066 185947 524100
rect 185981 524066 186039 524100
rect 186073 524066 186079 524100
rect 182569 524057 186079 524066
rect 186131 524100 186143 524109
rect 186131 524057 186143 524066
rect 186195 524057 186207 524109
rect 186259 524057 186271 524109
rect 186323 524100 186335 524109
rect 186387 524100 187482 524109
rect 186387 524066 186407 524100
rect 186441 524066 186499 524100
rect 186533 524066 186591 524100
rect 186625 524066 186683 524100
rect 186717 524066 186775 524100
rect 186809 524066 186867 524100
rect 186901 524066 186959 524100
rect 186993 524066 187051 524100
rect 187085 524066 187143 524100
rect 187177 524066 187235 524100
rect 187269 524066 187327 524100
rect 187361 524066 187419 524100
rect 187453 524066 187482 524100
rect 186323 524057 186335 524066
rect 186387 524057 187482 524066
rect 172210 524035 187482 524057
rect 193000 524000 195000 526000
rect 192430 523587 192630 523617
rect 172210 523565 192630 523587
rect 193000 523570 193130 524000
rect 172210 523556 173965 523565
rect 174017 523556 174029 523565
rect 174081 523556 174093 523565
rect 172210 523522 172239 523556
rect 172273 523522 172331 523556
rect 172365 523522 172423 523556
rect 172457 523522 172515 523556
rect 172549 523522 172607 523556
rect 172641 523522 172699 523556
rect 172733 523522 172791 523556
rect 172825 523522 172883 523556
rect 172917 523522 172975 523556
rect 173009 523522 173067 523556
rect 173101 523522 173159 523556
rect 173193 523522 173251 523556
rect 173285 523522 173343 523556
rect 173377 523522 173435 523556
rect 173469 523522 173527 523556
rect 173561 523522 173619 523556
rect 173653 523522 173711 523556
rect 173745 523522 173803 523556
rect 173837 523522 173895 523556
rect 173929 523522 173965 523556
rect 174021 523522 174029 523556
rect 172210 523513 173965 523522
rect 174017 523513 174029 523522
rect 174081 523513 174093 523522
rect 174145 523513 174157 523565
rect 174209 523513 174221 523565
rect 174273 523556 177783 523565
rect 174297 523522 174355 523556
rect 174389 523522 174447 523556
rect 174481 523522 174539 523556
rect 174573 523522 174631 523556
rect 174665 523522 174723 523556
rect 174757 523522 174815 523556
rect 174849 523522 174907 523556
rect 174941 523522 174999 523556
rect 175033 523522 175091 523556
rect 175125 523522 175183 523556
rect 175217 523522 175275 523556
rect 175309 523522 175367 523556
rect 175401 523522 175459 523556
rect 175493 523522 175551 523556
rect 175585 523522 175643 523556
rect 175677 523522 175735 523556
rect 175769 523522 175827 523556
rect 175861 523522 175919 523556
rect 175953 523522 176011 523556
rect 176045 523522 176103 523556
rect 176137 523522 176195 523556
rect 176229 523522 176287 523556
rect 176321 523522 176379 523556
rect 176413 523522 176471 523556
rect 176505 523522 176563 523556
rect 176597 523522 176655 523556
rect 176689 523522 176747 523556
rect 176781 523522 176839 523556
rect 176873 523522 176931 523556
rect 176965 523522 177023 523556
rect 177057 523522 177115 523556
rect 177149 523522 177207 523556
rect 177241 523522 177299 523556
rect 177333 523522 177391 523556
rect 177425 523522 177483 523556
rect 177517 523522 177575 523556
rect 177609 523522 177667 523556
rect 177701 523522 177759 523556
rect 174273 523513 177783 523522
rect 177835 523513 177847 523565
rect 177899 523513 177911 523565
rect 177963 523556 177975 523565
rect 178027 523556 178039 523565
rect 178091 523556 181601 523565
rect 181653 523556 181665 523565
rect 181717 523556 181729 523565
rect 178027 523522 178035 523556
rect 178091 523522 178127 523556
rect 178161 523522 178219 523556
rect 178253 523522 178311 523556
rect 178345 523522 178403 523556
rect 178437 523522 178495 523556
rect 178529 523522 178587 523556
rect 178621 523522 178679 523556
rect 178713 523522 178771 523556
rect 178805 523522 178863 523556
rect 178897 523522 178955 523556
rect 178989 523522 179047 523556
rect 179081 523522 179139 523556
rect 179173 523522 179231 523556
rect 179265 523522 179323 523556
rect 179357 523522 179415 523556
rect 179449 523522 179507 523556
rect 179541 523522 179599 523556
rect 179633 523522 179691 523556
rect 179725 523522 179783 523556
rect 179817 523522 179875 523556
rect 179909 523522 179967 523556
rect 180001 523522 180059 523556
rect 180093 523522 180151 523556
rect 180185 523522 180243 523556
rect 180277 523522 180335 523556
rect 180369 523522 180427 523556
rect 180461 523522 180519 523556
rect 180553 523522 180611 523556
rect 180645 523522 180703 523556
rect 180737 523522 180795 523556
rect 180829 523522 180887 523556
rect 180921 523522 180979 523556
rect 181013 523522 181071 523556
rect 181105 523522 181163 523556
rect 181197 523522 181255 523556
rect 181289 523522 181347 523556
rect 181381 523522 181439 523556
rect 181473 523522 181531 523556
rect 181565 523522 181601 523556
rect 181657 523522 181665 523556
rect 177963 523513 177975 523522
rect 178027 523513 178039 523522
rect 178091 523513 181601 523522
rect 181653 523513 181665 523522
rect 181717 523513 181729 523522
rect 181781 523513 181793 523565
rect 181845 523513 181857 523565
rect 181909 523556 185419 523565
rect 181933 523522 181991 523556
rect 182025 523522 182083 523556
rect 182117 523522 182175 523556
rect 182209 523522 182267 523556
rect 182301 523522 182359 523556
rect 182393 523522 182451 523556
rect 182485 523522 182543 523556
rect 182577 523522 182635 523556
rect 182669 523522 182727 523556
rect 182761 523522 182819 523556
rect 182853 523522 182911 523556
rect 182945 523522 183003 523556
rect 183037 523522 183095 523556
rect 183129 523522 183187 523556
rect 183221 523522 183279 523556
rect 183313 523522 183371 523556
rect 183405 523522 183463 523556
rect 183497 523522 183555 523556
rect 183589 523522 183647 523556
rect 183681 523522 183739 523556
rect 183773 523522 183831 523556
rect 183865 523522 183923 523556
rect 183957 523522 184015 523556
rect 184049 523522 184107 523556
rect 184141 523522 184199 523556
rect 184233 523522 184291 523556
rect 184325 523522 184383 523556
rect 184417 523522 184475 523556
rect 184509 523522 184567 523556
rect 184601 523522 184659 523556
rect 184693 523522 184751 523556
rect 184785 523522 184843 523556
rect 184877 523522 184935 523556
rect 184969 523522 185027 523556
rect 185061 523522 185119 523556
rect 185153 523522 185211 523556
rect 185245 523522 185303 523556
rect 185337 523522 185395 523556
rect 181909 523513 185419 523522
rect 185471 523513 185483 523565
rect 185535 523513 185547 523565
rect 185599 523556 185611 523565
rect 185663 523556 185675 523565
rect 185727 523556 192630 523565
rect 185663 523522 185671 523556
rect 185727 523522 185763 523556
rect 185797 523522 185855 523556
rect 185889 523522 185947 523556
rect 185981 523522 186039 523556
rect 186073 523522 186131 523556
rect 186165 523522 186223 523556
rect 186257 523522 186315 523556
rect 186349 523522 186407 523556
rect 186441 523522 186499 523556
rect 186533 523522 186591 523556
rect 186625 523522 186683 523556
rect 186717 523522 186775 523556
rect 186809 523522 186867 523556
rect 186901 523522 186959 523556
rect 186993 523522 187051 523556
rect 187085 523522 187143 523556
rect 187177 523522 187235 523556
rect 187269 523522 187327 523556
rect 187361 523522 187419 523556
rect 187453 523522 192630 523556
rect 185599 523513 185611 523522
rect 185663 523513 185675 523522
rect 185727 523513 192630 523522
rect 172210 523491 192630 523513
rect 187470 523487 192630 523491
rect 192430 523427 192630 523487
rect 192742 523450 193130 523570
rect 172210 523037 187482 523043
rect 192430 523037 192630 523097
rect 172210 523021 192110 523037
rect 172210 523012 174625 523021
rect 172210 522978 172239 523012
rect 172273 522978 172331 523012
rect 172365 522978 172423 523012
rect 172457 522978 172515 523012
rect 172549 522978 172607 523012
rect 172641 522978 172699 523012
rect 172733 522978 172791 523012
rect 172825 522978 172883 523012
rect 172917 522978 172975 523012
rect 173009 522978 173067 523012
rect 173101 522978 173159 523012
rect 173193 522978 173251 523012
rect 173285 522978 173343 523012
rect 173377 522978 173435 523012
rect 173469 522978 173527 523012
rect 173561 522978 173619 523012
rect 173653 522978 173711 523012
rect 173745 522978 173803 523012
rect 173837 522978 173895 523012
rect 173929 522978 173987 523012
rect 174021 522978 174079 523012
rect 174113 522978 174171 523012
rect 174205 522978 174263 523012
rect 174297 522978 174355 523012
rect 174389 522978 174447 523012
rect 174481 522978 174539 523012
rect 174573 522978 174625 523012
rect 172210 522969 174625 522978
rect 174677 522969 174689 523021
rect 174741 523012 174753 523021
rect 174805 523012 174817 523021
rect 174805 522978 174815 523012
rect 174741 522969 174753 522978
rect 174805 522969 174817 522978
rect 174869 522969 174881 523021
rect 174933 523012 178443 523021
rect 174941 522978 174999 523012
rect 175033 522978 175091 523012
rect 175125 522978 175183 523012
rect 175217 522978 175275 523012
rect 175309 522978 175367 523012
rect 175401 522978 175459 523012
rect 175493 522978 175551 523012
rect 175585 522978 175643 523012
rect 175677 522978 175735 523012
rect 175769 522978 175827 523012
rect 175861 522978 175919 523012
rect 175953 522978 176011 523012
rect 176045 522978 176103 523012
rect 176137 522978 176195 523012
rect 176229 522978 176287 523012
rect 176321 522978 176379 523012
rect 176413 522978 176471 523012
rect 176505 522978 176563 523012
rect 176597 522978 176655 523012
rect 176689 522978 176747 523012
rect 176781 522978 176839 523012
rect 176873 522978 176931 523012
rect 176965 522978 177023 523012
rect 177057 522978 177115 523012
rect 177149 522978 177207 523012
rect 177241 522978 177299 523012
rect 177333 522978 177391 523012
rect 177425 522978 177483 523012
rect 177517 522978 177575 523012
rect 177609 522978 177667 523012
rect 177701 522978 177759 523012
rect 177793 522978 177851 523012
rect 177885 522978 177943 523012
rect 177977 522978 178035 523012
rect 178069 522978 178127 523012
rect 178161 522978 178219 523012
rect 178253 522978 178311 523012
rect 178345 522978 178403 523012
rect 178437 522978 178443 523012
rect 174933 522969 178443 522978
rect 178495 523012 178507 523021
rect 178495 522969 178507 522978
rect 178559 522969 178571 523021
rect 178623 522969 178635 523021
rect 178687 523012 178699 523021
rect 178751 523012 182261 523021
rect 178751 522978 178771 523012
rect 178805 522978 178863 523012
rect 178897 522978 178955 523012
rect 178989 522978 179047 523012
rect 179081 522978 179139 523012
rect 179173 522978 179231 523012
rect 179265 522978 179323 523012
rect 179357 522978 179415 523012
rect 179449 522978 179507 523012
rect 179541 522978 179599 523012
rect 179633 522978 179691 523012
rect 179725 522978 179783 523012
rect 179817 522978 179875 523012
rect 179909 522978 179967 523012
rect 180001 522978 180059 523012
rect 180093 522978 180151 523012
rect 180185 522978 180243 523012
rect 180277 522978 180335 523012
rect 180369 522978 180427 523012
rect 180461 522978 180519 523012
rect 180553 522978 180611 523012
rect 180645 522978 180703 523012
rect 180737 522978 180795 523012
rect 180829 522978 180887 523012
rect 180921 522978 180979 523012
rect 181013 522978 181071 523012
rect 181105 522978 181163 523012
rect 181197 522978 181255 523012
rect 181289 522978 181347 523012
rect 181381 522978 181439 523012
rect 181473 522978 181531 523012
rect 181565 522978 181623 523012
rect 181657 522978 181715 523012
rect 181749 522978 181807 523012
rect 181841 522978 181899 523012
rect 181933 522978 181991 523012
rect 182025 522978 182083 523012
rect 182117 522978 182175 523012
rect 182209 522978 182261 523012
rect 178687 522969 178699 522978
rect 178751 522969 182261 522978
rect 182313 522969 182325 523021
rect 182377 523012 182389 523021
rect 182441 523012 182453 523021
rect 182441 522978 182451 523012
rect 182377 522969 182389 522978
rect 182441 522969 182453 522978
rect 182505 522969 182517 523021
rect 182569 523012 186079 523021
rect 182577 522978 182635 523012
rect 182669 522978 182727 523012
rect 182761 522978 182819 523012
rect 182853 522978 182911 523012
rect 182945 522978 183003 523012
rect 183037 522978 183095 523012
rect 183129 522978 183187 523012
rect 183221 522978 183279 523012
rect 183313 522978 183371 523012
rect 183405 522978 183463 523012
rect 183497 522978 183555 523012
rect 183589 522978 183647 523012
rect 183681 522978 183739 523012
rect 183773 522978 183831 523012
rect 183865 522978 183923 523012
rect 183957 522978 184015 523012
rect 184049 522978 184107 523012
rect 184141 522978 184199 523012
rect 184233 522978 184291 523012
rect 184325 522978 184383 523012
rect 184417 522978 184475 523012
rect 184509 522978 184567 523012
rect 184601 522978 184659 523012
rect 184693 522978 184751 523012
rect 184785 522978 184843 523012
rect 184877 522978 184935 523012
rect 184969 522978 185027 523012
rect 185061 522978 185119 523012
rect 185153 522978 185211 523012
rect 185245 522978 185303 523012
rect 185337 522978 185395 523012
rect 185429 522978 185487 523012
rect 185521 522978 185579 523012
rect 185613 522978 185671 523012
rect 185705 522978 185763 523012
rect 185797 522978 185855 523012
rect 185889 522978 185947 523012
rect 185981 522978 186039 523012
rect 186073 522978 186079 523012
rect 182569 522969 186079 522978
rect 186131 523012 186143 523021
rect 186131 522969 186143 522978
rect 186195 522969 186207 523021
rect 186259 522969 186271 523021
rect 186323 523012 186335 523021
rect 186387 523012 192110 523021
rect 186387 522978 186407 523012
rect 186441 522978 186499 523012
rect 186533 522978 186591 523012
rect 186625 522978 186683 523012
rect 186717 522978 186775 523012
rect 186809 522978 186867 523012
rect 186901 522978 186959 523012
rect 186993 522978 187051 523012
rect 187085 522978 187143 523012
rect 187177 522978 187235 523012
rect 187269 522978 187327 523012
rect 187361 522978 187419 523012
rect 187453 522978 192110 523012
rect 186323 522969 186335 522978
rect 186387 522969 192110 522978
rect 172210 522947 192110 522969
rect 192140 522947 192630 523037
rect 192430 522907 192630 522947
rect 192742 523000 193020 523010
rect 192742 522910 195000 523000
rect 172210 522477 187482 522499
rect 172210 522468 173965 522477
rect 174017 522468 174029 522477
rect 174081 522468 174093 522477
rect 172210 522434 172239 522468
rect 172273 522434 172331 522468
rect 172365 522434 172423 522468
rect 172457 522434 172515 522468
rect 172549 522434 172607 522468
rect 172641 522434 172699 522468
rect 172733 522434 172791 522468
rect 172825 522434 172883 522468
rect 172917 522434 172975 522468
rect 173009 522434 173067 522468
rect 173101 522434 173159 522468
rect 173193 522434 173251 522468
rect 173285 522434 173343 522468
rect 173377 522434 173435 522468
rect 173469 522434 173527 522468
rect 173561 522434 173619 522468
rect 173653 522434 173711 522468
rect 173745 522434 173803 522468
rect 173837 522434 173895 522468
rect 173929 522434 173965 522468
rect 174021 522434 174029 522468
rect 172210 522425 173965 522434
rect 174017 522425 174029 522434
rect 174081 522425 174093 522434
rect 174145 522425 174157 522477
rect 174209 522425 174221 522477
rect 174273 522468 177783 522477
rect 174297 522434 174355 522468
rect 174389 522434 174447 522468
rect 174481 522434 174539 522468
rect 174573 522434 174631 522468
rect 174665 522434 174723 522468
rect 174757 522434 174815 522468
rect 174849 522434 174907 522468
rect 174941 522434 174999 522468
rect 175033 522434 175091 522468
rect 175125 522434 175183 522468
rect 175217 522434 175275 522468
rect 175309 522434 175367 522468
rect 175401 522434 175459 522468
rect 175493 522434 175551 522468
rect 175585 522434 175643 522468
rect 175677 522434 175735 522468
rect 175769 522434 175827 522468
rect 175861 522434 175919 522468
rect 175953 522434 176011 522468
rect 176045 522434 176103 522468
rect 176137 522434 176195 522468
rect 176229 522434 176287 522468
rect 176321 522434 176379 522468
rect 176413 522434 176471 522468
rect 176505 522434 176563 522468
rect 176597 522434 176655 522468
rect 176689 522434 176747 522468
rect 176781 522434 176839 522468
rect 176873 522434 176931 522468
rect 176965 522434 177023 522468
rect 177057 522434 177115 522468
rect 177149 522434 177207 522468
rect 177241 522434 177299 522468
rect 177333 522434 177391 522468
rect 177425 522434 177483 522468
rect 177517 522434 177575 522468
rect 177609 522434 177667 522468
rect 177701 522434 177759 522468
rect 174273 522425 177783 522434
rect 177835 522425 177847 522477
rect 177899 522425 177911 522477
rect 177963 522468 177975 522477
rect 178027 522468 178039 522477
rect 178091 522468 181601 522477
rect 181653 522468 181665 522477
rect 181717 522468 181729 522477
rect 178027 522434 178035 522468
rect 178091 522434 178127 522468
rect 178161 522434 178219 522468
rect 178253 522434 178311 522468
rect 178345 522434 178403 522468
rect 178437 522434 178495 522468
rect 178529 522434 178587 522468
rect 178621 522434 178679 522468
rect 178713 522434 178771 522468
rect 178805 522434 178863 522468
rect 178897 522434 178955 522468
rect 178989 522434 179047 522468
rect 179081 522434 179139 522468
rect 179173 522434 179231 522468
rect 179265 522434 179323 522468
rect 179357 522434 179415 522468
rect 179449 522434 179507 522468
rect 179541 522434 179599 522468
rect 179633 522434 179691 522468
rect 179725 522434 179783 522468
rect 179817 522434 179875 522468
rect 179909 522434 179967 522468
rect 180001 522434 180059 522468
rect 180093 522434 180151 522468
rect 180185 522434 180243 522468
rect 180277 522434 180335 522468
rect 180369 522434 180427 522468
rect 180461 522434 180519 522468
rect 180553 522434 180611 522468
rect 180645 522434 180703 522468
rect 180737 522434 180795 522468
rect 180829 522434 180887 522468
rect 180921 522434 180979 522468
rect 181013 522434 181071 522468
rect 181105 522434 181163 522468
rect 181197 522434 181255 522468
rect 181289 522434 181347 522468
rect 181381 522434 181439 522468
rect 181473 522434 181531 522468
rect 181565 522434 181601 522468
rect 181657 522434 181665 522468
rect 177963 522425 177975 522434
rect 178027 522425 178039 522434
rect 178091 522425 181601 522434
rect 181653 522425 181665 522434
rect 181717 522425 181729 522434
rect 181781 522425 181793 522477
rect 181845 522425 181857 522477
rect 181909 522468 185419 522477
rect 181933 522434 181991 522468
rect 182025 522434 182083 522468
rect 182117 522434 182175 522468
rect 182209 522434 182267 522468
rect 182301 522434 182359 522468
rect 182393 522434 182451 522468
rect 182485 522434 182543 522468
rect 182577 522434 182635 522468
rect 182669 522434 182727 522468
rect 182761 522434 182819 522468
rect 182853 522434 182911 522468
rect 182945 522434 183003 522468
rect 183037 522434 183095 522468
rect 183129 522434 183187 522468
rect 183221 522434 183279 522468
rect 183313 522434 183371 522468
rect 183405 522434 183463 522468
rect 183497 522434 183555 522468
rect 183589 522434 183647 522468
rect 183681 522434 183739 522468
rect 183773 522434 183831 522468
rect 183865 522434 183923 522468
rect 183957 522434 184015 522468
rect 184049 522434 184107 522468
rect 184141 522434 184199 522468
rect 184233 522434 184291 522468
rect 184325 522434 184383 522468
rect 184417 522434 184475 522468
rect 184509 522434 184567 522468
rect 184601 522434 184659 522468
rect 184693 522434 184751 522468
rect 184785 522434 184843 522468
rect 184877 522434 184935 522468
rect 184969 522434 185027 522468
rect 185061 522434 185119 522468
rect 185153 522434 185211 522468
rect 185245 522434 185303 522468
rect 185337 522434 185395 522468
rect 181909 522425 185419 522434
rect 185471 522425 185483 522477
rect 185535 522425 185547 522477
rect 185599 522468 185611 522477
rect 185663 522468 185675 522477
rect 185727 522468 187482 522477
rect 185663 522434 185671 522468
rect 185727 522434 185763 522468
rect 185797 522434 185855 522468
rect 185889 522434 185947 522468
rect 185981 522434 186039 522468
rect 186073 522434 186131 522468
rect 186165 522434 186223 522468
rect 186257 522434 186315 522468
rect 186349 522434 186407 522468
rect 186441 522434 186499 522468
rect 186533 522434 186591 522468
rect 186625 522434 186683 522468
rect 186717 522434 186775 522468
rect 186809 522434 186867 522468
rect 186901 522434 186959 522468
rect 186993 522434 187051 522468
rect 187085 522434 187143 522468
rect 187177 522434 187235 522468
rect 187269 522434 187327 522468
rect 187361 522434 187419 522468
rect 187453 522434 187482 522468
rect 185599 522425 185611 522434
rect 185663 522425 185675 522434
rect 185727 522425 187482 522434
rect 172210 522403 187482 522425
rect 172210 521933 187482 521955
rect 172210 521924 174625 521933
rect 172210 521890 172239 521924
rect 172273 521890 172331 521924
rect 172365 521890 172423 521924
rect 172457 521890 172515 521924
rect 172549 521890 172607 521924
rect 172641 521890 172699 521924
rect 172733 521890 172791 521924
rect 172825 521890 172883 521924
rect 172917 521890 172975 521924
rect 173009 521890 173067 521924
rect 173101 521890 173159 521924
rect 173193 521890 173251 521924
rect 173285 521890 173343 521924
rect 173377 521890 173435 521924
rect 173469 521890 173527 521924
rect 173561 521890 173619 521924
rect 173653 521890 173711 521924
rect 173745 521890 173803 521924
rect 173837 521890 173895 521924
rect 173929 521890 173987 521924
rect 174021 521890 174079 521924
rect 174113 521890 174171 521924
rect 174205 521890 174263 521924
rect 174297 521890 174355 521924
rect 174389 521890 174447 521924
rect 174481 521890 174539 521924
rect 174573 521890 174625 521924
rect 172210 521881 174625 521890
rect 174677 521881 174689 521933
rect 174741 521924 174753 521933
rect 174805 521924 174817 521933
rect 174805 521890 174815 521924
rect 174741 521881 174753 521890
rect 174805 521881 174817 521890
rect 174869 521881 174881 521933
rect 174933 521924 178443 521933
rect 174941 521890 174999 521924
rect 175033 521890 175091 521924
rect 175125 521890 175183 521924
rect 175217 521890 175275 521924
rect 175309 521890 175367 521924
rect 175401 521890 175459 521924
rect 175493 521890 175551 521924
rect 175585 521890 175643 521924
rect 175677 521890 175735 521924
rect 175769 521890 175827 521924
rect 175861 521890 175919 521924
rect 175953 521890 176011 521924
rect 176045 521890 176103 521924
rect 176137 521890 176195 521924
rect 176229 521890 176287 521924
rect 176321 521890 176379 521924
rect 176413 521890 176471 521924
rect 176505 521890 176563 521924
rect 176597 521890 176655 521924
rect 176689 521890 176747 521924
rect 176781 521890 176839 521924
rect 176873 521890 176931 521924
rect 176965 521890 177023 521924
rect 177057 521890 177115 521924
rect 177149 521890 177207 521924
rect 177241 521890 177299 521924
rect 177333 521890 177391 521924
rect 177425 521890 177483 521924
rect 177517 521890 177575 521924
rect 177609 521890 177667 521924
rect 177701 521890 177759 521924
rect 177793 521890 177851 521924
rect 177885 521890 177943 521924
rect 177977 521890 178035 521924
rect 178069 521890 178127 521924
rect 178161 521890 178219 521924
rect 178253 521890 178311 521924
rect 178345 521890 178403 521924
rect 178437 521890 178443 521924
rect 174933 521881 178443 521890
rect 178495 521924 178507 521933
rect 178495 521881 178507 521890
rect 178559 521881 178571 521933
rect 178623 521881 178635 521933
rect 178687 521924 178699 521933
rect 178751 521924 182261 521933
rect 178751 521890 178771 521924
rect 178805 521890 178863 521924
rect 178897 521890 178955 521924
rect 178989 521890 179047 521924
rect 179081 521890 179139 521924
rect 179173 521890 179231 521924
rect 179265 521890 179323 521924
rect 179357 521890 179415 521924
rect 179449 521890 179507 521924
rect 179541 521890 179599 521924
rect 179633 521890 179691 521924
rect 179725 521890 179783 521924
rect 179817 521890 179875 521924
rect 179909 521890 179967 521924
rect 180001 521890 180059 521924
rect 180093 521890 180151 521924
rect 180185 521890 180243 521924
rect 180277 521890 180335 521924
rect 180369 521890 180427 521924
rect 180461 521890 180519 521924
rect 180553 521890 180611 521924
rect 180645 521890 180703 521924
rect 180737 521890 180795 521924
rect 180829 521890 180887 521924
rect 180921 521890 180979 521924
rect 181013 521890 181071 521924
rect 181105 521890 181163 521924
rect 181197 521890 181255 521924
rect 181289 521890 181347 521924
rect 181381 521890 181439 521924
rect 181473 521890 181531 521924
rect 181565 521890 181623 521924
rect 181657 521890 181715 521924
rect 181749 521890 181807 521924
rect 181841 521890 181899 521924
rect 181933 521890 181991 521924
rect 182025 521890 182083 521924
rect 182117 521890 182175 521924
rect 182209 521890 182261 521924
rect 178687 521881 178699 521890
rect 178751 521881 182261 521890
rect 182313 521881 182325 521933
rect 182377 521924 182389 521933
rect 182441 521924 182453 521933
rect 182441 521890 182451 521924
rect 182377 521881 182389 521890
rect 182441 521881 182453 521890
rect 182505 521881 182517 521933
rect 182569 521924 186079 521933
rect 182577 521890 182635 521924
rect 182669 521890 182727 521924
rect 182761 521890 182819 521924
rect 182853 521890 182911 521924
rect 182945 521890 183003 521924
rect 183037 521890 183095 521924
rect 183129 521890 183187 521924
rect 183221 521890 183279 521924
rect 183313 521890 183371 521924
rect 183405 521890 183463 521924
rect 183497 521890 183555 521924
rect 183589 521890 183647 521924
rect 183681 521890 183739 521924
rect 183773 521890 183831 521924
rect 183865 521890 183923 521924
rect 183957 521890 184015 521924
rect 184049 521890 184107 521924
rect 184141 521890 184199 521924
rect 184233 521890 184291 521924
rect 184325 521890 184383 521924
rect 184417 521890 184475 521924
rect 184509 521890 184567 521924
rect 184601 521890 184659 521924
rect 184693 521890 184751 521924
rect 184785 521890 184843 521924
rect 184877 521890 184935 521924
rect 184969 521890 185027 521924
rect 185061 521890 185119 521924
rect 185153 521890 185211 521924
rect 185245 521890 185303 521924
rect 185337 521890 185395 521924
rect 185429 521890 185487 521924
rect 185521 521890 185579 521924
rect 185613 521890 185671 521924
rect 185705 521890 185763 521924
rect 185797 521890 185855 521924
rect 185889 521890 185947 521924
rect 185981 521890 186039 521924
rect 186073 521890 186079 521924
rect 182569 521881 186079 521890
rect 186131 521924 186143 521933
rect 186131 521881 186143 521890
rect 186195 521881 186207 521933
rect 186259 521881 186271 521933
rect 186323 521924 186335 521933
rect 186387 521924 187482 521933
rect 186387 521890 186407 521924
rect 186441 521890 186499 521924
rect 186533 521890 186591 521924
rect 186625 521890 186683 521924
rect 186717 521890 186775 521924
rect 186809 521890 186867 521924
rect 186901 521890 186959 521924
rect 186993 521890 187051 521924
rect 187085 521890 187143 521924
rect 187177 521890 187235 521924
rect 187269 521890 187327 521924
rect 187361 521890 187419 521924
rect 187453 521890 187482 521924
rect 186323 521881 186335 521890
rect 186387 521881 187482 521890
rect 172210 521859 187482 521881
rect 172210 521389 187482 521411
rect 172210 521380 173965 521389
rect 174017 521380 174029 521389
rect 174081 521380 174093 521389
rect 172210 521346 172239 521380
rect 172273 521346 172331 521380
rect 172365 521346 172423 521380
rect 172457 521346 172515 521380
rect 172549 521346 172607 521380
rect 172641 521346 172699 521380
rect 172733 521346 172791 521380
rect 172825 521346 172883 521380
rect 172917 521346 172975 521380
rect 173009 521346 173067 521380
rect 173101 521346 173159 521380
rect 173193 521346 173251 521380
rect 173285 521346 173343 521380
rect 173377 521346 173435 521380
rect 173469 521346 173527 521380
rect 173561 521346 173619 521380
rect 173653 521346 173711 521380
rect 173745 521346 173803 521380
rect 173837 521346 173895 521380
rect 173929 521346 173965 521380
rect 174021 521346 174029 521380
rect 172210 521337 173965 521346
rect 174017 521337 174029 521346
rect 174081 521337 174093 521346
rect 174145 521337 174157 521389
rect 174209 521337 174221 521389
rect 174273 521380 177783 521389
rect 174297 521346 174355 521380
rect 174389 521346 174447 521380
rect 174481 521346 174539 521380
rect 174573 521346 174631 521380
rect 174665 521346 174723 521380
rect 174757 521346 174815 521380
rect 174849 521346 174907 521380
rect 174941 521346 174999 521380
rect 175033 521346 175091 521380
rect 175125 521346 175183 521380
rect 175217 521346 175275 521380
rect 175309 521346 175367 521380
rect 175401 521346 175459 521380
rect 175493 521346 175551 521380
rect 175585 521346 175643 521380
rect 175677 521346 175735 521380
rect 175769 521346 175827 521380
rect 175861 521346 175919 521380
rect 175953 521346 176011 521380
rect 176045 521346 176103 521380
rect 176137 521346 176195 521380
rect 176229 521346 176287 521380
rect 176321 521346 176379 521380
rect 176413 521346 176471 521380
rect 176505 521346 176563 521380
rect 176597 521346 176655 521380
rect 176689 521346 176747 521380
rect 176781 521346 176839 521380
rect 176873 521346 176931 521380
rect 176965 521346 177023 521380
rect 177057 521346 177115 521380
rect 177149 521346 177207 521380
rect 177241 521346 177299 521380
rect 177333 521346 177391 521380
rect 177425 521346 177483 521380
rect 177517 521346 177575 521380
rect 177609 521346 177667 521380
rect 177701 521346 177759 521380
rect 174273 521337 177783 521346
rect 177835 521337 177847 521389
rect 177899 521337 177911 521389
rect 177963 521380 177975 521389
rect 178027 521380 178039 521389
rect 178091 521380 181601 521389
rect 181653 521380 181665 521389
rect 181717 521380 181729 521389
rect 178027 521346 178035 521380
rect 178091 521346 178127 521380
rect 178161 521346 178219 521380
rect 178253 521346 178311 521380
rect 178345 521346 178403 521380
rect 178437 521346 178495 521380
rect 178529 521346 178587 521380
rect 178621 521346 178679 521380
rect 178713 521346 178771 521380
rect 178805 521346 178863 521380
rect 178897 521346 178955 521380
rect 178989 521346 179047 521380
rect 179081 521346 179139 521380
rect 179173 521346 179231 521380
rect 179265 521346 179323 521380
rect 179357 521346 179415 521380
rect 179449 521346 179507 521380
rect 179541 521346 179599 521380
rect 179633 521346 179691 521380
rect 179725 521346 179783 521380
rect 179817 521346 179875 521380
rect 179909 521346 179967 521380
rect 180001 521346 180059 521380
rect 180093 521346 180151 521380
rect 180185 521346 180243 521380
rect 180277 521346 180335 521380
rect 180369 521346 180427 521380
rect 180461 521346 180519 521380
rect 180553 521346 180611 521380
rect 180645 521346 180703 521380
rect 180737 521346 180795 521380
rect 180829 521346 180887 521380
rect 180921 521346 180979 521380
rect 181013 521346 181071 521380
rect 181105 521346 181163 521380
rect 181197 521346 181255 521380
rect 181289 521346 181347 521380
rect 181381 521346 181439 521380
rect 181473 521346 181531 521380
rect 181565 521346 181601 521380
rect 181657 521346 181665 521380
rect 177963 521337 177975 521346
rect 178027 521337 178039 521346
rect 178091 521337 181601 521346
rect 181653 521337 181665 521346
rect 181717 521337 181729 521346
rect 181781 521337 181793 521389
rect 181845 521337 181857 521389
rect 181909 521380 185419 521389
rect 181933 521346 181991 521380
rect 182025 521346 182083 521380
rect 182117 521346 182175 521380
rect 182209 521346 182267 521380
rect 182301 521346 182359 521380
rect 182393 521346 182451 521380
rect 182485 521346 182543 521380
rect 182577 521346 182635 521380
rect 182669 521346 182727 521380
rect 182761 521346 182819 521380
rect 182853 521346 182911 521380
rect 182945 521346 183003 521380
rect 183037 521346 183095 521380
rect 183129 521346 183187 521380
rect 183221 521346 183279 521380
rect 183313 521346 183371 521380
rect 183405 521346 183463 521380
rect 183497 521346 183555 521380
rect 183589 521346 183647 521380
rect 183681 521346 183739 521380
rect 183773 521346 183831 521380
rect 183865 521346 183923 521380
rect 183957 521346 184015 521380
rect 184049 521346 184107 521380
rect 184141 521346 184199 521380
rect 184233 521346 184291 521380
rect 184325 521346 184383 521380
rect 184417 521346 184475 521380
rect 184509 521346 184567 521380
rect 184601 521346 184659 521380
rect 184693 521346 184751 521380
rect 184785 521346 184843 521380
rect 184877 521346 184935 521380
rect 184969 521346 185027 521380
rect 185061 521346 185119 521380
rect 185153 521346 185211 521380
rect 185245 521346 185303 521380
rect 185337 521346 185395 521380
rect 181909 521337 185419 521346
rect 185471 521337 185483 521389
rect 185535 521337 185547 521389
rect 185599 521380 185611 521389
rect 185663 521380 185675 521389
rect 185727 521380 187482 521389
rect 185663 521346 185671 521380
rect 185727 521346 185763 521380
rect 185797 521346 185855 521380
rect 185889 521346 185947 521380
rect 185981 521346 186039 521380
rect 186073 521346 186131 521380
rect 186165 521346 186223 521380
rect 186257 521346 186315 521380
rect 186349 521346 186407 521380
rect 186441 521346 186499 521380
rect 186533 521346 186591 521380
rect 186625 521346 186683 521380
rect 186717 521346 186775 521380
rect 186809 521346 186867 521380
rect 186901 521346 186959 521380
rect 186993 521346 187051 521380
rect 187085 521346 187143 521380
rect 187177 521346 187235 521380
rect 187269 521346 187327 521380
rect 187361 521346 187419 521380
rect 187453 521346 187482 521380
rect 185599 521337 185611 521346
rect 185663 521337 185675 521346
rect 185727 521337 187482 521346
rect 172210 521315 187482 521337
rect 193000 521000 195000 522910
rect 172210 520845 187482 520867
rect 172210 520836 174625 520845
rect 172210 520802 172239 520836
rect 172273 520802 172331 520836
rect 172365 520802 172423 520836
rect 172457 520802 172515 520836
rect 172549 520802 172607 520836
rect 172641 520802 172699 520836
rect 172733 520802 172791 520836
rect 172825 520802 172883 520836
rect 172917 520802 172975 520836
rect 173009 520802 173067 520836
rect 173101 520802 173159 520836
rect 173193 520802 173251 520836
rect 173285 520802 173343 520836
rect 173377 520802 173435 520836
rect 173469 520802 173527 520836
rect 173561 520802 173619 520836
rect 173653 520802 173711 520836
rect 173745 520802 173803 520836
rect 173837 520802 173895 520836
rect 173929 520802 173987 520836
rect 174021 520802 174079 520836
rect 174113 520802 174171 520836
rect 174205 520802 174263 520836
rect 174297 520802 174355 520836
rect 174389 520802 174447 520836
rect 174481 520802 174539 520836
rect 174573 520802 174625 520836
rect 172210 520793 174625 520802
rect 174677 520793 174689 520845
rect 174741 520836 174753 520845
rect 174805 520836 174817 520845
rect 174805 520802 174815 520836
rect 174741 520793 174753 520802
rect 174805 520793 174817 520802
rect 174869 520793 174881 520845
rect 174933 520836 178443 520845
rect 174941 520802 174999 520836
rect 175033 520802 175091 520836
rect 175125 520802 175183 520836
rect 175217 520802 175275 520836
rect 175309 520802 175367 520836
rect 175401 520802 175459 520836
rect 175493 520802 175551 520836
rect 175585 520802 175643 520836
rect 175677 520802 175735 520836
rect 175769 520802 175827 520836
rect 175861 520802 175919 520836
rect 175953 520802 176011 520836
rect 176045 520802 176103 520836
rect 176137 520802 176195 520836
rect 176229 520802 176287 520836
rect 176321 520802 176379 520836
rect 176413 520802 176471 520836
rect 176505 520802 176563 520836
rect 176597 520802 176655 520836
rect 176689 520802 176747 520836
rect 176781 520802 176839 520836
rect 176873 520802 176931 520836
rect 176965 520802 177023 520836
rect 177057 520802 177115 520836
rect 177149 520802 177207 520836
rect 177241 520802 177299 520836
rect 177333 520802 177391 520836
rect 177425 520802 177483 520836
rect 177517 520802 177575 520836
rect 177609 520802 177667 520836
rect 177701 520802 177759 520836
rect 177793 520802 177851 520836
rect 177885 520802 177943 520836
rect 177977 520802 178035 520836
rect 178069 520802 178127 520836
rect 178161 520802 178219 520836
rect 178253 520802 178311 520836
rect 178345 520802 178403 520836
rect 178437 520802 178443 520836
rect 174933 520793 178443 520802
rect 178495 520836 178507 520845
rect 178495 520793 178507 520802
rect 178559 520793 178571 520845
rect 178623 520793 178635 520845
rect 178687 520836 178699 520845
rect 178751 520836 182261 520845
rect 178751 520802 178771 520836
rect 178805 520802 178863 520836
rect 178897 520802 178955 520836
rect 178989 520802 179047 520836
rect 179081 520802 179139 520836
rect 179173 520802 179231 520836
rect 179265 520802 179323 520836
rect 179357 520802 179415 520836
rect 179449 520802 179507 520836
rect 179541 520802 179599 520836
rect 179633 520802 179691 520836
rect 179725 520802 179783 520836
rect 179817 520802 179875 520836
rect 179909 520802 179967 520836
rect 180001 520802 180059 520836
rect 180093 520802 180151 520836
rect 180185 520802 180243 520836
rect 180277 520802 180335 520836
rect 180369 520802 180427 520836
rect 180461 520802 180519 520836
rect 180553 520802 180611 520836
rect 180645 520802 180703 520836
rect 180737 520802 180795 520836
rect 180829 520802 180887 520836
rect 180921 520802 180979 520836
rect 181013 520802 181071 520836
rect 181105 520802 181163 520836
rect 181197 520802 181255 520836
rect 181289 520802 181347 520836
rect 181381 520802 181439 520836
rect 181473 520802 181531 520836
rect 181565 520802 181623 520836
rect 181657 520802 181715 520836
rect 181749 520802 181807 520836
rect 181841 520802 181899 520836
rect 181933 520802 181991 520836
rect 182025 520802 182083 520836
rect 182117 520802 182175 520836
rect 182209 520802 182261 520836
rect 178687 520793 178699 520802
rect 178751 520793 182261 520802
rect 182313 520793 182325 520845
rect 182377 520836 182389 520845
rect 182441 520836 182453 520845
rect 182441 520802 182451 520836
rect 182377 520793 182389 520802
rect 182441 520793 182453 520802
rect 182505 520793 182517 520845
rect 182569 520836 186079 520845
rect 182577 520802 182635 520836
rect 182669 520802 182727 520836
rect 182761 520802 182819 520836
rect 182853 520802 182911 520836
rect 182945 520802 183003 520836
rect 183037 520802 183095 520836
rect 183129 520802 183187 520836
rect 183221 520802 183279 520836
rect 183313 520802 183371 520836
rect 183405 520802 183463 520836
rect 183497 520802 183555 520836
rect 183589 520802 183647 520836
rect 183681 520802 183739 520836
rect 183773 520802 183831 520836
rect 183865 520802 183923 520836
rect 183957 520802 184015 520836
rect 184049 520802 184107 520836
rect 184141 520802 184199 520836
rect 184233 520802 184291 520836
rect 184325 520802 184383 520836
rect 184417 520802 184475 520836
rect 184509 520802 184567 520836
rect 184601 520802 184659 520836
rect 184693 520802 184751 520836
rect 184785 520802 184843 520836
rect 184877 520802 184935 520836
rect 184969 520802 185027 520836
rect 185061 520802 185119 520836
rect 185153 520802 185211 520836
rect 185245 520802 185303 520836
rect 185337 520802 185395 520836
rect 185429 520802 185487 520836
rect 185521 520802 185579 520836
rect 185613 520802 185671 520836
rect 185705 520802 185763 520836
rect 185797 520802 185855 520836
rect 185889 520802 185947 520836
rect 185981 520802 186039 520836
rect 186073 520802 186079 520836
rect 182569 520793 186079 520802
rect 186131 520836 186143 520845
rect 186131 520793 186143 520802
rect 186195 520793 186207 520845
rect 186259 520793 186271 520845
rect 186323 520836 186335 520845
rect 186387 520836 187482 520845
rect 186387 520802 186407 520836
rect 186441 520802 186499 520836
rect 186533 520802 186591 520836
rect 186625 520802 186683 520836
rect 186717 520802 186775 520836
rect 186809 520802 186867 520836
rect 186901 520802 186959 520836
rect 186993 520802 187051 520836
rect 187085 520802 187143 520836
rect 187177 520802 187235 520836
rect 187269 520802 187327 520836
rect 187361 520802 187419 520836
rect 187453 520802 187482 520836
rect 186323 520793 186335 520802
rect 186387 520793 187482 520802
rect 172210 520771 187482 520793
rect 172210 520301 187482 520323
rect 172210 520292 173965 520301
rect 174017 520292 174029 520301
rect 174081 520292 174093 520301
rect 172210 520258 172239 520292
rect 172273 520258 172331 520292
rect 172365 520258 172423 520292
rect 172457 520258 172515 520292
rect 172549 520258 172607 520292
rect 172641 520258 172699 520292
rect 172733 520258 172791 520292
rect 172825 520258 172883 520292
rect 172917 520258 172975 520292
rect 173009 520258 173067 520292
rect 173101 520258 173159 520292
rect 173193 520258 173251 520292
rect 173285 520258 173343 520292
rect 173377 520258 173435 520292
rect 173469 520258 173527 520292
rect 173561 520258 173619 520292
rect 173653 520258 173711 520292
rect 173745 520258 173803 520292
rect 173837 520258 173895 520292
rect 173929 520258 173965 520292
rect 174021 520258 174029 520292
rect 172210 520249 173965 520258
rect 174017 520249 174029 520258
rect 174081 520249 174093 520258
rect 174145 520249 174157 520301
rect 174209 520249 174221 520301
rect 174273 520292 177783 520301
rect 174297 520258 174355 520292
rect 174389 520258 174447 520292
rect 174481 520258 174539 520292
rect 174573 520258 174631 520292
rect 174665 520258 174723 520292
rect 174757 520258 174815 520292
rect 174849 520258 174907 520292
rect 174941 520258 174999 520292
rect 175033 520258 175091 520292
rect 175125 520258 175183 520292
rect 175217 520258 175275 520292
rect 175309 520258 175367 520292
rect 175401 520258 175459 520292
rect 175493 520258 175551 520292
rect 175585 520258 175643 520292
rect 175677 520258 175735 520292
rect 175769 520258 175827 520292
rect 175861 520258 175919 520292
rect 175953 520258 176011 520292
rect 176045 520258 176103 520292
rect 176137 520258 176195 520292
rect 176229 520258 176287 520292
rect 176321 520258 176379 520292
rect 176413 520258 176471 520292
rect 176505 520258 176563 520292
rect 176597 520258 176655 520292
rect 176689 520258 176747 520292
rect 176781 520258 176839 520292
rect 176873 520258 176931 520292
rect 176965 520258 177023 520292
rect 177057 520258 177115 520292
rect 177149 520258 177207 520292
rect 177241 520258 177299 520292
rect 177333 520258 177391 520292
rect 177425 520258 177483 520292
rect 177517 520258 177575 520292
rect 177609 520258 177667 520292
rect 177701 520258 177759 520292
rect 174273 520249 177783 520258
rect 177835 520249 177847 520301
rect 177899 520249 177911 520301
rect 177963 520292 177975 520301
rect 178027 520292 178039 520301
rect 178091 520292 181601 520301
rect 181653 520292 181665 520301
rect 181717 520292 181729 520301
rect 178027 520258 178035 520292
rect 178091 520258 178127 520292
rect 178161 520258 178219 520292
rect 178253 520258 178311 520292
rect 178345 520258 178403 520292
rect 178437 520258 178495 520292
rect 178529 520258 178587 520292
rect 178621 520258 178679 520292
rect 178713 520258 178771 520292
rect 178805 520258 178863 520292
rect 178897 520258 178955 520292
rect 178989 520258 179047 520292
rect 179081 520258 179139 520292
rect 179173 520258 179231 520292
rect 179265 520258 179323 520292
rect 179357 520258 179415 520292
rect 179449 520258 179507 520292
rect 179541 520258 179599 520292
rect 179633 520258 179691 520292
rect 179725 520258 179783 520292
rect 179817 520258 179875 520292
rect 179909 520258 179967 520292
rect 180001 520258 180059 520292
rect 180093 520258 180151 520292
rect 180185 520258 180243 520292
rect 180277 520258 180335 520292
rect 180369 520258 180427 520292
rect 180461 520258 180519 520292
rect 180553 520258 180611 520292
rect 180645 520258 180703 520292
rect 180737 520258 180795 520292
rect 180829 520258 180887 520292
rect 180921 520258 180979 520292
rect 181013 520258 181071 520292
rect 181105 520258 181163 520292
rect 181197 520258 181255 520292
rect 181289 520258 181347 520292
rect 181381 520258 181439 520292
rect 181473 520258 181531 520292
rect 181565 520258 181601 520292
rect 181657 520258 181665 520292
rect 177963 520249 177975 520258
rect 178027 520249 178039 520258
rect 178091 520249 181601 520258
rect 181653 520249 181665 520258
rect 181717 520249 181729 520258
rect 181781 520249 181793 520301
rect 181845 520249 181857 520301
rect 181909 520292 185419 520301
rect 181933 520258 181991 520292
rect 182025 520258 182083 520292
rect 182117 520258 182175 520292
rect 182209 520258 182267 520292
rect 182301 520258 182359 520292
rect 182393 520258 182451 520292
rect 182485 520258 182543 520292
rect 182577 520258 182635 520292
rect 182669 520258 182727 520292
rect 182761 520258 182819 520292
rect 182853 520258 182911 520292
rect 182945 520258 183003 520292
rect 183037 520258 183095 520292
rect 183129 520258 183187 520292
rect 183221 520258 183279 520292
rect 183313 520258 183371 520292
rect 183405 520258 183463 520292
rect 183497 520258 183555 520292
rect 183589 520258 183647 520292
rect 183681 520258 183739 520292
rect 183773 520258 183831 520292
rect 183865 520258 183923 520292
rect 183957 520258 184015 520292
rect 184049 520258 184107 520292
rect 184141 520258 184199 520292
rect 184233 520258 184291 520292
rect 184325 520258 184383 520292
rect 184417 520258 184475 520292
rect 184509 520258 184567 520292
rect 184601 520258 184659 520292
rect 184693 520258 184751 520292
rect 184785 520258 184843 520292
rect 184877 520258 184935 520292
rect 184969 520258 185027 520292
rect 185061 520258 185119 520292
rect 185153 520258 185211 520292
rect 185245 520258 185303 520292
rect 185337 520258 185395 520292
rect 181909 520249 185419 520258
rect 185471 520249 185483 520301
rect 185535 520249 185547 520301
rect 185599 520292 185611 520301
rect 185663 520292 185675 520301
rect 185727 520292 187482 520301
rect 185663 520258 185671 520292
rect 185727 520258 185763 520292
rect 185797 520258 185855 520292
rect 185889 520258 185947 520292
rect 185981 520258 186039 520292
rect 186073 520258 186131 520292
rect 186165 520258 186223 520292
rect 186257 520258 186315 520292
rect 186349 520258 186407 520292
rect 186441 520258 186499 520292
rect 186533 520258 186591 520292
rect 186625 520258 186683 520292
rect 186717 520258 186775 520292
rect 186809 520258 186867 520292
rect 186901 520258 186959 520292
rect 186993 520258 187051 520292
rect 187085 520258 187143 520292
rect 187177 520258 187235 520292
rect 187269 520258 187327 520292
rect 187361 520258 187419 520292
rect 187453 520258 187482 520292
rect 185599 520249 185611 520258
rect 185663 520249 185675 520258
rect 185727 520249 187482 520258
rect 172210 520227 187482 520249
rect 172210 519757 187482 519779
rect 172210 519748 174625 519757
rect 172210 519714 172239 519748
rect 172273 519714 172331 519748
rect 172365 519714 172423 519748
rect 172457 519714 172515 519748
rect 172549 519714 172607 519748
rect 172641 519714 172699 519748
rect 172733 519714 172791 519748
rect 172825 519714 172883 519748
rect 172917 519714 172975 519748
rect 173009 519714 173067 519748
rect 173101 519714 173159 519748
rect 173193 519714 173251 519748
rect 173285 519714 173343 519748
rect 173377 519714 173435 519748
rect 173469 519714 173527 519748
rect 173561 519714 173619 519748
rect 173653 519714 173711 519748
rect 173745 519714 173803 519748
rect 173837 519714 173895 519748
rect 173929 519714 173987 519748
rect 174021 519714 174079 519748
rect 174113 519714 174171 519748
rect 174205 519714 174263 519748
rect 174297 519714 174355 519748
rect 174389 519714 174447 519748
rect 174481 519714 174539 519748
rect 174573 519714 174625 519748
rect 172210 519705 174625 519714
rect 174677 519705 174689 519757
rect 174741 519748 174753 519757
rect 174805 519748 174817 519757
rect 174805 519714 174815 519748
rect 174741 519705 174753 519714
rect 174805 519705 174817 519714
rect 174869 519705 174881 519757
rect 174933 519748 178443 519757
rect 174941 519714 174999 519748
rect 175033 519714 175091 519748
rect 175125 519714 175183 519748
rect 175217 519714 175275 519748
rect 175309 519714 175367 519748
rect 175401 519714 175459 519748
rect 175493 519714 175551 519748
rect 175585 519714 175643 519748
rect 175677 519714 175735 519748
rect 175769 519714 175827 519748
rect 175861 519714 175919 519748
rect 175953 519714 176011 519748
rect 176045 519714 176103 519748
rect 176137 519714 176195 519748
rect 176229 519714 176287 519748
rect 176321 519714 176379 519748
rect 176413 519714 176471 519748
rect 176505 519714 176563 519748
rect 176597 519714 176655 519748
rect 176689 519714 176747 519748
rect 176781 519714 176839 519748
rect 176873 519714 176931 519748
rect 176965 519714 177023 519748
rect 177057 519714 177115 519748
rect 177149 519714 177207 519748
rect 177241 519714 177299 519748
rect 177333 519714 177391 519748
rect 177425 519714 177483 519748
rect 177517 519714 177575 519748
rect 177609 519714 177667 519748
rect 177701 519714 177759 519748
rect 177793 519714 177851 519748
rect 177885 519714 177943 519748
rect 177977 519714 178035 519748
rect 178069 519714 178127 519748
rect 178161 519714 178219 519748
rect 178253 519714 178311 519748
rect 178345 519714 178403 519748
rect 178437 519714 178443 519748
rect 174933 519705 178443 519714
rect 178495 519748 178507 519757
rect 178495 519705 178507 519714
rect 178559 519705 178571 519757
rect 178623 519705 178635 519757
rect 178687 519748 178699 519757
rect 178751 519748 182261 519757
rect 178751 519714 178771 519748
rect 178805 519714 178863 519748
rect 178897 519714 178955 519748
rect 178989 519714 179047 519748
rect 179081 519714 179139 519748
rect 179173 519714 179231 519748
rect 179265 519714 179323 519748
rect 179357 519714 179415 519748
rect 179449 519714 179507 519748
rect 179541 519714 179599 519748
rect 179633 519714 179691 519748
rect 179725 519714 179783 519748
rect 179817 519714 179875 519748
rect 179909 519714 179967 519748
rect 180001 519714 180059 519748
rect 180093 519714 180151 519748
rect 180185 519714 180243 519748
rect 180277 519714 180335 519748
rect 180369 519714 180427 519748
rect 180461 519714 180519 519748
rect 180553 519714 180611 519748
rect 180645 519714 180703 519748
rect 180737 519714 180795 519748
rect 180829 519714 180887 519748
rect 180921 519714 180979 519748
rect 181013 519714 181071 519748
rect 181105 519714 181163 519748
rect 181197 519714 181255 519748
rect 181289 519714 181347 519748
rect 181381 519714 181439 519748
rect 181473 519714 181531 519748
rect 181565 519714 181623 519748
rect 181657 519714 181715 519748
rect 181749 519714 181807 519748
rect 181841 519714 181899 519748
rect 181933 519714 181991 519748
rect 182025 519714 182083 519748
rect 182117 519714 182175 519748
rect 182209 519714 182261 519748
rect 178687 519705 178699 519714
rect 178751 519705 182261 519714
rect 182313 519705 182325 519757
rect 182377 519748 182389 519757
rect 182441 519748 182453 519757
rect 182441 519714 182451 519748
rect 182377 519705 182389 519714
rect 182441 519705 182453 519714
rect 182505 519705 182517 519757
rect 182569 519748 186079 519757
rect 182577 519714 182635 519748
rect 182669 519714 182727 519748
rect 182761 519714 182819 519748
rect 182853 519714 182911 519748
rect 182945 519714 183003 519748
rect 183037 519714 183095 519748
rect 183129 519714 183187 519748
rect 183221 519714 183279 519748
rect 183313 519714 183371 519748
rect 183405 519714 183463 519748
rect 183497 519714 183555 519748
rect 183589 519714 183647 519748
rect 183681 519714 183739 519748
rect 183773 519714 183831 519748
rect 183865 519714 183923 519748
rect 183957 519714 184015 519748
rect 184049 519714 184107 519748
rect 184141 519714 184199 519748
rect 184233 519714 184291 519748
rect 184325 519714 184383 519748
rect 184417 519714 184475 519748
rect 184509 519714 184567 519748
rect 184601 519714 184659 519748
rect 184693 519714 184751 519748
rect 184785 519714 184843 519748
rect 184877 519714 184935 519748
rect 184969 519714 185027 519748
rect 185061 519714 185119 519748
rect 185153 519714 185211 519748
rect 185245 519714 185303 519748
rect 185337 519714 185395 519748
rect 185429 519714 185487 519748
rect 185521 519714 185579 519748
rect 185613 519714 185671 519748
rect 185705 519714 185763 519748
rect 185797 519714 185855 519748
rect 185889 519714 185947 519748
rect 185981 519714 186039 519748
rect 186073 519714 186079 519748
rect 182569 519705 186079 519714
rect 186131 519748 186143 519757
rect 186131 519705 186143 519714
rect 186195 519705 186207 519757
rect 186259 519705 186271 519757
rect 186323 519748 186335 519757
rect 186387 519748 187482 519757
rect 186387 519714 186407 519748
rect 186441 519714 186499 519748
rect 186533 519714 186591 519748
rect 186625 519714 186683 519748
rect 186717 519714 186775 519748
rect 186809 519714 186867 519748
rect 186901 519714 186959 519748
rect 186993 519714 187051 519748
rect 187085 519714 187143 519748
rect 187177 519714 187235 519748
rect 187269 519714 187327 519748
rect 187361 519714 187419 519748
rect 187453 519714 187482 519748
rect 186323 519705 186335 519714
rect 186387 519705 187482 519714
rect 172210 519683 187482 519705
rect 172210 519213 187482 519235
rect 172210 519204 173965 519213
rect 174017 519204 174029 519213
rect 174081 519204 174093 519213
rect 172210 519170 172239 519204
rect 172273 519170 172331 519204
rect 172365 519170 172423 519204
rect 172457 519170 172515 519204
rect 172549 519170 172607 519204
rect 172641 519170 172699 519204
rect 172733 519170 172791 519204
rect 172825 519170 172883 519204
rect 172917 519170 172975 519204
rect 173009 519170 173067 519204
rect 173101 519170 173159 519204
rect 173193 519170 173251 519204
rect 173285 519170 173343 519204
rect 173377 519170 173435 519204
rect 173469 519170 173527 519204
rect 173561 519170 173619 519204
rect 173653 519170 173711 519204
rect 173745 519170 173803 519204
rect 173837 519170 173895 519204
rect 173929 519170 173965 519204
rect 174021 519170 174029 519204
rect 172210 519161 173965 519170
rect 174017 519161 174029 519170
rect 174081 519161 174093 519170
rect 174145 519161 174157 519213
rect 174209 519161 174221 519213
rect 174273 519204 177783 519213
rect 174297 519170 174355 519204
rect 174389 519170 174447 519204
rect 174481 519170 174539 519204
rect 174573 519170 174631 519204
rect 174665 519170 174723 519204
rect 174757 519170 174815 519204
rect 174849 519170 174907 519204
rect 174941 519170 174999 519204
rect 175033 519170 175091 519204
rect 175125 519170 175183 519204
rect 175217 519170 175275 519204
rect 175309 519170 175367 519204
rect 175401 519170 175459 519204
rect 175493 519170 175551 519204
rect 175585 519170 175643 519204
rect 175677 519170 175735 519204
rect 175769 519170 175827 519204
rect 175861 519170 175919 519204
rect 175953 519170 176011 519204
rect 176045 519170 176103 519204
rect 176137 519170 176195 519204
rect 176229 519170 176287 519204
rect 176321 519170 176379 519204
rect 176413 519170 176471 519204
rect 176505 519170 176563 519204
rect 176597 519170 176655 519204
rect 176689 519170 176747 519204
rect 176781 519170 176839 519204
rect 176873 519170 176931 519204
rect 176965 519170 177023 519204
rect 177057 519170 177115 519204
rect 177149 519170 177207 519204
rect 177241 519170 177299 519204
rect 177333 519170 177391 519204
rect 177425 519170 177483 519204
rect 177517 519170 177575 519204
rect 177609 519170 177667 519204
rect 177701 519170 177759 519204
rect 174273 519161 177783 519170
rect 177835 519161 177847 519213
rect 177899 519161 177911 519213
rect 177963 519204 177975 519213
rect 178027 519204 178039 519213
rect 178091 519204 181601 519213
rect 181653 519204 181665 519213
rect 181717 519204 181729 519213
rect 178027 519170 178035 519204
rect 178091 519170 178127 519204
rect 178161 519170 178219 519204
rect 178253 519170 178311 519204
rect 178345 519170 178403 519204
rect 178437 519170 178495 519204
rect 178529 519170 178587 519204
rect 178621 519170 178679 519204
rect 178713 519170 178771 519204
rect 178805 519170 178863 519204
rect 178897 519170 178955 519204
rect 178989 519170 179047 519204
rect 179081 519170 179139 519204
rect 179173 519170 179231 519204
rect 179265 519170 179323 519204
rect 179357 519170 179415 519204
rect 179449 519170 179507 519204
rect 179541 519170 179599 519204
rect 179633 519170 179691 519204
rect 179725 519170 179783 519204
rect 179817 519170 179875 519204
rect 179909 519170 179967 519204
rect 180001 519170 180059 519204
rect 180093 519170 180151 519204
rect 180185 519170 180243 519204
rect 180277 519170 180335 519204
rect 180369 519170 180427 519204
rect 180461 519170 180519 519204
rect 180553 519170 180611 519204
rect 180645 519170 180703 519204
rect 180737 519170 180795 519204
rect 180829 519170 180887 519204
rect 180921 519170 180979 519204
rect 181013 519170 181071 519204
rect 181105 519170 181163 519204
rect 181197 519170 181255 519204
rect 181289 519170 181347 519204
rect 181381 519170 181439 519204
rect 181473 519170 181531 519204
rect 181565 519170 181601 519204
rect 181657 519170 181665 519204
rect 177963 519161 177975 519170
rect 178027 519161 178039 519170
rect 178091 519161 181601 519170
rect 181653 519161 181665 519170
rect 181717 519161 181729 519170
rect 181781 519161 181793 519213
rect 181845 519161 181857 519213
rect 181909 519204 185419 519213
rect 181933 519170 181991 519204
rect 182025 519170 182083 519204
rect 182117 519170 182175 519204
rect 182209 519170 182267 519204
rect 182301 519170 182359 519204
rect 182393 519170 182451 519204
rect 182485 519170 182543 519204
rect 182577 519170 182635 519204
rect 182669 519170 182727 519204
rect 182761 519170 182819 519204
rect 182853 519170 182911 519204
rect 182945 519170 183003 519204
rect 183037 519170 183095 519204
rect 183129 519170 183187 519204
rect 183221 519170 183279 519204
rect 183313 519170 183371 519204
rect 183405 519170 183463 519204
rect 183497 519170 183555 519204
rect 183589 519170 183647 519204
rect 183681 519170 183739 519204
rect 183773 519170 183831 519204
rect 183865 519170 183923 519204
rect 183957 519170 184015 519204
rect 184049 519170 184107 519204
rect 184141 519170 184199 519204
rect 184233 519170 184291 519204
rect 184325 519170 184383 519204
rect 184417 519170 184475 519204
rect 184509 519170 184567 519204
rect 184601 519170 184659 519204
rect 184693 519170 184751 519204
rect 184785 519170 184843 519204
rect 184877 519170 184935 519204
rect 184969 519170 185027 519204
rect 185061 519170 185119 519204
rect 185153 519170 185211 519204
rect 185245 519170 185303 519204
rect 185337 519170 185395 519204
rect 181909 519161 185419 519170
rect 185471 519161 185483 519213
rect 185535 519161 185547 519213
rect 185599 519204 185611 519213
rect 185663 519204 185675 519213
rect 185727 519204 187482 519213
rect 185663 519170 185671 519204
rect 185727 519170 185763 519204
rect 185797 519170 185855 519204
rect 185889 519170 185947 519204
rect 185981 519170 186039 519204
rect 186073 519170 186131 519204
rect 186165 519170 186223 519204
rect 186257 519170 186315 519204
rect 186349 519170 186407 519204
rect 186441 519170 186499 519204
rect 186533 519170 186591 519204
rect 186625 519170 186683 519204
rect 186717 519170 186775 519204
rect 186809 519170 186867 519204
rect 186901 519170 186959 519204
rect 186993 519170 187051 519204
rect 187085 519170 187143 519204
rect 187177 519170 187235 519204
rect 187269 519170 187327 519204
rect 187361 519170 187419 519204
rect 187453 519170 187482 519204
rect 185599 519161 185611 519170
rect 185663 519161 185675 519170
rect 185727 519161 187482 519170
rect 172210 519139 187482 519161
rect 172210 518669 187482 518691
rect 172210 518660 174625 518669
rect 172210 518626 172239 518660
rect 172273 518626 172331 518660
rect 172365 518626 172423 518660
rect 172457 518626 172515 518660
rect 172549 518626 172607 518660
rect 172641 518626 172699 518660
rect 172733 518626 172791 518660
rect 172825 518626 172883 518660
rect 172917 518626 172975 518660
rect 173009 518626 173067 518660
rect 173101 518626 173159 518660
rect 173193 518626 173251 518660
rect 173285 518626 173343 518660
rect 173377 518626 173435 518660
rect 173469 518626 173527 518660
rect 173561 518626 173619 518660
rect 173653 518626 173711 518660
rect 173745 518626 173803 518660
rect 173837 518626 173895 518660
rect 173929 518626 173987 518660
rect 174021 518626 174079 518660
rect 174113 518626 174171 518660
rect 174205 518626 174263 518660
rect 174297 518626 174355 518660
rect 174389 518626 174447 518660
rect 174481 518626 174539 518660
rect 174573 518626 174625 518660
rect 172210 518617 174625 518626
rect 174677 518617 174689 518669
rect 174741 518660 174753 518669
rect 174805 518660 174817 518669
rect 174805 518626 174815 518660
rect 174741 518617 174753 518626
rect 174805 518617 174817 518626
rect 174869 518617 174881 518669
rect 174933 518660 178443 518669
rect 174941 518626 174999 518660
rect 175033 518626 175091 518660
rect 175125 518626 175183 518660
rect 175217 518626 175275 518660
rect 175309 518626 175367 518660
rect 175401 518626 175459 518660
rect 175493 518626 175551 518660
rect 175585 518626 175643 518660
rect 175677 518626 175735 518660
rect 175769 518626 175827 518660
rect 175861 518626 175919 518660
rect 175953 518626 176011 518660
rect 176045 518626 176103 518660
rect 176137 518626 176195 518660
rect 176229 518626 176287 518660
rect 176321 518626 176379 518660
rect 176413 518626 176471 518660
rect 176505 518626 176563 518660
rect 176597 518626 176655 518660
rect 176689 518626 176747 518660
rect 176781 518626 176839 518660
rect 176873 518626 176931 518660
rect 176965 518626 177023 518660
rect 177057 518626 177115 518660
rect 177149 518626 177207 518660
rect 177241 518626 177299 518660
rect 177333 518626 177391 518660
rect 177425 518626 177483 518660
rect 177517 518626 177575 518660
rect 177609 518626 177667 518660
rect 177701 518626 177759 518660
rect 177793 518626 177851 518660
rect 177885 518626 177943 518660
rect 177977 518626 178035 518660
rect 178069 518626 178127 518660
rect 178161 518626 178219 518660
rect 178253 518626 178311 518660
rect 178345 518626 178403 518660
rect 178437 518626 178443 518660
rect 174933 518617 178443 518626
rect 178495 518660 178507 518669
rect 178495 518617 178507 518626
rect 178559 518617 178571 518669
rect 178623 518617 178635 518669
rect 178687 518660 178699 518669
rect 178751 518660 182261 518669
rect 178751 518626 178771 518660
rect 178805 518626 178863 518660
rect 178897 518626 178955 518660
rect 178989 518626 179047 518660
rect 179081 518626 179139 518660
rect 179173 518626 179231 518660
rect 179265 518626 179323 518660
rect 179357 518626 179415 518660
rect 179449 518626 179507 518660
rect 179541 518626 179599 518660
rect 179633 518626 179691 518660
rect 179725 518626 179783 518660
rect 179817 518626 179875 518660
rect 179909 518626 179967 518660
rect 180001 518626 180059 518660
rect 180093 518626 180151 518660
rect 180185 518626 180243 518660
rect 180277 518626 180335 518660
rect 180369 518626 180427 518660
rect 180461 518626 180519 518660
rect 180553 518626 180611 518660
rect 180645 518626 180703 518660
rect 180737 518626 180795 518660
rect 180829 518626 180887 518660
rect 180921 518626 180979 518660
rect 181013 518626 181071 518660
rect 181105 518626 181163 518660
rect 181197 518626 181255 518660
rect 181289 518626 181347 518660
rect 181381 518626 181439 518660
rect 181473 518626 181531 518660
rect 181565 518626 181623 518660
rect 181657 518626 181715 518660
rect 181749 518626 181807 518660
rect 181841 518626 181899 518660
rect 181933 518626 181991 518660
rect 182025 518626 182083 518660
rect 182117 518626 182175 518660
rect 182209 518626 182261 518660
rect 178687 518617 178699 518626
rect 178751 518617 182261 518626
rect 182313 518617 182325 518669
rect 182377 518660 182389 518669
rect 182441 518660 182453 518669
rect 182441 518626 182451 518660
rect 182377 518617 182389 518626
rect 182441 518617 182453 518626
rect 182505 518617 182517 518669
rect 182569 518660 186079 518669
rect 182577 518626 182635 518660
rect 182669 518626 182727 518660
rect 182761 518626 182819 518660
rect 182853 518626 182911 518660
rect 182945 518626 183003 518660
rect 183037 518626 183095 518660
rect 183129 518626 183187 518660
rect 183221 518626 183279 518660
rect 183313 518626 183371 518660
rect 183405 518626 183463 518660
rect 183497 518626 183555 518660
rect 183589 518626 183647 518660
rect 183681 518626 183739 518660
rect 183773 518626 183831 518660
rect 183865 518626 183923 518660
rect 183957 518626 184015 518660
rect 184049 518626 184107 518660
rect 184141 518626 184199 518660
rect 184233 518626 184291 518660
rect 184325 518626 184383 518660
rect 184417 518626 184475 518660
rect 184509 518626 184567 518660
rect 184601 518626 184659 518660
rect 184693 518626 184751 518660
rect 184785 518626 184843 518660
rect 184877 518626 184935 518660
rect 184969 518626 185027 518660
rect 185061 518626 185119 518660
rect 185153 518626 185211 518660
rect 185245 518626 185303 518660
rect 185337 518626 185395 518660
rect 185429 518626 185487 518660
rect 185521 518626 185579 518660
rect 185613 518626 185671 518660
rect 185705 518626 185763 518660
rect 185797 518626 185855 518660
rect 185889 518626 185947 518660
rect 185981 518626 186039 518660
rect 186073 518626 186079 518660
rect 182569 518617 186079 518626
rect 186131 518660 186143 518669
rect 186131 518617 186143 518626
rect 186195 518617 186207 518669
rect 186259 518617 186271 518669
rect 186323 518660 186335 518669
rect 186387 518660 187482 518669
rect 186387 518626 186407 518660
rect 186441 518626 186499 518660
rect 186533 518626 186591 518660
rect 186625 518626 186683 518660
rect 186717 518626 186775 518660
rect 186809 518626 186867 518660
rect 186901 518626 186959 518660
rect 186993 518626 187051 518660
rect 187085 518626 187143 518660
rect 187177 518626 187235 518660
rect 187269 518626 187327 518660
rect 187361 518626 187419 518660
rect 187453 518626 187482 518660
rect 186323 518617 186335 518626
rect 186387 518617 187482 518626
rect 172210 518595 187482 518617
rect 172210 518125 187482 518147
rect 172210 518116 173965 518125
rect 174017 518116 174029 518125
rect 174081 518116 174093 518125
rect 172210 518082 172239 518116
rect 172273 518082 172331 518116
rect 172365 518082 172423 518116
rect 172457 518082 172515 518116
rect 172549 518082 172607 518116
rect 172641 518082 172699 518116
rect 172733 518082 172791 518116
rect 172825 518082 172883 518116
rect 172917 518082 172975 518116
rect 173009 518082 173067 518116
rect 173101 518082 173159 518116
rect 173193 518082 173251 518116
rect 173285 518082 173343 518116
rect 173377 518082 173435 518116
rect 173469 518082 173527 518116
rect 173561 518082 173619 518116
rect 173653 518082 173711 518116
rect 173745 518082 173803 518116
rect 173837 518082 173895 518116
rect 173929 518082 173965 518116
rect 174021 518082 174029 518116
rect 172210 518073 173965 518082
rect 174017 518073 174029 518082
rect 174081 518073 174093 518082
rect 174145 518073 174157 518125
rect 174209 518073 174221 518125
rect 174273 518116 177783 518125
rect 174297 518082 174355 518116
rect 174389 518082 174447 518116
rect 174481 518082 174539 518116
rect 174573 518082 174631 518116
rect 174665 518082 174723 518116
rect 174757 518082 174815 518116
rect 174849 518082 174907 518116
rect 174941 518082 174999 518116
rect 175033 518082 175091 518116
rect 175125 518082 175183 518116
rect 175217 518082 175275 518116
rect 175309 518082 175367 518116
rect 175401 518082 175459 518116
rect 175493 518082 175551 518116
rect 175585 518082 175643 518116
rect 175677 518082 175735 518116
rect 175769 518082 175827 518116
rect 175861 518082 175919 518116
rect 175953 518082 176011 518116
rect 176045 518082 176103 518116
rect 176137 518082 176195 518116
rect 176229 518082 176287 518116
rect 176321 518082 176379 518116
rect 176413 518082 176471 518116
rect 176505 518082 176563 518116
rect 176597 518082 176655 518116
rect 176689 518082 176747 518116
rect 176781 518082 176839 518116
rect 176873 518082 176931 518116
rect 176965 518082 177023 518116
rect 177057 518082 177115 518116
rect 177149 518082 177207 518116
rect 177241 518082 177299 518116
rect 177333 518082 177391 518116
rect 177425 518082 177483 518116
rect 177517 518082 177575 518116
rect 177609 518082 177667 518116
rect 177701 518082 177759 518116
rect 174273 518073 177783 518082
rect 177835 518073 177847 518125
rect 177899 518073 177911 518125
rect 177963 518116 177975 518125
rect 178027 518116 178039 518125
rect 178091 518116 181601 518125
rect 181653 518116 181665 518125
rect 181717 518116 181729 518125
rect 178027 518082 178035 518116
rect 178091 518082 178127 518116
rect 178161 518082 178219 518116
rect 178253 518082 178311 518116
rect 178345 518082 178403 518116
rect 178437 518082 178495 518116
rect 178529 518082 178587 518116
rect 178621 518082 178679 518116
rect 178713 518082 178771 518116
rect 178805 518082 178863 518116
rect 178897 518082 178955 518116
rect 178989 518082 179047 518116
rect 179081 518082 179139 518116
rect 179173 518082 179231 518116
rect 179265 518082 179323 518116
rect 179357 518082 179415 518116
rect 179449 518082 179507 518116
rect 179541 518082 179599 518116
rect 179633 518082 179691 518116
rect 179725 518082 179783 518116
rect 179817 518082 179875 518116
rect 179909 518082 179967 518116
rect 180001 518082 180059 518116
rect 180093 518082 180151 518116
rect 180185 518082 180243 518116
rect 180277 518082 180335 518116
rect 180369 518082 180427 518116
rect 180461 518082 180519 518116
rect 180553 518082 180611 518116
rect 180645 518082 180703 518116
rect 180737 518082 180795 518116
rect 180829 518082 180887 518116
rect 180921 518082 180979 518116
rect 181013 518082 181071 518116
rect 181105 518082 181163 518116
rect 181197 518082 181255 518116
rect 181289 518082 181347 518116
rect 181381 518082 181439 518116
rect 181473 518082 181531 518116
rect 181565 518082 181601 518116
rect 181657 518082 181665 518116
rect 177963 518073 177975 518082
rect 178027 518073 178039 518082
rect 178091 518073 181601 518082
rect 181653 518073 181665 518082
rect 181717 518073 181729 518082
rect 181781 518073 181793 518125
rect 181845 518073 181857 518125
rect 181909 518116 185419 518125
rect 181933 518082 181991 518116
rect 182025 518082 182083 518116
rect 182117 518082 182175 518116
rect 182209 518082 182267 518116
rect 182301 518082 182359 518116
rect 182393 518082 182451 518116
rect 182485 518082 182543 518116
rect 182577 518082 182635 518116
rect 182669 518082 182727 518116
rect 182761 518082 182819 518116
rect 182853 518082 182911 518116
rect 182945 518082 183003 518116
rect 183037 518082 183095 518116
rect 183129 518082 183187 518116
rect 183221 518082 183279 518116
rect 183313 518082 183371 518116
rect 183405 518082 183463 518116
rect 183497 518082 183555 518116
rect 183589 518082 183647 518116
rect 183681 518082 183739 518116
rect 183773 518082 183831 518116
rect 183865 518082 183923 518116
rect 183957 518082 184015 518116
rect 184049 518082 184107 518116
rect 184141 518082 184199 518116
rect 184233 518082 184291 518116
rect 184325 518082 184383 518116
rect 184417 518082 184475 518116
rect 184509 518082 184567 518116
rect 184601 518082 184659 518116
rect 184693 518082 184751 518116
rect 184785 518082 184843 518116
rect 184877 518082 184935 518116
rect 184969 518082 185027 518116
rect 185061 518082 185119 518116
rect 185153 518082 185211 518116
rect 185245 518082 185303 518116
rect 185337 518082 185395 518116
rect 181909 518073 185419 518082
rect 185471 518073 185483 518125
rect 185535 518073 185547 518125
rect 185599 518116 185611 518125
rect 185663 518116 185675 518125
rect 185727 518116 187482 518125
rect 185663 518082 185671 518116
rect 185727 518082 185763 518116
rect 185797 518082 185855 518116
rect 185889 518082 185947 518116
rect 185981 518082 186039 518116
rect 186073 518082 186131 518116
rect 186165 518082 186223 518116
rect 186257 518082 186315 518116
rect 186349 518082 186407 518116
rect 186441 518082 186499 518116
rect 186533 518082 186591 518116
rect 186625 518082 186683 518116
rect 186717 518082 186775 518116
rect 186809 518082 186867 518116
rect 186901 518082 186959 518116
rect 186993 518082 187051 518116
rect 187085 518082 187143 518116
rect 187177 518082 187235 518116
rect 187269 518082 187327 518116
rect 187361 518082 187419 518116
rect 187453 518082 187482 518116
rect 185599 518073 185611 518082
rect 185663 518073 185675 518082
rect 185727 518073 187482 518082
rect 172210 518051 187482 518073
rect 172210 517581 187482 517603
rect 172210 517572 174625 517581
rect 172210 517538 172239 517572
rect 172273 517538 172331 517572
rect 172365 517538 172423 517572
rect 172457 517538 172515 517572
rect 172549 517538 172607 517572
rect 172641 517538 172699 517572
rect 172733 517538 172791 517572
rect 172825 517538 172883 517572
rect 172917 517538 172975 517572
rect 173009 517538 173067 517572
rect 173101 517538 173159 517572
rect 173193 517538 173251 517572
rect 173285 517538 173343 517572
rect 173377 517538 173435 517572
rect 173469 517538 173527 517572
rect 173561 517538 173619 517572
rect 173653 517538 173711 517572
rect 173745 517538 173803 517572
rect 173837 517538 173895 517572
rect 173929 517538 173987 517572
rect 174021 517538 174079 517572
rect 174113 517538 174171 517572
rect 174205 517538 174263 517572
rect 174297 517538 174355 517572
rect 174389 517538 174447 517572
rect 174481 517538 174539 517572
rect 174573 517538 174625 517572
rect 172210 517529 174625 517538
rect 174677 517529 174689 517581
rect 174741 517572 174753 517581
rect 174805 517572 174817 517581
rect 174805 517538 174815 517572
rect 174741 517529 174753 517538
rect 174805 517529 174817 517538
rect 174869 517529 174881 517581
rect 174933 517572 178443 517581
rect 174941 517538 174999 517572
rect 175033 517538 175091 517572
rect 175125 517538 175183 517572
rect 175217 517538 175275 517572
rect 175309 517538 175367 517572
rect 175401 517538 175459 517572
rect 175493 517538 175551 517572
rect 175585 517538 175643 517572
rect 175677 517538 175735 517572
rect 175769 517538 175827 517572
rect 175861 517538 175919 517572
rect 175953 517538 176011 517572
rect 176045 517538 176103 517572
rect 176137 517538 176195 517572
rect 176229 517538 176287 517572
rect 176321 517538 176379 517572
rect 176413 517538 176471 517572
rect 176505 517538 176563 517572
rect 176597 517538 176655 517572
rect 176689 517538 176747 517572
rect 176781 517538 176839 517572
rect 176873 517538 176931 517572
rect 176965 517538 177023 517572
rect 177057 517538 177115 517572
rect 177149 517538 177207 517572
rect 177241 517538 177299 517572
rect 177333 517538 177391 517572
rect 177425 517538 177483 517572
rect 177517 517538 177575 517572
rect 177609 517538 177667 517572
rect 177701 517538 177759 517572
rect 177793 517538 177851 517572
rect 177885 517538 177943 517572
rect 177977 517538 178035 517572
rect 178069 517538 178127 517572
rect 178161 517538 178219 517572
rect 178253 517538 178311 517572
rect 178345 517538 178403 517572
rect 178437 517538 178443 517572
rect 174933 517529 178443 517538
rect 178495 517572 178507 517581
rect 178495 517529 178507 517538
rect 178559 517529 178571 517581
rect 178623 517529 178635 517581
rect 178687 517572 178699 517581
rect 178751 517572 182261 517581
rect 178751 517538 178771 517572
rect 178805 517538 178863 517572
rect 178897 517538 178955 517572
rect 178989 517538 179047 517572
rect 179081 517538 179139 517572
rect 179173 517538 179231 517572
rect 179265 517538 179323 517572
rect 179357 517538 179415 517572
rect 179449 517538 179507 517572
rect 179541 517538 179599 517572
rect 179633 517538 179691 517572
rect 179725 517538 179783 517572
rect 179817 517538 179875 517572
rect 179909 517538 179967 517572
rect 180001 517538 180059 517572
rect 180093 517538 180151 517572
rect 180185 517538 180243 517572
rect 180277 517538 180335 517572
rect 180369 517538 180427 517572
rect 180461 517538 180519 517572
rect 180553 517538 180611 517572
rect 180645 517538 180703 517572
rect 180737 517538 180795 517572
rect 180829 517538 180887 517572
rect 180921 517538 180979 517572
rect 181013 517538 181071 517572
rect 181105 517538 181163 517572
rect 181197 517538 181255 517572
rect 181289 517538 181347 517572
rect 181381 517538 181439 517572
rect 181473 517538 181531 517572
rect 181565 517538 181623 517572
rect 181657 517538 181715 517572
rect 181749 517538 181807 517572
rect 181841 517538 181899 517572
rect 181933 517538 181991 517572
rect 182025 517538 182083 517572
rect 182117 517538 182175 517572
rect 182209 517538 182261 517572
rect 178687 517529 178699 517538
rect 178751 517529 182261 517538
rect 182313 517529 182325 517581
rect 182377 517572 182389 517581
rect 182441 517572 182453 517581
rect 182441 517538 182451 517572
rect 182377 517529 182389 517538
rect 182441 517529 182453 517538
rect 182505 517529 182517 517581
rect 182569 517572 186079 517581
rect 182577 517538 182635 517572
rect 182669 517538 182727 517572
rect 182761 517538 182819 517572
rect 182853 517538 182911 517572
rect 182945 517538 183003 517572
rect 183037 517538 183095 517572
rect 183129 517538 183187 517572
rect 183221 517538 183279 517572
rect 183313 517538 183371 517572
rect 183405 517538 183463 517572
rect 183497 517538 183555 517572
rect 183589 517538 183647 517572
rect 183681 517538 183739 517572
rect 183773 517538 183831 517572
rect 183865 517538 183923 517572
rect 183957 517538 184015 517572
rect 184049 517538 184107 517572
rect 184141 517538 184199 517572
rect 184233 517538 184291 517572
rect 184325 517538 184383 517572
rect 184417 517538 184475 517572
rect 184509 517538 184567 517572
rect 184601 517538 184659 517572
rect 184693 517538 184751 517572
rect 184785 517538 184843 517572
rect 184877 517538 184935 517572
rect 184969 517538 185027 517572
rect 185061 517538 185119 517572
rect 185153 517538 185211 517572
rect 185245 517538 185303 517572
rect 185337 517538 185395 517572
rect 185429 517538 185487 517572
rect 185521 517538 185579 517572
rect 185613 517538 185671 517572
rect 185705 517538 185763 517572
rect 185797 517538 185855 517572
rect 185889 517538 185947 517572
rect 185981 517538 186039 517572
rect 186073 517538 186079 517572
rect 182569 517529 186079 517538
rect 186131 517572 186143 517581
rect 186131 517529 186143 517538
rect 186195 517529 186207 517581
rect 186259 517529 186271 517581
rect 186323 517572 186335 517581
rect 186387 517572 187482 517581
rect 186387 517538 186407 517572
rect 186441 517538 186499 517572
rect 186533 517538 186591 517572
rect 186625 517538 186683 517572
rect 186717 517538 186775 517572
rect 186809 517538 186867 517572
rect 186901 517538 186959 517572
rect 186993 517538 187051 517572
rect 187085 517538 187143 517572
rect 187177 517538 187235 517572
rect 187269 517538 187327 517572
rect 187361 517538 187419 517572
rect 187453 517538 187482 517572
rect 186323 517529 186335 517538
rect 186387 517529 187482 517538
rect 172210 517507 187482 517529
rect 177652 517427 177658 517479
rect 177710 517467 177716 517479
rect 178296 517467 178302 517479
rect 177710 517439 178302 517467
rect 177710 517427 177716 517439
rect 178296 517427 178302 517439
rect 178354 517427 178360 517479
rect 172210 517037 187482 517059
rect 172210 517028 173965 517037
rect 174017 517028 174029 517037
rect 174081 517028 174093 517037
rect 172210 516994 172239 517028
rect 172273 516994 172331 517028
rect 172365 516994 172423 517028
rect 172457 516994 172515 517028
rect 172549 516994 172607 517028
rect 172641 516994 172699 517028
rect 172733 516994 172791 517028
rect 172825 516994 172883 517028
rect 172917 516994 172975 517028
rect 173009 516994 173067 517028
rect 173101 516994 173159 517028
rect 173193 516994 173251 517028
rect 173285 516994 173343 517028
rect 173377 516994 173435 517028
rect 173469 516994 173527 517028
rect 173561 516994 173619 517028
rect 173653 516994 173711 517028
rect 173745 516994 173803 517028
rect 173837 516994 173895 517028
rect 173929 516994 173965 517028
rect 174021 516994 174029 517028
rect 172210 516985 173965 516994
rect 174017 516985 174029 516994
rect 174081 516985 174093 516994
rect 174145 516985 174157 517037
rect 174209 516985 174221 517037
rect 174273 517028 177783 517037
rect 174297 516994 174355 517028
rect 174389 516994 174447 517028
rect 174481 516994 174539 517028
rect 174573 516994 174631 517028
rect 174665 516994 174723 517028
rect 174757 516994 174815 517028
rect 174849 516994 174907 517028
rect 174941 516994 174999 517028
rect 175033 516994 175091 517028
rect 175125 516994 175183 517028
rect 175217 516994 175275 517028
rect 175309 516994 175367 517028
rect 175401 516994 175459 517028
rect 175493 516994 175551 517028
rect 175585 516994 175643 517028
rect 175677 516994 175735 517028
rect 175769 516994 175827 517028
rect 175861 516994 175919 517028
rect 175953 516994 176011 517028
rect 176045 516994 176103 517028
rect 176137 516994 176195 517028
rect 176229 516994 176287 517028
rect 176321 516994 176379 517028
rect 176413 516994 176471 517028
rect 176505 516994 176563 517028
rect 176597 516994 176655 517028
rect 176689 516994 176747 517028
rect 176781 516994 176839 517028
rect 176873 516994 176931 517028
rect 176965 516994 177023 517028
rect 177057 516994 177115 517028
rect 177149 516994 177207 517028
rect 177241 516994 177299 517028
rect 177333 516994 177391 517028
rect 177425 516994 177483 517028
rect 177517 516994 177575 517028
rect 177609 516994 177667 517028
rect 177701 516994 177759 517028
rect 174273 516985 177783 516994
rect 177835 516985 177847 517037
rect 177899 516985 177911 517037
rect 177963 517028 177975 517037
rect 178027 517028 178039 517037
rect 178091 517028 181601 517037
rect 181653 517028 181665 517037
rect 181717 517028 181729 517037
rect 178027 516994 178035 517028
rect 178091 516994 178127 517028
rect 178161 516994 178219 517028
rect 178253 516994 178311 517028
rect 178345 516994 178403 517028
rect 178437 516994 178495 517028
rect 178529 516994 178587 517028
rect 178621 516994 178679 517028
rect 178713 516994 178771 517028
rect 178805 516994 178863 517028
rect 178897 516994 178955 517028
rect 178989 516994 179047 517028
rect 179081 516994 179139 517028
rect 179173 516994 179231 517028
rect 179265 516994 179323 517028
rect 179357 516994 179415 517028
rect 179449 516994 179507 517028
rect 179541 516994 179599 517028
rect 179633 516994 179691 517028
rect 179725 516994 179783 517028
rect 179817 516994 179875 517028
rect 179909 516994 179967 517028
rect 180001 516994 180059 517028
rect 180093 516994 180151 517028
rect 180185 516994 180243 517028
rect 180277 516994 180335 517028
rect 180369 516994 180427 517028
rect 180461 516994 180519 517028
rect 180553 516994 180611 517028
rect 180645 516994 180703 517028
rect 180737 516994 180795 517028
rect 180829 516994 180887 517028
rect 180921 516994 180979 517028
rect 181013 516994 181071 517028
rect 181105 516994 181163 517028
rect 181197 516994 181255 517028
rect 181289 516994 181347 517028
rect 181381 516994 181439 517028
rect 181473 516994 181531 517028
rect 181565 516994 181601 517028
rect 181657 516994 181665 517028
rect 177963 516985 177975 516994
rect 178027 516985 178039 516994
rect 178091 516985 181601 516994
rect 181653 516985 181665 516994
rect 181717 516985 181729 516994
rect 181781 516985 181793 517037
rect 181845 516985 181857 517037
rect 181909 517028 185419 517037
rect 181933 516994 181991 517028
rect 182025 516994 182083 517028
rect 182117 516994 182175 517028
rect 182209 516994 182267 517028
rect 182301 516994 182359 517028
rect 182393 516994 182451 517028
rect 182485 516994 182543 517028
rect 182577 516994 182635 517028
rect 182669 516994 182727 517028
rect 182761 516994 182819 517028
rect 182853 516994 182911 517028
rect 182945 516994 183003 517028
rect 183037 516994 183095 517028
rect 183129 516994 183187 517028
rect 183221 516994 183279 517028
rect 183313 516994 183371 517028
rect 183405 516994 183463 517028
rect 183497 516994 183555 517028
rect 183589 516994 183647 517028
rect 183681 516994 183739 517028
rect 183773 516994 183831 517028
rect 183865 516994 183923 517028
rect 183957 516994 184015 517028
rect 184049 516994 184107 517028
rect 184141 516994 184199 517028
rect 184233 516994 184291 517028
rect 184325 516994 184383 517028
rect 184417 516994 184475 517028
rect 184509 516994 184567 517028
rect 184601 516994 184659 517028
rect 184693 516994 184751 517028
rect 184785 516994 184843 517028
rect 184877 516994 184935 517028
rect 184969 516994 185027 517028
rect 185061 516994 185119 517028
rect 185153 516994 185211 517028
rect 185245 516994 185303 517028
rect 185337 516994 185395 517028
rect 181909 516985 185419 516994
rect 185471 516985 185483 517037
rect 185535 516985 185547 517037
rect 185599 517028 185611 517037
rect 185663 517028 185675 517037
rect 185727 517028 187482 517037
rect 185663 516994 185671 517028
rect 185727 516994 185763 517028
rect 185797 516994 185855 517028
rect 185889 516994 185947 517028
rect 185981 516994 186039 517028
rect 186073 516994 186131 517028
rect 186165 516994 186223 517028
rect 186257 516994 186315 517028
rect 186349 516994 186407 517028
rect 186441 516994 186499 517028
rect 186533 516994 186591 517028
rect 186625 516994 186683 517028
rect 186717 516994 186775 517028
rect 186809 516994 186867 517028
rect 186901 516994 186959 517028
rect 186993 516994 187051 517028
rect 187085 516994 187143 517028
rect 187177 516994 187235 517028
rect 187269 516994 187327 517028
rect 187361 516994 187419 517028
rect 187453 516994 187482 517028
rect 185599 516985 185611 516994
rect 185663 516985 185675 516994
rect 185727 516985 187482 516994
rect 172210 516963 187482 516985
rect 172210 516493 187482 516515
rect 172210 516484 174625 516493
rect 172210 516450 172239 516484
rect 172273 516450 172331 516484
rect 172365 516450 172423 516484
rect 172457 516450 172515 516484
rect 172549 516450 172607 516484
rect 172641 516450 172699 516484
rect 172733 516450 172791 516484
rect 172825 516450 172883 516484
rect 172917 516450 172975 516484
rect 173009 516450 173067 516484
rect 173101 516450 173159 516484
rect 173193 516450 173251 516484
rect 173285 516450 173343 516484
rect 173377 516450 173435 516484
rect 173469 516450 173527 516484
rect 173561 516450 173619 516484
rect 173653 516450 173711 516484
rect 173745 516450 173803 516484
rect 173837 516450 173895 516484
rect 173929 516450 173987 516484
rect 174021 516450 174079 516484
rect 174113 516450 174171 516484
rect 174205 516450 174263 516484
rect 174297 516450 174355 516484
rect 174389 516450 174447 516484
rect 174481 516450 174539 516484
rect 174573 516450 174625 516484
rect 172210 516441 174625 516450
rect 174677 516441 174689 516493
rect 174741 516484 174753 516493
rect 174805 516484 174817 516493
rect 174805 516450 174815 516484
rect 174741 516441 174753 516450
rect 174805 516441 174817 516450
rect 174869 516441 174881 516493
rect 174933 516484 178443 516493
rect 174941 516450 174999 516484
rect 175033 516450 175091 516484
rect 175125 516450 175183 516484
rect 175217 516450 175275 516484
rect 175309 516450 175367 516484
rect 175401 516450 175459 516484
rect 175493 516450 175551 516484
rect 175585 516450 175643 516484
rect 175677 516450 175735 516484
rect 175769 516450 175827 516484
rect 175861 516450 175919 516484
rect 175953 516450 176011 516484
rect 176045 516450 176103 516484
rect 176137 516450 176195 516484
rect 176229 516450 176287 516484
rect 176321 516450 176379 516484
rect 176413 516450 176471 516484
rect 176505 516450 176563 516484
rect 176597 516450 176655 516484
rect 176689 516450 176747 516484
rect 176781 516450 176839 516484
rect 176873 516450 176931 516484
rect 176965 516450 177023 516484
rect 177057 516450 177115 516484
rect 177149 516450 177207 516484
rect 177241 516450 177299 516484
rect 177333 516450 177391 516484
rect 177425 516450 177483 516484
rect 177517 516450 177575 516484
rect 177609 516450 177667 516484
rect 177701 516450 177759 516484
rect 177793 516450 177851 516484
rect 177885 516450 177943 516484
rect 177977 516450 178035 516484
rect 178069 516450 178127 516484
rect 178161 516450 178219 516484
rect 178253 516450 178311 516484
rect 178345 516450 178403 516484
rect 178437 516450 178443 516484
rect 174933 516441 178443 516450
rect 178495 516484 178507 516493
rect 178495 516441 178507 516450
rect 178559 516441 178571 516493
rect 178623 516441 178635 516493
rect 178687 516484 178699 516493
rect 178751 516484 182261 516493
rect 178751 516450 178771 516484
rect 178805 516450 178863 516484
rect 178897 516450 178955 516484
rect 178989 516450 179047 516484
rect 179081 516450 179139 516484
rect 179173 516450 179231 516484
rect 179265 516450 179323 516484
rect 179357 516450 179415 516484
rect 179449 516450 179507 516484
rect 179541 516450 179599 516484
rect 179633 516450 179691 516484
rect 179725 516450 179783 516484
rect 179817 516450 179875 516484
rect 179909 516450 179967 516484
rect 180001 516450 180059 516484
rect 180093 516450 180151 516484
rect 180185 516450 180243 516484
rect 180277 516450 180335 516484
rect 180369 516450 180427 516484
rect 180461 516450 180519 516484
rect 180553 516450 180611 516484
rect 180645 516450 180703 516484
rect 180737 516450 180795 516484
rect 180829 516450 180887 516484
rect 180921 516450 180979 516484
rect 181013 516450 181071 516484
rect 181105 516450 181163 516484
rect 181197 516450 181255 516484
rect 181289 516450 181347 516484
rect 181381 516450 181439 516484
rect 181473 516450 181531 516484
rect 181565 516450 181623 516484
rect 181657 516450 181715 516484
rect 181749 516450 181807 516484
rect 181841 516450 181899 516484
rect 181933 516450 181991 516484
rect 182025 516450 182083 516484
rect 182117 516450 182175 516484
rect 182209 516450 182261 516484
rect 178687 516441 178699 516450
rect 178751 516441 182261 516450
rect 182313 516441 182325 516493
rect 182377 516484 182389 516493
rect 182441 516484 182453 516493
rect 182441 516450 182451 516484
rect 182377 516441 182389 516450
rect 182441 516441 182453 516450
rect 182505 516441 182517 516493
rect 182569 516484 186079 516493
rect 182577 516450 182635 516484
rect 182669 516450 182727 516484
rect 182761 516450 182819 516484
rect 182853 516450 182911 516484
rect 182945 516450 183003 516484
rect 183037 516450 183095 516484
rect 183129 516450 183187 516484
rect 183221 516450 183279 516484
rect 183313 516450 183371 516484
rect 183405 516450 183463 516484
rect 183497 516450 183555 516484
rect 183589 516450 183647 516484
rect 183681 516450 183739 516484
rect 183773 516450 183831 516484
rect 183865 516450 183923 516484
rect 183957 516450 184015 516484
rect 184049 516450 184107 516484
rect 184141 516450 184199 516484
rect 184233 516450 184291 516484
rect 184325 516450 184383 516484
rect 184417 516450 184475 516484
rect 184509 516450 184567 516484
rect 184601 516450 184659 516484
rect 184693 516450 184751 516484
rect 184785 516450 184843 516484
rect 184877 516450 184935 516484
rect 184969 516450 185027 516484
rect 185061 516450 185119 516484
rect 185153 516450 185211 516484
rect 185245 516450 185303 516484
rect 185337 516450 185395 516484
rect 185429 516450 185487 516484
rect 185521 516450 185579 516484
rect 185613 516450 185671 516484
rect 185705 516450 185763 516484
rect 185797 516450 185855 516484
rect 185889 516450 185947 516484
rect 185981 516450 186039 516484
rect 186073 516450 186079 516484
rect 182569 516441 186079 516450
rect 186131 516484 186143 516493
rect 186131 516441 186143 516450
rect 186195 516441 186207 516493
rect 186259 516441 186271 516493
rect 186323 516484 186335 516493
rect 186387 516484 187482 516493
rect 186387 516450 186407 516484
rect 186441 516450 186499 516484
rect 186533 516450 186591 516484
rect 186625 516450 186683 516484
rect 186717 516450 186775 516484
rect 186809 516450 186867 516484
rect 186901 516450 186959 516484
rect 186993 516450 187051 516484
rect 187085 516450 187143 516484
rect 187177 516450 187235 516484
rect 187269 516450 187327 516484
rect 187361 516450 187419 516484
rect 187453 516450 187482 516484
rect 186323 516441 186335 516450
rect 186387 516441 187482 516450
rect 172210 516419 187482 516441
rect 172210 515949 187482 515971
rect 172210 515940 173965 515949
rect 174017 515940 174029 515949
rect 174081 515940 174093 515949
rect 172210 515906 172239 515940
rect 172273 515906 172331 515940
rect 172365 515906 172423 515940
rect 172457 515906 172515 515940
rect 172549 515906 172607 515940
rect 172641 515906 172699 515940
rect 172733 515906 172791 515940
rect 172825 515906 172883 515940
rect 172917 515906 172975 515940
rect 173009 515906 173067 515940
rect 173101 515906 173159 515940
rect 173193 515906 173251 515940
rect 173285 515906 173343 515940
rect 173377 515906 173435 515940
rect 173469 515906 173527 515940
rect 173561 515906 173619 515940
rect 173653 515906 173711 515940
rect 173745 515906 173803 515940
rect 173837 515906 173895 515940
rect 173929 515906 173965 515940
rect 174021 515906 174029 515940
rect 172210 515897 173965 515906
rect 174017 515897 174029 515906
rect 174081 515897 174093 515906
rect 174145 515897 174157 515949
rect 174209 515897 174221 515949
rect 174273 515940 177783 515949
rect 174297 515906 174355 515940
rect 174389 515906 174447 515940
rect 174481 515906 174539 515940
rect 174573 515906 174631 515940
rect 174665 515906 174723 515940
rect 174757 515906 174815 515940
rect 174849 515906 174907 515940
rect 174941 515906 174999 515940
rect 175033 515906 175091 515940
rect 175125 515906 175183 515940
rect 175217 515906 175275 515940
rect 175309 515906 175367 515940
rect 175401 515906 175459 515940
rect 175493 515906 175551 515940
rect 175585 515906 175643 515940
rect 175677 515906 175735 515940
rect 175769 515906 175827 515940
rect 175861 515906 175919 515940
rect 175953 515906 176011 515940
rect 176045 515906 176103 515940
rect 176137 515906 176195 515940
rect 176229 515906 176287 515940
rect 176321 515906 176379 515940
rect 176413 515906 176471 515940
rect 176505 515906 176563 515940
rect 176597 515906 176655 515940
rect 176689 515906 176747 515940
rect 176781 515906 176839 515940
rect 176873 515906 176931 515940
rect 176965 515906 177023 515940
rect 177057 515906 177115 515940
rect 177149 515906 177207 515940
rect 177241 515906 177299 515940
rect 177333 515906 177391 515940
rect 177425 515906 177483 515940
rect 177517 515906 177575 515940
rect 177609 515906 177667 515940
rect 177701 515906 177759 515940
rect 174273 515897 177783 515906
rect 177835 515897 177847 515949
rect 177899 515897 177911 515949
rect 177963 515940 177975 515949
rect 178027 515940 178039 515949
rect 178091 515940 181601 515949
rect 181653 515940 181665 515949
rect 181717 515940 181729 515949
rect 178027 515906 178035 515940
rect 178091 515906 178127 515940
rect 178161 515906 178219 515940
rect 178253 515906 178311 515940
rect 178345 515906 178403 515940
rect 178437 515906 178495 515940
rect 178529 515906 178587 515940
rect 178621 515906 178679 515940
rect 178713 515906 178771 515940
rect 178805 515906 178863 515940
rect 178897 515906 178955 515940
rect 178989 515906 179047 515940
rect 179081 515906 179139 515940
rect 179173 515906 179231 515940
rect 179265 515906 179323 515940
rect 179357 515906 179415 515940
rect 179449 515906 179507 515940
rect 179541 515906 179599 515940
rect 179633 515906 179691 515940
rect 179725 515906 179783 515940
rect 179817 515906 179875 515940
rect 179909 515906 179967 515940
rect 180001 515906 180059 515940
rect 180093 515906 180151 515940
rect 180185 515906 180243 515940
rect 180277 515906 180335 515940
rect 180369 515906 180427 515940
rect 180461 515906 180519 515940
rect 180553 515906 180611 515940
rect 180645 515906 180703 515940
rect 180737 515906 180795 515940
rect 180829 515906 180887 515940
rect 180921 515906 180979 515940
rect 181013 515906 181071 515940
rect 181105 515906 181163 515940
rect 181197 515906 181255 515940
rect 181289 515906 181347 515940
rect 181381 515906 181439 515940
rect 181473 515906 181531 515940
rect 181565 515906 181601 515940
rect 181657 515906 181665 515940
rect 177963 515897 177975 515906
rect 178027 515897 178039 515906
rect 178091 515897 181601 515906
rect 181653 515897 181665 515906
rect 181717 515897 181729 515906
rect 181781 515897 181793 515949
rect 181845 515897 181857 515949
rect 181909 515940 185419 515949
rect 181933 515906 181991 515940
rect 182025 515906 182083 515940
rect 182117 515906 182175 515940
rect 182209 515906 182267 515940
rect 182301 515906 182359 515940
rect 182393 515906 182451 515940
rect 182485 515906 182543 515940
rect 182577 515906 182635 515940
rect 182669 515906 182727 515940
rect 182761 515906 182819 515940
rect 182853 515906 182911 515940
rect 182945 515906 183003 515940
rect 183037 515906 183095 515940
rect 183129 515906 183187 515940
rect 183221 515906 183279 515940
rect 183313 515906 183371 515940
rect 183405 515906 183463 515940
rect 183497 515906 183555 515940
rect 183589 515906 183647 515940
rect 183681 515906 183739 515940
rect 183773 515906 183831 515940
rect 183865 515906 183923 515940
rect 183957 515906 184015 515940
rect 184049 515906 184107 515940
rect 184141 515906 184199 515940
rect 184233 515906 184291 515940
rect 184325 515906 184383 515940
rect 184417 515906 184475 515940
rect 184509 515906 184567 515940
rect 184601 515906 184659 515940
rect 184693 515906 184751 515940
rect 184785 515906 184843 515940
rect 184877 515906 184935 515940
rect 184969 515906 185027 515940
rect 185061 515906 185119 515940
rect 185153 515906 185211 515940
rect 185245 515906 185303 515940
rect 185337 515906 185395 515940
rect 181909 515897 185419 515906
rect 185471 515897 185483 515949
rect 185535 515897 185547 515949
rect 185599 515940 185611 515949
rect 185663 515940 185675 515949
rect 185727 515940 187482 515949
rect 185663 515906 185671 515940
rect 185727 515906 185763 515940
rect 185797 515906 185855 515940
rect 185889 515906 185947 515940
rect 185981 515906 186039 515940
rect 186073 515906 186131 515940
rect 186165 515906 186223 515940
rect 186257 515906 186315 515940
rect 186349 515906 186407 515940
rect 186441 515906 186499 515940
rect 186533 515906 186591 515940
rect 186625 515906 186683 515940
rect 186717 515906 186775 515940
rect 186809 515906 186867 515940
rect 186901 515906 186959 515940
rect 186993 515906 187051 515940
rect 187085 515906 187143 515940
rect 187177 515906 187235 515940
rect 187269 515906 187327 515940
rect 187361 515906 187419 515940
rect 187453 515906 187482 515940
rect 185599 515897 185611 515906
rect 185663 515897 185675 515906
rect 185727 515897 187482 515906
rect 172210 515875 187482 515897
rect 173604 515795 173610 515847
rect 173662 515795 173668 515847
rect 181332 515795 181338 515847
rect 181390 515835 181396 515847
rect 182071 515838 182129 515844
rect 182071 515835 182083 515838
rect 181390 515807 182083 515835
rect 181390 515795 181396 515807
rect 182071 515804 182083 515807
rect 182117 515804 182129 515838
rect 182071 515798 182129 515804
rect 186576 515795 186582 515847
rect 186634 515795 186640 515847
rect 182255 515634 182313 515640
rect 182255 515631 182267 515634
rect 182178 515603 182267 515631
rect 173328 515523 173334 515575
rect 173386 515563 173392 515575
rect 173515 515566 173573 515572
rect 173515 515563 173527 515566
rect 173386 515535 173527 515563
rect 173386 515523 173392 515535
rect 173515 515532 173527 515535
rect 173561 515532 173573 515566
rect 173515 515526 173573 515532
rect 182178 515507 182206 515603
rect 182255 515600 182267 515603
rect 182301 515600 182313 515634
rect 182255 515594 182313 515600
rect 186484 515523 186490 515575
rect 186542 515523 186548 515575
rect 182160 515455 182166 515507
rect 182218 515455 182224 515507
rect 172210 515405 187482 515427
rect 172210 515396 174625 515405
rect 172210 515362 172239 515396
rect 172273 515362 172331 515396
rect 172365 515362 172423 515396
rect 172457 515362 172515 515396
rect 172549 515362 172607 515396
rect 172641 515362 172699 515396
rect 172733 515362 172791 515396
rect 172825 515362 172883 515396
rect 172917 515362 172975 515396
rect 173009 515362 173067 515396
rect 173101 515362 173159 515396
rect 173193 515362 173251 515396
rect 173285 515362 173343 515396
rect 173377 515362 173435 515396
rect 173469 515362 173527 515396
rect 173561 515362 173619 515396
rect 173653 515362 173711 515396
rect 173745 515362 173803 515396
rect 173837 515362 173895 515396
rect 173929 515362 173987 515396
rect 174021 515362 174079 515396
rect 174113 515362 174171 515396
rect 174205 515362 174263 515396
rect 174297 515362 174355 515396
rect 174389 515362 174447 515396
rect 174481 515362 174539 515396
rect 174573 515362 174625 515396
rect 172210 515353 174625 515362
rect 174677 515353 174689 515405
rect 174741 515396 174753 515405
rect 174805 515396 174817 515405
rect 174805 515362 174815 515396
rect 174741 515353 174753 515362
rect 174805 515353 174817 515362
rect 174869 515353 174881 515405
rect 174933 515396 178443 515405
rect 174941 515362 174999 515396
rect 175033 515362 175091 515396
rect 175125 515362 175183 515396
rect 175217 515362 175275 515396
rect 175309 515362 175367 515396
rect 175401 515362 175459 515396
rect 175493 515362 175551 515396
rect 175585 515362 175643 515396
rect 175677 515362 175735 515396
rect 175769 515362 175827 515396
rect 175861 515362 175919 515396
rect 175953 515362 176011 515396
rect 176045 515362 176103 515396
rect 176137 515362 176195 515396
rect 176229 515362 176287 515396
rect 176321 515362 176379 515396
rect 176413 515362 176471 515396
rect 176505 515362 176563 515396
rect 176597 515362 176655 515396
rect 176689 515362 176747 515396
rect 176781 515362 176839 515396
rect 176873 515362 176931 515396
rect 176965 515362 177023 515396
rect 177057 515362 177115 515396
rect 177149 515362 177207 515396
rect 177241 515362 177299 515396
rect 177333 515362 177391 515396
rect 177425 515362 177483 515396
rect 177517 515362 177575 515396
rect 177609 515362 177667 515396
rect 177701 515362 177759 515396
rect 177793 515362 177851 515396
rect 177885 515362 177943 515396
rect 177977 515362 178035 515396
rect 178069 515362 178127 515396
rect 178161 515362 178219 515396
rect 178253 515362 178311 515396
rect 178345 515362 178403 515396
rect 178437 515362 178443 515396
rect 174933 515353 178443 515362
rect 178495 515396 178507 515405
rect 178495 515353 178507 515362
rect 178559 515353 178571 515405
rect 178623 515353 178635 515405
rect 178687 515396 178699 515405
rect 178751 515396 182261 515405
rect 178751 515362 178771 515396
rect 178805 515362 178863 515396
rect 178897 515362 178955 515396
rect 178989 515362 179047 515396
rect 179081 515362 179139 515396
rect 179173 515362 179231 515396
rect 179265 515362 179323 515396
rect 179357 515362 179415 515396
rect 179449 515362 179507 515396
rect 179541 515362 179599 515396
rect 179633 515362 179691 515396
rect 179725 515362 179783 515396
rect 179817 515362 179875 515396
rect 179909 515362 179967 515396
rect 180001 515362 180059 515396
rect 180093 515362 180151 515396
rect 180185 515362 180243 515396
rect 180277 515362 180335 515396
rect 180369 515362 180427 515396
rect 180461 515362 180519 515396
rect 180553 515362 180611 515396
rect 180645 515362 180703 515396
rect 180737 515362 180795 515396
rect 180829 515362 180887 515396
rect 180921 515362 180979 515396
rect 181013 515362 181071 515396
rect 181105 515362 181163 515396
rect 181197 515362 181255 515396
rect 181289 515362 181347 515396
rect 181381 515362 181439 515396
rect 181473 515362 181531 515396
rect 181565 515362 181623 515396
rect 181657 515362 181715 515396
rect 181749 515362 181807 515396
rect 181841 515362 181899 515396
rect 181933 515362 181991 515396
rect 182025 515362 182083 515396
rect 182117 515362 182175 515396
rect 182209 515362 182261 515396
rect 178687 515353 178699 515362
rect 178751 515353 182261 515362
rect 182313 515353 182325 515405
rect 182377 515396 182389 515405
rect 182441 515396 182453 515405
rect 182441 515362 182451 515396
rect 182377 515353 182389 515362
rect 182441 515353 182453 515362
rect 182505 515353 182517 515405
rect 182569 515396 186079 515405
rect 182577 515362 182635 515396
rect 182669 515362 182727 515396
rect 182761 515362 182819 515396
rect 182853 515362 182911 515396
rect 182945 515362 183003 515396
rect 183037 515362 183095 515396
rect 183129 515362 183187 515396
rect 183221 515362 183279 515396
rect 183313 515362 183371 515396
rect 183405 515362 183463 515396
rect 183497 515362 183555 515396
rect 183589 515362 183647 515396
rect 183681 515362 183739 515396
rect 183773 515362 183831 515396
rect 183865 515362 183923 515396
rect 183957 515362 184015 515396
rect 184049 515362 184107 515396
rect 184141 515362 184199 515396
rect 184233 515362 184291 515396
rect 184325 515362 184383 515396
rect 184417 515362 184475 515396
rect 184509 515362 184567 515396
rect 184601 515362 184659 515396
rect 184693 515362 184751 515396
rect 184785 515362 184843 515396
rect 184877 515362 184935 515396
rect 184969 515362 185027 515396
rect 185061 515362 185119 515396
rect 185153 515362 185211 515396
rect 185245 515362 185303 515396
rect 185337 515362 185395 515396
rect 185429 515362 185487 515396
rect 185521 515362 185579 515396
rect 185613 515362 185671 515396
rect 185705 515362 185763 515396
rect 185797 515362 185855 515396
rect 185889 515362 185947 515396
rect 185981 515362 186039 515396
rect 186073 515362 186079 515396
rect 182569 515353 186079 515362
rect 186131 515396 186143 515405
rect 186131 515353 186143 515362
rect 186195 515353 186207 515405
rect 186259 515353 186271 515405
rect 186323 515396 186335 515405
rect 186387 515396 187482 515405
rect 186387 515362 186407 515396
rect 186441 515362 186499 515396
rect 186533 515362 186591 515396
rect 186625 515362 186683 515396
rect 186717 515362 186775 515396
rect 186809 515362 186867 515396
rect 186901 515362 186959 515396
rect 186993 515362 187051 515396
rect 187085 515362 187143 515396
rect 187177 515362 187235 515396
rect 187269 515362 187327 515396
rect 187361 515362 187419 515396
rect 187453 515362 187482 515396
rect 186323 515353 186335 515362
rect 186387 515353 187482 515362
rect 172210 515331 187482 515353
rect 173000 512810 173250 513000
rect 173450 512810 175000 513000
rect 173000 509000 175000 512810
rect 1990 507000 2000 509000
rect 4000 507000 175000 509000
rect 177000 512810 177580 513000
rect 177780 512810 179000 513000
rect 177000 506000 179000 512810
rect 5000 504000 179000 506000
rect 181000 512810 181910 513000
rect 182110 512810 183000 513000
rect 5000 466000 7000 504000
rect 181000 503000 183000 512810
rect 1990 464000 2000 466000
rect 4000 464000 7000 466000
rect 8000 501000 183000 503000
rect 185000 512810 186230 513000
rect 186430 512810 187000 513000
rect 8000 423000 10000 501000
rect 185000 500000 187000 512810
rect 1990 421000 2000 423000
rect 4000 421000 10000 423000
rect 11000 498000 187000 500000
rect 11000 380000 13000 498000
rect 1990 378000 2000 380000
rect 4000 378000 13000 380000
<< rmetal1 >>
rect 192110 522947 192140 523037
<< via1 >>
rect 18000 699000 20000 701000
rect 70000 699000 72000 701000
rect 122000 699000 124000 701000
rect 3000 682000 5000 684000
rect 146000 626000 148000 628000
rect 154000 551000 156000 553000
rect 146000 544000 148000 546000
rect 154000 538000 156000 540000
rect 161390 538577 161510 538697
rect 163030 538697 163330 538897
rect 159400 538247 159480 538327
rect 165890 540927 165945 541027
rect 165945 540927 165979 541027
rect 165979 540927 166000 541027
rect 165890 540807 165945 540907
rect 165945 540807 165979 540907
rect 165979 540807 166000 540907
rect 165890 540687 165945 540787
rect 165945 540687 165979 540787
rect 165979 540687 166000 540787
rect 166690 540097 166870 540277
rect 161690 537738 161750 537767
rect 161690 537707 161700 537738
rect 161700 537707 161734 537738
rect 161734 537707 161750 537738
rect 162880 537917 162940 537977
rect 165900 538737 166040 538837
rect 166690 539157 166870 539337
rect 157420 536877 157510 536957
rect 161790 536857 161850 536937
rect 158480 536427 158580 536587
rect 161090 536497 161170 536577
rect 160200 535467 160350 535607
rect 163840 535937 164050 536267
rect 166930 536077 167260 536297
rect 166720 535457 166850 535587
rect 166900 535447 167030 535577
rect 167080 535427 167210 535557
rect 166700 535267 166830 535397
rect 166890 535257 167020 535387
rect 167090 535247 167220 535377
rect 169690 540927 169745 541027
rect 169745 540927 169779 541027
rect 169779 540927 169800 541027
rect 169690 540807 169745 540907
rect 169745 540807 169779 540907
rect 169779 540807 169800 540907
rect 169690 540687 169745 540787
rect 169745 540687 169779 540787
rect 169779 540687 169800 540787
rect 170490 540097 170670 540277
rect 169700 538737 169840 538837
rect 170490 539157 170670 539337
rect 169570 536007 169870 536287
rect 173390 540927 173445 541027
rect 173445 540927 173479 541027
rect 173479 540927 173500 541027
rect 173390 540807 173445 540907
rect 173445 540807 173479 540907
rect 173479 540807 173500 540907
rect 173390 540687 173445 540787
rect 173445 540687 173479 540787
rect 173479 540687 173500 540787
rect 174190 540107 174370 540287
rect 173400 538737 173540 538837
rect 174190 539157 174370 539337
rect 172610 536007 172940 536297
rect 176890 540927 176945 541027
rect 176945 540927 176979 541027
rect 176979 540927 177000 541027
rect 176890 540807 176945 540907
rect 176945 540807 176979 540907
rect 176979 540807 177000 540907
rect 176890 540687 176945 540787
rect 176945 540687 176979 540787
rect 176979 540687 177000 540787
rect 177700 540097 177880 540277
rect 176900 538737 177040 538837
rect 177690 539157 177870 539337
rect 175280 536051 175360 536287
rect 175360 536051 175398 536287
rect 175398 536051 175500 536287
rect 175280 535977 175500 536051
rect 172360 532597 172490 532767
rect 174490 532607 174620 532777
rect 176580 532597 176710 532767
rect 180490 540927 180545 541027
rect 180545 540927 180579 541027
rect 180579 540927 180600 541027
rect 180490 540807 180545 540907
rect 180545 540807 180579 540907
rect 180579 540807 180600 540907
rect 180490 540687 180545 540787
rect 180545 540687 180579 540787
rect 180579 540687 180600 540787
rect 181290 540097 181470 540277
rect 180500 538737 180640 538837
rect 181290 539157 181470 539337
rect 178870 535997 179070 536307
rect 183790 540927 183845 541027
rect 183845 540927 183879 541027
rect 183879 540927 183900 541027
rect 183790 540807 183845 540907
rect 183845 540807 183879 540907
rect 183879 540807 183900 540907
rect 183790 540687 183845 540787
rect 183845 540687 183879 540787
rect 183879 540687 183900 540787
rect 184590 540097 184770 540277
rect 183800 538737 183940 538837
rect 184590 539157 184770 539337
rect 182190 536057 182390 536317
rect 187090 540927 187145 541027
rect 187145 540927 187179 541027
rect 187179 540927 187200 541027
rect 187090 540807 187145 540907
rect 187145 540807 187179 540907
rect 187179 540807 187200 540907
rect 187090 540687 187145 540787
rect 187145 540687 187179 540787
rect 187179 540687 187200 540787
rect 187900 540097 188080 540277
rect 187100 538737 187240 538837
rect 187890 539157 188070 539337
rect 185490 536177 185700 536297
rect 178700 532597 178830 532767
rect 180870 532597 181000 532767
rect 190390 540927 190445 541027
rect 190445 540927 190479 541027
rect 190479 540927 190500 541027
rect 190390 540807 190445 540907
rect 190445 540807 190479 540907
rect 190479 540807 190500 540907
rect 190390 540687 190445 540787
rect 190445 540687 190479 540787
rect 190479 540687 190500 540787
rect 191190 540097 191370 540277
rect 190400 538737 190540 538837
rect 191200 539167 191380 539347
rect 188780 536067 189000 536307
rect 182960 532597 183090 532767
rect 185060 532637 185190 532807
rect 191810 540097 191990 540277
rect 191820 539157 192000 539337
rect 187170 532627 187270 532767
rect 174625 530628 174677 530637
rect 174625 530594 174631 530628
rect 174631 530594 174665 530628
rect 174665 530594 174677 530628
rect 174625 530585 174677 530594
rect 174689 530628 174741 530637
rect 174753 530628 174805 530637
rect 174817 530628 174869 530637
rect 174689 530594 174723 530628
rect 174723 530594 174741 530628
rect 174753 530594 174757 530628
rect 174757 530594 174805 530628
rect 174817 530594 174849 530628
rect 174849 530594 174869 530628
rect 174689 530585 174741 530594
rect 174753 530585 174805 530594
rect 174817 530585 174869 530594
rect 174881 530628 174933 530637
rect 174881 530594 174907 530628
rect 174907 530594 174933 530628
rect 174881 530585 174933 530594
rect 178443 530585 178495 530637
rect 178507 530628 178559 530637
rect 178507 530594 178529 530628
rect 178529 530594 178559 530628
rect 178507 530585 178559 530594
rect 178571 530628 178623 530637
rect 178571 530594 178587 530628
rect 178587 530594 178621 530628
rect 178621 530594 178623 530628
rect 178571 530585 178623 530594
rect 178635 530628 178687 530637
rect 178699 530628 178751 530637
rect 182261 530628 182313 530637
rect 178635 530594 178679 530628
rect 178679 530594 178687 530628
rect 178699 530594 178713 530628
rect 178713 530594 178751 530628
rect 182261 530594 182267 530628
rect 182267 530594 182301 530628
rect 182301 530594 182313 530628
rect 178635 530585 178687 530594
rect 178699 530585 178751 530594
rect 182261 530585 182313 530594
rect 182325 530628 182377 530637
rect 182389 530628 182441 530637
rect 182453 530628 182505 530637
rect 182325 530594 182359 530628
rect 182359 530594 182377 530628
rect 182389 530594 182393 530628
rect 182393 530594 182441 530628
rect 182453 530594 182485 530628
rect 182485 530594 182505 530628
rect 182325 530585 182377 530594
rect 182389 530585 182441 530594
rect 182453 530585 182505 530594
rect 182517 530628 182569 530637
rect 182517 530594 182543 530628
rect 182543 530594 182569 530628
rect 182517 530585 182569 530594
rect 186079 530585 186131 530637
rect 186143 530628 186195 530637
rect 186143 530594 186165 530628
rect 186165 530594 186195 530628
rect 186143 530585 186195 530594
rect 186207 530628 186259 530637
rect 186207 530594 186223 530628
rect 186223 530594 186257 530628
rect 186257 530594 186259 530628
rect 186207 530585 186259 530594
rect 186271 530628 186323 530637
rect 186335 530628 186387 530637
rect 186271 530594 186315 530628
rect 186315 530594 186323 530628
rect 186335 530594 186349 530628
rect 186349 530594 186387 530628
rect 186271 530585 186323 530594
rect 186335 530585 186387 530594
rect 172414 530415 172466 530467
rect 174530 530415 174582 530467
rect 176830 530483 176882 530535
rect 178762 530526 178814 530535
rect 178762 530492 178771 530526
rect 178771 530492 178805 530526
rect 178805 530492 178814 530526
rect 178762 530483 178814 530492
rect 174806 530347 174858 530399
rect 175450 530347 175502 530399
rect 176738 530415 176790 530467
rect 179498 530483 179550 530535
rect 182994 530483 183046 530535
rect 185110 530483 185162 530535
rect 178946 530347 178998 530399
rect 179222 530347 179274 530399
rect 176646 530279 176698 530331
rect 177290 530322 177342 530331
rect 177290 530288 177299 530322
rect 177299 530288 177333 530322
rect 177333 530288 177342 530322
rect 177290 530279 177342 530288
rect 178210 530322 178262 530331
rect 178210 530288 178219 530322
rect 178219 530288 178253 530322
rect 178253 530288 178262 530322
rect 178210 530279 178262 530288
rect 180694 530279 180746 530331
rect 182258 530347 182310 530399
rect 183178 530390 183230 530399
rect 183178 530356 183187 530390
rect 183187 530356 183221 530390
rect 183221 530356 183230 530390
rect 183178 530347 183230 530356
rect 187134 530390 187186 530399
rect 187134 530356 187143 530390
rect 187143 530356 187177 530390
rect 187177 530356 187186 530390
rect 187134 530347 187186 530356
rect 182626 530279 182678 530331
rect 177658 530186 177710 530195
rect 177658 530152 177667 530186
rect 177667 530152 177701 530186
rect 177701 530152 177710 530186
rect 177658 530143 177710 530152
rect 178302 530143 178354 530195
rect 179682 530143 179734 530195
rect 182166 530186 182218 530195
rect 182166 530152 182175 530186
rect 182175 530152 182209 530186
rect 182209 530152 182218 530186
rect 182166 530143 182218 530152
rect 182718 530143 182770 530195
rect 173965 530084 174017 530093
rect 174029 530084 174081 530093
rect 174093 530084 174145 530093
rect 173965 530050 173987 530084
rect 173987 530050 174017 530084
rect 174029 530050 174079 530084
rect 174079 530050 174081 530084
rect 174093 530050 174113 530084
rect 174113 530050 174145 530084
rect 173965 530041 174017 530050
rect 174029 530041 174081 530050
rect 174093 530041 174145 530050
rect 174157 530084 174209 530093
rect 174157 530050 174171 530084
rect 174171 530050 174205 530084
rect 174205 530050 174209 530084
rect 174157 530041 174209 530050
rect 174221 530084 174273 530093
rect 177783 530084 177835 530093
rect 174221 530050 174263 530084
rect 174263 530050 174273 530084
rect 177783 530050 177793 530084
rect 177793 530050 177835 530084
rect 174221 530041 174273 530050
rect 177783 530041 177835 530050
rect 177847 530084 177899 530093
rect 177847 530050 177851 530084
rect 177851 530050 177885 530084
rect 177885 530050 177899 530084
rect 177847 530041 177899 530050
rect 177911 530084 177963 530093
rect 177975 530084 178027 530093
rect 178039 530084 178091 530093
rect 181601 530084 181653 530093
rect 181665 530084 181717 530093
rect 181729 530084 181781 530093
rect 177911 530050 177943 530084
rect 177943 530050 177963 530084
rect 177975 530050 177977 530084
rect 177977 530050 178027 530084
rect 178039 530050 178069 530084
rect 178069 530050 178091 530084
rect 181601 530050 181623 530084
rect 181623 530050 181653 530084
rect 181665 530050 181715 530084
rect 181715 530050 181717 530084
rect 181729 530050 181749 530084
rect 181749 530050 181781 530084
rect 177911 530041 177963 530050
rect 177975 530041 178027 530050
rect 178039 530041 178091 530050
rect 181601 530041 181653 530050
rect 181665 530041 181717 530050
rect 181729 530041 181781 530050
rect 181793 530084 181845 530093
rect 181793 530050 181807 530084
rect 181807 530050 181841 530084
rect 181841 530050 181845 530084
rect 181793 530041 181845 530050
rect 181857 530084 181909 530093
rect 185419 530084 185471 530093
rect 181857 530050 181899 530084
rect 181899 530050 181909 530084
rect 185419 530050 185429 530084
rect 185429 530050 185471 530084
rect 181857 530041 181909 530050
rect 185419 530041 185471 530050
rect 185483 530084 185535 530093
rect 185483 530050 185487 530084
rect 185487 530050 185521 530084
rect 185521 530050 185535 530084
rect 185483 530041 185535 530050
rect 185547 530084 185599 530093
rect 185611 530084 185663 530093
rect 185675 530084 185727 530093
rect 185547 530050 185579 530084
rect 185579 530050 185599 530084
rect 185611 530050 185613 530084
rect 185613 530050 185663 530084
rect 185675 530050 185705 530084
rect 185705 530050 185727 530084
rect 185547 530041 185599 530050
rect 185611 530041 185663 530050
rect 185675 530041 185727 530050
rect 178210 529939 178262 529991
rect 179498 529939 179550 529991
rect 180878 529939 180930 529991
rect 182166 529939 182218 529991
rect 182626 529982 182678 529991
rect 182626 529948 182635 529982
rect 182635 529948 182669 529982
rect 182669 529948 182678 529982
rect 182626 529939 182678 529948
rect 178118 529871 178170 529923
rect 174806 529846 174858 529855
rect 174806 529812 174815 529846
rect 174815 529812 174849 529846
rect 174849 529812 174858 529846
rect 174806 529803 174858 529812
rect 176830 529735 176882 529787
rect 179314 529803 179366 529855
rect 179866 529846 179918 529855
rect 179866 529812 179875 529846
rect 179875 529812 179909 529846
rect 179909 529812 179918 529846
rect 179866 529803 179918 529812
rect 175358 529599 175410 529651
rect 176094 529599 176146 529651
rect 177382 529667 177434 529719
rect 177566 529667 177618 529719
rect 177658 529667 177710 529719
rect 177934 529599 177986 529651
rect 181522 529667 181574 529719
rect 183178 529846 183230 529855
rect 183178 529812 183187 529846
rect 183187 529812 183221 529846
rect 183221 529812 183230 529846
rect 183178 529803 183230 529812
rect 180510 529599 180562 529651
rect 181798 529599 181850 529651
rect 174625 529540 174677 529549
rect 174625 529506 174631 529540
rect 174631 529506 174665 529540
rect 174665 529506 174677 529540
rect 174625 529497 174677 529506
rect 174689 529540 174741 529549
rect 174753 529540 174805 529549
rect 174817 529540 174869 529549
rect 174689 529506 174723 529540
rect 174723 529506 174741 529540
rect 174753 529506 174757 529540
rect 174757 529506 174805 529540
rect 174817 529506 174849 529540
rect 174849 529506 174869 529540
rect 174689 529497 174741 529506
rect 174753 529497 174805 529506
rect 174817 529497 174869 529506
rect 174881 529540 174933 529549
rect 174881 529506 174907 529540
rect 174907 529506 174933 529540
rect 174881 529497 174933 529506
rect 178443 529497 178495 529549
rect 178507 529540 178559 529549
rect 178507 529506 178529 529540
rect 178529 529506 178559 529540
rect 178507 529497 178559 529506
rect 178571 529540 178623 529549
rect 178571 529506 178587 529540
rect 178587 529506 178621 529540
rect 178621 529506 178623 529540
rect 178571 529497 178623 529506
rect 178635 529540 178687 529549
rect 178699 529540 178751 529549
rect 182261 529540 182313 529549
rect 178635 529506 178679 529540
rect 178679 529506 178687 529540
rect 178699 529506 178713 529540
rect 178713 529506 178751 529540
rect 182261 529506 182267 529540
rect 182267 529506 182301 529540
rect 182301 529506 182313 529540
rect 178635 529497 178687 529506
rect 178699 529497 178751 529506
rect 182261 529497 182313 529506
rect 182325 529540 182377 529549
rect 182389 529540 182441 529549
rect 182453 529540 182505 529549
rect 182325 529506 182359 529540
rect 182359 529506 182377 529540
rect 182389 529506 182393 529540
rect 182393 529506 182441 529540
rect 182453 529506 182485 529540
rect 182485 529506 182505 529540
rect 182325 529497 182377 529506
rect 182389 529497 182441 529506
rect 182453 529497 182505 529506
rect 182517 529540 182569 529549
rect 182517 529506 182543 529540
rect 182543 529506 182569 529540
rect 182517 529497 182569 529506
rect 186079 529497 186131 529549
rect 186143 529540 186195 529549
rect 186143 529506 186165 529540
rect 186165 529506 186195 529540
rect 186143 529497 186195 529506
rect 186207 529540 186259 529549
rect 186207 529506 186223 529540
rect 186223 529506 186257 529540
rect 186257 529506 186259 529540
rect 186207 529497 186259 529506
rect 186271 529540 186323 529549
rect 186335 529540 186387 529549
rect 186271 529506 186315 529540
rect 186315 529506 186323 529540
rect 186335 529506 186349 529540
rect 186349 529506 186387 529540
rect 186271 529497 186323 529506
rect 186335 529497 186387 529506
rect 175358 529438 175410 529447
rect 175358 529404 175367 529438
rect 175367 529404 175401 529438
rect 175401 529404 175410 529438
rect 175358 529395 175410 529404
rect 177934 529395 177986 529447
rect 178302 529327 178354 529379
rect 179866 529438 179918 529447
rect 179866 529404 179875 529438
rect 179875 529404 179909 529438
rect 179909 529404 179918 529438
rect 179866 529395 179918 529404
rect 181798 529395 181850 529447
rect 175450 529302 175502 529311
rect 175450 529268 175459 529302
rect 175459 529268 175493 529302
rect 175493 529268 175502 529302
rect 175450 529259 175502 529268
rect 176738 529259 176790 529311
rect 177658 529302 177710 529311
rect 177658 529268 177667 529302
rect 177667 529268 177701 529302
rect 177701 529268 177710 529302
rect 177658 529259 177710 529268
rect 179682 529302 179734 529311
rect 179682 529268 179691 529302
rect 179691 529268 179725 529302
rect 179725 529268 179734 529302
rect 179682 529259 179734 529268
rect 173610 529191 173662 529243
rect 175266 529234 175318 529243
rect 175266 529200 175275 529234
rect 175275 529200 175309 529234
rect 175309 529200 175318 529234
rect 175266 529191 175318 529200
rect 175910 529055 175962 529107
rect 176094 529055 176146 529107
rect 177290 529191 177342 529243
rect 181522 529259 181574 529311
rect 182718 529302 182770 529311
rect 182718 529268 182727 529302
rect 182727 529268 182761 529302
rect 182761 529268 182770 529302
rect 182718 529259 182770 529268
rect 179314 529055 179366 529107
rect 179682 529055 179734 529107
rect 180510 529055 180562 529107
rect 173965 528996 174017 529005
rect 174029 528996 174081 529005
rect 174093 528996 174145 529005
rect 173965 528962 173987 528996
rect 173987 528962 174017 528996
rect 174029 528962 174079 528996
rect 174079 528962 174081 528996
rect 174093 528962 174113 528996
rect 174113 528962 174145 528996
rect 173965 528953 174017 528962
rect 174029 528953 174081 528962
rect 174093 528953 174145 528962
rect 174157 528996 174209 529005
rect 174157 528962 174171 528996
rect 174171 528962 174205 528996
rect 174205 528962 174209 528996
rect 174157 528953 174209 528962
rect 174221 528996 174273 529005
rect 177783 528996 177835 529005
rect 174221 528962 174263 528996
rect 174263 528962 174273 528996
rect 177783 528962 177793 528996
rect 177793 528962 177835 528996
rect 174221 528953 174273 528962
rect 177783 528953 177835 528962
rect 177847 528996 177899 529005
rect 177847 528962 177851 528996
rect 177851 528962 177885 528996
rect 177885 528962 177899 528996
rect 177847 528953 177899 528962
rect 177911 528996 177963 529005
rect 177975 528996 178027 529005
rect 178039 528996 178091 529005
rect 181601 528996 181653 529005
rect 181665 528996 181717 529005
rect 181729 528996 181781 529005
rect 177911 528962 177943 528996
rect 177943 528962 177963 528996
rect 177975 528962 177977 528996
rect 177977 528962 178027 528996
rect 178039 528962 178069 528996
rect 178069 528962 178091 528996
rect 181601 528962 181623 528996
rect 181623 528962 181653 528996
rect 181665 528962 181715 528996
rect 181715 528962 181717 528996
rect 181729 528962 181749 528996
rect 181749 528962 181781 528996
rect 177911 528953 177963 528962
rect 177975 528953 178027 528962
rect 178039 528953 178091 528962
rect 181601 528953 181653 528962
rect 181665 528953 181717 528962
rect 181729 528953 181781 528962
rect 181793 528996 181845 529005
rect 181793 528962 181807 528996
rect 181807 528962 181841 528996
rect 181841 528962 181845 528996
rect 181793 528953 181845 528962
rect 181857 528996 181909 529005
rect 185419 528996 185471 529005
rect 181857 528962 181899 528996
rect 181899 528962 181909 528996
rect 185419 528962 185429 528996
rect 185429 528962 185471 528996
rect 181857 528953 181909 528962
rect 185419 528953 185471 528962
rect 185483 528996 185535 529005
rect 185483 528962 185487 528996
rect 185487 528962 185521 528996
rect 185521 528962 185535 528996
rect 185483 528953 185535 528962
rect 185547 528996 185599 529005
rect 185611 528996 185663 529005
rect 185675 528996 185727 529005
rect 185547 528962 185579 528996
rect 185579 528962 185599 528996
rect 185611 528962 185613 528996
rect 185613 528962 185663 528996
rect 185675 528962 185705 528996
rect 185705 528962 185727 528996
rect 185547 528953 185599 528962
rect 185611 528953 185663 528962
rect 185675 528953 185727 528962
rect 175266 528851 175318 528903
rect 176646 528851 176698 528903
rect 177658 528851 177710 528903
rect 179682 528894 179734 528903
rect 179682 528860 179691 528894
rect 179691 528860 179725 528894
rect 179725 528860 179734 528894
rect 179682 528851 179734 528860
rect 177566 528715 177618 528767
rect 178026 528715 178078 528767
rect 178210 528715 178262 528767
rect 180510 528758 180562 528767
rect 180510 528724 180519 528758
rect 180519 528724 180553 528758
rect 180553 528724 180562 528758
rect 180510 528715 180562 528724
rect 182166 528851 182218 528903
rect 181522 528715 181574 528767
rect 175910 528690 175962 528699
rect 175910 528656 175919 528690
rect 175919 528656 175953 528690
rect 175953 528656 175962 528690
rect 175910 528647 175962 528656
rect 178394 528622 178446 528631
rect 178394 528588 178403 528622
rect 178403 528588 178437 528622
rect 178437 528588 178446 528622
rect 178394 528579 178446 528588
rect 186582 528579 186634 528631
rect 176278 528511 176330 528563
rect 176370 528554 176422 528563
rect 176370 528520 176379 528554
rect 176379 528520 176413 528554
rect 176413 528520 176422 528554
rect 176370 528511 176422 528520
rect 176738 528554 176790 528563
rect 176738 528520 176747 528554
rect 176747 528520 176781 528554
rect 176781 528520 176790 528554
rect 176738 528511 176790 528520
rect 177014 528511 177066 528563
rect 180970 528511 181022 528563
rect 174625 528452 174677 528461
rect 174625 528418 174631 528452
rect 174631 528418 174665 528452
rect 174665 528418 174677 528452
rect 174625 528409 174677 528418
rect 174689 528452 174741 528461
rect 174753 528452 174805 528461
rect 174817 528452 174869 528461
rect 174689 528418 174723 528452
rect 174723 528418 174741 528452
rect 174753 528418 174757 528452
rect 174757 528418 174805 528452
rect 174817 528418 174849 528452
rect 174849 528418 174869 528452
rect 174689 528409 174741 528418
rect 174753 528409 174805 528418
rect 174817 528409 174869 528418
rect 174881 528452 174933 528461
rect 174881 528418 174907 528452
rect 174907 528418 174933 528452
rect 174881 528409 174933 528418
rect 178443 528409 178495 528461
rect 178507 528452 178559 528461
rect 178507 528418 178529 528452
rect 178529 528418 178559 528452
rect 178507 528409 178559 528418
rect 178571 528452 178623 528461
rect 178571 528418 178587 528452
rect 178587 528418 178621 528452
rect 178621 528418 178623 528452
rect 178571 528409 178623 528418
rect 178635 528452 178687 528461
rect 178699 528452 178751 528461
rect 182261 528452 182313 528461
rect 178635 528418 178679 528452
rect 178679 528418 178687 528452
rect 178699 528418 178713 528452
rect 178713 528418 178751 528452
rect 182261 528418 182267 528452
rect 182267 528418 182301 528452
rect 182301 528418 182313 528452
rect 178635 528409 178687 528418
rect 178699 528409 178751 528418
rect 182261 528409 182313 528418
rect 182325 528452 182377 528461
rect 182389 528452 182441 528461
rect 182453 528452 182505 528461
rect 182325 528418 182359 528452
rect 182359 528418 182377 528452
rect 182389 528418 182393 528452
rect 182393 528418 182441 528452
rect 182453 528418 182485 528452
rect 182485 528418 182505 528452
rect 182325 528409 182377 528418
rect 182389 528409 182441 528418
rect 182453 528409 182505 528418
rect 182517 528452 182569 528461
rect 182517 528418 182543 528452
rect 182543 528418 182569 528452
rect 182517 528409 182569 528418
rect 186079 528409 186131 528461
rect 186143 528452 186195 528461
rect 186143 528418 186165 528452
rect 186165 528418 186195 528452
rect 186143 528409 186195 528418
rect 186207 528452 186259 528461
rect 186207 528418 186223 528452
rect 186223 528418 186257 528452
rect 186257 528418 186259 528452
rect 186207 528409 186259 528418
rect 186271 528452 186323 528461
rect 186335 528452 186387 528461
rect 186271 528418 186315 528452
rect 186315 528418 186323 528452
rect 186335 528418 186349 528452
rect 186349 528418 186387 528452
rect 186271 528409 186323 528418
rect 186335 528409 186387 528418
rect 176738 528307 176790 528359
rect 178026 528307 178078 528359
rect 178946 528350 178998 528359
rect 178946 528316 178955 528350
rect 178955 528316 178989 528350
rect 178989 528316 178998 528350
rect 178946 528307 178998 528316
rect 179314 528307 179366 528359
rect 180970 528350 181022 528359
rect 180970 528316 180979 528350
rect 180979 528316 181013 528350
rect 181013 528316 181022 528350
rect 180970 528307 181022 528316
rect 182166 528307 182218 528359
rect 176370 528282 176422 528291
rect 176370 528248 176379 528282
rect 176379 528248 176413 528282
rect 176413 528248 176422 528282
rect 176370 528239 176422 528248
rect 176830 528282 176882 528291
rect 176830 528248 176835 528282
rect 176835 528248 176869 528282
rect 176869 528248 176882 528282
rect 176830 528239 176882 528248
rect 176094 528214 176146 528223
rect 176094 528180 176103 528214
rect 176103 528180 176137 528214
rect 176137 528180 176146 528214
rect 176094 528171 176146 528180
rect 178118 528214 178170 528223
rect 178118 528180 178127 528214
rect 178127 528180 178161 528214
rect 178161 528180 178170 528214
rect 178118 528171 178170 528180
rect 177382 528035 177434 528087
rect 178946 527967 178998 528019
rect 181338 528214 181390 528223
rect 181338 528180 181347 528214
rect 181347 528180 181381 528214
rect 181381 528180 181390 528214
rect 181338 528171 181390 528180
rect 180694 528103 180746 528155
rect 173965 527908 174017 527917
rect 174029 527908 174081 527917
rect 174093 527908 174145 527917
rect 173965 527874 173987 527908
rect 173987 527874 174017 527908
rect 174029 527874 174079 527908
rect 174079 527874 174081 527908
rect 174093 527874 174113 527908
rect 174113 527874 174145 527908
rect 173965 527865 174017 527874
rect 174029 527865 174081 527874
rect 174093 527865 174145 527874
rect 174157 527908 174209 527917
rect 174157 527874 174171 527908
rect 174171 527874 174205 527908
rect 174205 527874 174209 527908
rect 174157 527865 174209 527874
rect 174221 527908 174273 527917
rect 177783 527908 177835 527917
rect 174221 527874 174263 527908
rect 174263 527874 174273 527908
rect 177783 527874 177793 527908
rect 177793 527874 177835 527908
rect 174221 527865 174273 527874
rect 177783 527865 177835 527874
rect 177847 527908 177899 527917
rect 177847 527874 177851 527908
rect 177851 527874 177885 527908
rect 177885 527874 177899 527908
rect 177847 527865 177899 527874
rect 177911 527908 177963 527917
rect 177975 527908 178027 527917
rect 178039 527908 178091 527917
rect 181601 527908 181653 527917
rect 181665 527908 181717 527917
rect 181729 527908 181781 527917
rect 177911 527874 177943 527908
rect 177943 527874 177963 527908
rect 177975 527874 177977 527908
rect 177977 527874 178027 527908
rect 178039 527874 178069 527908
rect 178069 527874 178091 527908
rect 181601 527874 181623 527908
rect 181623 527874 181653 527908
rect 181665 527874 181715 527908
rect 181715 527874 181717 527908
rect 181729 527874 181749 527908
rect 181749 527874 181781 527908
rect 177911 527865 177963 527874
rect 177975 527865 178027 527874
rect 178039 527865 178091 527874
rect 181601 527865 181653 527874
rect 181665 527865 181717 527874
rect 181729 527865 181781 527874
rect 181793 527908 181845 527917
rect 181793 527874 181807 527908
rect 181807 527874 181841 527908
rect 181841 527874 181845 527908
rect 181793 527865 181845 527874
rect 181857 527908 181909 527917
rect 185419 527908 185471 527917
rect 181857 527874 181899 527908
rect 181899 527874 181909 527908
rect 185419 527874 185429 527908
rect 185429 527874 185471 527908
rect 181857 527865 181909 527874
rect 185419 527865 185471 527874
rect 185483 527908 185535 527917
rect 185483 527874 185487 527908
rect 185487 527874 185521 527908
rect 185521 527874 185535 527908
rect 185483 527865 185535 527874
rect 185547 527908 185599 527917
rect 185611 527908 185663 527917
rect 185675 527908 185727 527917
rect 185547 527874 185579 527908
rect 185579 527874 185599 527908
rect 185611 527874 185613 527908
rect 185613 527874 185663 527908
rect 185675 527874 185705 527908
rect 185705 527874 185727 527908
rect 185547 527865 185599 527874
rect 185611 527865 185663 527874
rect 185675 527865 185727 527874
rect 176278 527763 176330 527815
rect 178946 527806 178998 527815
rect 178946 527772 178955 527806
rect 178955 527772 178989 527806
rect 178989 527772 178998 527806
rect 178946 527763 178998 527772
rect 177014 527670 177066 527679
rect 177014 527636 177023 527670
rect 177023 527636 177057 527670
rect 177057 527636 177066 527670
rect 177014 527627 177066 527636
rect 179498 527670 179550 527679
rect 179498 527636 179507 527670
rect 179507 527636 179541 527670
rect 179541 527636 179550 527670
rect 179498 527627 179550 527636
rect 174625 527364 174677 527373
rect 174625 527330 174631 527364
rect 174631 527330 174665 527364
rect 174665 527330 174677 527364
rect 174625 527321 174677 527330
rect 174689 527364 174741 527373
rect 174753 527364 174805 527373
rect 174817 527364 174869 527373
rect 174689 527330 174723 527364
rect 174723 527330 174741 527364
rect 174753 527330 174757 527364
rect 174757 527330 174805 527364
rect 174817 527330 174849 527364
rect 174849 527330 174869 527364
rect 174689 527321 174741 527330
rect 174753 527321 174805 527330
rect 174817 527321 174869 527330
rect 174881 527364 174933 527373
rect 174881 527330 174907 527364
rect 174907 527330 174933 527364
rect 174881 527321 174933 527330
rect 178443 527321 178495 527373
rect 178507 527364 178559 527373
rect 178507 527330 178529 527364
rect 178529 527330 178559 527364
rect 178507 527321 178559 527330
rect 178571 527364 178623 527373
rect 178571 527330 178587 527364
rect 178587 527330 178621 527364
rect 178621 527330 178623 527364
rect 178571 527321 178623 527330
rect 178635 527364 178687 527373
rect 178699 527364 178751 527373
rect 182261 527364 182313 527373
rect 178635 527330 178679 527364
rect 178679 527330 178687 527364
rect 178699 527330 178713 527364
rect 178713 527330 178751 527364
rect 182261 527330 182267 527364
rect 182267 527330 182301 527364
rect 182301 527330 182313 527364
rect 178635 527321 178687 527330
rect 178699 527321 178751 527330
rect 182261 527321 182313 527330
rect 182325 527364 182377 527373
rect 182389 527364 182441 527373
rect 182453 527364 182505 527373
rect 182325 527330 182359 527364
rect 182359 527330 182377 527364
rect 182389 527330 182393 527364
rect 182393 527330 182441 527364
rect 182453 527330 182485 527364
rect 182485 527330 182505 527364
rect 182325 527321 182377 527330
rect 182389 527321 182441 527330
rect 182453 527321 182505 527330
rect 182517 527364 182569 527373
rect 182517 527330 182543 527364
rect 182543 527330 182569 527364
rect 182517 527321 182569 527330
rect 186079 527321 186131 527373
rect 186143 527364 186195 527373
rect 186143 527330 186165 527364
rect 186165 527330 186195 527364
rect 186143 527321 186195 527330
rect 186207 527364 186259 527373
rect 186207 527330 186223 527364
rect 186223 527330 186257 527364
rect 186257 527330 186259 527364
rect 186207 527321 186259 527330
rect 186271 527364 186323 527373
rect 186335 527364 186387 527373
rect 186271 527330 186315 527364
rect 186315 527330 186323 527364
rect 186335 527330 186349 527364
rect 186349 527330 186387 527364
rect 186271 527321 186323 527330
rect 186335 527321 186387 527330
rect 173965 526820 174017 526829
rect 174029 526820 174081 526829
rect 174093 526820 174145 526829
rect 173965 526786 173987 526820
rect 173987 526786 174017 526820
rect 174029 526786 174079 526820
rect 174079 526786 174081 526820
rect 174093 526786 174113 526820
rect 174113 526786 174145 526820
rect 173965 526777 174017 526786
rect 174029 526777 174081 526786
rect 174093 526777 174145 526786
rect 174157 526820 174209 526829
rect 174157 526786 174171 526820
rect 174171 526786 174205 526820
rect 174205 526786 174209 526820
rect 174157 526777 174209 526786
rect 174221 526820 174273 526829
rect 177783 526820 177835 526829
rect 174221 526786 174263 526820
rect 174263 526786 174273 526820
rect 177783 526786 177793 526820
rect 177793 526786 177835 526820
rect 174221 526777 174273 526786
rect 177783 526777 177835 526786
rect 177847 526820 177899 526829
rect 177847 526786 177851 526820
rect 177851 526786 177885 526820
rect 177885 526786 177899 526820
rect 177847 526777 177899 526786
rect 177911 526820 177963 526829
rect 177975 526820 178027 526829
rect 178039 526820 178091 526829
rect 181601 526820 181653 526829
rect 181665 526820 181717 526829
rect 181729 526820 181781 526829
rect 177911 526786 177943 526820
rect 177943 526786 177963 526820
rect 177975 526786 177977 526820
rect 177977 526786 178027 526820
rect 178039 526786 178069 526820
rect 178069 526786 178091 526820
rect 181601 526786 181623 526820
rect 181623 526786 181653 526820
rect 181665 526786 181715 526820
rect 181715 526786 181717 526820
rect 181729 526786 181749 526820
rect 181749 526786 181781 526820
rect 177911 526777 177963 526786
rect 177975 526777 178027 526786
rect 178039 526777 178091 526786
rect 181601 526777 181653 526786
rect 181665 526777 181717 526786
rect 181729 526777 181781 526786
rect 181793 526820 181845 526829
rect 181793 526786 181807 526820
rect 181807 526786 181841 526820
rect 181841 526786 181845 526820
rect 181793 526777 181845 526786
rect 181857 526820 181909 526829
rect 185419 526820 185471 526829
rect 181857 526786 181899 526820
rect 181899 526786 181909 526820
rect 185419 526786 185429 526820
rect 185429 526786 185471 526820
rect 181857 526777 181909 526786
rect 185419 526777 185471 526786
rect 185483 526820 185535 526829
rect 185483 526786 185487 526820
rect 185487 526786 185521 526820
rect 185521 526786 185535 526820
rect 185483 526777 185535 526786
rect 185547 526820 185599 526829
rect 185611 526820 185663 526829
rect 185675 526820 185727 526829
rect 185547 526786 185579 526820
rect 185579 526786 185599 526820
rect 185611 526786 185613 526820
rect 185613 526786 185663 526820
rect 185675 526786 185705 526820
rect 185705 526786 185727 526820
rect 185547 526777 185599 526786
rect 185611 526777 185663 526786
rect 185675 526777 185727 526786
rect 174625 526276 174677 526285
rect 174625 526242 174631 526276
rect 174631 526242 174665 526276
rect 174665 526242 174677 526276
rect 174625 526233 174677 526242
rect 174689 526276 174741 526285
rect 174753 526276 174805 526285
rect 174817 526276 174869 526285
rect 174689 526242 174723 526276
rect 174723 526242 174741 526276
rect 174753 526242 174757 526276
rect 174757 526242 174805 526276
rect 174817 526242 174849 526276
rect 174849 526242 174869 526276
rect 174689 526233 174741 526242
rect 174753 526233 174805 526242
rect 174817 526233 174869 526242
rect 174881 526276 174933 526285
rect 174881 526242 174907 526276
rect 174907 526242 174933 526276
rect 174881 526233 174933 526242
rect 178443 526233 178495 526285
rect 178507 526276 178559 526285
rect 178507 526242 178529 526276
rect 178529 526242 178559 526276
rect 178507 526233 178559 526242
rect 178571 526276 178623 526285
rect 178571 526242 178587 526276
rect 178587 526242 178621 526276
rect 178621 526242 178623 526276
rect 178571 526233 178623 526242
rect 178635 526276 178687 526285
rect 178699 526276 178751 526285
rect 182261 526276 182313 526285
rect 178635 526242 178679 526276
rect 178679 526242 178687 526276
rect 178699 526242 178713 526276
rect 178713 526242 178751 526276
rect 182261 526242 182267 526276
rect 182267 526242 182301 526276
rect 182301 526242 182313 526276
rect 178635 526233 178687 526242
rect 178699 526233 178751 526242
rect 182261 526233 182313 526242
rect 182325 526276 182377 526285
rect 182389 526276 182441 526285
rect 182453 526276 182505 526285
rect 182325 526242 182359 526276
rect 182359 526242 182377 526276
rect 182389 526242 182393 526276
rect 182393 526242 182441 526276
rect 182453 526242 182485 526276
rect 182485 526242 182505 526276
rect 182325 526233 182377 526242
rect 182389 526233 182441 526242
rect 182453 526233 182505 526242
rect 182517 526276 182569 526285
rect 182517 526242 182543 526276
rect 182543 526242 182569 526276
rect 182517 526233 182569 526242
rect 186079 526233 186131 526285
rect 186143 526276 186195 526285
rect 186143 526242 186165 526276
rect 186165 526242 186195 526276
rect 186143 526233 186195 526242
rect 186207 526276 186259 526285
rect 186207 526242 186223 526276
rect 186223 526242 186257 526276
rect 186257 526242 186259 526276
rect 186207 526233 186259 526242
rect 186271 526276 186323 526285
rect 186335 526276 186387 526285
rect 186271 526242 186315 526276
rect 186315 526242 186323 526276
rect 186335 526242 186349 526276
rect 186349 526242 186387 526276
rect 186271 526233 186323 526242
rect 186335 526233 186387 526242
rect 173965 525732 174017 525741
rect 174029 525732 174081 525741
rect 174093 525732 174145 525741
rect 173965 525698 173987 525732
rect 173987 525698 174017 525732
rect 174029 525698 174079 525732
rect 174079 525698 174081 525732
rect 174093 525698 174113 525732
rect 174113 525698 174145 525732
rect 173965 525689 174017 525698
rect 174029 525689 174081 525698
rect 174093 525689 174145 525698
rect 174157 525732 174209 525741
rect 174157 525698 174171 525732
rect 174171 525698 174205 525732
rect 174205 525698 174209 525732
rect 174157 525689 174209 525698
rect 174221 525732 174273 525741
rect 177783 525732 177835 525741
rect 174221 525698 174263 525732
rect 174263 525698 174273 525732
rect 177783 525698 177793 525732
rect 177793 525698 177835 525732
rect 174221 525689 174273 525698
rect 177783 525689 177835 525698
rect 177847 525732 177899 525741
rect 177847 525698 177851 525732
rect 177851 525698 177885 525732
rect 177885 525698 177899 525732
rect 177847 525689 177899 525698
rect 177911 525732 177963 525741
rect 177975 525732 178027 525741
rect 178039 525732 178091 525741
rect 181601 525732 181653 525741
rect 181665 525732 181717 525741
rect 181729 525732 181781 525741
rect 177911 525698 177943 525732
rect 177943 525698 177963 525732
rect 177975 525698 177977 525732
rect 177977 525698 178027 525732
rect 178039 525698 178069 525732
rect 178069 525698 178091 525732
rect 181601 525698 181623 525732
rect 181623 525698 181653 525732
rect 181665 525698 181715 525732
rect 181715 525698 181717 525732
rect 181729 525698 181749 525732
rect 181749 525698 181781 525732
rect 177911 525689 177963 525698
rect 177975 525689 178027 525698
rect 178039 525689 178091 525698
rect 181601 525689 181653 525698
rect 181665 525689 181717 525698
rect 181729 525689 181781 525698
rect 181793 525732 181845 525741
rect 181793 525698 181807 525732
rect 181807 525698 181841 525732
rect 181841 525698 181845 525732
rect 181793 525689 181845 525698
rect 181857 525732 181909 525741
rect 185419 525732 185471 525741
rect 181857 525698 181899 525732
rect 181899 525698 181909 525732
rect 185419 525698 185429 525732
rect 185429 525698 185471 525732
rect 181857 525689 181909 525698
rect 185419 525689 185471 525698
rect 185483 525732 185535 525741
rect 185483 525698 185487 525732
rect 185487 525698 185521 525732
rect 185521 525698 185535 525732
rect 185483 525689 185535 525698
rect 185547 525732 185599 525741
rect 185611 525732 185663 525741
rect 185675 525732 185727 525741
rect 185547 525698 185579 525732
rect 185579 525698 185599 525732
rect 185611 525698 185613 525732
rect 185613 525698 185663 525732
rect 185675 525698 185705 525732
rect 185705 525698 185727 525732
rect 185547 525689 185599 525698
rect 185611 525689 185663 525698
rect 185675 525689 185727 525698
rect 174625 525188 174677 525197
rect 174625 525154 174631 525188
rect 174631 525154 174665 525188
rect 174665 525154 174677 525188
rect 174625 525145 174677 525154
rect 174689 525188 174741 525197
rect 174753 525188 174805 525197
rect 174817 525188 174869 525197
rect 174689 525154 174723 525188
rect 174723 525154 174741 525188
rect 174753 525154 174757 525188
rect 174757 525154 174805 525188
rect 174817 525154 174849 525188
rect 174849 525154 174869 525188
rect 174689 525145 174741 525154
rect 174753 525145 174805 525154
rect 174817 525145 174869 525154
rect 174881 525188 174933 525197
rect 174881 525154 174907 525188
rect 174907 525154 174933 525188
rect 174881 525145 174933 525154
rect 178443 525145 178495 525197
rect 178507 525188 178559 525197
rect 178507 525154 178529 525188
rect 178529 525154 178559 525188
rect 178507 525145 178559 525154
rect 178571 525188 178623 525197
rect 178571 525154 178587 525188
rect 178587 525154 178621 525188
rect 178621 525154 178623 525188
rect 178571 525145 178623 525154
rect 178635 525188 178687 525197
rect 178699 525188 178751 525197
rect 182261 525188 182313 525197
rect 178635 525154 178679 525188
rect 178679 525154 178687 525188
rect 178699 525154 178713 525188
rect 178713 525154 178751 525188
rect 182261 525154 182267 525188
rect 182267 525154 182301 525188
rect 182301 525154 182313 525188
rect 178635 525145 178687 525154
rect 178699 525145 178751 525154
rect 182261 525145 182313 525154
rect 182325 525188 182377 525197
rect 182389 525188 182441 525197
rect 182453 525188 182505 525197
rect 182325 525154 182359 525188
rect 182359 525154 182377 525188
rect 182389 525154 182393 525188
rect 182393 525154 182441 525188
rect 182453 525154 182485 525188
rect 182485 525154 182505 525188
rect 182325 525145 182377 525154
rect 182389 525145 182441 525154
rect 182453 525145 182505 525154
rect 182517 525188 182569 525197
rect 182517 525154 182543 525188
rect 182543 525154 182569 525188
rect 182517 525145 182569 525154
rect 186079 525145 186131 525197
rect 186143 525188 186195 525197
rect 186143 525154 186165 525188
rect 186165 525154 186195 525188
rect 186143 525145 186195 525154
rect 186207 525188 186259 525197
rect 186207 525154 186223 525188
rect 186223 525154 186257 525188
rect 186257 525154 186259 525188
rect 186207 525145 186259 525154
rect 186271 525188 186323 525197
rect 186335 525188 186387 525197
rect 186271 525154 186315 525188
rect 186315 525154 186323 525188
rect 186335 525154 186349 525188
rect 186349 525154 186387 525188
rect 186271 525145 186323 525154
rect 186335 525145 186387 525154
rect 173965 524644 174017 524653
rect 174029 524644 174081 524653
rect 174093 524644 174145 524653
rect 173965 524610 173987 524644
rect 173987 524610 174017 524644
rect 174029 524610 174079 524644
rect 174079 524610 174081 524644
rect 174093 524610 174113 524644
rect 174113 524610 174145 524644
rect 173965 524601 174017 524610
rect 174029 524601 174081 524610
rect 174093 524601 174145 524610
rect 174157 524644 174209 524653
rect 174157 524610 174171 524644
rect 174171 524610 174205 524644
rect 174205 524610 174209 524644
rect 174157 524601 174209 524610
rect 174221 524644 174273 524653
rect 177783 524644 177835 524653
rect 174221 524610 174263 524644
rect 174263 524610 174273 524644
rect 177783 524610 177793 524644
rect 177793 524610 177835 524644
rect 174221 524601 174273 524610
rect 177783 524601 177835 524610
rect 177847 524644 177899 524653
rect 177847 524610 177851 524644
rect 177851 524610 177885 524644
rect 177885 524610 177899 524644
rect 177847 524601 177899 524610
rect 177911 524644 177963 524653
rect 177975 524644 178027 524653
rect 178039 524644 178091 524653
rect 181601 524644 181653 524653
rect 181665 524644 181717 524653
rect 181729 524644 181781 524653
rect 177911 524610 177943 524644
rect 177943 524610 177963 524644
rect 177975 524610 177977 524644
rect 177977 524610 178027 524644
rect 178039 524610 178069 524644
rect 178069 524610 178091 524644
rect 181601 524610 181623 524644
rect 181623 524610 181653 524644
rect 181665 524610 181715 524644
rect 181715 524610 181717 524644
rect 181729 524610 181749 524644
rect 181749 524610 181781 524644
rect 177911 524601 177963 524610
rect 177975 524601 178027 524610
rect 178039 524601 178091 524610
rect 181601 524601 181653 524610
rect 181665 524601 181717 524610
rect 181729 524601 181781 524610
rect 181793 524644 181845 524653
rect 181793 524610 181807 524644
rect 181807 524610 181841 524644
rect 181841 524610 181845 524644
rect 181793 524601 181845 524610
rect 181857 524644 181909 524653
rect 185419 524644 185471 524653
rect 181857 524610 181899 524644
rect 181899 524610 181909 524644
rect 185419 524610 185429 524644
rect 185429 524610 185471 524644
rect 181857 524601 181909 524610
rect 185419 524601 185471 524610
rect 185483 524644 185535 524653
rect 185483 524610 185487 524644
rect 185487 524610 185521 524644
rect 185521 524610 185535 524644
rect 185483 524601 185535 524610
rect 185547 524644 185599 524653
rect 185611 524644 185663 524653
rect 185675 524644 185727 524653
rect 185547 524610 185579 524644
rect 185579 524610 185599 524644
rect 185611 524610 185613 524644
rect 185613 524610 185663 524644
rect 185675 524610 185705 524644
rect 185705 524610 185727 524644
rect 185547 524601 185599 524610
rect 185611 524601 185663 524610
rect 185675 524601 185727 524610
rect 174625 524100 174677 524109
rect 174625 524066 174631 524100
rect 174631 524066 174665 524100
rect 174665 524066 174677 524100
rect 174625 524057 174677 524066
rect 174689 524100 174741 524109
rect 174753 524100 174805 524109
rect 174817 524100 174869 524109
rect 174689 524066 174723 524100
rect 174723 524066 174741 524100
rect 174753 524066 174757 524100
rect 174757 524066 174805 524100
rect 174817 524066 174849 524100
rect 174849 524066 174869 524100
rect 174689 524057 174741 524066
rect 174753 524057 174805 524066
rect 174817 524057 174869 524066
rect 174881 524100 174933 524109
rect 174881 524066 174907 524100
rect 174907 524066 174933 524100
rect 174881 524057 174933 524066
rect 178443 524057 178495 524109
rect 178507 524100 178559 524109
rect 178507 524066 178529 524100
rect 178529 524066 178559 524100
rect 178507 524057 178559 524066
rect 178571 524100 178623 524109
rect 178571 524066 178587 524100
rect 178587 524066 178621 524100
rect 178621 524066 178623 524100
rect 178571 524057 178623 524066
rect 178635 524100 178687 524109
rect 178699 524100 178751 524109
rect 182261 524100 182313 524109
rect 178635 524066 178679 524100
rect 178679 524066 178687 524100
rect 178699 524066 178713 524100
rect 178713 524066 178751 524100
rect 182261 524066 182267 524100
rect 182267 524066 182301 524100
rect 182301 524066 182313 524100
rect 178635 524057 178687 524066
rect 178699 524057 178751 524066
rect 182261 524057 182313 524066
rect 182325 524100 182377 524109
rect 182389 524100 182441 524109
rect 182453 524100 182505 524109
rect 182325 524066 182359 524100
rect 182359 524066 182377 524100
rect 182389 524066 182393 524100
rect 182393 524066 182441 524100
rect 182453 524066 182485 524100
rect 182485 524066 182505 524100
rect 182325 524057 182377 524066
rect 182389 524057 182441 524066
rect 182453 524057 182505 524066
rect 182517 524100 182569 524109
rect 182517 524066 182543 524100
rect 182543 524066 182569 524100
rect 182517 524057 182569 524066
rect 186079 524057 186131 524109
rect 186143 524100 186195 524109
rect 186143 524066 186165 524100
rect 186165 524066 186195 524100
rect 186143 524057 186195 524066
rect 186207 524100 186259 524109
rect 186207 524066 186223 524100
rect 186223 524066 186257 524100
rect 186257 524066 186259 524100
rect 186207 524057 186259 524066
rect 186271 524100 186323 524109
rect 186335 524100 186387 524109
rect 186271 524066 186315 524100
rect 186315 524066 186323 524100
rect 186335 524066 186349 524100
rect 186349 524066 186387 524100
rect 186271 524057 186323 524066
rect 186335 524057 186387 524066
rect 173965 523556 174017 523565
rect 174029 523556 174081 523565
rect 174093 523556 174145 523565
rect 173965 523522 173987 523556
rect 173987 523522 174017 523556
rect 174029 523522 174079 523556
rect 174079 523522 174081 523556
rect 174093 523522 174113 523556
rect 174113 523522 174145 523556
rect 173965 523513 174017 523522
rect 174029 523513 174081 523522
rect 174093 523513 174145 523522
rect 174157 523556 174209 523565
rect 174157 523522 174171 523556
rect 174171 523522 174205 523556
rect 174205 523522 174209 523556
rect 174157 523513 174209 523522
rect 174221 523556 174273 523565
rect 177783 523556 177835 523565
rect 174221 523522 174263 523556
rect 174263 523522 174273 523556
rect 177783 523522 177793 523556
rect 177793 523522 177835 523556
rect 174221 523513 174273 523522
rect 177783 523513 177835 523522
rect 177847 523556 177899 523565
rect 177847 523522 177851 523556
rect 177851 523522 177885 523556
rect 177885 523522 177899 523556
rect 177847 523513 177899 523522
rect 177911 523556 177963 523565
rect 177975 523556 178027 523565
rect 178039 523556 178091 523565
rect 181601 523556 181653 523565
rect 181665 523556 181717 523565
rect 181729 523556 181781 523565
rect 177911 523522 177943 523556
rect 177943 523522 177963 523556
rect 177975 523522 177977 523556
rect 177977 523522 178027 523556
rect 178039 523522 178069 523556
rect 178069 523522 178091 523556
rect 181601 523522 181623 523556
rect 181623 523522 181653 523556
rect 181665 523522 181715 523556
rect 181715 523522 181717 523556
rect 181729 523522 181749 523556
rect 181749 523522 181781 523556
rect 177911 523513 177963 523522
rect 177975 523513 178027 523522
rect 178039 523513 178091 523522
rect 181601 523513 181653 523522
rect 181665 523513 181717 523522
rect 181729 523513 181781 523522
rect 181793 523556 181845 523565
rect 181793 523522 181807 523556
rect 181807 523522 181841 523556
rect 181841 523522 181845 523556
rect 181793 523513 181845 523522
rect 181857 523556 181909 523565
rect 185419 523556 185471 523565
rect 181857 523522 181899 523556
rect 181899 523522 181909 523556
rect 185419 523522 185429 523556
rect 185429 523522 185471 523556
rect 181857 523513 181909 523522
rect 185419 523513 185471 523522
rect 185483 523556 185535 523565
rect 185483 523522 185487 523556
rect 185487 523522 185521 523556
rect 185521 523522 185535 523556
rect 185483 523513 185535 523522
rect 185547 523556 185599 523565
rect 185611 523556 185663 523565
rect 185675 523556 185727 523565
rect 185547 523522 185579 523556
rect 185579 523522 185599 523556
rect 185611 523522 185613 523556
rect 185613 523522 185663 523556
rect 185675 523522 185705 523556
rect 185705 523522 185727 523556
rect 185547 523513 185599 523522
rect 185611 523513 185663 523522
rect 185675 523513 185727 523522
rect 174625 523012 174677 523021
rect 174625 522978 174631 523012
rect 174631 522978 174665 523012
rect 174665 522978 174677 523012
rect 174625 522969 174677 522978
rect 174689 523012 174741 523021
rect 174753 523012 174805 523021
rect 174817 523012 174869 523021
rect 174689 522978 174723 523012
rect 174723 522978 174741 523012
rect 174753 522978 174757 523012
rect 174757 522978 174805 523012
rect 174817 522978 174849 523012
rect 174849 522978 174869 523012
rect 174689 522969 174741 522978
rect 174753 522969 174805 522978
rect 174817 522969 174869 522978
rect 174881 523012 174933 523021
rect 174881 522978 174907 523012
rect 174907 522978 174933 523012
rect 174881 522969 174933 522978
rect 178443 522969 178495 523021
rect 178507 523012 178559 523021
rect 178507 522978 178529 523012
rect 178529 522978 178559 523012
rect 178507 522969 178559 522978
rect 178571 523012 178623 523021
rect 178571 522978 178587 523012
rect 178587 522978 178621 523012
rect 178621 522978 178623 523012
rect 178571 522969 178623 522978
rect 178635 523012 178687 523021
rect 178699 523012 178751 523021
rect 182261 523012 182313 523021
rect 178635 522978 178679 523012
rect 178679 522978 178687 523012
rect 178699 522978 178713 523012
rect 178713 522978 178751 523012
rect 182261 522978 182267 523012
rect 182267 522978 182301 523012
rect 182301 522978 182313 523012
rect 178635 522969 178687 522978
rect 178699 522969 178751 522978
rect 182261 522969 182313 522978
rect 182325 523012 182377 523021
rect 182389 523012 182441 523021
rect 182453 523012 182505 523021
rect 182325 522978 182359 523012
rect 182359 522978 182377 523012
rect 182389 522978 182393 523012
rect 182393 522978 182441 523012
rect 182453 522978 182485 523012
rect 182485 522978 182505 523012
rect 182325 522969 182377 522978
rect 182389 522969 182441 522978
rect 182453 522969 182505 522978
rect 182517 523012 182569 523021
rect 182517 522978 182543 523012
rect 182543 522978 182569 523012
rect 182517 522969 182569 522978
rect 186079 522969 186131 523021
rect 186143 523012 186195 523021
rect 186143 522978 186165 523012
rect 186165 522978 186195 523012
rect 186143 522969 186195 522978
rect 186207 523012 186259 523021
rect 186207 522978 186223 523012
rect 186223 522978 186257 523012
rect 186257 522978 186259 523012
rect 186207 522969 186259 522978
rect 186271 523012 186323 523021
rect 186335 523012 186387 523021
rect 186271 522978 186315 523012
rect 186315 522978 186323 523012
rect 186335 522978 186349 523012
rect 186349 522978 186387 523012
rect 186271 522969 186323 522978
rect 186335 522969 186387 522978
rect 173965 522468 174017 522477
rect 174029 522468 174081 522477
rect 174093 522468 174145 522477
rect 173965 522434 173987 522468
rect 173987 522434 174017 522468
rect 174029 522434 174079 522468
rect 174079 522434 174081 522468
rect 174093 522434 174113 522468
rect 174113 522434 174145 522468
rect 173965 522425 174017 522434
rect 174029 522425 174081 522434
rect 174093 522425 174145 522434
rect 174157 522468 174209 522477
rect 174157 522434 174171 522468
rect 174171 522434 174205 522468
rect 174205 522434 174209 522468
rect 174157 522425 174209 522434
rect 174221 522468 174273 522477
rect 177783 522468 177835 522477
rect 174221 522434 174263 522468
rect 174263 522434 174273 522468
rect 177783 522434 177793 522468
rect 177793 522434 177835 522468
rect 174221 522425 174273 522434
rect 177783 522425 177835 522434
rect 177847 522468 177899 522477
rect 177847 522434 177851 522468
rect 177851 522434 177885 522468
rect 177885 522434 177899 522468
rect 177847 522425 177899 522434
rect 177911 522468 177963 522477
rect 177975 522468 178027 522477
rect 178039 522468 178091 522477
rect 181601 522468 181653 522477
rect 181665 522468 181717 522477
rect 181729 522468 181781 522477
rect 177911 522434 177943 522468
rect 177943 522434 177963 522468
rect 177975 522434 177977 522468
rect 177977 522434 178027 522468
rect 178039 522434 178069 522468
rect 178069 522434 178091 522468
rect 181601 522434 181623 522468
rect 181623 522434 181653 522468
rect 181665 522434 181715 522468
rect 181715 522434 181717 522468
rect 181729 522434 181749 522468
rect 181749 522434 181781 522468
rect 177911 522425 177963 522434
rect 177975 522425 178027 522434
rect 178039 522425 178091 522434
rect 181601 522425 181653 522434
rect 181665 522425 181717 522434
rect 181729 522425 181781 522434
rect 181793 522468 181845 522477
rect 181793 522434 181807 522468
rect 181807 522434 181841 522468
rect 181841 522434 181845 522468
rect 181793 522425 181845 522434
rect 181857 522468 181909 522477
rect 185419 522468 185471 522477
rect 181857 522434 181899 522468
rect 181899 522434 181909 522468
rect 185419 522434 185429 522468
rect 185429 522434 185471 522468
rect 181857 522425 181909 522434
rect 185419 522425 185471 522434
rect 185483 522468 185535 522477
rect 185483 522434 185487 522468
rect 185487 522434 185521 522468
rect 185521 522434 185535 522468
rect 185483 522425 185535 522434
rect 185547 522468 185599 522477
rect 185611 522468 185663 522477
rect 185675 522468 185727 522477
rect 185547 522434 185579 522468
rect 185579 522434 185599 522468
rect 185611 522434 185613 522468
rect 185613 522434 185663 522468
rect 185675 522434 185705 522468
rect 185705 522434 185727 522468
rect 185547 522425 185599 522434
rect 185611 522425 185663 522434
rect 185675 522425 185727 522434
rect 174625 521924 174677 521933
rect 174625 521890 174631 521924
rect 174631 521890 174665 521924
rect 174665 521890 174677 521924
rect 174625 521881 174677 521890
rect 174689 521924 174741 521933
rect 174753 521924 174805 521933
rect 174817 521924 174869 521933
rect 174689 521890 174723 521924
rect 174723 521890 174741 521924
rect 174753 521890 174757 521924
rect 174757 521890 174805 521924
rect 174817 521890 174849 521924
rect 174849 521890 174869 521924
rect 174689 521881 174741 521890
rect 174753 521881 174805 521890
rect 174817 521881 174869 521890
rect 174881 521924 174933 521933
rect 174881 521890 174907 521924
rect 174907 521890 174933 521924
rect 174881 521881 174933 521890
rect 178443 521881 178495 521933
rect 178507 521924 178559 521933
rect 178507 521890 178529 521924
rect 178529 521890 178559 521924
rect 178507 521881 178559 521890
rect 178571 521924 178623 521933
rect 178571 521890 178587 521924
rect 178587 521890 178621 521924
rect 178621 521890 178623 521924
rect 178571 521881 178623 521890
rect 178635 521924 178687 521933
rect 178699 521924 178751 521933
rect 182261 521924 182313 521933
rect 178635 521890 178679 521924
rect 178679 521890 178687 521924
rect 178699 521890 178713 521924
rect 178713 521890 178751 521924
rect 182261 521890 182267 521924
rect 182267 521890 182301 521924
rect 182301 521890 182313 521924
rect 178635 521881 178687 521890
rect 178699 521881 178751 521890
rect 182261 521881 182313 521890
rect 182325 521924 182377 521933
rect 182389 521924 182441 521933
rect 182453 521924 182505 521933
rect 182325 521890 182359 521924
rect 182359 521890 182377 521924
rect 182389 521890 182393 521924
rect 182393 521890 182441 521924
rect 182453 521890 182485 521924
rect 182485 521890 182505 521924
rect 182325 521881 182377 521890
rect 182389 521881 182441 521890
rect 182453 521881 182505 521890
rect 182517 521924 182569 521933
rect 182517 521890 182543 521924
rect 182543 521890 182569 521924
rect 182517 521881 182569 521890
rect 186079 521881 186131 521933
rect 186143 521924 186195 521933
rect 186143 521890 186165 521924
rect 186165 521890 186195 521924
rect 186143 521881 186195 521890
rect 186207 521924 186259 521933
rect 186207 521890 186223 521924
rect 186223 521890 186257 521924
rect 186257 521890 186259 521924
rect 186207 521881 186259 521890
rect 186271 521924 186323 521933
rect 186335 521924 186387 521933
rect 186271 521890 186315 521924
rect 186315 521890 186323 521924
rect 186335 521890 186349 521924
rect 186349 521890 186387 521924
rect 186271 521881 186323 521890
rect 186335 521881 186387 521890
rect 173965 521380 174017 521389
rect 174029 521380 174081 521389
rect 174093 521380 174145 521389
rect 173965 521346 173987 521380
rect 173987 521346 174017 521380
rect 174029 521346 174079 521380
rect 174079 521346 174081 521380
rect 174093 521346 174113 521380
rect 174113 521346 174145 521380
rect 173965 521337 174017 521346
rect 174029 521337 174081 521346
rect 174093 521337 174145 521346
rect 174157 521380 174209 521389
rect 174157 521346 174171 521380
rect 174171 521346 174205 521380
rect 174205 521346 174209 521380
rect 174157 521337 174209 521346
rect 174221 521380 174273 521389
rect 177783 521380 177835 521389
rect 174221 521346 174263 521380
rect 174263 521346 174273 521380
rect 177783 521346 177793 521380
rect 177793 521346 177835 521380
rect 174221 521337 174273 521346
rect 177783 521337 177835 521346
rect 177847 521380 177899 521389
rect 177847 521346 177851 521380
rect 177851 521346 177885 521380
rect 177885 521346 177899 521380
rect 177847 521337 177899 521346
rect 177911 521380 177963 521389
rect 177975 521380 178027 521389
rect 178039 521380 178091 521389
rect 181601 521380 181653 521389
rect 181665 521380 181717 521389
rect 181729 521380 181781 521389
rect 177911 521346 177943 521380
rect 177943 521346 177963 521380
rect 177975 521346 177977 521380
rect 177977 521346 178027 521380
rect 178039 521346 178069 521380
rect 178069 521346 178091 521380
rect 181601 521346 181623 521380
rect 181623 521346 181653 521380
rect 181665 521346 181715 521380
rect 181715 521346 181717 521380
rect 181729 521346 181749 521380
rect 181749 521346 181781 521380
rect 177911 521337 177963 521346
rect 177975 521337 178027 521346
rect 178039 521337 178091 521346
rect 181601 521337 181653 521346
rect 181665 521337 181717 521346
rect 181729 521337 181781 521346
rect 181793 521380 181845 521389
rect 181793 521346 181807 521380
rect 181807 521346 181841 521380
rect 181841 521346 181845 521380
rect 181793 521337 181845 521346
rect 181857 521380 181909 521389
rect 185419 521380 185471 521389
rect 181857 521346 181899 521380
rect 181899 521346 181909 521380
rect 185419 521346 185429 521380
rect 185429 521346 185471 521380
rect 181857 521337 181909 521346
rect 185419 521337 185471 521346
rect 185483 521380 185535 521389
rect 185483 521346 185487 521380
rect 185487 521346 185521 521380
rect 185521 521346 185535 521380
rect 185483 521337 185535 521346
rect 185547 521380 185599 521389
rect 185611 521380 185663 521389
rect 185675 521380 185727 521389
rect 185547 521346 185579 521380
rect 185579 521346 185599 521380
rect 185611 521346 185613 521380
rect 185613 521346 185663 521380
rect 185675 521346 185705 521380
rect 185705 521346 185727 521380
rect 185547 521337 185599 521346
rect 185611 521337 185663 521346
rect 185675 521337 185727 521346
rect 174625 520836 174677 520845
rect 174625 520802 174631 520836
rect 174631 520802 174665 520836
rect 174665 520802 174677 520836
rect 174625 520793 174677 520802
rect 174689 520836 174741 520845
rect 174753 520836 174805 520845
rect 174817 520836 174869 520845
rect 174689 520802 174723 520836
rect 174723 520802 174741 520836
rect 174753 520802 174757 520836
rect 174757 520802 174805 520836
rect 174817 520802 174849 520836
rect 174849 520802 174869 520836
rect 174689 520793 174741 520802
rect 174753 520793 174805 520802
rect 174817 520793 174869 520802
rect 174881 520836 174933 520845
rect 174881 520802 174907 520836
rect 174907 520802 174933 520836
rect 174881 520793 174933 520802
rect 178443 520793 178495 520845
rect 178507 520836 178559 520845
rect 178507 520802 178529 520836
rect 178529 520802 178559 520836
rect 178507 520793 178559 520802
rect 178571 520836 178623 520845
rect 178571 520802 178587 520836
rect 178587 520802 178621 520836
rect 178621 520802 178623 520836
rect 178571 520793 178623 520802
rect 178635 520836 178687 520845
rect 178699 520836 178751 520845
rect 182261 520836 182313 520845
rect 178635 520802 178679 520836
rect 178679 520802 178687 520836
rect 178699 520802 178713 520836
rect 178713 520802 178751 520836
rect 182261 520802 182267 520836
rect 182267 520802 182301 520836
rect 182301 520802 182313 520836
rect 178635 520793 178687 520802
rect 178699 520793 178751 520802
rect 182261 520793 182313 520802
rect 182325 520836 182377 520845
rect 182389 520836 182441 520845
rect 182453 520836 182505 520845
rect 182325 520802 182359 520836
rect 182359 520802 182377 520836
rect 182389 520802 182393 520836
rect 182393 520802 182441 520836
rect 182453 520802 182485 520836
rect 182485 520802 182505 520836
rect 182325 520793 182377 520802
rect 182389 520793 182441 520802
rect 182453 520793 182505 520802
rect 182517 520836 182569 520845
rect 182517 520802 182543 520836
rect 182543 520802 182569 520836
rect 182517 520793 182569 520802
rect 186079 520793 186131 520845
rect 186143 520836 186195 520845
rect 186143 520802 186165 520836
rect 186165 520802 186195 520836
rect 186143 520793 186195 520802
rect 186207 520836 186259 520845
rect 186207 520802 186223 520836
rect 186223 520802 186257 520836
rect 186257 520802 186259 520836
rect 186207 520793 186259 520802
rect 186271 520836 186323 520845
rect 186335 520836 186387 520845
rect 186271 520802 186315 520836
rect 186315 520802 186323 520836
rect 186335 520802 186349 520836
rect 186349 520802 186387 520836
rect 186271 520793 186323 520802
rect 186335 520793 186387 520802
rect 173965 520292 174017 520301
rect 174029 520292 174081 520301
rect 174093 520292 174145 520301
rect 173965 520258 173987 520292
rect 173987 520258 174017 520292
rect 174029 520258 174079 520292
rect 174079 520258 174081 520292
rect 174093 520258 174113 520292
rect 174113 520258 174145 520292
rect 173965 520249 174017 520258
rect 174029 520249 174081 520258
rect 174093 520249 174145 520258
rect 174157 520292 174209 520301
rect 174157 520258 174171 520292
rect 174171 520258 174205 520292
rect 174205 520258 174209 520292
rect 174157 520249 174209 520258
rect 174221 520292 174273 520301
rect 177783 520292 177835 520301
rect 174221 520258 174263 520292
rect 174263 520258 174273 520292
rect 177783 520258 177793 520292
rect 177793 520258 177835 520292
rect 174221 520249 174273 520258
rect 177783 520249 177835 520258
rect 177847 520292 177899 520301
rect 177847 520258 177851 520292
rect 177851 520258 177885 520292
rect 177885 520258 177899 520292
rect 177847 520249 177899 520258
rect 177911 520292 177963 520301
rect 177975 520292 178027 520301
rect 178039 520292 178091 520301
rect 181601 520292 181653 520301
rect 181665 520292 181717 520301
rect 181729 520292 181781 520301
rect 177911 520258 177943 520292
rect 177943 520258 177963 520292
rect 177975 520258 177977 520292
rect 177977 520258 178027 520292
rect 178039 520258 178069 520292
rect 178069 520258 178091 520292
rect 181601 520258 181623 520292
rect 181623 520258 181653 520292
rect 181665 520258 181715 520292
rect 181715 520258 181717 520292
rect 181729 520258 181749 520292
rect 181749 520258 181781 520292
rect 177911 520249 177963 520258
rect 177975 520249 178027 520258
rect 178039 520249 178091 520258
rect 181601 520249 181653 520258
rect 181665 520249 181717 520258
rect 181729 520249 181781 520258
rect 181793 520292 181845 520301
rect 181793 520258 181807 520292
rect 181807 520258 181841 520292
rect 181841 520258 181845 520292
rect 181793 520249 181845 520258
rect 181857 520292 181909 520301
rect 185419 520292 185471 520301
rect 181857 520258 181899 520292
rect 181899 520258 181909 520292
rect 185419 520258 185429 520292
rect 185429 520258 185471 520292
rect 181857 520249 181909 520258
rect 185419 520249 185471 520258
rect 185483 520292 185535 520301
rect 185483 520258 185487 520292
rect 185487 520258 185521 520292
rect 185521 520258 185535 520292
rect 185483 520249 185535 520258
rect 185547 520292 185599 520301
rect 185611 520292 185663 520301
rect 185675 520292 185727 520301
rect 185547 520258 185579 520292
rect 185579 520258 185599 520292
rect 185611 520258 185613 520292
rect 185613 520258 185663 520292
rect 185675 520258 185705 520292
rect 185705 520258 185727 520292
rect 185547 520249 185599 520258
rect 185611 520249 185663 520258
rect 185675 520249 185727 520258
rect 174625 519748 174677 519757
rect 174625 519714 174631 519748
rect 174631 519714 174665 519748
rect 174665 519714 174677 519748
rect 174625 519705 174677 519714
rect 174689 519748 174741 519757
rect 174753 519748 174805 519757
rect 174817 519748 174869 519757
rect 174689 519714 174723 519748
rect 174723 519714 174741 519748
rect 174753 519714 174757 519748
rect 174757 519714 174805 519748
rect 174817 519714 174849 519748
rect 174849 519714 174869 519748
rect 174689 519705 174741 519714
rect 174753 519705 174805 519714
rect 174817 519705 174869 519714
rect 174881 519748 174933 519757
rect 174881 519714 174907 519748
rect 174907 519714 174933 519748
rect 174881 519705 174933 519714
rect 178443 519705 178495 519757
rect 178507 519748 178559 519757
rect 178507 519714 178529 519748
rect 178529 519714 178559 519748
rect 178507 519705 178559 519714
rect 178571 519748 178623 519757
rect 178571 519714 178587 519748
rect 178587 519714 178621 519748
rect 178621 519714 178623 519748
rect 178571 519705 178623 519714
rect 178635 519748 178687 519757
rect 178699 519748 178751 519757
rect 182261 519748 182313 519757
rect 178635 519714 178679 519748
rect 178679 519714 178687 519748
rect 178699 519714 178713 519748
rect 178713 519714 178751 519748
rect 182261 519714 182267 519748
rect 182267 519714 182301 519748
rect 182301 519714 182313 519748
rect 178635 519705 178687 519714
rect 178699 519705 178751 519714
rect 182261 519705 182313 519714
rect 182325 519748 182377 519757
rect 182389 519748 182441 519757
rect 182453 519748 182505 519757
rect 182325 519714 182359 519748
rect 182359 519714 182377 519748
rect 182389 519714 182393 519748
rect 182393 519714 182441 519748
rect 182453 519714 182485 519748
rect 182485 519714 182505 519748
rect 182325 519705 182377 519714
rect 182389 519705 182441 519714
rect 182453 519705 182505 519714
rect 182517 519748 182569 519757
rect 182517 519714 182543 519748
rect 182543 519714 182569 519748
rect 182517 519705 182569 519714
rect 186079 519705 186131 519757
rect 186143 519748 186195 519757
rect 186143 519714 186165 519748
rect 186165 519714 186195 519748
rect 186143 519705 186195 519714
rect 186207 519748 186259 519757
rect 186207 519714 186223 519748
rect 186223 519714 186257 519748
rect 186257 519714 186259 519748
rect 186207 519705 186259 519714
rect 186271 519748 186323 519757
rect 186335 519748 186387 519757
rect 186271 519714 186315 519748
rect 186315 519714 186323 519748
rect 186335 519714 186349 519748
rect 186349 519714 186387 519748
rect 186271 519705 186323 519714
rect 186335 519705 186387 519714
rect 173965 519204 174017 519213
rect 174029 519204 174081 519213
rect 174093 519204 174145 519213
rect 173965 519170 173987 519204
rect 173987 519170 174017 519204
rect 174029 519170 174079 519204
rect 174079 519170 174081 519204
rect 174093 519170 174113 519204
rect 174113 519170 174145 519204
rect 173965 519161 174017 519170
rect 174029 519161 174081 519170
rect 174093 519161 174145 519170
rect 174157 519204 174209 519213
rect 174157 519170 174171 519204
rect 174171 519170 174205 519204
rect 174205 519170 174209 519204
rect 174157 519161 174209 519170
rect 174221 519204 174273 519213
rect 177783 519204 177835 519213
rect 174221 519170 174263 519204
rect 174263 519170 174273 519204
rect 177783 519170 177793 519204
rect 177793 519170 177835 519204
rect 174221 519161 174273 519170
rect 177783 519161 177835 519170
rect 177847 519204 177899 519213
rect 177847 519170 177851 519204
rect 177851 519170 177885 519204
rect 177885 519170 177899 519204
rect 177847 519161 177899 519170
rect 177911 519204 177963 519213
rect 177975 519204 178027 519213
rect 178039 519204 178091 519213
rect 181601 519204 181653 519213
rect 181665 519204 181717 519213
rect 181729 519204 181781 519213
rect 177911 519170 177943 519204
rect 177943 519170 177963 519204
rect 177975 519170 177977 519204
rect 177977 519170 178027 519204
rect 178039 519170 178069 519204
rect 178069 519170 178091 519204
rect 181601 519170 181623 519204
rect 181623 519170 181653 519204
rect 181665 519170 181715 519204
rect 181715 519170 181717 519204
rect 181729 519170 181749 519204
rect 181749 519170 181781 519204
rect 177911 519161 177963 519170
rect 177975 519161 178027 519170
rect 178039 519161 178091 519170
rect 181601 519161 181653 519170
rect 181665 519161 181717 519170
rect 181729 519161 181781 519170
rect 181793 519204 181845 519213
rect 181793 519170 181807 519204
rect 181807 519170 181841 519204
rect 181841 519170 181845 519204
rect 181793 519161 181845 519170
rect 181857 519204 181909 519213
rect 185419 519204 185471 519213
rect 181857 519170 181899 519204
rect 181899 519170 181909 519204
rect 185419 519170 185429 519204
rect 185429 519170 185471 519204
rect 181857 519161 181909 519170
rect 185419 519161 185471 519170
rect 185483 519204 185535 519213
rect 185483 519170 185487 519204
rect 185487 519170 185521 519204
rect 185521 519170 185535 519204
rect 185483 519161 185535 519170
rect 185547 519204 185599 519213
rect 185611 519204 185663 519213
rect 185675 519204 185727 519213
rect 185547 519170 185579 519204
rect 185579 519170 185599 519204
rect 185611 519170 185613 519204
rect 185613 519170 185663 519204
rect 185675 519170 185705 519204
rect 185705 519170 185727 519204
rect 185547 519161 185599 519170
rect 185611 519161 185663 519170
rect 185675 519161 185727 519170
rect 174625 518660 174677 518669
rect 174625 518626 174631 518660
rect 174631 518626 174665 518660
rect 174665 518626 174677 518660
rect 174625 518617 174677 518626
rect 174689 518660 174741 518669
rect 174753 518660 174805 518669
rect 174817 518660 174869 518669
rect 174689 518626 174723 518660
rect 174723 518626 174741 518660
rect 174753 518626 174757 518660
rect 174757 518626 174805 518660
rect 174817 518626 174849 518660
rect 174849 518626 174869 518660
rect 174689 518617 174741 518626
rect 174753 518617 174805 518626
rect 174817 518617 174869 518626
rect 174881 518660 174933 518669
rect 174881 518626 174907 518660
rect 174907 518626 174933 518660
rect 174881 518617 174933 518626
rect 178443 518617 178495 518669
rect 178507 518660 178559 518669
rect 178507 518626 178529 518660
rect 178529 518626 178559 518660
rect 178507 518617 178559 518626
rect 178571 518660 178623 518669
rect 178571 518626 178587 518660
rect 178587 518626 178621 518660
rect 178621 518626 178623 518660
rect 178571 518617 178623 518626
rect 178635 518660 178687 518669
rect 178699 518660 178751 518669
rect 182261 518660 182313 518669
rect 178635 518626 178679 518660
rect 178679 518626 178687 518660
rect 178699 518626 178713 518660
rect 178713 518626 178751 518660
rect 182261 518626 182267 518660
rect 182267 518626 182301 518660
rect 182301 518626 182313 518660
rect 178635 518617 178687 518626
rect 178699 518617 178751 518626
rect 182261 518617 182313 518626
rect 182325 518660 182377 518669
rect 182389 518660 182441 518669
rect 182453 518660 182505 518669
rect 182325 518626 182359 518660
rect 182359 518626 182377 518660
rect 182389 518626 182393 518660
rect 182393 518626 182441 518660
rect 182453 518626 182485 518660
rect 182485 518626 182505 518660
rect 182325 518617 182377 518626
rect 182389 518617 182441 518626
rect 182453 518617 182505 518626
rect 182517 518660 182569 518669
rect 182517 518626 182543 518660
rect 182543 518626 182569 518660
rect 182517 518617 182569 518626
rect 186079 518617 186131 518669
rect 186143 518660 186195 518669
rect 186143 518626 186165 518660
rect 186165 518626 186195 518660
rect 186143 518617 186195 518626
rect 186207 518660 186259 518669
rect 186207 518626 186223 518660
rect 186223 518626 186257 518660
rect 186257 518626 186259 518660
rect 186207 518617 186259 518626
rect 186271 518660 186323 518669
rect 186335 518660 186387 518669
rect 186271 518626 186315 518660
rect 186315 518626 186323 518660
rect 186335 518626 186349 518660
rect 186349 518626 186387 518660
rect 186271 518617 186323 518626
rect 186335 518617 186387 518626
rect 173965 518116 174017 518125
rect 174029 518116 174081 518125
rect 174093 518116 174145 518125
rect 173965 518082 173987 518116
rect 173987 518082 174017 518116
rect 174029 518082 174079 518116
rect 174079 518082 174081 518116
rect 174093 518082 174113 518116
rect 174113 518082 174145 518116
rect 173965 518073 174017 518082
rect 174029 518073 174081 518082
rect 174093 518073 174145 518082
rect 174157 518116 174209 518125
rect 174157 518082 174171 518116
rect 174171 518082 174205 518116
rect 174205 518082 174209 518116
rect 174157 518073 174209 518082
rect 174221 518116 174273 518125
rect 177783 518116 177835 518125
rect 174221 518082 174263 518116
rect 174263 518082 174273 518116
rect 177783 518082 177793 518116
rect 177793 518082 177835 518116
rect 174221 518073 174273 518082
rect 177783 518073 177835 518082
rect 177847 518116 177899 518125
rect 177847 518082 177851 518116
rect 177851 518082 177885 518116
rect 177885 518082 177899 518116
rect 177847 518073 177899 518082
rect 177911 518116 177963 518125
rect 177975 518116 178027 518125
rect 178039 518116 178091 518125
rect 181601 518116 181653 518125
rect 181665 518116 181717 518125
rect 181729 518116 181781 518125
rect 177911 518082 177943 518116
rect 177943 518082 177963 518116
rect 177975 518082 177977 518116
rect 177977 518082 178027 518116
rect 178039 518082 178069 518116
rect 178069 518082 178091 518116
rect 181601 518082 181623 518116
rect 181623 518082 181653 518116
rect 181665 518082 181715 518116
rect 181715 518082 181717 518116
rect 181729 518082 181749 518116
rect 181749 518082 181781 518116
rect 177911 518073 177963 518082
rect 177975 518073 178027 518082
rect 178039 518073 178091 518082
rect 181601 518073 181653 518082
rect 181665 518073 181717 518082
rect 181729 518073 181781 518082
rect 181793 518116 181845 518125
rect 181793 518082 181807 518116
rect 181807 518082 181841 518116
rect 181841 518082 181845 518116
rect 181793 518073 181845 518082
rect 181857 518116 181909 518125
rect 185419 518116 185471 518125
rect 181857 518082 181899 518116
rect 181899 518082 181909 518116
rect 185419 518082 185429 518116
rect 185429 518082 185471 518116
rect 181857 518073 181909 518082
rect 185419 518073 185471 518082
rect 185483 518116 185535 518125
rect 185483 518082 185487 518116
rect 185487 518082 185521 518116
rect 185521 518082 185535 518116
rect 185483 518073 185535 518082
rect 185547 518116 185599 518125
rect 185611 518116 185663 518125
rect 185675 518116 185727 518125
rect 185547 518082 185579 518116
rect 185579 518082 185599 518116
rect 185611 518082 185613 518116
rect 185613 518082 185663 518116
rect 185675 518082 185705 518116
rect 185705 518082 185727 518116
rect 185547 518073 185599 518082
rect 185611 518073 185663 518082
rect 185675 518073 185727 518082
rect 174625 517572 174677 517581
rect 174625 517538 174631 517572
rect 174631 517538 174665 517572
rect 174665 517538 174677 517572
rect 174625 517529 174677 517538
rect 174689 517572 174741 517581
rect 174753 517572 174805 517581
rect 174817 517572 174869 517581
rect 174689 517538 174723 517572
rect 174723 517538 174741 517572
rect 174753 517538 174757 517572
rect 174757 517538 174805 517572
rect 174817 517538 174849 517572
rect 174849 517538 174869 517572
rect 174689 517529 174741 517538
rect 174753 517529 174805 517538
rect 174817 517529 174869 517538
rect 174881 517572 174933 517581
rect 174881 517538 174907 517572
rect 174907 517538 174933 517572
rect 174881 517529 174933 517538
rect 178443 517529 178495 517581
rect 178507 517572 178559 517581
rect 178507 517538 178529 517572
rect 178529 517538 178559 517572
rect 178507 517529 178559 517538
rect 178571 517572 178623 517581
rect 178571 517538 178587 517572
rect 178587 517538 178621 517572
rect 178621 517538 178623 517572
rect 178571 517529 178623 517538
rect 178635 517572 178687 517581
rect 178699 517572 178751 517581
rect 182261 517572 182313 517581
rect 178635 517538 178679 517572
rect 178679 517538 178687 517572
rect 178699 517538 178713 517572
rect 178713 517538 178751 517572
rect 182261 517538 182267 517572
rect 182267 517538 182301 517572
rect 182301 517538 182313 517572
rect 178635 517529 178687 517538
rect 178699 517529 178751 517538
rect 182261 517529 182313 517538
rect 182325 517572 182377 517581
rect 182389 517572 182441 517581
rect 182453 517572 182505 517581
rect 182325 517538 182359 517572
rect 182359 517538 182377 517572
rect 182389 517538 182393 517572
rect 182393 517538 182441 517572
rect 182453 517538 182485 517572
rect 182485 517538 182505 517572
rect 182325 517529 182377 517538
rect 182389 517529 182441 517538
rect 182453 517529 182505 517538
rect 182517 517572 182569 517581
rect 182517 517538 182543 517572
rect 182543 517538 182569 517572
rect 182517 517529 182569 517538
rect 186079 517529 186131 517581
rect 186143 517572 186195 517581
rect 186143 517538 186165 517572
rect 186165 517538 186195 517572
rect 186143 517529 186195 517538
rect 186207 517572 186259 517581
rect 186207 517538 186223 517572
rect 186223 517538 186257 517572
rect 186257 517538 186259 517572
rect 186207 517529 186259 517538
rect 186271 517572 186323 517581
rect 186335 517572 186387 517581
rect 186271 517538 186315 517572
rect 186315 517538 186323 517572
rect 186335 517538 186349 517572
rect 186349 517538 186387 517572
rect 186271 517529 186323 517538
rect 186335 517529 186387 517538
rect 177658 517427 177710 517479
rect 178302 517427 178354 517479
rect 173965 517028 174017 517037
rect 174029 517028 174081 517037
rect 174093 517028 174145 517037
rect 173965 516994 173987 517028
rect 173987 516994 174017 517028
rect 174029 516994 174079 517028
rect 174079 516994 174081 517028
rect 174093 516994 174113 517028
rect 174113 516994 174145 517028
rect 173965 516985 174017 516994
rect 174029 516985 174081 516994
rect 174093 516985 174145 516994
rect 174157 517028 174209 517037
rect 174157 516994 174171 517028
rect 174171 516994 174205 517028
rect 174205 516994 174209 517028
rect 174157 516985 174209 516994
rect 174221 517028 174273 517037
rect 177783 517028 177835 517037
rect 174221 516994 174263 517028
rect 174263 516994 174273 517028
rect 177783 516994 177793 517028
rect 177793 516994 177835 517028
rect 174221 516985 174273 516994
rect 177783 516985 177835 516994
rect 177847 517028 177899 517037
rect 177847 516994 177851 517028
rect 177851 516994 177885 517028
rect 177885 516994 177899 517028
rect 177847 516985 177899 516994
rect 177911 517028 177963 517037
rect 177975 517028 178027 517037
rect 178039 517028 178091 517037
rect 181601 517028 181653 517037
rect 181665 517028 181717 517037
rect 181729 517028 181781 517037
rect 177911 516994 177943 517028
rect 177943 516994 177963 517028
rect 177975 516994 177977 517028
rect 177977 516994 178027 517028
rect 178039 516994 178069 517028
rect 178069 516994 178091 517028
rect 181601 516994 181623 517028
rect 181623 516994 181653 517028
rect 181665 516994 181715 517028
rect 181715 516994 181717 517028
rect 181729 516994 181749 517028
rect 181749 516994 181781 517028
rect 177911 516985 177963 516994
rect 177975 516985 178027 516994
rect 178039 516985 178091 516994
rect 181601 516985 181653 516994
rect 181665 516985 181717 516994
rect 181729 516985 181781 516994
rect 181793 517028 181845 517037
rect 181793 516994 181807 517028
rect 181807 516994 181841 517028
rect 181841 516994 181845 517028
rect 181793 516985 181845 516994
rect 181857 517028 181909 517037
rect 185419 517028 185471 517037
rect 181857 516994 181899 517028
rect 181899 516994 181909 517028
rect 185419 516994 185429 517028
rect 185429 516994 185471 517028
rect 181857 516985 181909 516994
rect 185419 516985 185471 516994
rect 185483 517028 185535 517037
rect 185483 516994 185487 517028
rect 185487 516994 185521 517028
rect 185521 516994 185535 517028
rect 185483 516985 185535 516994
rect 185547 517028 185599 517037
rect 185611 517028 185663 517037
rect 185675 517028 185727 517037
rect 185547 516994 185579 517028
rect 185579 516994 185599 517028
rect 185611 516994 185613 517028
rect 185613 516994 185663 517028
rect 185675 516994 185705 517028
rect 185705 516994 185727 517028
rect 185547 516985 185599 516994
rect 185611 516985 185663 516994
rect 185675 516985 185727 516994
rect 174625 516484 174677 516493
rect 174625 516450 174631 516484
rect 174631 516450 174665 516484
rect 174665 516450 174677 516484
rect 174625 516441 174677 516450
rect 174689 516484 174741 516493
rect 174753 516484 174805 516493
rect 174817 516484 174869 516493
rect 174689 516450 174723 516484
rect 174723 516450 174741 516484
rect 174753 516450 174757 516484
rect 174757 516450 174805 516484
rect 174817 516450 174849 516484
rect 174849 516450 174869 516484
rect 174689 516441 174741 516450
rect 174753 516441 174805 516450
rect 174817 516441 174869 516450
rect 174881 516484 174933 516493
rect 174881 516450 174907 516484
rect 174907 516450 174933 516484
rect 174881 516441 174933 516450
rect 178443 516441 178495 516493
rect 178507 516484 178559 516493
rect 178507 516450 178529 516484
rect 178529 516450 178559 516484
rect 178507 516441 178559 516450
rect 178571 516484 178623 516493
rect 178571 516450 178587 516484
rect 178587 516450 178621 516484
rect 178621 516450 178623 516484
rect 178571 516441 178623 516450
rect 178635 516484 178687 516493
rect 178699 516484 178751 516493
rect 182261 516484 182313 516493
rect 178635 516450 178679 516484
rect 178679 516450 178687 516484
rect 178699 516450 178713 516484
rect 178713 516450 178751 516484
rect 182261 516450 182267 516484
rect 182267 516450 182301 516484
rect 182301 516450 182313 516484
rect 178635 516441 178687 516450
rect 178699 516441 178751 516450
rect 182261 516441 182313 516450
rect 182325 516484 182377 516493
rect 182389 516484 182441 516493
rect 182453 516484 182505 516493
rect 182325 516450 182359 516484
rect 182359 516450 182377 516484
rect 182389 516450 182393 516484
rect 182393 516450 182441 516484
rect 182453 516450 182485 516484
rect 182485 516450 182505 516484
rect 182325 516441 182377 516450
rect 182389 516441 182441 516450
rect 182453 516441 182505 516450
rect 182517 516484 182569 516493
rect 182517 516450 182543 516484
rect 182543 516450 182569 516484
rect 182517 516441 182569 516450
rect 186079 516441 186131 516493
rect 186143 516484 186195 516493
rect 186143 516450 186165 516484
rect 186165 516450 186195 516484
rect 186143 516441 186195 516450
rect 186207 516484 186259 516493
rect 186207 516450 186223 516484
rect 186223 516450 186257 516484
rect 186257 516450 186259 516484
rect 186207 516441 186259 516450
rect 186271 516484 186323 516493
rect 186335 516484 186387 516493
rect 186271 516450 186315 516484
rect 186315 516450 186323 516484
rect 186335 516450 186349 516484
rect 186349 516450 186387 516484
rect 186271 516441 186323 516450
rect 186335 516441 186387 516450
rect 173965 515940 174017 515949
rect 174029 515940 174081 515949
rect 174093 515940 174145 515949
rect 173965 515906 173987 515940
rect 173987 515906 174017 515940
rect 174029 515906 174079 515940
rect 174079 515906 174081 515940
rect 174093 515906 174113 515940
rect 174113 515906 174145 515940
rect 173965 515897 174017 515906
rect 174029 515897 174081 515906
rect 174093 515897 174145 515906
rect 174157 515940 174209 515949
rect 174157 515906 174171 515940
rect 174171 515906 174205 515940
rect 174205 515906 174209 515940
rect 174157 515897 174209 515906
rect 174221 515940 174273 515949
rect 177783 515940 177835 515949
rect 174221 515906 174263 515940
rect 174263 515906 174273 515940
rect 177783 515906 177793 515940
rect 177793 515906 177835 515940
rect 174221 515897 174273 515906
rect 177783 515897 177835 515906
rect 177847 515940 177899 515949
rect 177847 515906 177851 515940
rect 177851 515906 177885 515940
rect 177885 515906 177899 515940
rect 177847 515897 177899 515906
rect 177911 515940 177963 515949
rect 177975 515940 178027 515949
rect 178039 515940 178091 515949
rect 181601 515940 181653 515949
rect 181665 515940 181717 515949
rect 181729 515940 181781 515949
rect 177911 515906 177943 515940
rect 177943 515906 177963 515940
rect 177975 515906 177977 515940
rect 177977 515906 178027 515940
rect 178039 515906 178069 515940
rect 178069 515906 178091 515940
rect 181601 515906 181623 515940
rect 181623 515906 181653 515940
rect 181665 515906 181715 515940
rect 181715 515906 181717 515940
rect 181729 515906 181749 515940
rect 181749 515906 181781 515940
rect 177911 515897 177963 515906
rect 177975 515897 178027 515906
rect 178039 515897 178091 515906
rect 181601 515897 181653 515906
rect 181665 515897 181717 515906
rect 181729 515897 181781 515906
rect 181793 515940 181845 515949
rect 181793 515906 181807 515940
rect 181807 515906 181841 515940
rect 181841 515906 181845 515940
rect 181793 515897 181845 515906
rect 181857 515940 181909 515949
rect 185419 515940 185471 515949
rect 181857 515906 181899 515940
rect 181899 515906 181909 515940
rect 185419 515906 185429 515940
rect 185429 515906 185471 515940
rect 181857 515897 181909 515906
rect 185419 515897 185471 515906
rect 185483 515940 185535 515949
rect 185483 515906 185487 515940
rect 185487 515906 185521 515940
rect 185521 515906 185535 515940
rect 185483 515897 185535 515906
rect 185547 515940 185599 515949
rect 185611 515940 185663 515949
rect 185675 515940 185727 515949
rect 185547 515906 185579 515940
rect 185579 515906 185599 515940
rect 185611 515906 185613 515940
rect 185613 515906 185663 515940
rect 185675 515906 185705 515940
rect 185705 515906 185727 515940
rect 185547 515897 185599 515906
rect 185611 515897 185663 515906
rect 185675 515897 185727 515906
rect 173610 515838 173662 515847
rect 173610 515804 173619 515838
rect 173619 515804 173653 515838
rect 173653 515804 173662 515838
rect 173610 515795 173662 515804
rect 181338 515795 181390 515847
rect 186582 515838 186634 515847
rect 186582 515804 186591 515838
rect 186591 515804 186625 515838
rect 186625 515804 186634 515838
rect 186582 515795 186634 515804
rect 173334 515523 173386 515575
rect 186490 515566 186542 515575
rect 186490 515532 186499 515566
rect 186499 515532 186533 515566
rect 186533 515532 186542 515566
rect 186490 515523 186542 515532
rect 182166 515455 182218 515507
rect 174625 515396 174677 515405
rect 174625 515362 174631 515396
rect 174631 515362 174665 515396
rect 174665 515362 174677 515396
rect 174625 515353 174677 515362
rect 174689 515396 174741 515405
rect 174753 515396 174805 515405
rect 174817 515396 174869 515405
rect 174689 515362 174723 515396
rect 174723 515362 174741 515396
rect 174753 515362 174757 515396
rect 174757 515362 174805 515396
rect 174817 515362 174849 515396
rect 174849 515362 174869 515396
rect 174689 515353 174741 515362
rect 174753 515353 174805 515362
rect 174817 515353 174869 515362
rect 174881 515396 174933 515405
rect 174881 515362 174907 515396
rect 174907 515362 174933 515396
rect 174881 515353 174933 515362
rect 178443 515353 178495 515405
rect 178507 515396 178559 515405
rect 178507 515362 178529 515396
rect 178529 515362 178559 515396
rect 178507 515353 178559 515362
rect 178571 515396 178623 515405
rect 178571 515362 178587 515396
rect 178587 515362 178621 515396
rect 178621 515362 178623 515396
rect 178571 515353 178623 515362
rect 178635 515396 178687 515405
rect 178699 515396 178751 515405
rect 182261 515396 182313 515405
rect 178635 515362 178679 515396
rect 178679 515362 178687 515396
rect 178699 515362 178713 515396
rect 178713 515362 178751 515396
rect 182261 515362 182267 515396
rect 182267 515362 182301 515396
rect 182301 515362 182313 515396
rect 178635 515353 178687 515362
rect 178699 515353 178751 515362
rect 182261 515353 182313 515362
rect 182325 515396 182377 515405
rect 182389 515396 182441 515405
rect 182453 515396 182505 515405
rect 182325 515362 182359 515396
rect 182359 515362 182377 515396
rect 182389 515362 182393 515396
rect 182393 515362 182441 515396
rect 182453 515362 182485 515396
rect 182485 515362 182505 515396
rect 182325 515353 182377 515362
rect 182389 515353 182441 515362
rect 182453 515353 182505 515362
rect 182517 515396 182569 515405
rect 182517 515362 182543 515396
rect 182543 515362 182569 515396
rect 182517 515353 182569 515362
rect 186079 515353 186131 515405
rect 186143 515396 186195 515405
rect 186143 515362 186165 515396
rect 186165 515362 186195 515396
rect 186143 515353 186195 515362
rect 186207 515396 186259 515405
rect 186207 515362 186223 515396
rect 186223 515362 186257 515396
rect 186257 515362 186259 515396
rect 186207 515353 186259 515362
rect 186271 515396 186323 515405
rect 186335 515396 186387 515405
rect 186271 515362 186315 515396
rect 186315 515362 186323 515396
rect 186335 515362 186349 515396
rect 186349 515362 186387 515396
rect 186271 515353 186323 515362
rect 186335 515353 186387 515362
rect 173250 512810 173450 513000
rect 2000 507000 4000 509000
rect 177580 512810 177780 513000
rect 181910 512810 182110 513000
rect 2000 464000 4000 466000
rect 186230 512810 186430 513000
rect 2000 421000 4000 423000
rect 2000 378000 4000 380000
<< metal2 >>
rect 18000 701000 20000 701010
rect 18000 698990 20000 699000
rect 70000 701000 72000 701010
rect 70000 698990 72000 699000
rect 122000 701000 124000 701010
rect 122000 698990 124000 699000
rect 3000 684000 5000 684010
rect 3000 681990 5000 682000
rect 146000 628000 148000 628010
rect 146000 546000 148000 626000
rect 146000 543990 148000 544000
rect 154000 553000 156000 553010
rect 154000 540000 156000 551000
rect 165880 541027 166010 541057
rect 165880 540927 165890 541027
rect 166000 540927 166010 541027
rect 165880 540907 166010 540927
rect 165880 540807 165890 540907
rect 166000 540807 166010 540907
rect 165880 540787 166010 540807
rect 165880 540687 165890 540787
rect 166000 540687 166010 540787
rect 165880 540667 166010 540687
rect 169680 541027 169810 541057
rect 169680 540927 169690 541027
rect 169800 540927 169810 541027
rect 169680 540907 169810 540927
rect 169680 540807 169690 540907
rect 169800 540807 169810 540907
rect 169680 540787 169810 540807
rect 169680 540687 169690 540787
rect 169800 540687 169810 540787
rect 169680 540667 169810 540687
rect 173380 541027 173510 541057
rect 173380 540927 173390 541027
rect 173500 540927 173510 541027
rect 173380 540907 173510 540927
rect 173380 540807 173390 540907
rect 173500 540807 173510 540907
rect 173380 540787 173510 540807
rect 173380 540687 173390 540787
rect 173500 540687 173510 540787
rect 173380 540667 173510 540687
rect 176880 541027 177010 541057
rect 176880 540927 176890 541027
rect 177000 540927 177010 541027
rect 176880 540907 177010 540927
rect 176880 540807 176890 540907
rect 177000 540807 177010 540907
rect 176880 540787 177010 540807
rect 176880 540687 176890 540787
rect 177000 540687 177010 540787
rect 176880 540667 177010 540687
rect 180480 541027 180610 541057
rect 180480 540927 180490 541027
rect 180600 540927 180610 541027
rect 180480 540907 180610 540927
rect 180480 540807 180490 540907
rect 180600 540807 180610 540907
rect 180480 540787 180610 540807
rect 180480 540687 180490 540787
rect 180600 540687 180610 540787
rect 180480 540667 180610 540687
rect 183780 541027 183910 541057
rect 183780 540927 183790 541027
rect 183900 540927 183910 541027
rect 183780 540907 183910 540927
rect 183780 540807 183790 540907
rect 183900 540807 183910 540907
rect 183780 540787 183910 540807
rect 183780 540687 183790 540787
rect 183900 540687 183910 540787
rect 183780 540667 183910 540687
rect 187080 541027 187210 541057
rect 187080 540927 187090 541027
rect 187200 540927 187210 541027
rect 187080 540907 187210 540927
rect 187080 540807 187090 540907
rect 187200 540807 187210 540907
rect 187080 540787 187210 540807
rect 187080 540687 187090 540787
rect 187200 540687 187210 540787
rect 187080 540667 187210 540687
rect 190380 541027 190510 541057
rect 190380 540927 190390 541027
rect 190500 540927 190510 541027
rect 190380 540907 190510 540927
rect 190380 540807 190390 540907
rect 190500 540807 190510 540907
rect 190380 540787 190510 540807
rect 190380 540687 190390 540787
rect 190500 540687 190510 540787
rect 190380 540667 190510 540687
rect 163030 538897 163330 538907
rect 161380 538697 161530 538707
rect 159390 538687 159490 538697
rect 159390 538587 159400 538687
rect 159480 538587 159490 538687
rect 159390 538372 159490 538587
rect 161380 538577 161390 538697
rect 161510 538577 161530 538697
rect 165930 538847 166010 540667
rect 166680 540277 166880 540287
rect 166680 540097 166690 540277
rect 166870 540097 166880 540277
rect 166680 540087 166880 540097
rect 166680 539337 166880 539347
rect 166680 539157 166690 539337
rect 166870 539157 166880 539337
rect 166680 539147 166880 539157
rect 169730 538847 169810 540667
rect 170480 540277 170680 540287
rect 170480 540097 170490 540277
rect 170670 540097 170680 540277
rect 170480 540087 170680 540097
rect 170480 539337 170680 539347
rect 170480 539157 170490 539337
rect 170670 539157 170680 539337
rect 170480 539147 170680 539157
rect 173430 538847 173510 540667
rect 174180 540287 174380 540297
rect 174180 540107 174190 540287
rect 174370 540107 174380 540287
rect 174180 540097 174380 540107
rect 174180 539337 174380 539347
rect 174180 539157 174190 539337
rect 174370 539157 174380 539337
rect 174180 539147 174380 539157
rect 176930 538847 177010 540667
rect 177690 540277 177890 540287
rect 177690 540097 177700 540277
rect 177880 540097 177890 540277
rect 177690 540087 177890 540097
rect 177680 539337 177880 539347
rect 177680 539157 177690 539337
rect 177870 539157 177880 539337
rect 177680 539147 177880 539157
rect 180530 538847 180610 540667
rect 181280 540277 181480 540287
rect 181280 540097 181290 540277
rect 181470 540097 181480 540277
rect 181280 540087 181480 540097
rect 181280 539337 181480 539347
rect 181280 539157 181290 539337
rect 181470 539157 181480 539337
rect 181280 539147 181480 539157
rect 183830 538847 183910 540667
rect 184580 540277 184780 540287
rect 184580 540097 184590 540277
rect 184770 540097 184780 540277
rect 184580 540087 184780 540097
rect 184580 539337 184780 539347
rect 184580 539157 184590 539337
rect 184770 539157 184780 539337
rect 184580 539147 184780 539157
rect 187130 538847 187210 540667
rect 187890 540277 188090 540287
rect 187890 540097 187900 540277
rect 188080 540097 188090 540277
rect 187890 540087 188090 540097
rect 187880 539337 188080 539347
rect 187880 539157 187890 539337
rect 188070 539157 188080 539337
rect 187880 539147 188080 539157
rect 190430 538847 190510 540667
rect 191180 540277 191380 540287
rect 191180 540097 191190 540277
rect 191370 540097 191380 540277
rect 191180 540087 191380 540097
rect 191780 540277 192000 540287
rect 191780 540097 191810 540277
rect 191990 540097 192000 540277
rect 191780 540087 192000 540097
rect 191190 539347 191390 539357
rect 191190 539167 191200 539347
rect 191380 539167 191390 539347
rect 191190 539157 191390 539167
rect 191810 539337 192010 539347
rect 191810 539157 191820 539337
rect 192000 539157 192010 539337
rect 191810 539147 192010 539157
rect 165880 538837 166060 538847
rect 165880 538737 165900 538837
rect 166040 538737 166060 538837
rect 165880 538727 166060 538737
rect 169680 538837 169860 538847
rect 169680 538737 169700 538837
rect 169840 538737 169860 538837
rect 169680 538727 169860 538737
rect 173380 538837 173560 538847
rect 173380 538737 173400 538837
rect 173540 538737 173560 538837
rect 173380 538727 173560 538737
rect 176880 538837 177060 538847
rect 176880 538737 176900 538837
rect 177040 538737 177060 538837
rect 176880 538727 177060 538737
rect 180480 538837 180660 538847
rect 180480 538737 180500 538837
rect 180640 538737 180660 538837
rect 180480 538727 180660 538737
rect 183780 538837 183960 538847
rect 183780 538737 183800 538837
rect 183940 538737 183960 538837
rect 183780 538727 183960 538737
rect 187080 538837 187260 538847
rect 187080 538737 187100 538837
rect 187240 538737 187260 538837
rect 187080 538727 187260 538737
rect 190380 538837 190560 538847
rect 190380 538737 190400 538837
rect 190540 538737 190560 538837
rect 190380 538727 190560 538737
rect 163030 538687 163330 538697
rect 161380 538567 161530 538577
rect 154000 537990 156000 538000
rect 159385 538327 159495 538372
rect 159385 538247 159400 538327
rect 159480 538247 159495 538327
rect 159385 536967 159495 538247
rect 162870 537977 162950 537987
rect 162870 537967 162880 537977
rect 161690 537917 162880 537967
rect 162940 537917 162950 537977
rect 161690 537777 161740 537917
rect 162870 537907 162950 537917
rect 161680 537767 161760 537777
rect 161680 537707 161690 537767
rect 161750 537707 161760 537767
rect 161680 537697 161760 537707
rect 157415 536957 159495 536967
rect 157415 536877 157420 536957
rect 157510 536877 159495 536957
rect 161770 536937 161870 536957
rect 161770 536917 161790 536937
rect 157415 536857 159495 536877
rect 161090 536857 161790 536917
rect 161850 536857 161870 536937
rect 157420 535007 157500 536857
rect 158480 536597 158590 536857
rect 161090 536837 161870 536857
rect 161090 536597 161170 536837
rect 158470 536587 158600 536597
rect 158470 536427 158480 536587
rect 158580 536427 158600 536587
rect 161070 536577 161190 536597
rect 161070 536497 161090 536577
rect 161170 536497 161190 536577
rect 161070 536477 161190 536497
rect 158470 536407 158600 536427
rect 163820 536317 189030 536327
rect 163820 536307 182190 536317
rect 163820 536297 178870 536307
rect 163820 536267 166930 536297
rect 163820 535937 163840 536267
rect 164050 536077 166930 536267
rect 167260 536287 172610 536297
rect 167260 536077 169570 536287
rect 164050 536007 169570 536077
rect 169870 536007 172610 536287
rect 172940 536287 178870 536297
rect 172940 536007 175280 536287
rect 164050 535977 175280 536007
rect 175500 535997 178870 536287
rect 179070 536057 182190 536307
rect 182390 536307 189030 536317
rect 182390 536297 188780 536307
rect 182390 536177 185490 536297
rect 185700 536177 188780 536297
rect 182390 536067 188780 536177
rect 189000 536067 189030 536307
rect 182390 536057 189030 536067
rect 179070 535997 189030 536057
rect 175500 535977 189030 535997
rect 164050 535937 189030 535977
rect 163820 535907 189030 535937
rect 160170 535607 160370 535637
rect 163530 535607 167240 535637
rect 160170 535467 160200 535607
rect 160350 535597 160370 535607
rect 160170 535457 160210 535467
rect 160360 535457 160370 535597
rect 160170 535447 160370 535457
rect 163480 535587 167240 535607
rect 163480 535457 166720 535587
rect 166850 535577 167240 535587
rect 166850 535457 166900 535577
rect 163480 535447 166900 535457
rect 167030 535557 167240 535577
rect 167030 535447 167080 535557
rect 163480 535427 167080 535447
rect 167210 535427 167240 535557
rect 163480 535397 167240 535427
rect 163480 535267 166700 535397
rect 166830 535387 167240 535397
rect 166830 535267 166890 535387
rect 163480 535257 166890 535267
rect 167020 535377 167240 535387
rect 167020 535257 167090 535377
rect 163480 535247 167090 535257
rect 167220 535247 167240 535377
rect 163480 535217 167240 535247
rect 163480 535007 163900 535217
rect 157420 534587 163900 535007
rect 185060 532807 185190 532817
rect 172412 532777 172468 532787
rect 174490 532777 174620 532787
rect 176644 532777 176700 532787
rect 178760 532777 178816 532787
rect 180876 532777 180932 532787
rect 182992 532777 183048 532787
rect 172360 532767 172490 532777
rect 174490 532597 174620 532607
rect 176580 532767 176710 532777
rect 172360 532587 172490 532597
rect 172412 531987 172468 532587
rect 174528 531987 174584 532597
rect 176580 532587 176710 532597
rect 178700 532767 178830 532777
rect 178700 532587 178830 532597
rect 180870 532767 181000 532777
rect 180870 532587 181000 532597
rect 182960 532767 183090 532777
rect 187224 532777 187280 532787
rect 185060 532627 185190 532637
rect 187170 532767 187290 532777
rect 187270 532627 187290 532767
rect 182960 532587 183090 532597
rect 176644 531987 176700 532587
rect 178760 531987 178816 532587
rect 180876 531987 180932 532587
rect 182992 531987 183048 532587
rect 185108 531987 185164 532627
rect 187170 532607 187290 532627
rect 187224 531987 187280 532607
rect 172426 530473 172454 531987
rect 174542 530473 174570 531987
rect 176658 531645 176686 531987
rect 178774 531645 178802 531987
rect 176658 531617 176778 531645
rect 178774 531617 178894 531645
rect 174625 530639 174933 530648
rect 174625 530637 174631 530639
rect 174687 530637 174711 530639
rect 174767 530637 174791 530639
rect 174847 530637 174871 530639
rect 174927 530637 174933 530639
rect 174687 530585 174689 530637
rect 174869 530585 174871 530637
rect 174625 530583 174631 530585
rect 174687 530583 174711 530585
rect 174767 530583 174791 530585
rect 174847 530583 174871 530585
rect 174927 530583 174933 530585
rect 174625 530574 174933 530583
rect 176750 530473 176778 531617
rect 178443 530639 178751 530648
rect 178443 530637 178449 530639
rect 178505 530637 178529 530639
rect 178585 530637 178609 530639
rect 178665 530637 178689 530639
rect 178745 530637 178751 530639
rect 178505 530585 178507 530637
rect 178687 530585 178689 530637
rect 178443 530583 178449 530585
rect 178505 530583 178529 530585
rect 178585 530583 178609 530585
rect 178665 530583 178689 530585
rect 178745 530583 178751 530585
rect 178443 530574 178751 530583
rect 178866 530557 178894 531617
rect 178774 530541 178894 530557
rect 176830 530535 176882 530541
rect 176830 530477 176882 530483
rect 178762 530535 178894 530541
rect 178814 530529 178894 530535
rect 179498 530535 179550 530541
rect 178762 530477 178814 530483
rect 179498 530477 179550 530483
rect 172414 530467 172466 530473
rect 172414 530409 172466 530415
rect 174530 530467 174582 530473
rect 174530 530409 174582 530415
rect 176738 530467 176790 530473
rect 176738 530409 176790 530415
rect 174806 530399 174858 530405
rect 174806 530341 174858 530347
rect 175450 530399 175502 530405
rect 175450 530341 175502 530347
rect 173965 530095 174273 530104
rect 173965 530093 173971 530095
rect 174027 530093 174051 530095
rect 174107 530093 174131 530095
rect 174187 530093 174211 530095
rect 174267 530093 174273 530095
rect 174027 530041 174029 530093
rect 174209 530041 174211 530093
rect 173965 530039 173971 530041
rect 174027 530039 174051 530041
rect 174107 530039 174131 530041
rect 174187 530039 174211 530041
rect 174267 530039 174273 530041
rect 173965 530030 174273 530039
rect 174818 529861 174846 530341
rect 174806 529855 174858 529861
rect 174806 529797 174858 529803
rect 175358 529651 175410 529657
rect 175358 529593 175410 529599
rect 174625 529551 174933 529560
rect 174625 529549 174631 529551
rect 174687 529549 174711 529551
rect 174767 529549 174791 529551
rect 174847 529549 174871 529551
rect 174927 529549 174933 529551
rect 174687 529497 174689 529549
rect 174869 529497 174871 529549
rect 174625 529495 174631 529497
rect 174687 529495 174711 529497
rect 174767 529495 174791 529497
rect 174847 529495 174871 529497
rect 174927 529495 174933 529497
rect 174625 529486 174933 529495
rect 175370 529453 175398 529593
rect 175358 529447 175410 529453
rect 175358 529389 175410 529395
rect 175462 529317 175490 530341
rect 176646 530331 176698 530337
rect 176646 530273 176698 530279
rect 176094 529651 176146 529657
rect 176094 529593 176146 529599
rect 175450 529311 175502 529317
rect 175450 529253 175502 529259
rect 173610 529243 173662 529249
rect 173610 529185 173662 529191
rect 175266 529243 175318 529249
rect 175266 529185 175318 529191
rect 173622 515853 173650 529185
rect 173965 529007 174273 529016
rect 173965 529005 173971 529007
rect 174027 529005 174051 529007
rect 174107 529005 174131 529007
rect 174187 529005 174211 529007
rect 174267 529005 174273 529007
rect 174027 528953 174029 529005
rect 174209 528953 174211 529005
rect 173965 528951 173971 528953
rect 174027 528951 174051 528953
rect 174107 528951 174131 528953
rect 174187 528951 174211 528953
rect 174267 528951 174273 528953
rect 173965 528942 174273 528951
rect 175278 528909 175306 529185
rect 176106 529113 176134 529593
rect 175910 529107 175962 529113
rect 175910 529049 175962 529055
rect 176094 529107 176146 529113
rect 176094 529049 176146 529055
rect 175266 528903 175318 528909
rect 175266 528845 175318 528851
rect 175922 528705 175950 529049
rect 175910 528699 175962 528705
rect 175910 528641 175962 528647
rect 174625 528463 174933 528472
rect 174625 528461 174631 528463
rect 174687 528461 174711 528463
rect 174767 528461 174791 528463
rect 174847 528461 174871 528463
rect 174927 528461 174933 528463
rect 174687 528409 174689 528461
rect 174869 528409 174871 528461
rect 174625 528407 174631 528409
rect 174687 528407 174711 528409
rect 174767 528407 174791 528409
rect 174847 528407 174871 528409
rect 174927 528407 174933 528409
rect 174625 528398 174933 528407
rect 176106 528229 176134 529049
rect 176658 528909 176686 530273
rect 176842 529793 176870 530477
rect 178946 530399 178998 530405
rect 178946 530341 178998 530347
rect 179222 530399 179274 530405
rect 179222 530341 179274 530347
rect 177290 530331 177342 530337
rect 177290 530273 177342 530279
rect 178210 530331 178262 530337
rect 178210 530273 178262 530279
rect 176830 529787 176882 529793
rect 176830 529729 176882 529735
rect 176738 529311 176790 529317
rect 176738 529253 176790 529259
rect 176646 528903 176698 528909
rect 176646 528845 176698 528851
rect 176750 528569 176778 529253
rect 176278 528563 176330 528569
rect 176278 528505 176330 528511
rect 176370 528563 176422 528569
rect 176370 528505 176422 528511
rect 176738 528563 176790 528569
rect 176738 528505 176790 528511
rect 176094 528223 176146 528229
rect 176094 528165 176146 528171
rect 173965 527919 174273 527928
rect 173965 527917 173971 527919
rect 174027 527917 174051 527919
rect 174107 527917 174131 527919
rect 174187 527917 174211 527919
rect 174267 527917 174273 527919
rect 174027 527865 174029 527917
rect 174209 527865 174211 527917
rect 173965 527863 173971 527865
rect 174027 527863 174051 527865
rect 174107 527863 174131 527865
rect 174187 527863 174211 527865
rect 174267 527863 174273 527865
rect 173965 527854 174273 527863
rect 176290 527821 176318 528505
rect 176382 528297 176410 528505
rect 176750 528365 176778 528505
rect 176738 528359 176790 528365
rect 176738 528301 176790 528307
rect 176842 528297 176870 529729
rect 177302 529249 177330 530273
rect 177658 530195 177710 530201
rect 177658 530137 177710 530143
rect 177670 529725 177698 530137
rect 177783 530095 178091 530104
rect 177783 530093 177789 530095
rect 177845 530093 177869 530095
rect 177925 530093 177949 530095
rect 178005 530093 178029 530095
rect 178085 530093 178091 530095
rect 177845 530041 177847 530093
rect 178027 530041 178029 530093
rect 177783 530039 177789 530041
rect 177845 530039 177869 530041
rect 177925 530039 177949 530041
rect 178005 530039 178029 530041
rect 178085 530039 178091 530041
rect 177783 530030 178091 530039
rect 178222 529997 178250 530273
rect 178302 530195 178354 530201
rect 178302 530137 178354 530143
rect 178210 529991 178262 529997
rect 178210 529933 178262 529939
rect 178118 529923 178170 529929
rect 178118 529865 178170 529871
rect 177382 529719 177434 529725
rect 177382 529661 177434 529667
rect 177566 529719 177618 529725
rect 177566 529661 177618 529667
rect 177658 529719 177710 529725
rect 177658 529661 177710 529667
rect 177290 529243 177342 529249
rect 177290 529185 177342 529191
rect 177014 528563 177066 528569
rect 177014 528505 177066 528511
rect 176370 528291 176422 528297
rect 176370 528233 176422 528239
rect 176830 528291 176882 528297
rect 176830 528233 176882 528239
rect 176278 527815 176330 527821
rect 176278 527757 176330 527763
rect 177026 527685 177054 528505
rect 177394 528093 177422 529661
rect 177578 528773 177606 529661
rect 177934 529651 177986 529657
rect 177934 529593 177986 529599
rect 177946 529453 177974 529593
rect 177934 529447 177986 529453
rect 177934 529389 177986 529395
rect 177658 529311 177710 529317
rect 177658 529253 177710 529259
rect 177670 528909 177698 529253
rect 177783 529007 178091 529016
rect 177783 529005 177789 529007
rect 177845 529005 177869 529007
rect 177925 529005 177949 529007
rect 178005 529005 178029 529007
rect 178085 529005 178091 529007
rect 177845 528953 177847 529005
rect 178027 528953 178029 529005
rect 177783 528951 177789 528953
rect 177845 528951 177869 528953
rect 177925 528951 177949 528953
rect 178005 528951 178029 528953
rect 178085 528951 178091 528953
rect 177783 528942 178091 528951
rect 177658 528903 177710 528909
rect 177658 528845 177710 528851
rect 177566 528767 177618 528773
rect 177566 528709 177618 528715
rect 178026 528767 178078 528773
rect 178026 528709 178078 528715
rect 178038 528365 178066 528709
rect 178026 528359 178078 528365
rect 178026 528301 178078 528307
rect 178130 528229 178158 529865
rect 178222 528773 178250 529933
rect 178314 529385 178342 530137
rect 178443 529551 178751 529560
rect 178443 529549 178449 529551
rect 178505 529549 178529 529551
rect 178585 529549 178609 529551
rect 178665 529549 178689 529551
rect 178745 529549 178751 529551
rect 178505 529497 178507 529549
rect 178687 529497 178689 529549
rect 178443 529495 178449 529497
rect 178505 529495 178529 529497
rect 178585 529495 178609 529497
rect 178665 529495 178689 529497
rect 178745 529495 178751 529497
rect 178443 529486 178751 529495
rect 178302 529379 178354 529385
rect 178302 529321 178354 529327
rect 178210 528767 178262 528773
rect 178210 528709 178262 528715
rect 178314 528637 178434 528653
rect 178314 528631 178446 528637
rect 178314 528625 178394 528631
rect 178118 528223 178170 528229
rect 178118 528165 178170 528171
rect 177382 528087 177434 528093
rect 177382 528029 177434 528035
rect 177783 527919 178091 527928
rect 177783 527917 177789 527919
rect 177845 527917 177869 527919
rect 177925 527917 177949 527919
rect 178005 527917 178029 527919
rect 178085 527917 178091 527919
rect 177845 527865 177847 527917
rect 178027 527865 178029 527917
rect 177783 527863 177789 527865
rect 177845 527863 177869 527865
rect 177925 527863 177949 527865
rect 178005 527863 178029 527865
rect 178085 527863 178091 527865
rect 177783 527854 178091 527863
rect 177014 527679 177066 527685
rect 177014 527621 177066 527627
rect 174625 527375 174933 527384
rect 174625 527373 174631 527375
rect 174687 527373 174711 527375
rect 174767 527373 174791 527375
rect 174847 527373 174871 527375
rect 174927 527373 174933 527375
rect 174687 527321 174689 527373
rect 174869 527321 174871 527373
rect 174625 527319 174631 527321
rect 174687 527319 174711 527321
rect 174767 527319 174791 527321
rect 174847 527319 174871 527321
rect 174927 527319 174933 527321
rect 174625 527310 174933 527319
rect 173965 526831 174273 526840
rect 173965 526829 173971 526831
rect 174027 526829 174051 526831
rect 174107 526829 174131 526831
rect 174187 526829 174211 526831
rect 174267 526829 174273 526831
rect 174027 526777 174029 526829
rect 174209 526777 174211 526829
rect 173965 526775 173971 526777
rect 174027 526775 174051 526777
rect 174107 526775 174131 526777
rect 174187 526775 174211 526777
rect 174267 526775 174273 526777
rect 173965 526766 174273 526775
rect 177783 526831 178091 526840
rect 177783 526829 177789 526831
rect 177845 526829 177869 526831
rect 177925 526829 177949 526831
rect 178005 526829 178029 526831
rect 178085 526829 178091 526831
rect 177845 526777 177847 526829
rect 178027 526777 178029 526829
rect 177783 526775 177789 526777
rect 177845 526775 177869 526777
rect 177925 526775 177949 526777
rect 178005 526775 178029 526777
rect 178085 526775 178091 526777
rect 177783 526766 178091 526775
rect 174625 526287 174933 526296
rect 174625 526285 174631 526287
rect 174687 526285 174711 526287
rect 174767 526285 174791 526287
rect 174847 526285 174871 526287
rect 174927 526285 174933 526287
rect 174687 526233 174689 526285
rect 174869 526233 174871 526285
rect 174625 526231 174631 526233
rect 174687 526231 174711 526233
rect 174767 526231 174791 526233
rect 174847 526231 174871 526233
rect 174927 526231 174933 526233
rect 174625 526222 174933 526231
rect 173965 525743 174273 525752
rect 173965 525741 173971 525743
rect 174027 525741 174051 525743
rect 174107 525741 174131 525743
rect 174187 525741 174211 525743
rect 174267 525741 174273 525743
rect 174027 525689 174029 525741
rect 174209 525689 174211 525741
rect 173965 525687 173971 525689
rect 174027 525687 174051 525689
rect 174107 525687 174131 525689
rect 174187 525687 174211 525689
rect 174267 525687 174273 525689
rect 173965 525678 174273 525687
rect 177783 525743 178091 525752
rect 177783 525741 177789 525743
rect 177845 525741 177869 525743
rect 177925 525741 177949 525743
rect 178005 525741 178029 525743
rect 178085 525741 178091 525743
rect 177845 525689 177847 525741
rect 178027 525689 178029 525741
rect 177783 525687 177789 525689
rect 177845 525687 177869 525689
rect 177925 525687 177949 525689
rect 178005 525687 178029 525689
rect 178085 525687 178091 525689
rect 177783 525678 178091 525687
rect 174625 525199 174933 525208
rect 174625 525197 174631 525199
rect 174687 525197 174711 525199
rect 174767 525197 174791 525199
rect 174847 525197 174871 525199
rect 174927 525197 174933 525199
rect 174687 525145 174689 525197
rect 174869 525145 174871 525197
rect 174625 525143 174631 525145
rect 174687 525143 174711 525145
rect 174767 525143 174791 525145
rect 174847 525143 174871 525145
rect 174927 525143 174933 525145
rect 174625 525134 174933 525143
rect 173965 524655 174273 524664
rect 173965 524653 173971 524655
rect 174027 524653 174051 524655
rect 174107 524653 174131 524655
rect 174187 524653 174211 524655
rect 174267 524653 174273 524655
rect 174027 524601 174029 524653
rect 174209 524601 174211 524653
rect 173965 524599 173971 524601
rect 174027 524599 174051 524601
rect 174107 524599 174131 524601
rect 174187 524599 174211 524601
rect 174267 524599 174273 524601
rect 173965 524590 174273 524599
rect 177783 524655 178091 524664
rect 177783 524653 177789 524655
rect 177845 524653 177869 524655
rect 177925 524653 177949 524655
rect 178005 524653 178029 524655
rect 178085 524653 178091 524655
rect 177845 524601 177847 524653
rect 178027 524601 178029 524653
rect 177783 524599 177789 524601
rect 177845 524599 177869 524601
rect 177925 524599 177949 524601
rect 178005 524599 178029 524601
rect 178085 524599 178091 524601
rect 177783 524590 178091 524599
rect 174625 524111 174933 524120
rect 174625 524109 174631 524111
rect 174687 524109 174711 524111
rect 174767 524109 174791 524111
rect 174847 524109 174871 524111
rect 174927 524109 174933 524111
rect 174687 524057 174689 524109
rect 174869 524057 174871 524109
rect 174625 524055 174631 524057
rect 174687 524055 174711 524057
rect 174767 524055 174791 524057
rect 174847 524055 174871 524057
rect 174927 524055 174933 524057
rect 174625 524046 174933 524055
rect 173965 523567 174273 523576
rect 173965 523565 173971 523567
rect 174027 523565 174051 523567
rect 174107 523565 174131 523567
rect 174187 523565 174211 523567
rect 174267 523565 174273 523567
rect 174027 523513 174029 523565
rect 174209 523513 174211 523565
rect 173965 523511 173971 523513
rect 174027 523511 174051 523513
rect 174107 523511 174131 523513
rect 174187 523511 174211 523513
rect 174267 523511 174273 523513
rect 173965 523502 174273 523511
rect 177783 523567 178091 523576
rect 177783 523565 177789 523567
rect 177845 523565 177869 523567
rect 177925 523565 177949 523567
rect 178005 523565 178029 523567
rect 178085 523565 178091 523567
rect 177845 523513 177847 523565
rect 178027 523513 178029 523565
rect 177783 523511 177789 523513
rect 177845 523511 177869 523513
rect 177925 523511 177949 523513
rect 178005 523511 178029 523513
rect 178085 523511 178091 523513
rect 177783 523502 178091 523511
rect 174625 523023 174933 523032
rect 174625 523021 174631 523023
rect 174687 523021 174711 523023
rect 174767 523021 174791 523023
rect 174847 523021 174871 523023
rect 174927 523021 174933 523023
rect 174687 522969 174689 523021
rect 174869 522969 174871 523021
rect 174625 522967 174631 522969
rect 174687 522967 174711 522969
rect 174767 522967 174791 522969
rect 174847 522967 174871 522969
rect 174927 522967 174933 522969
rect 174625 522958 174933 522967
rect 173965 522479 174273 522488
rect 173965 522477 173971 522479
rect 174027 522477 174051 522479
rect 174107 522477 174131 522479
rect 174187 522477 174211 522479
rect 174267 522477 174273 522479
rect 174027 522425 174029 522477
rect 174209 522425 174211 522477
rect 173965 522423 173971 522425
rect 174027 522423 174051 522425
rect 174107 522423 174131 522425
rect 174187 522423 174211 522425
rect 174267 522423 174273 522425
rect 173965 522414 174273 522423
rect 177783 522479 178091 522488
rect 177783 522477 177789 522479
rect 177845 522477 177869 522479
rect 177925 522477 177949 522479
rect 178005 522477 178029 522479
rect 178085 522477 178091 522479
rect 177845 522425 177847 522477
rect 178027 522425 178029 522477
rect 177783 522423 177789 522425
rect 177845 522423 177869 522425
rect 177925 522423 177949 522425
rect 178005 522423 178029 522425
rect 178085 522423 178091 522425
rect 177783 522414 178091 522423
rect 174625 521935 174933 521944
rect 174625 521933 174631 521935
rect 174687 521933 174711 521935
rect 174767 521933 174791 521935
rect 174847 521933 174871 521935
rect 174927 521933 174933 521935
rect 174687 521881 174689 521933
rect 174869 521881 174871 521933
rect 174625 521879 174631 521881
rect 174687 521879 174711 521881
rect 174767 521879 174791 521881
rect 174847 521879 174871 521881
rect 174927 521879 174933 521881
rect 174625 521870 174933 521879
rect 173965 521391 174273 521400
rect 173965 521389 173971 521391
rect 174027 521389 174051 521391
rect 174107 521389 174131 521391
rect 174187 521389 174211 521391
rect 174267 521389 174273 521391
rect 174027 521337 174029 521389
rect 174209 521337 174211 521389
rect 173965 521335 173971 521337
rect 174027 521335 174051 521337
rect 174107 521335 174131 521337
rect 174187 521335 174211 521337
rect 174267 521335 174273 521337
rect 173965 521326 174273 521335
rect 177783 521391 178091 521400
rect 177783 521389 177789 521391
rect 177845 521389 177869 521391
rect 177925 521389 177949 521391
rect 178005 521389 178029 521391
rect 178085 521389 178091 521391
rect 177845 521337 177847 521389
rect 178027 521337 178029 521389
rect 177783 521335 177789 521337
rect 177845 521335 177869 521337
rect 177925 521335 177949 521337
rect 178005 521335 178029 521337
rect 178085 521335 178091 521337
rect 177783 521326 178091 521335
rect 174625 520847 174933 520856
rect 174625 520845 174631 520847
rect 174687 520845 174711 520847
rect 174767 520845 174791 520847
rect 174847 520845 174871 520847
rect 174927 520845 174933 520847
rect 174687 520793 174689 520845
rect 174869 520793 174871 520845
rect 174625 520791 174631 520793
rect 174687 520791 174711 520793
rect 174767 520791 174791 520793
rect 174847 520791 174871 520793
rect 174927 520791 174933 520793
rect 174625 520782 174933 520791
rect 173965 520303 174273 520312
rect 173965 520301 173971 520303
rect 174027 520301 174051 520303
rect 174107 520301 174131 520303
rect 174187 520301 174211 520303
rect 174267 520301 174273 520303
rect 174027 520249 174029 520301
rect 174209 520249 174211 520301
rect 173965 520247 173971 520249
rect 174027 520247 174051 520249
rect 174107 520247 174131 520249
rect 174187 520247 174211 520249
rect 174267 520247 174273 520249
rect 173965 520238 174273 520247
rect 177783 520303 178091 520312
rect 177783 520301 177789 520303
rect 177845 520301 177869 520303
rect 177925 520301 177949 520303
rect 178005 520301 178029 520303
rect 178085 520301 178091 520303
rect 177845 520249 177847 520301
rect 178027 520249 178029 520301
rect 177783 520247 177789 520249
rect 177845 520247 177869 520249
rect 177925 520247 177949 520249
rect 178005 520247 178029 520249
rect 178085 520247 178091 520249
rect 177783 520238 178091 520247
rect 174625 519759 174933 519768
rect 174625 519757 174631 519759
rect 174687 519757 174711 519759
rect 174767 519757 174791 519759
rect 174847 519757 174871 519759
rect 174927 519757 174933 519759
rect 174687 519705 174689 519757
rect 174869 519705 174871 519757
rect 174625 519703 174631 519705
rect 174687 519703 174711 519705
rect 174767 519703 174791 519705
rect 174847 519703 174871 519705
rect 174927 519703 174933 519705
rect 174625 519694 174933 519703
rect 173965 519215 174273 519224
rect 173965 519213 173971 519215
rect 174027 519213 174051 519215
rect 174107 519213 174131 519215
rect 174187 519213 174211 519215
rect 174267 519213 174273 519215
rect 174027 519161 174029 519213
rect 174209 519161 174211 519213
rect 173965 519159 173971 519161
rect 174027 519159 174051 519161
rect 174107 519159 174131 519161
rect 174187 519159 174211 519161
rect 174267 519159 174273 519161
rect 173965 519150 174273 519159
rect 177783 519215 178091 519224
rect 177783 519213 177789 519215
rect 177845 519213 177869 519215
rect 177925 519213 177949 519215
rect 178005 519213 178029 519215
rect 178085 519213 178091 519215
rect 177845 519161 177847 519213
rect 178027 519161 178029 519213
rect 177783 519159 177789 519161
rect 177845 519159 177869 519161
rect 177925 519159 177949 519161
rect 178005 519159 178029 519161
rect 178085 519159 178091 519161
rect 177783 519150 178091 519159
rect 174625 518671 174933 518680
rect 174625 518669 174631 518671
rect 174687 518669 174711 518671
rect 174767 518669 174791 518671
rect 174847 518669 174871 518671
rect 174927 518669 174933 518671
rect 174687 518617 174689 518669
rect 174869 518617 174871 518669
rect 174625 518615 174631 518617
rect 174687 518615 174711 518617
rect 174767 518615 174791 518617
rect 174847 518615 174871 518617
rect 174927 518615 174933 518617
rect 174625 518606 174933 518615
rect 173965 518127 174273 518136
rect 173965 518125 173971 518127
rect 174027 518125 174051 518127
rect 174107 518125 174131 518127
rect 174187 518125 174211 518127
rect 174267 518125 174273 518127
rect 174027 518073 174029 518125
rect 174209 518073 174211 518125
rect 173965 518071 173971 518073
rect 174027 518071 174051 518073
rect 174107 518071 174131 518073
rect 174187 518071 174211 518073
rect 174267 518071 174273 518073
rect 173965 518062 174273 518071
rect 177783 518127 178091 518136
rect 177783 518125 177789 518127
rect 177845 518125 177869 518127
rect 177925 518125 177949 518127
rect 178005 518125 178029 518127
rect 178085 518125 178091 518127
rect 177845 518073 177847 518125
rect 178027 518073 178029 518125
rect 177783 518071 177789 518073
rect 177845 518071 177869 518073
rect 177925 518071 177949 518073
rect 178005 518071 178029 518073
rect 178085 518071 178091 518073
rect 177783 518062 178091 518071
rect 174625 517583 174933 517592
rect 174625 517581 174631 517583
rect 174687 517581 174711 517583
rect 174767 517581 174791 517583
rect 174847 517581 174871 517583
rect 174927 517581 174933 517583
rect 174687 517529 174689 517581
rect 174869 517529 174871 517581
rect 174625 517527 174631 517529
rect 174687 517527 174711 517529
rect 174767 517527 174791 517529
rect 174847 517527 174871 517529
rect 174927 517527 174933 517529
rect 174625 517518 174933 517527
rect 178314 517485 178342 528625
rect 178394 528573 178446 528579
rect 178443 528463 178751 528472
rect 178443 528461 178449 528463
rect 178505 528461 178529 528463
rect 178585 528461 178609 528463
rect 178665 528461 178689 528463
rect 178745 528461 178751 528463
rect 178505 528409 178507 528461
rect 178687 528409 178689 528461
rect 178443 528407 178449 528409
rect 178505 528407 178529 528409
rect 178585 528407 178609 528409
rect 178665 528407 178689 528409
rect 178745 528407 178751 528409
rect 178443 528398 178751 528407
rect 178958 528365 178986 530341
rect 179234 530285 179262 530341
rect 179234 530257 179354 530285
rect 179326 529861 179354 530257
rect 179510 529997 179538 530477
rect 180694 530331 180746 530337
rect 180694 530273 180746 530279
rect 179682 530195 179734 530201
rect 179682 530137 179734 530143
rect 179498 529991 179550 529997
rect 179498 529933 179550 529939
rect 179314 529855 179366 529861
rect 179314 529797 179366 529803
rect 179326 529113 179354 529797
rect 179314 529107 179366 529113
rect 179314 529049 179366 529055
rect 179326 528365 179354 529049
rect 178946 528359 178998 528365
rect 178946 528301 178998 528307
rect 179314 528359 179366 528365
rect 179314 528301 179366 528307
rect 178946 528019 178998 528025
rect 178946 527961 178998 527967
rect 178958 527821 178986 527961
rect 178946 527815 178998 527821
rect 178946 527757 178998 527763
rect 179510 527685 179538 529933
rect 179694 529317 179722 530137
rect 179866 529855 179918 529861
rect 179866 529797 179918 529803
rect 179878 529453 179906 529797
rect 180510 529651 180562 529657
rect 180510 529593 180562 529599
rect 179866 529447 179918 529453
rect 179866 529389 179918 529395
rect 179682 529311 179734 529317
rect 179682 529253 179734 529259
rect 180522 529113 180550 529593
rect 179682 529107 179734 529113
rect 179682 529049 179734 529055
rect 180510 529107 180562 529113
rect 180510 529049 180562 529055
rect 179694 528909 179722 529049
rect 179682 528903 179734 528909
rect 179682 528845 179734 528851
rect 180522 528773 180550 529049
rect 180510 528767 180562 528773
rect 180510 528709 180562 528715
rect 180706 528161 180734 530273
rect 180890 529997 180918 531987
rect 182261 530639 182569 530648
rect 182261 530637 182267 530639
rect 182323 530637 182347 530639
rect 182403 530637 182427 530639
rect 182483 530637 182507 530639
rect 182563 530637 182569 530639
rect 182323 530585 182325 530637
rect 182505 530585 182507 530637
rect 182261 530583 182267 530585
rect 182323 530583 182347 530585
rect 182403 530583 182427 530585
rect 182483 530583 182507 530585
rect 182563 530583 182569 530585
rect 182261 530574 182569 530583
rect 183006 530541 183034 531987
rect 185122 530541 185150 531987
rect 187238 531509 187266 531987
rect 187146 531481 187266 531509
rect 186079 530639 186387 530648
rect 186079 530637 186085 530639
rect 186141 530637 186165 530639
rect 186221 530637 186245 530639
rect 186301 530637 186325 530639
rect 186381 530637 186387 530639
rect 186141 530585 186143 530637
rect 186323 530585 186325 530637
rect 186079 530583 186085 530585
rect 186141 530583 186165 530585
rect 186221 530583 186245 530585
rect 186301 530583 186325 530585
rect 186381 530583 186387 530585
rect 186079 530574 186387 530583
rect 182994 530535 183046 530541
rect 182994 530477 183046 530483
rect 185110 530535 185162 530541
rect 185110 530477 185162 530483
rect 187146 530405 187174 531481
rect 182258 530399 182310 530405
rect 182258 530341 182310 530347
rect 183178 530399 183230 530405
rect 183178 530341 183230 530347
rect 187134 530399 187186 530405
rect 187134 530341 187186 530347
rect 182166 530195 182218 530201
rect 182166 530137 182218 530143
rect 181601 530095 181909 530104
rect 181601 530093 181607 530095
rect 181663 530093 181687 530095
rect 181743 530093 181767 530095
rect 181823 530093 181847 530095
rect 181903 530093 181909 530095
rect 181663 530041 181665 530093
rect 181845 530041 181847 530093
rect 181601 530039 181607 530041
rect 181663 530039 181687 530041
rect 181743 530039 181767 530041
rect 181823 530039 181847 530041
rect 181903 530039 181909 530041
rect 181601 530030 181909 530039
rect 182178 529997 182206 530137
rect 180878 529991 180930 529997
rect 180878 529933 180930 529939
rect 182166 529991 182218 529997
rect 182166 529933 182218 529939
rect 181522 529719 181574 529725
rect 181522 529661 181574 529667
rect 181534 529317 181562 529661
rect 181798 529651 181850 529657
rect 182270 529639 182298 530341
rect 182626 530331 182678 530337
rect 182626 530273 182678 530279
rect 182638 529997 182666 530273
rect 182718 530195 182770 530201
rect 182718 530137 182770 530143
rect 182626 529991 182678 529997
rect 182626 529933 182678 529939
rect 181798 529593 181850 529599
rect 182178 529611 182298 529639
rect 181810 529453 181838 529593
rect 181798 529447 181850 529453
rect 181798 529389 181850 529395
rect 181522 529311 181574 529317
rect 181522 529253 181574 529259
rect 181534 528773 181562 529253
rect 181601 529007 181909 529016
rect 181601 529005 181607 529007
rect 181663 529005 181687 529007
rect 181743 529005 181767 529007
rect 181823 529005 181847 529007
rect 181903 529005 181909 529007
rect 181663 528953 181665 529005
rect 181845 528953 181847 529005
rect 181601 528951 181607 528953
rect 181663 528951 181687 528953
rect 181743 528951 181767 528953
rect 181823 528951 181847 528953
rect 181903 528951 181909 528953
rect 181601 528942 181909 528951
rect 182178 528909 182206 529611
rect 182261 529551 182569 529560
rect 182261 529549 182267 529551
rect 182323 529549 182347 529551
rect 182403 529549 182427 529551
rect 182483 529549 182507 529551
rect 182563 529549 182569 529551
rect 182323 529497 182325 529549
rect 182505 529497 182507 529549
rect 182261 529495 182267 529497
rect 182323 529495 182347 529497
rect 182403 529495 182427 529497
rect 182483 529495 182507 529497
rect 182563 529495 182569 529497
rect 182261 529486 182569 529495
rect 182730 529317 182758 530137
rect 183190 529861 183218 530341
rect 185419 530095 185727 530104
rect 185419 530093 185425 530095
rect 185481 530093 185505 530095
rect 185561 530093 185585 530095
rect 185641 530093 185665 530095
rect 185721 530093 185727 530095
rect 185481 530041 185483 530093
rect 185663 530041 185665 530093
rect 185419 530039 185425 530041
rect 185481 530039 185505 530041
rect 185561 530039 185585 530041
rect 185641 530039 185665 530041
rect 185721 530039 185727 530041
rect 185419 530030 185727 530039
rect 183178 529855 183230 529861
rect 183178 529797 183230 529803
rect 186079 529551 186387 529560
rect 186079 529549 186085 529551
rect 186141 529549 186165 529551
rect 186221 529549 186245 529551
rect 186301 529549 186325 529551
rect 186381 529549 186387 529551
rect 186141 529497 186143 529549
rect 186323 529497 186325 529549
rect 186079 529495 186085 529497
rect 186141 529495 186165 529497
rect 186221 529495 186245 529497
rect 186301 529495 186325 529497
rect 186381 529495 186387 529497
rect 186079 529486 186387 529495
rect 182718 529311 182770 529317
rect 182718 529253 182770 529259
rect 185419 529007 185727 529016
rect 185419 529005 185425 529007
rect 185481 529005 185505 529007
rect 185561 529005 185585 529007
rect 185641 529005 185665 529007
rect 185721 529005 185727 529007
rect 185481 528953 185483 529005
rect 185663 528953 185665 529005
rect 185419 528951 185425 528953
rect 185481 528951 185505 528953
rect 185561 528951 185585 528953
rect 185641 528951 185665 528953
rect 185721 528951 185727 528953
rect 185419 528942 185727 528951
rect 182166 528903 182218 528909
rect 182166 528845 182218 528851
rect 181522 528767 181574 528773
rect 181522 528709 181574 528715
rect 180970 528563 181022 528569
rect 180970 528505 181022 528511
rect 180982 528365 181010 528505
rect 182178 528365 182206 528845
rect 186582 528631 186634 528637
rect 186582 528573 186634 528579
rect 182261 528463 182569 528472
rect 182261 528461 182267 528463
rect 182323 528461 182347 528463
rect 182403 528461 182427 528463
rect 182483 528461 182507 528463
rect 182563 528461 182569 528463
rect 182323 528409 182325 528461
rect 182505 528409 182507 528461
rect 182261 528407 182267 528409
rect 182323 528407 182347 528409
rect 182403 528407 182427 528409
rect 182483 528407 182507 528409
rect 182563 528407 182569 528409
rect 182261 528398 182569 528407
rect 186079 528463 186387 528472
rect 186079 528461 186085 528463
rect 186141 528461 186165 528463
rect 186221 528461 186245 528463
rect 186301 528461 186325 528463
rect 186381 528461 186387 528463
rect 186141 528409 186143 528461
rect 186323 528409 186325 528461
rect 186079 528407 186085 528409
rect 186141 528407 186165 528409
rect 186221 528407 186245 528409
rect 186301 528407 186325 528409
rect 186381 528407 186387 528409
rect 186079 528398 186387 528407
rect 180970 528359 181022 528365
rect 180970 528301 181022 528307
rect 182166 528359 182218 528365
rect 182166 528301 182218 528307
rect 181338 528223 181390 528229
rect 181338 528165 181390 528171
rect 180694 528155 180746 528161
rect 180694 528097 180746 528103
rect 179498 527679 179550 527685
rect 179498 527621 179550 527627
rect 178443 527375 178751 527384
rect 178443 527373 178449 527375
rect 178505 527373 178529 527375
rect 178585 527373 178609 527375
rect 178665 527373 178689 527375
rect 178745 527373 178751 527375
rect 178505 527321 178507 527373
rect 178687 527321 178689 527373
rect 178443 527319 178449 527321
rect 178505 527319 178529 527321
rect 178585 527319 178609 527321
rect 178665 527319 178689 527321
rect 178745 527319 178751 527321
rect 178443 527310 178751 527319
rect 178443 526287 178751 526296
rect 178443 526285 178449 526287
rect 178505 526285 178529 526287
rect 178585 526285 178609 526287
rect 178665 526285 178689 526287
rect 178745 526285 178751 526287
rect 178505 526233 178507 526285
rect 178687 526233 178689 526285
rect 178443 526231 178449 526233
rect 178505 526231 178529 526233
rect 178585 526231 178609 526233
rect 178665 526231 178689 526233
rect 178745 526231 178751 526233
rect 178443 526222 178751 526231
rect 178443 525199 178751 525208
rect 178443 525197 178449 525199
rect 178505 525197 178529 525199
rect 178585 525197 178609 525199
rect 178665 525197 178689 525199
rect 178745 525197 178751 525199
rect 178505 525145 178507 525197
rect 178687 525145 178689 525197
rect 178443 525143 178449 525145
rect 178505 525143 178529 525145
rect 178585 525143 178609 525145
rect 178665 525143 178689 525145
rect 178745 525143 178751 525145
rect 178443 525134 178751 525143
rect 178443 524111 178751 524120
rect 178443 524109 178449 524111
rect 178505 524109 178529 524111
rect 178585 524109 178609 524111
rect 178665 524109 178689 524111
rect 178745 524109 178751 524111
rect 178505 524057 178507 524109
rect 178687 524057 178689 524109
rect 178443 524055 178449 524057
rect 178505 524055 178529 524057
rect 178585 524055 178609 524057
rect 178665 524055 178689 524057
rect 178745 524055 178751 524057
rect 178443 524046 178751 524055
rect 178443 523023 178751 523032
rect 178443 523021 178449 523023
rect 178505 523021 178529 523023
rect 178585 523021 178609 523023
rect 178665 523021 178689 523023
rect 178745 523021 178751 523023
rect 178505 522969 178507 523021
rect 178687 522969 178689 523021
rect 178443 522967 178449 522969
rect 178505 522967 178529 522969
rect 178585 522967 178609 522969
rect 178665 522967 178689 522969
rect 178745 522967 178751 522969
rect 178443 522958 178751 522967
rect 178443 521935 178751 521944
rect 178443 521933 178449 521935
rect 178505 521933 178529 521935
rect 178585 521933 178609 521935
rect 178665 521933 178689 521935
rect 178745 521933 178751 521935
rect 178505 521881 178507 521933
rect 178687 521881 178689 521933
rect 178443 521879 178449 521881
rect 178505 521879 178529 521881
rect 178585 521879 178609 521881
rect 178665 521879 178689 521881
rect 178745 521879 178751 521881
rect 178443 521870 178751 521879
rect 178443 520847 178751 520856
rect 178443 520845 178449 520847
rect 178505 520845 178529 520847
rect 178585 520845 178609 520847
rect 178665 520845 178689 520847
rect 178745 520845 178751 520847
rect 178505 520793 178507 520845
rect 178687 520793 178689 520845
rect 178443 520791 178449 520793
rect 178505 520791 178529 520793
rect 178585 520791 178609 520793
rect 178665 520791 178689 520793
rect 178745 520791 178751 520793
rect 178443 520782 178751 520791
rect 178443 519759 178751 519768
rect 178443 519757 178449 519759
rect 178505 519757 178529 519759
rect 178585 519757 178609 519759
rect 178665 519757 178689 519759
rect 178745 519757 178751 519759
rect 178505 519705 178507 519757
rect 178687 519705 178689 519757
rect 178443 519703 178449 519705
rect 178505 519703 178529 519705
rect 178585 519703 178609 519705
rect 178665 519703 178689 519705
rect 178745 519703 178751 519705
rect 178443 519694 178751 519703
rect 178443 518671 178751 518680
rect 178443 518669 178449 518671
rect 178505 518669 178529 518671
rect 178585 518669 178609 518671
rect 178665 518669 178689 518671
rect 178745 518669 178751 518671
rect 178505 518617 178507 518669
rect 178687 518617 178689 518669
rect 178443 518615 178449 518617
rect 178505 518615 178529 518617
rect 178585 518615 178609 518617
rect 178665 518615 178689 518617
rect 178745 518615 178751 518617
rect 178443 518606 178751 518615
rect 178443 517583 178751 517592
rect 178443 517581 178449 517583
rect 178505 517581 178529 517583
rect 178585 517581 178609 517583
rect 178665 517581 178689 517583
rect 178745 517581 178751 517583
rect 178505 517529 178507 517581
rect 178687 517529 178689 517581
rect 178443 517527 178449 517529
rect 178505 517527 178529 517529
rect 178585 517527 178609 517529
rect 178665 517527 178689 517529
rect 178745 517527 178751 517529
rect 178443 517518 178751 517527
rect 177658 517479 177710 517485
rect 177658 517421 177710 517427
rect 178302 517479 178354 517485
rect 178302 517421 178354 517427
rect 173965 517039 174273 517048
rect 173965 517037 173971 517039
rect 174027 517037 174051 517039
rect 174107 517037 174131 517039
rect 174187 517037 174211 517039
rect 174267 517037 174273 517039
rect 174027 516985 174029 517037
rect 174209 516985 174211 517037
rect 173965 516983 173971 516985
rect 174027 516983 174051 516985
rect 174107 516983 174131 516985
rect 174187 516983 174211 516985
rect 174267 516983 174273 516985
rect 173965 516974 174273 516983
rect 174625 516495 174933 516504
rect 174625 516493 174631 516495
rect 174687 516493 174711 516495
rect 174767 516493 174791 516495
rect 174847 516493 174871 516495
rect 174927 516493 174933 516495
rect 174687 516441 174689 516493
rect 174869 516441 174871 516493
rect 174625 516439 174631 516441
rect 174687 516439 174711 516441
rect 174767 516439 174791 516441
rect 174847 516439 174871 516441
rect 174927 516439 174933 516441
rect 174625 516430 174933 516439
rect 173965 515951 174273 515960
rect 173965 515949 173971 515951
rect 174027 515949 174051 515951
rect 174107 515949 174131 515951
rect 174187 515949 174211 515951
rect 174267 515949 174273 515951
rect 174027 515897 174029 515949
rect 174209 515897 174211 515949
rect 173965 515895 173971 515897
rect 174027 515895 174051 515897
rect 174107 515895 174131 515897
rect 174187 515895 174211 515897
rect 174267 515895 174273 515897
rect 173965 515886 174273 515895
rect 173610 515847 173662 515853
rect 173610 515789 173662 515795
rect 173334 515575 173386 515581
rect 173334 515517 173386 515523
rect 173346 513931 173374 515517
rect 174625 515407 174933 515416
rect 174625 515405 174631 515407
rect 174687 515405 174711 515407
rect 174767 515405 174791 515407
rect 174847 515405 174871 515407
rect 174927 515405 174933 515407
rect 174687 515353 174689 515405
rect 174869 515353 174871 515405
rect 174625 515351 174631 515353
rect 174687 515351 174711 515353
rect 174767 515351 174791 515353
rect 174847 515351 174871 515353
rect 174927 515351 174933 515353
rect 174625 515342 174933 515351
rect 177670 513931 177698 517421
rect 177783 517039 178091 517048
rect 177783 517037 177789 517039
rect 177845 517037 177869 517039
rect 177925 517037 177949 517039
rect 178005 517037 178029 517039
rect 178085 517037 178091 517039
rect 177845 516985 177847 517037
rect 178027 516985 178029 517037
rect 177783 516983 177789 516985
rect 177845 516983 177869 516985
rect 177925 516983 177949 516985
rect 178005 516983 178029 516985
rect 178085 516983 178091 516985
rect 177783 516974 178091 516983
rect 178443 516495 178751 516504
rect 178443 516493 178449 516495
rect 178505 516493 178529 516495
rect 178585 516493 178609 516495
rect 178665 516493 178689 516495
rect 178745 516493 178751 516495
rect 178505 516441 178507 516493
rect 178687 516441 178689 516493
rect 178443 516439 178449 516441
rect 178505 516439 178529 516441
rect 178585 516439 178609 516441
rect 178665 516439 178689 516441
rect 178745 516439 178751 516441
rect 178443 516430 178751 516439
rect 177783 515951 178091 515960
rect 177783 515949 177789 515951
rect 177845 515949 177869 515951
rect 177925 515949 177949 515951
rect 178005 515949 178029 515951
rect 178085 515949 178091 515951
rect 177845 515897 177847 515949
rect 178027 515897 178029 515949
rect 177783 515895 177789 515897
rect 177845 515895 177869 515897
rect 177925 515895 177949 515897
rect 178005 515895 178029 515897
rect 178085 515895 178091 515897
rect 177783 515886 178091 515895
rect 181350 515853 181378 528165
rect 181601 527919 181909 527928
rect 181601 527917 181607 527919
rect 181663 527917 181687 527919
rect 181743 527917 181767 527919
rect 181823 527917 181847 527919
rect 181903 527917 181909 527919
rect 181663 527865 181665 527917
rect 181845 527865 181847 527917
rect 181601 527863 181607 527865
rect 181663 527863 181687 527865
rect 181743 527863 181767 527865
rect 181823 527863 181847 527865
rect 181903 527863 181909 527865
rect 181601 527854 181909 527863
rect 185419 527919 185727 527928
rect 185419 527917 185425 527919
rect 185481 527917 185505 527919
rect 185561 527917 185585 527919
rect 185641 527917 185665 527919
rect 185721 527917 185727 527919
rect 185481 527865 185483 527917
rect 185663 527865 185665 527917
rect 185419 527863 185425 527865
rect 185481 527863 185505 527865
rect 185561 527863 185585 527865
rect 185641 527863 185665 527865
rect 185721 527863 185727 527865
rect 185419 527854 185727 527863
rect 182261 527375 182569 527384
rect 182261 527373 182267 527375
rect 182323 527373 182347 527375
rect 182403 527373 182427 527375
rect 182483 527373 182507 527375
rect 182563 527373 182569 527375
rect 182323 527321 182325 527373
rect 182505 527321 182507 527373
rect 182261 527319 182267 527321
rect 182323 527319 182347 527321
rect 182403 527319 182427 527321
rect 182483 527319 182507 527321
rect 182563 527319 182569 527321
rect 182261 527310 182569 527319
rect 186079 527375 186387 527384
rect 186079 527373 186085 527375
rect 186141 527373 186165 527375
rect 186221 527373 186245 527375
rect 186301 527373 186325 527375
rect 186381 527373 186387 527375
rect 186141 527321 186143 527373
rect 186323 527321 186325 527373
rect 186079 527319 186085 527321
rect 186141 527319 186165 527321
rect 186221 527319 186245 527321
rect 186301 527319 186325 527321
rect 186381 527319 186387 527321
rect 186079 527310 186387 527319
rect 181601 526831 181909 526840
rect 181601 526829 181607 526831
rect 181663 526829 181687 526831
rect 181743 526829 181767 526831
rect 181823 526829 181847 526831
rect 181903 526829 181909 526831
rect 181663 526777 181665 526829
rect 181845 526777 181847 526829
rect 181601 526775 181607 526777
rect 181663 526775 181687 526777
rect 181743 526775 181767 526777
rect 181823 526775 181847 526777
rect 181903 526775 181909 526777
rect 181601 526766 181909 526775
rect 185419 526831 185727 526840
rect 185419 526829 185425 526831
rect 185481 526829 185505 526831
rect 185561 526829 185585 526831
rect 185641 526829 185665 526831
rect 185721 526829 185727 526831
rect 185481 526777 185483 526829
rect 185663 526777 185665 526829
rect 185419 526775 185425 526777
rect 185481 526775 185505 526777
rect 185561 526775 185585 526777
rect 185641 526775 185665 526777
rect 185721 526775 185727 526777
rect 185419 526766 185727 526775
rect 182261 526287 182569 526296
rect 182261 526285 182267 526287
rect 182323 526285 182347 526287
rect 182403 526285 182427 526287
rect 182483 526285 182507 526287
rect 182563 526285 182569 526287
rect 182323 526233 182325 526285
rect 182505 526233 182507 526285
rect 182261 526231 182267 526233
rect 182323 526231 182347 526233
rect 182403 526231 182427 526233
rect 182483 526231 182507 526233
rect 182563 526231 182569 526233
rect 182261 526222 182569 526231
rect 186079 526287 186387 526296
rect 186079 526285 186085 526287
rect 186141 526285 186165 526287
rect 186221 526285 186245 526287
rect 186301 526285 186325 526287
rect 186381 526285 186387 526287
rect 186141 526233 186143 526285
rect 186323 526233 186325 526285
rect 186079 526231 186085 526233
rect 186141 526231 186165 526233
rect 186221 526231 186245 526233
rect 186301 526231 186325 526233
rect 186381 526231 186387 526233
rect 186079 526222 186387 526231
rect 181601 525743 181909 525752
rect 181601 525741 181607 525743
rect 181663 525741 181687 525743
rect 181743 525741 181767 525743
rect 181823 525741 181847 525743
rect 181903 525741 181909 525743
rect 181663 525689 181665 525741
rect 181845 525689 181847 525741
rect 181601 525687 181607 525689
rect 181663 525687 181687 525689
rect 181743 525687 181767 525689
rect 181823 525687 181847 525689
rect 181903 525687 181909 525689
rect 181601 525678 181909 525687
rect 185419 525743 185727 525752
rect 185419 525741 185425 525743
rect 185481 525741 185505 525743
rect 185561 525741 185585 525743
rect 185641 525741 185665 525743
rect 185721 525741 185727 525743
rect 185481 525689 185483 525741
rect 185663 525689 185665 525741
rect 185419 525687 185425 525689
rect 185481 525687 185505 525689
rect 185561 525687 185585 525689
rect 185641 525687 185665 525689
rect 185721 525687 185727 525689
rect 185419 525678 185727 525687
rect 182261 525199 182569 525208
rect 182261 525197 182267 525199
rect 182323 525197 182347 525199
rect 182403 525197 182427 525199
rect 182483 525197 182507 525199
rect 182563 525197 182569 525199
rect 182323 525145 182325 525197
rect 182505 525145 182507 525197
rect 182261 525143 182267 525145
rect 182323 525143 182347 525145
rect 182403 525143 182427 525145
rect 182483 525143 182507 525145
rect 182563 525143 182569 525145
rect 182261 525134 182569 525143
rect 186079 525199 186387 525208
rect 186079 525197 186085 525199
rect 186141 525197 186165 525199
rect 186221 525197 186245 525199
rect 186301 525197 186325 525199
rect 186381 525197 186387 525199
rect 186141 525145 186143 525197
rect 186323 525145 186325 525197
rect 186079 525143 186085 525145
rect 186141 525143 186165 525145
rect 186221 525143 186245 525145
rect 186301 525143 186325 525145
rect 186381 525143 186387 525145
rect 186079 525134 186387 525143
rect 181601 524655 181909 524664
rect 181601 524653 181607 524655
rect 181663 524653 181687 524655
rect 181743 524653 181767 524655
rect 181823 524653 181847 524655
rect 181903 524653 181909 524655
rect 181663 524601 181665 524653
rect 181845 524601 181847 524653
rect 181601 524599 181607 524601
rect 181663 524599 181687 524601
rect 181743 524599 181767 524601
rect 181823 524599 181847 524601
rect 181903 524599 181909 524601
rect 181601 524590 181909 524599
rect 185419 524655 185727 524664
rect 185419 524653 185425 524655
rect 185481 524653 185505 524655
rect 185561 524653 185585 524655
rect 185641 524653 185665 524655
rect 185721 524653 185727 524655
rect 185481 524601 185483 524653
rect 185663 524601 185665 524653
rect 185419 524599 185425 524601
rect 185481 524599 185505 524601
rect 185561 524599 185585 524601
rect 185641 524599 185665 524601
rect 185721 524599 185727 524601
rect 185419 524590 185727 524599
rect 182261 524111 182569 524120
rect 182261 524109 182267 524111
rect 182323 524109 182347 524111
rect 182403 524109 182427 524111
rect 182483 524109 182507 524111
rect 182563 524109 182569 524111
rect 182323 524057 182325 524109
rect 182505 524057 182507 524109
rect 182261 524055 182267 524057
rect 182323 524055 182347 524057
rect 182403 524055 182427 524057
rect 182483 524055 182507 524057
rect 182563 524055 182569 524057
rect 182261 524046 182569 524055
rect 186079 524111 186387 524120
rect 186079 524109 186085 524111
rect 186141 524109 186165 524111
rect 186221 524109 186245 524111
rect 186301 524109 186325 524111
rect 186381 524109 186387 524111
rect 186141 524057 186143 524109
rect 186323 524057 186325 524109
rect 186079 524055 186085 524057
rect 186141 524055 186165 524057
rect 186221 524055 186245 524057
rect 186301 524055 186325 524057
rect 186381 524055 186387 524057
rect 186079 524046 186387 524055
rect 181601 523567 181909 523576
rect 181601 523565 181607 523567
rect 181663 523565 181687 523567
rect 181743 523565 181767 523567
rect 181823 523565 181847 523567
rect 181903 523565 181909 523567
rect 181663 523513 181665 523565
rect 181845 523513 181847 523565
rect 181601 523511 181607 523513
rect 181663 523511 181687 523513
rect 181743 523511 181767 523513
rect 181823 523511 181847 523513
rect 181903 523511 181909 523513
rect 181601 523502 181909 523511
rect 185419 523567 185727 523576
rect 185419 523565 185425 523567
rect 185481 523565 185505 523567
rect 185561 523565 185585 523567
rect 185641 523565 185665 523567
rect 185721 523565 185727 523567
rect 185481 523513 185483 523565
rect 185663 523513 185665 523565
rect 185419 523511 185425 523513
rect 185481 523511 185505 523513
rect 185561 523511 185585 523513
rect 185641 523511 185665 523513
rect 185721 523511 185727 523513
rect 185419 523502 185727 523511
rect 182261 523023 182569 523032
rect 182261 523021 182267 523023
rect 182323 523021 182347 523023
rect 182403 523021 182427 523023
rect 182483 523021 182507 523023
rect 182563 523021 182569 523023
rect 182323 522969 182325 523021
rect 182505 522969 182507 523021
rect 182261 522967 182267 522969
rect 182323 522967 182347 522969
rect 182403 522967 182427 522969
rect 182483 522967 182507 522969
rect 182563 522967 182569 522969
rect 182261 522958 182569 522967
rect 186079 523023 186387 523032
rect 186079 523021 186085 523023
rect 186141 523021 186165 523023
rect 186221 523021 186245 523023
rect 186301 523021 186325 523023
rect 186381 523021 186387 523023
rect 186141 522969 186143 523021
rect 186323 522969 186325 523021
rect 186079 522967 186085 522969
rect 186141 522967 186165 522969
rect 186221 522967 186245 522969
rect 186301 522967 186325 522969
rect 186381 522967 186387 522969
rect 186079 522958 186387 522967
rect 181601 522479 181909 522488
rect 181601 522477 181607 522479
rect 181663 522477 181687 522479
rect 181743 522477 181767 522479
rect 181823 522477 181847 522479
rect 181903 522477 181909 522479
rect 181663 522425 181665 522477
rect 181845 522425 181847 522477
rect 181601 522423 181607 522425
rect 181663 522423 181687 522425
rect 181743 522423 181767 522425
rect 181823 522423 181847 522425
rect 181903 522423 181909 522425
rect 181601 522414 181909 522423
rect 185419 522479 185727 522488
rect 185419 522477 185425 522479
rect 185481 522477 185505 522479
rect 185561 522477 185585 522479
rect 185641 522477 185665 522479
rect 185721 522477 185727 522479
rect 185481 522425 185483 522477
rect 185663 522425 185665 522477
rect 185419 522423 185425 522425
rect 185481 522423 185505 522425
rect 185561 522423 185585 522425
rect 185641 522423 185665 522425
rect 185721 522423 185727 522425
rect 185419 522414 185727 522423
rect 182261 521935 182569 521944
rect 182261 521933 182267 521935
rect 182323 521933 182347 521935
rect 182403 521933 182427 521935
rect 182483 521933 182507 521935
rect 182563 521933 182569 521935
rect 182323 521881 182325 521933
rect 182505 521881 182507 521933
rect 182261 521879 182267 521881
rect 182323 521879 182347 521881
rect 182403 521879 182427 521881
rect 182483 521879 182507 521881
rect 182563 521879 182569 521881
rect 182261 521870 182569 521879
rect 186079 521935 186387 521944
rect 186079 521933 186085 521935
rect 186141 521933 186165 521935
rect 186221 521933 186245 521935
rect 186301 521933 186325 521935
rect 186381 521933 186387 521935
rect 186141 521881 186143 521933
rect 186323 521881 186325 521933
rect 186079 521879 186085 521881
rect 186141 521879 186165 521881
rect 186221 521879 186245 521881
rect 186301 521879 186325 521881
rect 186381 521879 186387 521881
rect 186079 521870 186387 521879
rect 181601 521391 181909 521400
rect 181601 521389 181607 521391
rect 181663 521389 181687 521391
rect 181743 521389 181767 521391
rect 181823 521389 181847 521391
rect 181903 521389 181909 521391
rect 181663 521337 181665 521389
rect 181845 521337 181847 521389
rect 181601 521335 181607 521337
rect 181663 521335 181687 521337
rect 181743 521335 181767 521337
rect 181823 521335 181847 521337
rect 181903 521335 181909 521337
rect 181601 521326 181909 521335
rect 185419 521391 185727 521400
rect 185419 521389 185425 521391
rect 185481 521389 185505 521391
rect 185561 521389 185585 521391
rect 185641 521389 185665 521391
rect 185721 521389 185727 521391
rect 185481 521337 185483 521389
rect 185663 521337 185665 521389
rect 185419 521335 185425 521337
rect 185481 521335 185505 521337
rect 185561 521335 185585 521337
rect 185641 521335 185665 521337
rect 185721 521335 185727 521337
rect 185419 521326 185727 521335
rect 182261 520847 182569 520856
rect 182261 520845 182267 520847
rect 182323 520845 182347 520847
rect 182403 520845 182427 520847
rect 182483 520845 182507 520847
rect 182563 520845 182569 520847
rect 182323 520793 182325 520845
rect 182505 520793 182507 520845
rect 182261 520791 182267 520793
rect 182323 520791 182347 520793
rect 182403 520791 182427 520793
rect 182483 520791 182507 520793
rect 182563 520791 182569 520793
rect 182261 520782 182569 520791
rect 186079 520847 186387 520856
rect 186079 520845 186085 520847
rect 186141 520845 186165 520847
rect 186221 520845 186245 520847
rect 186301 520845 186325 520847
rect 186381 520845 186387 520847
rect 186141 520793 186143 520845
rect 186323 520793 186325 520845
rect 186079 520791 186085 520793
rect 186141 520791 186165 520793
rect 186221 520791 186245 520793
rect 186301 520791 186325 520793
rect 186381 520791 186387 520793
rect 186079 520782 186387 520791
rect 181601 520303 181909 520312
rect 181601 520301 181607 520303
rect 181663 520301 181687 520303
rect 181743 520301 181767 520303
rect 181823 520301 181847 520303
rect 181903 520301 181909 520303
rect 181663 520249 181665 520301
rect 181845 520249 181847 520301
rect 181601 520247 181607 520249
rect 181663 520247 181687 520249
rect 181743 520247 181767 520249
rect 181823 520247 181847 520249
rect 181903 520247 181909 520249
rect 181601 520238 181909 520247
rect 185419 520303 185727 520312
rect 185419 520301 185425 520303
rect 185481 520301 185505 520303
rect 185561 520301 185585 520303
rect 185641 520301 185665 520303
rect 185721 520301 185727 520303
rect 185481 520249 185483 520301
rect 185663 520249 185665 520301
rect 185419 520247 185425 520249
rect 185481 520247 185505 520249
rect 185561 520247 185585 520249
rect 185641 520247 185665 520249
rect 185721 520247 185727 520249
rect 185419 520238 185727 520247
rect 182261 519759 182569 519768
rect 182261 519757 182267 519759
rect 182323 519757 182347 519759
rect 182403 519757 182427 519759
rect 182483 519757 182507 519759
rect 182563 519757 182569 519759
rect 182323 519705 182325 519757
rect 182505 519705 182507 519757
rect 182261 519703 182267 519705
rect 182323 519703 182347 519705
rect 182403 519703 182427 519705
rect 182483 519703 182507 519705
rect 182563 519703 182569 519705
rect 182261 519694 182569 519703
rect 186079 519759 186387 519768
rect 186079 519757 186085 519759
rect 186141 519757 186165 519759
rect 186221 519757 186245 519759
rect 186301 519757 186325 519759
rect 186381 519757 186387 519759
rect 186141 519705 186143 519757
rect 186323 519705 186325 519757
rect 186079 519703 186085 519705
rect 186141 519703 186165 519705
rect 186221 519703 186245 519705
rect 186301 519703 186325 519705
rect 186381 519703 186387 519705
rect 186079 519694 186387 519703
rect 181601 519215 181909 519224
rect 181601 519213 181607 519215
rect 181663 519213 181687 519215
rect 181743 519213 181767 519215
rect 181823 519213 181847 519215
rect 181903 519213 181909 519215
rect 181663 519161 181665 519213
rect 181845 519161 181847 519213
rect 181601 519159 181607 519161
rect 181663 519159 181687 519161
rect 181743 519159 181767 519161
rect 181823 519159 181847 519161
rect 181903 519159 181909 519161
rect 181601 519150 181909 519159
rect 185419 519215 185727 519224
rect 185419 519213 185425 519215
rect 185481 519213 185505 519215
rect 185561 519213 185585 519215
rect 185641 519213 185665 519215
rect 185721 519213 185727 519215
rect 185481 519161 185483 519213
rect 185663 519161 185665 519213
rect 185419 519159 185425 519161
rect 185481 519159 185505 519161
rect 185561 519159 185585 519161
rect 185641 519159 185665 519161
rect 185721 519159 185727 519161
rect 185419 519150 185727 519159
rect 182261 518671 182569 518680
rect 182261 518669 182267 518671
rect 182323 518669 182347 518671
rect 182403 518669 182427 518671
rect 182483 518669 182507 518671
rect 182563 518669 182569 518671
rect 182323 518617 182325 518669
rect 182505 518617 182507 518669
rect 182261 518615 182267 518617
rect 182323 518615 182347 518617
rect 182403 518615 182427 518617
rect 182483 518615 182507 518617
rect 182563 518615 182569 518617
rect 182261 518606 182569 518615
rect 186079 518671 186387 518680
rect 186079 518669 186085 518671
rect 186141 518669 186165 518671
rect 186221 518669 186245 518671
rect 186301 518669 186325 518671
rect 186381 518669 186387 518671
rect 186141 518617 186143 518669
rect 186323 518617 186325 518669
rect 186079 518615 186085 518617
rect 186141 518615 186165 518617
rect 186221 518615 186245 518617
rect 186301 518615 186325 518617
rect 186381 518615 186387 518617
rect 186079 518606 186387 518615
rect 181601 518127 181909 518136
rect 181601 518125 181607 518127
rect 181663 518125 181687 518127
rect 181743 518125 181767 518127
rect 181823 518125 181847 518127
rect 181903 518125 181909 518127
rect 181663 518073 181665 518125
rect 181845 518073 181847 518125
rect 181601 518071 181607 518073
rect 181663 518071 181687 518073
rect 181743 518071 181767 518073
rect 181823 518071 181847 518073
rect 181903 518071 181909 518073
rect 181601 518062 181909 518071
rect 185419 518127 185727 518136
rect 185419 518125 185425 518127
rect 185481 518125 185505 518127
rect 185561 518125 185585 518127
rect 185641 518125 185665 518127
rect 185721 518125 185727 518127
rect 185481 518073 185483 518125
rect 185663 518073 185665 518125
rect 185419 518071 185425 518073
rect 185481 518071 185505 518073
rect 185561 518071 185585 518073
rect 185641 518071 185665 518073
rect 185721 518071 185727 518073
rect 185419 518062 185727 518071
rect 182261 517583 182569 517592
rect 182261 517581 182267 517583
rect 182323 517581 182347 517583
rect 182403 517581 182427 517583
rect 182483 517581 182507 517583
rect 182563 517581 182569 517583
rect 182323 517529 182325 517581
rect 182505 517529 182507 517581
rect 182261 517527 182267 517529
rect 182323 517527 182347 517529
rect 182403 517527 182427 517529
rect 182483 517527 182507 517529
rect 182563 517527 182569 517529
rect 182261 517518 182569 517527
rect 186079 517583 186387 517592
rect 186079 517581 186085 517583
rect 186141 517581 186165 517583
rect 186221 517581 186245 517583
rect 186301 517581 186325 517583
rect 186381 517581 186387 517583
rect 186141 517529 186143 517581
rect 186323 517529 186325 517581
rect 186079 517527 186085 517529
rect 186141 517527 186165 517529
rect 186221 517527 186245 517529
rect 186301 517527 186325 517529
rect 186381 517527 186387 517529
rect 186079 517518 186387 517527
rect 181601 517039 181909 517048
rect 181601 517037 181607 517039
rect 181663 517037 181687 517039
rect 181743 517037 181767 517039
rect 181823 517037 181847 517039
rect 181903 517037 181909 517039
rect 181663 516985 181665 517037
rect 181845 516985 181847 517037
rect 181601 516983 181607 516985
rect 181663 516983 181687 516985
rect 181743 516983 181767 516985
rect 181823 516983 181847 516985
rect 181903 516983 181909 516985
rect 181601 516974 181909 516983
rect 185419 517039 185727 517048
rect 185419 517037 185425 517039
rect 185481 517037 185505 517039
rect 185561 517037 185585 517039
rect 185641 517037 185665 517039
rect 185721 517037 185727 517039
rect 185481 516985 185483 517037
rect 185663 516985 185665 517037
rect 185419 516983 185425 516985
rect 185481 516983 185505 516985
rect 185561 516983 185585 516985
rect 185641 516983 185665 516985
rect 185721 516983 185727 516985
rect 185419 516974 185727 516983
rect 182261 516495 182569 516504
rect 182261 516493 182267 516495
rect 182323 516493 182347 516495
rect 182403 516493 182427 516495
rect 182483 516493 182507 516495
rect 182563 516493 182569 516495
rect 182323 516441 182325 516493
rect 182505 516441 182507 516493
rect 182261 516439 182267 516441
rect 182323 516439 182347 516441
rect 182403 516439 182427 516441
rect 182483 516439 182507 516441
rect 182563 516439 182569 516441
rect 182261 516430 182569 516439
rect 186079 516495 186387 516504
rect 186079 516493 186085 516495
rect 186141 516493 186165 516495
rect 186221 516493 186245 516495
rect 186301 516493 186325 516495
rect 186381 516493 186387 516495
rect 186141 516441 186143 516493
rect 186323 516441 186325 516493
rect 186079 516439 186085 516441
rect 186141 516439 186165 516441
rect 186221 516439 186245 516441
rect 186301 516439 186325 516441
rect 186381 516439 186387 516441
rect 186079 516430 186387 516439
rect 181601 515951 181909 515960
rect 181601 515949 181607 515951
rect 181663 515949 181687 515951
rect 181743 515949 181767 515951
rect 181823 515949 181847 515951
rect 181903 515949 181909 515951
rect 181663 515897 181665 515949
rect 181845 515897 181847 515949
rect 181601 515895 181607 515897
rect 181663 515895 181687 515897
rect 181743 515895 181767 515897
rect 181823 515895 181847 515897
rect 181903 515895 181909 515897
rect 181601 515886 181909 515895
rect 185419 515951 185727 515960
rect 185419 515949 185425 515951
rect 185481 515949 185505 515951
rect 185561 515949 185585 515951
rect 185641 515949 185665 515951
rect 185721 515949 185727 515951
rect 185481 515897 185483 515949
rect 185663 515897 185665 515949
rect 185419 515895 185425 515897
rect 185481 515895 185505 515897
rect 185561 515895 185585 515897
rect 185641 515895 185665 515897
rect 185721 515895 185727 515897
rect 185419 515886 185727 515895
rect 186594 515853 186622 528573
rect 181338 515847 181390 515853
rect 181338 515789 181390 515795
rect 186582 515847 186634 515853
rect 186582 515789 186634 515795
rect 186490 515575 186542 515581
rect 186490 515517 186542 515523
rect 182166 515507 182218 515513
rect 182086 515455 182166 515461
rect 182086 515449 182218 515455
rect 182086 515433 182206 515449
rect 178443 515407 178751 515416
rect 178443 515405 178449 515407
rect 178505 515405 178529 515407
rect 178585 515405 178609 515407
rect 178665 515405 178689 515407
rect 178745 515405 178751 515407
rect 178505 515353 178507 515405
rect 178687 515353 178689 515405
rect 178443 515351 178449 515353
rect 178505 515351 178529 515353
rect 178585 515351 178609 515353
rect 178665 515351 178689 515353
rect 178745 515351 178751 515353
rect 178443 515342 178751 515351
rect 173332 513317 173388 513931
rect 177656 513367 177712 513931
rect 181980 513829 182036 513931
rect 182086 513829 182114 515433
rect 182261 515407 182569 515416
rect 182261 515405 182267 515407
rect 182323 515405 182347 515407
rect 182403 515405 182427 515407
rect 182483 515405 182507 515407
rect 182563 515405 182569 515407
rect 182323 515353 182325 515405
rect 182505 515353 182507 515405
rect 182261 515351 182267 515353
rect 182323 515351 182347 515353
rect 182403 515351 182427 515353
rect 182483 515351 182507 515353
rect 182563 515351 182569 515353
rect 182261 515342 182569 515351
rect 186079 515407 186387 515416
rect 186079 515405 186085 515407
rect 186141 515405 186165 515407
rect 186221 515405 186245 515407
rect 186301 515405 186325 515407
rect 186381 515405 186387 515407
rect 186141 515353 186143 515405
rect 186323 515353 186325 515405
rect 186079 515351 186085 515353
rect 186141 515351 186165 515353
rect 186221 515351 186245 515353
rect 186301 515351 186325 515353
rect 186381 515351 186387 515353
rect 186079 515342 186387 515351
rect 181980 513801 182114 513829
rect 186304 513829 186360 513931
rect 186502 513829 186530 515517
rect 186304 513801 186530 513829
rect 173250 513000 173450 513317
rect 173250 512800 173450 512810
rect 177580 513000 177780 513367
rect 181980 513317 182036 513801
rect 177580 512800 177780 512810
rect 181910 513000 182110 513317
rect 186304 513277 186360 513801
rect 181910 512800 182110 512810
rect 186230 513000 186430 513277
rect 186230 512800 186430 512810
rect 2000 509000 4000 509010
rect 2000 506990 4000 507000
rect 2000 466000 4000 466010
rect 2000 463990 4000 464000
rect 2000 423000 4000 423010
rect 2000 420990 4000 421000
rect 2000 380000 4000 380010
rect 2000 377990 4000 378000
<< via2 >>
rect 18000 699000 20000 701000
rect 70000 699000 72000 701000
rect 122000 699000 124000 701000
rect 3000 682000 5000 684000
rect 159400 538587 159480 538687
rect 161390 538577 161510 538697
rect 163030 538697 163330 538897
rect 166690 540097 166870 540277
rect 166690 539157 166870 539337
rect 170490 540097 170670 540277
rect 170490 539157 170670 539337
rect 174190 540107 174370 540287
rect 174190 539157 174370 539337
rect 177700 540097 177880 540277
rect 177690 539157 177870 539337
rect 181290 540097 181470 540277
rect 181290 539157 181470 539337
rect 184590 540097 184770 540277
rect 184590 539157 184770 539337
rect 187900 540097 188080 540277
rect 187890 539157 188070 539337
rect 191190 540097 191370 540277
rect 191810 540097 191990 540277
rect 191200 539167 191380 539347
rect 191820 539157 192000 539337
rect 160210 535467 160350 535597
rect 160350 535467 160360 535597
rect 160210 535457 160360 535467
rect 174631 530637 174687 530639
rect 174711 530637 174767 530639
rect 174791 530637 174847 530639
rect 174871 530637 174927 530639
rect 174631 530585 174677 530637
rect 174677 530585 174687 530637
rect 174711 530585 174741 530637
rect 174741 530585 174753 530637
rect 174753 530585 174767 530637
rect 174791 530585 174805 530637
rect 174805 530585 174817 530637
rect 174817 530585 174847 530637
rect 174871 530585 174881 530637
rect 174881 530585 174927 530637
rect 174631 530583 174687 530585
rect 174711 530583 174767 530585
rect 174791 530583 174847 530585
rect 174871 530583 174927 530585
rect 178449 530637 178505 530639
rect 178529 530637 178585 530639
rect 178609 530637 178665 530639
rect 178689 530637 178745 530639
rect 178449 530585 178495 530637
rect 178495 530585 178505 530637
rect 178529 530585 178559 530637
rect 178559 530585 178571 530637
rect 178571 530585 178585 530637
rect 178609 530585 178623 530637
rect 178623 530585 178635 530637
rect 178635 530585 178665 530637
rect 178689 530585 178699 530637
rect 178699 530585 178745 530637
rect 178449 530583 178505 530585
rect 178529 530583 178585 530585
rect 178609 530583 178665 530585
rect 178689 530583 178745 530585
rect 173971 530093 174027 530095
rect 174051 530093 174107 530095
rect 174131 530093 174187 530095
rect 174211 530093 174267 530095
rect 173971 530041 174017 530093
rect 174017 530041 174027 530093
rect 174051 530041 174081 530093
rect 174081 530041 174093 530093
rect 174093 530041 174107 530093
rect 174131 530041 174145 530093
rect 174145 530041 174157 530093
rect 174157 530041 174187 530093
rect 174211 530041 174221 530093
rect 174221 530041 174267 530093
rect 173971 530039 174027 530041
rect 174051 530039 174107 530041
rect 174131 530039 174187 530041
rect 174211 530039 174267 530041
rect 174631 529549 174687 529551
rect 174711 529549 174767 529551
rect 174791 529549 174847 529551
rect 174871 529549 174927 529551
rect 174631 529497 174677 529549
rect 174677 529497 174687 529549
rect 174711 529497 174741 529549
rect 174741 529497 174753 529549
rect 174753 529497 174767 529549
rect 174791 529497 174805 529549
rect 174805 529497 174817 529549
rect 174817 529497 174847 529549
rect 174871 529497 174881 529549
rect 174881 529497 174927 529549
rect 174631 529495 174687 529497
rect 174711 529495 174767 529497
rect 174791 529495 174847 529497
rect 174871 529495 174927 529497
rect 173971 529005 174027 529007
rect 174051 529005 174107 529007
rect 174131 529005 174187 529007
rect 174211 529005 174267 529007
rect 173971 528953 174017 529005
rect 174017 528953 174027 529005
rect 174051 528953 174081 529005
rect 174081 528953 174093 529005
rect 174093 528953 174107 529005
rect 174131 528953 174145 529005
rect 174145 528953 174157 529005
rect 174157 528953 174187 529005
rect 174211 528953 174221 529005
rect 174221 528953 174267 529005
rect 173971 528951 174027 528953
rect 174051 528951 174107 528953
rect 174131 528951 174187 528953
rect 174211 528951 174267 528953
rect 174631 528461 174687 528463
rect 174711 528461 174767 528463
rect 174791 528461 174847 528463
rect 174871 528461 174927 528463
rect 174631 528409 174677 528461
rect 174677 528409 174687 528461
rect 174711 528409 174741 528461
rect 174741 528409 174753 528461
rect 174753 528409 174767 528461
rect 174791 528409 174805 528461
rect 174805 528409 174817 528461
rect 174817 528409 174847 528461
rect 174871 528409 174881 528461
rect 174881 528409 174927 528461
rect 174631 528407 174687 528409
rect 174711 528407 174767 528409
rect 174791 528407 174847 528409
rect 174871 528407 174927 528409
rect 173971 527917 174027 527919
rect 174051 527917 174107 527919
rect 174131 527917 174187 527919
rect 174211 527917 174267 527919
rect 173971 527865 174017 527917
rect 174017 527865 174027 527917
rect 174051 527865 174081 527917
rect 174081 527865 174093 527917
rect 174093 527865 174107 527917
rect 174131 527865 174145 527917
rect 174145 527865 174157 527917
rect 174157 527865 174187 527917
rect 174211 527865 174221 527917
rect 174221 527865 174267 527917
rect 173971 527863 174027 527865
rect 174051 527863 174107 527865
rect 174131 527863 174187 527865
rect 174211 527863 174267 527865
rect 177789 530093 177845 530095
rect 177869 530093 177925 530095
rect 177949 530093 178005 530095
rect 178029 530093 178085 530095
rect 177789 530041 177835 530093
rect 177835 530041 177845 530093
rect 177869 530041 177899 530093
rect 177899 530041 177911 530093
rect 177911 530041 177925 530093
rect 177949 530041 177963 530093
rect 177963 530041 177975 530093
rect 177975 530041 178005 530093
rect 178029 530041 178039 530093
rect 178039 530041 178085 530093
rect 177789 530039 177845 530041
rect 177869 530039 177925 530041
rect 177949 530039 178005 530041
rect 178029 530039 178085 530041
rect 177789 529005 177845 529007
rect 177869 529005 177925 529007
rect 177949 529005 178005 529007
rect 178029 529005 178085 529007
rect 177789 528953 177835 529005
rect 177835 528953 177845 529005
rect 177869 528953 177899 529005
rect 177899 528953 177911 529005
rect 177911 528953 177925 529005
rect 177949 528953 177963 529005
rect 177963 528953 177975 529005
rect 177975 528953 178005 529005
rect 178029 528953 178039 529005
rect 178039 528953 178085 529005
rect 177789 528951 177845 528953
rect 177869 528951 177925 528953
rect 177949 528951 178005 528953
rect 178029 528951 178085 528953
rect 178449 529549 178505 529551
rect 178529 529549 178585 529551
rect 178609 529549 178665 529551
rect 178689 529549 178745 529551
rect 178449 529497 178495 529549
rect 178495 529497 178505 529549
rect 178529 529497 178559 529549
rect 178559 529497 178571 529549
rect 178571 529497 178585 529549
rect 178609 529497 178623 529549
rect 178623 529497 178635 529549
rect 178635 529497 178665 529549
rect 178689 529497 178699 529549
rect 178699 529497 178745 529549
rect 178449 529495 178505 529497
rect 178529 529495 178585 529497
rect 178609 529495 178665 529497
rect 178689 529495 178745 529497
rect 177789 527917 177845 527919
rect 177869 527917 177925 527919
rect 177949 527917 178005 527919
rect 178029 527917 178085 527919
rect 177789 527865 177835 527917
rect 177835 527865 177845 527917
rect 177869 527865 177899 527917
rect 177899 527865 177911 527917
rect 177911 527865 177925 527917
rect 177949 527865 177963 527917
rect 177963 527865 177975 527917
rect 177975 527865 178005 527917
rect 178029 527865 178039 527917
rect 178039 527865 178085 527917
rect 177789 527863 177845 527865
rect 177869 527863 177925 527865
rect 177949 527863 178005 527865
rect 178029 527863 178085 527865
rect 174631 527373 174687 527375
rect 174711 527373 174767 527375
rect 174791 527373 174847 527375
rect 174871 527373 174927 527375
rect 174631 527321 174677 527373
rect 174677 527321 174687 527373
rect 174711 527321 174741 527373
rect 174741 527321 174753 527373
rect 174753 527321 174767 527373
rect 174791 527321 174805 527373
rect 174805 527321 174817 527373
rect 174817 527321 174847 527373
rect 174871 527321 174881 527373
rect 174881 527321 174927 527373
rect 174631 527319 174687 527321
rect 174711 527319 174767 527321
rect 174791 527319 174847 527321
rect 174871 527319 174927 527321
rect 173971 526829 174027 526831
rect 174051 526829 174107 526831
rect 174131 526829 174187 526831
rect 174211 526829 174267 526831
rect 173971 526777 174017 526829
rect 174017 526777 174027 526829
rect 174051 526777 174081 526829
rect 174081 526777 174093 526829
rect 174093 526777 174107 526829
rect 174131 526777 174145 526829
rect 174145 526777 174157 526829
rect 174157 526777 174187 526829
rect 174211 526777 174221 526829
rect 174221 526777 174267 526829
rect 173971 526775 174027 526777
rect 174051 526775 174107 526777
rect 174131 526775 174187 526777
rect 174211 526775 174267 526777
rect 177789 526829 177845 526831
rect 177869 526829 177925 526831
rect 177949 526829 178005 526831
rect 178029 526829 178085 526831
rect 177789 526777 177835 526829
rect 177835 526777 177845 526829
rect 177869 526777 177899 526829
rect 177899 526777 177911 526829
rect 177911 526777 177925 526829
rect 177949 526777 177963 526829
rect 177963 526777 177975 526829
rect 177975 526777 178005 526829
rect 178029 526777 178039 526829
rect 178039 526777 178085 526829
rect 177789 526775 177845 526777
rect 177869 526775 177925 526777
rect 177949 526775 178005 526777
rect 178029 526775 178085 526777
rect 174631 526285 174687 526287
rect 174711 526285 174767 526287
rect 174791 526285 174847 526287
rect 174871 526285 174927 526287
rect 174631 526233 174677 526285
rect 174677 526233 174687 526285
rect 174711 526233 174741 526285
rect 174741 526233 174753 526285
rect 174753 526233 174767 526285
rect 174791 526233 174805 526285
rect 174805 526233 174817 526285
rect 174817 526233 174847 526285
rect 174871 526233 174881 526285
rect 174881 526233 174927 526285
rect 174631 526231 174687 526233
rect 174711 526231 174767 526233
rect 174791 526231 174847 526233
rect 174871 526231 174927 526233
rect 173971 525741 174027 525743
rect 174051 525741 174107 525743
rect 174131 525741 174187 525743
rect 174211 525741 174267 525743
rect 173971 525689 174017 525741
rect 174017 525689 174027 525741
rect 174051 525689 174081 525741
rect 174081 525689 174093 525741
rect 174093 525689 174107 525741
rect 174131 525689 174145 525741
rect 174145 525689 174157 525741
rect 174157 525689 174187 525741
rect 174211 525689 174221 525741
rect 174221 525689 174267 525741
rect 173971 525687 174027 525689
rect 174051 525687 174107 525689
rect 174131 525687 174187 525689
rect 174211 525687 174267 525689
rect 177789 525741 177845 525743
rect 177869 525741 177925 525743
rect 177949 525741 178005 525743
rect 178029 525741 178085 525743
rect 177789 525689 177835 525741
rect 177835 525689 177845 525741
rect 177869 525689 177899 525741
rect 177899 525689 177911 525741
rect 177911 525689 177925 525741
rect 177949 525689 177963 525741
rect 177963 525689 177975 525741
rect 177975 525689 178005 525741
rect 178029 525689 178039 525741
rect 178039 525689 178085 525741
rect 177789 525687 177845 525689
rect 177869 525687 177925 525689
rect 177949 525687 178005 525689
rect 178029 525687 178085 525689
rect 174631 525197 174687 525199
rect 174711 525197 174767 525199
rect 174791 525197 174847 525199
rect 174871 525197 174927 525199
rect 174631 525145 174677 525197
rect 174677 525145 174687 525197
rect 174711 525145 174741 525197
rect 174741 525145 174753 525197
rect 174753 525145 174767 525197
rect 174791 525145 174805 525197
rect 174805 525145 174817 525197
rect 174817 525145 174847 525197
rect 174871 525145 174881 525197
rect 174881 525145 174927 525197
rect 174631 525143 174687 525145
rect 174711 525143 174767 525145
rect 174791 525143 174847 525145
rect 174871 525143 174927 525145
rect 173971 524653 174027 524655
rect 174051 524653 174107 524655
rect 174131 524653 174187 524655
rect 174211 524653 174267 524655
rect 173971 524601 174017 524653
rect 174017 524601 174027 524653
rect 174051 524601 174081 524653
rect 174081 524601 174093 524653
rect 174093 524601 174107 524653
rect 174131 524601 174145 524653
rect 174145 524601 174157 524653
rect 174157 524601 174187 524653
rect 174211 524601 174221 524653
rect 174221 524601 174267 524653
rect 173971 524599 174027 524601
rect 174051 524599 174107 524601
rect 174131 524599 174187 524601
rect 174211 524599 174267 524601
rect 177789 524653 177845 524655
rect 177869 524653 177925 524655
rect 177949 524653 178005 524655
rect 178029 524653 178085 524655
rect 177789 524601 177835 524653
rect 177835 524601 177845 524653
rect 177869 524601 177899 524653
rect 177899 524601 177911 524653
rect 177911 524601 177925 524653
rect 177949 524601 177963 524653
rect 177963 524601 177975 524653
rect 177975 524601 178005 524653
rect 178029 524601 178039 524653
rect 178039 524601 178085 524653
rect 177789 524599 177845 524601
rect 177869 524599 177925 524601
rect 177949 524599 178005 524601
rect 178029 524599 178085 524601
rect 174631 524109 174687 524111
rect 174711 524109 174767 524111
rect 174791 524109 174847 524111
rect 174871 524109 174927 524111
rect 174631 524057 174677 524109
rect 174677 524057 174687 524109
rect 174711 524057 174741 524109
rect 174741 524057 174753 524109
rect 174753 524057 174767 524109
rect 174791 524057 174805 524109
rect 174805 524057 174817 524109
rect 174817 524057 174847 524109
rect 174871 524057 174881 524109
rect 174881 524057 174927 524109
rect 174631 524055 174687 524057
rect 174711 524055 174767 524057
rect 174791 524055 174847 524057
rect 174871 524055 174927 524057
rect 173971 523565 174027 523567
rect 174051 523565 174107 523567
rect 174131 523565 174187 523567
rect 174211 523565 174267 523567
rect 173971 523513 174017 523565
rect 174017 523513 174027 523565
rect 174051 523513 174081 523565
rect 174081 523513 174093 523565
rect 174093 523513 174107 523565
rect 174131 523513 174145 523565
rect 174145 523513 174157 523565
rect 174157 523513 174187 523565
rect 174211 523513 174221 523565
rect 174221 523513 174267 523565
rect 173971 523511 174027 523513
rect 174051 523511 174107 523513
rect 174131 523511 174187 523513
rect 174211 523511 174267 523513
rect 177789 523565 177845 523567
rect 177869 523565 177925 523567
rect 177949 523565 178005 523567
rect 178029 523565 178085 523567
rect 177789 523513 177835 523565
rect 177835 523513 177845 523565
rect 177869 523513 177899 523565
rect 177899 523513 177911 523565
rect 177911 523513 177925 523565
rect 177949 523513 177963 523565
rect 177963 523513 177975 523565
rect 177975 523513 178005 523565
rect 178029 523513 178039 523565
rect 178039 523513 178085 523565
rect 177789 523511 177845 523513
rect 177869 523511 177925 523513
rect 177949 523511 178005 523513
rect 178029 523511 178085 523513
rect 174631 523021 174687 523023
rect 174711 523021 174767 523023
rect 174791 523021 174847 523023
rect 174871 523021 174927 523023
rect 174631 522969 174677 523021
rect 174677 522969 174687 523021
rect 174711 522969 174741 523021
rect 174741 522969 174753 523021
rect 174753 522969 174767 523021
rect 174791 522969 174805 523021
rect 174805 522969 174817 523021
rect 174817 522969 174847 523021
rect 174871 522969 174881 523021
rect 174881 522969 174927 523021
rect 174631 522967 174687 522969
rect 174711 522967 174767 522969
rect 174791 522967 174847 522969
rect 174871 522967 174927 522969
rect 173971 522477 174027 522479
rect 174051 522477 174107 522479
rect 174131 522477 174187 522479
rect 174211 522477 174267 522479
rect 173971 522425 174017 522477
rect 174017 522425 174027 522477
rect 174051 522425 174081 522477
rect 174081 522425 174093 522477
rect 174093 522425 174107 522477
rect 174131 522425 174145 522477
rect 174145 522425 174157 522477
rect 174157 522425 174187 522477
rect 174211 522425 174221 522477
rect 174221 522425 174267 522477
rect 173971 522423 174027 522425
rect 174051 522423 174107 522425
rect 174131 522423 174187 522425
rect 174211 522423 174267 522425
rect 177789 522477 177845 522479
rect 177869 522477 177925 522479
rect 177949 522477 178005 522479
rect 178029 522477 178085 522479
rect 177789 522425 177835 522477
rect 177835 522425 177845 522477
rect 177869 522425 177899 522477
rect 177899 522425 177911 522477
rect 177911 522425 177925 522477
rect 177949 522425 177963 522477
rect 177963 522425 177975 522477
rect 177975 522425 178005 522477
rect 178029 522425 178039 522477
rect 178039 522425 178085 522477
rect 177789 522423 177845 522425
rect 177869 522423 177925 522425
rect 177949 522423 178005 522425
rect 178029 522423 178085 522425
rect 174631 521933 174687 521935
rect 174711 521933 174767 521935
rect 174791 521933 174847 521935
rect 174871 521933 174927 521935
rect 174631 521881 174677 521933
rect 174677 521881 174687 521933
rect 174711 521881 174741 521933
rect 174741 521881 174753 521933
rect 174753 521881 174767 521933
rect 174791 521881 174805 521933
rect 174805 521881 174817 521933
rect 174817 521881 174847 521933
rect 174871 521881 174881 521933
rect 174881 521881 174927 521933
rect 174631 521879 174687 521881
rect 174711 521879 174767 521881
rect 174791 521879 174847 521881
rect 174871 521879 174927 521881
rect 173971 521389 174027 521391
rect 174051 521389 174107 521391
rect 174131 521389 174187 521391
rect 174211 521389 174267 521391
rect 173971 521337 174017 521389
rect 174017 521337 174027 521389
rect 174051 521337 174081 521389
rect 174081 521337 174093 521389
rect 174093 521337 174107 521389
rect 174131 521337 174145 521389
rect 174145 521337 174157 521389
rect 174157 521337 174187 521389
rect 174211 521337 174221 521389
rect 174221 521337 174267 521389
rect 173971 521335 174027 521337
rect 174051 521335 174107 521337
rect 174131 521335 174187 521337
rect 174211 521335 174267 521337
rect 177789 521389 177845 521391
rect 177869 521389 177925 521391
rect 177949 521389 178005 521391
rect 178029 521389 178085 521391
rect 177789 521337 177835 521389
rect 177835 521337 177845 521389
rect 177869 521337 177899 521389
rect 177899 521337 177911 521389
rect 177911 521337 177925 521389
rect 177949 521337 177963 521389
rect 177963 521337 177975 521389
rect 177975 521337 178005 521389
rect 178029 521337 178039 521389
rect 178039 521337 178085 521389
rect 177789 521335 177845 521337
rect 177869 521335 177925 521337
rect 177949 521335 178005 521337
rect 178029 521335 178085 521337
rect 174631 520845 174687 520847
rect 174711 520845 174767 520847
rect 174791 520845 174847 520847
rect 174871 520845 174927 520847
rect 174631 520793 174677 520845
rect 174677 520793 174687 520845
rect 174711 520793 174741 520845
rect 174741 520793 174753 520845
rect 174753 520793 174767 520845
rect 174791 520793 174805 520845
rect 174805 520793 174817 520845
rect 174817 520793 174847 520845
rect 174871 520793 174881 520845
rect 174881 520793 174927 520845
rect 174631 520791 174687 520793
rect 174711 520791 174767 520793
rect 174791 520791 174847 520793
rect 174871 520791 174927 520793
rect 173971 520301 174027 520303
rect 174051 520301 174107 520303
rect 174131 520301 174187 520303
rect 174211 520301 174267 520303
rect 173971 520249 174017 520301
rect 174017 520249 174027 520301
rect 174051 520249 174081 520301
rect 174081 520249 174093 520301
rect 174093 520249 174107 520301
rect 174131 520249 174145 520301
rect 174145 520249 174157 520301
rect 174157 520249 174187 520301
rect 174211 520249 174221 520301
rect 174221 520249 174267 520301
rect 173971 520247 174027 520249
rect 174051 520247 174107 520249
rect 174131 520247 174187 520249
rect 174211 520247 174267 520249
rect 177789 520301 177845 520303
rect 177869 520301 177925 520303
rect 177949 520301 178005 520303
rect 178029 520301 178085 520303
rect 177789 520249 177835 520301
rect 177835 520249 177845 520301
rect 177869 520249 177899 520301
rect 177899 520249 177911 520301
rect 177911 520249 177925 520301
rect 177949 520249 177963 520301
rect 177963 520249 177975 520301
rect 177975 520249 178005 520301
rect 178029 520249 178039 520301
rect 178039 520249 178085 520301
rect 177789 520247 177845 520249
rect 177869 520247 177925 520249
rect 177949 520247 178005 520249
rect 178029 520247 178085 520249
rect 174631 519757 174687 519759
rect 174711 519757 174767 519759
rect 174791 519757 174847 519759
rect 174871 519757 174927 519759
rect 174631 519705 174677 519757
rect 174677 519705 174687 519757
rect 174711 519705 174741 519757
rect 174741 519705 174753 519757
rect 174753 519705 174767 519757
rect 174791 519705 174805 519757
rect 174805 519705 174817 519757
rect 174817 519705 174847 519757
rect 174871 519705 174881 519757
rect 174881 519705 174927 519757
rect 174631 519703 174687 519705
rect 174711 519703 174767 519705
rect 174791 519703 174847 519705
rect 174871 519703 174927 519705
rect 173971 519213 174027 519215
rect 174051 519213 174107 519215
rect 174131 519213 174187 519215
rect 174211 519213 174267 519215
rect 173971 519161 174017 519213
rect 174017 519161 174027 519213
rect 174051 519161 174081 519213
rect 174081 519161 174093 519213
rect 174093 519161 174107 519213
rect 174131 519161 174145 519213
rect 174145 519161 174157 519213
rect 174157 519161 174187 519213
rect 174211 519161 174221 519213
rect 174221 519161 174267 519213
rect 173971 519159 174027 519161
rect 174051 519159 174107 519161
rect 174131 519159 174187 519161
rect 174211 519159 174267 519161
rect 177789 519213 177845 519215
rect 177869 519213 177925 519215
rect 177949 519213 178005 519215
rect 178029 519213 178085 519215
rect 177789 519161 177835 519213
rect 177835 519161 177845 519213
rect 177869 519161 177899 519213
rect 177899 519161 177911 519213
rect 177911 519161 177925 519213
rect 177949 519161 177963 519213
rect 177963 519161 177975 519213
rect 177975 519161 178005 519213
rect 178029 519161 178039 519213
rect 178039 519161 178085 519213
rect 177789 519159 177845 519161
rect 177869 519159 177925 519161
rect 177949 519159 178005 519161
rect 178029 519159 178085 519161
rect 174631 518669 174687 518671
rect 174711 518669 174767 518671
rect 174791 518669 174847 518671
rect 174871 518669 174927 518671
rect 174631 518617 174677 518669
rect 174677 518617 174687 518669
rect 174711 518617 174741 518669
rect 174741 518617 174753 518669
rect 174753 518617 174767 518669
rect 174791 518617 174805 518669
rect 174805 518617 174817 518669
rect 174817 518617 174847 518669
rect 174871 518617 174881 518669
rect 174881 518617 174927 518669
rect 174631 518615 174687 518617
rect 174711 518615 174767 518617
rect 174791 518615 174847 518617
rect 174871 518615 174927 518617
rect 173971 518125 174027 518127
rect 174051 518125 174107 518127
rect 174131 518125 174187 518127
rect 174211 518125 174267 518127
rect 173971 518073 174017 518125
rect 174017 518073 174027 518125
rect 174051 518073 174081 518125
rect 174081 518073 174093 518125
rect 174093 518073 174107 518125
rect 174131 518073 174145 518125
rect 174145 518073 174157 518125
rect 174157 518073 174187 518125
rect 174211 518073 174221 518125
rect 174221 518073 174267 518125
rect 173971 518071 174027 518073
rect 174051 518071 174107 518073
rect 174131 518071 174187 518073
rect 174211 518071 174267 518073
rect 177789 518125 177845 518127
rect 177869 518125 177925 518127
rect 177949 518125 178005 518127
rect 178029 518125 178085 518127
rect 177789 518073 177835 518125
rect 177835 518073 177845 518125
rect 177869 518073 177899 518125
rect 177899 518073 177911 518125
rect 177911 518073 177925 518125
rect 177949 518073 177963 518125
rect 177963 518073 177975 518125
rect 177975 518073 178005 518125
rect 178029 518073 178039 518125
rect 178039 518073 178085 518125
rect 177789 518071 177845 518073
rect 177869 518071 177925 518073
rect 177949 518071 178005 518073
rect 178029 518071 178085 518073
rect 174631 517581 174687 517583
rect 174711 517581 174767 517583
rect 174791 517581 174847 517583
rect 174871 517581 174927 517583
rect 174631 517529 174677 517581
rect 174677 517529 174687 517581
rect 174711 517529 174741 517581
rect 174741 517529 174753 517581
rect 174753 517529 174767 517581
rect 174791 517529 174805 517581
rect 174805 517529 174817 517581
rect 174817 517529 174847 517581
rect 174871 517529 174881 517581
rect 174881 517529 174927 517581
rect 174631 517527 174687 517529
rect 174711 517527 174767 517529
rect 174791 517527 174847 517529
rect 174871 517527 174927 517529
rect 178449 528461 178505 528463
rect 178529 528461 178585 528463
rect 178609 528461 178665 528463
rect 178689 528461 178745 528463
rect 178449 528409 178495 528461
rect 178495 528409 178505 528461
rect 178529 528409 178559 528461
rect 178559 528409 178571 528461
rect 178571 528409 178585 528461
rect 178609 528409 178623 528461
rect 178623 528409 178635 528461
rect 178635 528409 178665 528461
rect 178689 528409 178699 528461
rect 178699 528409 178745 528461
rect 178449 528407 178505 528409
rect 178529 528407 178585 528409
rect 178609 528407 178665 528409
rect 178689 528407 178745 528409
rect 182267 530637 182323 530639
rect 182347 530637 182403 530639
rect 182427 530637 182483 530639
rect 182507 530637 182563 530639
rect 182267 530585 182313 530637
rect 182313 530585 182323 530637
rect 182347 530585 182377 530637
rect 182377 530585 182389 530637
rect 182389 530585 182403 530637
rect 182427 530585 182441 530637
rect 182441 530585 182453 530637
rect 182453 530585 182483 530637
rect 182507 530585 182517 530637
rect 182517 530585 182563 530637
rect 182267 530583 182323 530585
rect 182347 530583 182403 530585
rect 182427 530583 182483 530585
rect 182507 530583 182563 530585
rect 186085 530637 186141 530639
rect 186165 530637 186221 530639
rect 186245 530637 186301 530639
rect 186325 530637 186381 530639
rect 186085 530585 186131 530637
rect 186131 530585 186141 530637
rect 186165 530585 186195 530637
rect 186195 530585 186207 530637
rect 186207 530585 186221 530637
rect 186245 530585 186259 530637
rect 186259 530585 186271 530637
rect 186271 530585 186301 530637
rect 186325 530585 186335 530637
rect 186335 530585 186381 530637
rect 186085 530583 186141 530585
rect 186165 530583 186221 530585
rect 186245 530583 186301 530585
rect 186325 530583 186381 530585
rect 181607 530093 181663 530095
rect 181687 530093 181743 530095
rect 181767 530093 181823 530095
rect 181847 530093 181903 530095
rect 181607 530041 181653 530093
rect 181653 530041 181663 530093
rect 181687 530041 181717 530093
rect 181717 530041 181729 530093
rect 181729 530041 181743 530093
rect 181767 530041 181781 530093
rect 181781 530041 181793 530093
rect 181793 530041 181823 530093
rect 181847 530041 181857 530093
rect 181857 530041 181903 530093
rect 181607 530039 181663 530041
rect 181687 530039 181743 530041
rect 181767 530039 181823 530041
rect 181847 530039 181903 530041
rect 181607 529005 181663 529007
rect 181687 529005 181743 529007
rect 181767 529005 181823 529007
rect 181847 529005 181903 529007
rect 181607 528953 181653 529005
rect 181653 528953 181663 529005
rect 181687 528953 181717 529005
rect 181717 528953 181729 529005
rect 181729 528953 181743 529005
rect 181767 528953 181781 529005
rect 181781 528953 181793 529005
rect 181793 528953 181823 529005
rect 181847 528953 181857 529005
rect 181857 528953 181903 529005
rect 181607 528951 181663 528953
rect 181687 528951 181743 528953
rect 181767 528951 181823 528953
rect 181847 528951 181903 528953
rect 182267 529549 182323 529551
rect 182347 529549 182403 529551
rect 182427 529549 182483 529551
rect 182507 529549 182563 529551
rect 182267 529497 182313 529549
rect 182313 529497 182323 529549
rect 182347 529497 182377 529549
rect 182377 529497 182389 529549
rect 182389 529497 182403 529549
rect 182427 529497 182441 529549
rect 182441 529497 182453 529549
rect 182453 529497 182483 529549
rect 182507 529497 182517 529549
rect 182517 529497 182563 529549
rect 182267 529495 182323 529497
rect 182347 529495 182403 529497
rect 182427 529495 182483 529497
rect 182507 529495 182563 529497
rect 185425 530093 185481 530095
rect 185505 530093 185561 530095
rect 185585 530093 185641 530095
rect 185665 530093 185721 530095
rect 185425 530041 185471 530093
rect 185471 530041 185481 530093
rect 185505 530041 185535 530093
rect 185535 530041 185547 530093
rect 185547 530041 185561 530093
rect 185585 530041 185599 530093
rect 185599 530041 185611 530093
rect 185611 530041 185641 530093
rect 185665 530041 185675 530093
rect 185675 530041 185721 530093
rect 185425 530039 185481 530041
rect 185505 530039 185561 530041
rect 185585 530039 185641 530041
rect 185665 530039 185721 530041
rect 186085 529549 186141 529551
rect 186165 529549 186221 529551
rect 186245 529549 186301 529551
rect 186325 529549 186381 529551
rect 186085 529497 186131 529549
rect 186131 529497 186141 529549
rect 186165 529497 186195 529549
rect 186195 529497 186207 529549
rect 186207 529497 186221 529549
rect 186245 529497 186259 529549
rect 186259 529497 186271 529549
rect 186271 529497 186301 529549
rect 186325 529497 186335 529549
rect 186335 529497 186381 529549
rect 186085 529495 186141 529497
rect 186165 529495 186221 529497
rect 186245 529495 186301 529497
rect 186325 529495 186381 529497
rect 185425 529005 185481 529007
rect 185505 529005 185561 529007
rect 185585 529005 185641 529007
rect 185665 529005 185721 529007
rect 185425 528953 185471 529005
rect 185471 528953 185481 529005
rect 185505 528953 185535 529005
rect 185535 528953 185547 529005
rect 185547 528953 185561 529005
rect 185585 528953 185599 529005
rect 185599 528953 185611 529005
rect 185611 528953 185641 529005
rect 185665 528953 185675 529005
rect 185675 528953 185721 529005
rect 185425 528951 185481 528953
rect 185505 528951 185561 528953
rect 185585 528951 185641 528953
rect 185665 528951 185721 528953
rect 182267 528461 182323 528463
rect 182347 528461 182403 528463
rect 182427 528461 182483 528463
rect 182507 528461 182563 528463
rect 182267 528409 182313 528461
rect 182313 528409 182323 528461
rect 182347 528409 182377 528461
rect 182377 528409 182389 528461
rect 182389 528409 182403 528461
rect 182427 528409 182441 528461
rect 182441 528409 182453 528461
rect 182453 528409 182483 528461
rect 182507 528409 182517 528461
rect 182517 528409 182563 528461
rect 182267 528407 182323 528409
rect 182347 528407 182403 528409
rect 182427 528407 182483 528409
rect 182507 528407 182563 528409
rect 186085 528461 186141 528463
rect 186165 528461 186221 528463
rect 186245 528461 186301 528463
rect 186325 528461 186381 528463
rect 186085 528409 186131 528461
rect 186131 528409 186141 528461
rect 186165 528409 186195 528461
rect 186195 528409 186207 528461
rect 186207 528409 186221 528461
rect 186245 528409 186259 528461
rect 186259 528409 186271 528461
rect 186271 528409 186301 528461
rect 186325 528409 186335 528461
rect 186335 528409 186381 528461
rect 186085 528407 186141 528409
rect 186165 528407 186221 528409
rect 186245 528407 186301 528409
rect 186325 528407 186381 528409
rect 178449 527373 178505 527375
rect 178529 527373 178585 527375
rect 178609 527373 178665 527375
rect 178689 527373 178745 527375
rect 178449 527321 178495 527373
rect 178495 527321 178505 527373
rect 178529 527321 178559 527373
rect 178559 527321 178571 527373
rect 178571 527321 178585 527373
rect 178609 527321 178623 527373
rect 178623 527321 178635 527373
rect 178635 527321 178665 527373
rect 178689 527321 178699 527373
rect 178699 527321 178745 527373
rect 178449 527319 178505 527321
rect 178529 527319 178585 527321
rect 178609 527319 178665 527321
rect 178689 527319 178745 527321
rect 178449 526285 178505 526287
rect 178529 526285 178585 526287
rect 178609 526285 178665 526287
rect 178689 526285 178745 526287
rect 178449 526233 178495 526285
rect 178495 526233 178505 526285
rect 178529 526233 178559 526285
rect 178559 526233 178571 526285
rect 178571 526233 178585 526285
rect 178609 526233 178623 526285
rect 178623 526233 178635 526285
rect 178635 526233 178665 526285
rect 178689 526233 178699 526285
rect 178699 526233 178745 526285
rect 178449 526231 178505 526233
rect 178529 526231 178585 526233
rect 178609 526231 178665 526233
rect 178689 526231 178745 526233
rect 178449 525197 178505 525199
rect 178529 525197 178585 525199
rect 178609 525197 178665 525199
rect 178689 525197 178745 525199
rect 178449 525145 178495 525197
rect 178495 525145 178505 525197
rect 178529 525145 178559 525197
rect 178559 525145 178571 525197
rect 178571 525145 178585 525197
rect 178609 525145 178623 525197
rect 178623 525145 178635 525197
rect 178635 525145 178665 525197
rect 178689 525145 178699 525197
rect 178699 525145 178745 525197
rect 178449 525143 178505 525145
rect 178529 525143 178585 525145
rect 178609 525143 178665 525145
rect 178689 525143 178745 525145
rect 178449 524109 178505 524111
rect 178529 524109 178585 524111
rect 178609 524109 178665 524111
rect 178689 524109 178745 524111
rect 178449 524057 178495 524109
rect 178495 524057 178505 524109
rect 178529 524057 178559 524109
rect 178559 524057 178571 524109
rect 178571 524057 178585 524109
rect 178609 524057 178623 524109
rect 178623 524057 178635 524109
rect 178635 524057 178665 524109
rect 178689 524057 178699 524109
rect 178699 524057 178745 524109
rect 178449 524055 178505 524057
rect 178529 524055 178585 524057
rect 178609 524055 178665 524057
rect 178689 524055 178745 524057
rect 178449 523021 178505 523023
rect 178529 523021 178585 523023
rect 178609 523021 178665 523023
rect 178689 523021 178745 523023
rect 178449 522969 178495 523021
rect 178495 522969 178505 523021
rect 178529 522969 178559 523021
rect 178559 522969 178571 523021
rect 178571 522969 178585 523021
rect 178609 522969 178623 523021
rect 178623 522969 178635 523021
rect 178635 522969 178665 523021
rect 178689 522969 178699 523021
rect 178699 522969 178745 523021
rect 178449 522967 178505 522969
rect 178529 522967 178585 522969
rect 178609 522967 178665 522969
rect 178689 522967 178745 522969
rect 178449 521933 178505 521935
rect 178529 521933 178585 521935
rect 178609 521933 178665 521935
rect 178689 521933 178745 521935
rect 178449 521881 178495 521933
rect 178495 521881 178505 521933
rect 178529 521881 178559 521933
rect 178559 521881 178571 521933
rect 178571 521881 178585 521933
rect 178609 521881 178623 521933
rect 178623 521881 178635 521933
rect 178635 521881 178665 521933
rect 178689 521881 178699 521933
rect 178699 521881 178745 521933
rect 178449 521879 178505 521881
rect 178529 521879 178585 521881
rect 178609 521879 178665 521881
rect 178689 521879 178745 521881
rect 178449 520845 178505 520847
rect 178529 520845 178585 520847
rect 178609 520845 178665 520847
rect 178689 520845 178745 520847
rect 178449 520793 178495 520845
rect 178495 520793 178505 520845
rect 178529 520793 178559 520845
rect 178559 520793 178571 520845
rect 178571 520793 178585 520845
rect 178609 520793 178623 520845
rect 178623 520793 178635 520845
rect 178635 520793 178665 520845
rect 178689 520793 178699 520845
rect 178699 520793 178745 520845
rect 178449 520791 178505 520793
rect 178529 520791 178585 520793
rect 178609 520791 178665 520793
rect 178689 520791 178745 520793
rect 178449 519757 178505 519759
rect 178529 519757 178585 519759
rect 178609 519757 178665 519759
rect 178689 519757 178745 519759
rect 178449 519705 178495 519757
rect 178495 519705 178505 519757
rect 178529 519705 178559 519757
rect 178559 519705 178571 519757
rect 178571 519705 178585 519757
rect 178609 519705 178623 519757
rect 178623 519705 178635 519757
rect 178635 519705 178665 519757
rect 178689 519705 178699 519757
rect 178699 519705 178745 519757
rect 178449 519703 178505 519705
rect 178529 519703 178585 519705
rect 178609 519703 178665 519705
rect 178689 519703 178745 519705
rect 178449 518669 178505 518671
rect 178529 518669 178585 518671
rect 178609 518669 178665 518671
rect 178689 518669 178745 518671
rect 178449 518617 178495 518669
rect 178495 518617 178505 518669
rect 178529 518617 178559 518669
rect 178559 518617 178571 518669
rect 178571 518617 178585 518669
rect 178609 518617 178623 518669
rect 178623 518617 178635 518669
rect 178635 518617 178665 518669
rect 178689 518617 178699 518669
rect 178699 518617 178745 518669
rect 178449 518615 178505 518617
rect 178529 518615 178585 518617
rect 178609 518615 178665 518617
rect 178689 518615 178745 518617
rect 178449 517581 178505 517583
rect 178529 517581 178585 517583
rect 178609 517581 178665 517583
rect 178689 517581 178745 517583
rect 178449 517529 178495 517581
rect 178495 517529 178505 517581
rect 178529 517529 178559 517581
rect 178559 517529 178571 517581
rect 178571 517529 178585 517581
rect 178609 517529 178623 517581
rect 178623 517529 178635 517581
rect 178635 517529 178665 517581
rect 178689 517529 178699 517581
rect 178699 517529 178745 517581
rect 178449 517527 178505 517529
rect 178529 517527 178585 517529
rect 178609 517527 178665 517529
rect 178689 517527 178745 517529
rect 173971 517037 174027 517039
rect 174051 517037 174107 517039
rect 174131 517037 174187 517039
rect 174211 517037 174267 517039
rect 173971 516985 174017 517037
rect 174017 516985 174027 517037
rect 174051 516985 174081 517037
rect 174081 516985 174093 517037
rect 174093 516985 174107 517037
rect 174131 516985 174145 517037
rect 174145 516985 174157 517037
rect 174157 516985 174187 517037
rect 174211 516985 174221 517037
rect 174221 516985 174267 517037
rect 173971 516983 174027 516985
rect 174051 516983 174107 516985
rect 174131 516983 174187 516985
rect 174211 516983 174267 516985
rect 174631 516493 174687 516495
rect 174711 516493 174767 516495
rect 174791 516493 174847 516495
rect 174871 516493 174927 516495
rect 174631 516441 174677 516493
rect 174677 516441 174687 516493
rect 174711 516441 174741 516493
rect 174741 516441 174753 516493
rect 174753 516441 174767 516493
rect 174791 516441 174805 516493
rect 174805 516441 174817 516493
rect 174817 516441 174847 516493
rect 174871 516441 174881 516493
rect 174881 516441 174927 516493
rect 174631 516439 174687 516441
rect 174711 516439 174767 516441
rect 174791 516439 174847 516441
rect 174871 516439 174927 516441
rect 173971 515949 174027 515951
rect 174051 515949 174107 515951
rect 174131 515949 174187 515951
rect 174211 515949 174267 515951
rect 173971 515897 174017 515949
rect 174017 515897 174027 515949
rect 174051 515897 174081 515949
rect 174081 515897 174093 515949
rect 174093 515897 174107 515949
rect 174131 515897 174145 515949
rect 174145 515897 174157 515949
rect 174157 515897 174187 515949
rect 174211 515897 174221 515949
rect 174221 515897 174267 515949
rect 173971 515895 174027 515897
rect 174051 515895 174107 515897
rect 174131 515895 174187 515897
rect 174211 515895 174267 515897
rect 174631 515405 174687 515407
rect 174711 515405 174767 515407
rect 174791 515405 174847 515407
rect 174871 515405 174927 515407
rect 174631 515353 174677 515405
rect 174677 515353 174687 515405
rect 174711 515353 174741 515405
rect 174741 515353 174753 515405
rect 174753 515353 174767 515405
rect 174791 515353 174805 515405
rect 174805 515353 174817 515405
rect 174817 515353 174847 515405
rect 174871 515353 174881 515405
rect 174881 515353 174927 515405
rect 174631 515351 174687 515353
rect 174711 515351 174767 515353
rect 174791 515351 174847 515353
rect 174871 515351 174927 515353
rect 177789 517037 177845 517039
rect 177869 517037 177925 517039
rect 177949 517037 178005 517039
rect 178029 517037 178085 517039
rect 177789 516985 177835 517037
rect 177835 516985 177845 517037
rect 177869 516985 177899 517037
rect 177899 516985 177911 517037
rect 177911 516985 177925 517037
rect 177949 516985 177963 517037
rect 177963 516985 177975 517037
rect 177975 516985 178005 517037
rect 178029 516985 178039 517037
rect 178039 516985 178085 517037
rect 177789 516983 177845 516985
rect 177869 516983 177925 516985
rect 177949 516983 178005 516985
rect 178029 516983 178085 516985
rect 178449 516493 178505 516495
rect 178529 516493 178585 516495
rect 178609 516493 178665 516495
rect 178689 516493 178745 516495
rect 178449 516441 178495 516493
rect 178495 516441 178505 516493
rect 178529 516441 178559 516493
rect 178559 516441 178571 516493
rect 178571 516441 178585 516493
rect 178609 516441 178623 516493
rect 178623 516441 178635 516493
rect 178635 516441 178665 516493
rect 178689 516441 178699 516493
rect 178699 516441 178745 516493
rect 178449 516439 178505 516441
rect 178529 516439 178585 516441
rect 178609 516439 178665 516441
rect 178689 516439 178745 516441
rect 177789 515949 177845 515951
rect 177869 515949 177925 515951
rect 177949 515949 178005 515951
rect 178029 515949 178085 515951
rect 177789 515897 177835 515949
rect 177835 515897 177845 515949
rect 177869 515897 177899 515949
rect 177899 515897 177911 515949
rect 177911 515897 177925 515949
rect 177949 515897 177963 515949
rect 177963 515897 177975 515949
rect 177975 515897 178005 515949
rect 178029 515897 178039 515949
rect 178039 515897 178085 515949
rect 177789 515895 177845 515897
rect 177869 515895 177925 515897
rect 177949 515895 178005 515897
rect 178029 515895 178085 515897
rect 181607 527917 181663 527919
rect 181687 527917 181743 527919
rect 181767 527917 181823 527919
rect 181847 527917 181903 527919
rect 181607 527865 181653 527917
rect 181653 527865 181663 527917
rect 181687 527865 181717 527917
rect 181717 527865 181729 527917
rect 181729 527865 181743 527917
rect 181767 527865 181781 527917
rect 181781 527865 181793 527917
rect 181793 527865 181823 527917
rect 181847 527865 181857 527917
rect 181857 527865 181903 527917
rect 181607 527863 181663 527865
rect 181687 527863 181743 527865
rect 181767 527863 181823 527865
rect 181847 527863 181903 527865
rect 185425 527917 185481 527919
rect 185505 527917 185561 527919
rect 185585 527917 185641 527919
rect 185665 527917 185721 527919
rect 185425 527865 185471 527917
rect 185471 527865 185481 527917
rect 185505 527865 185535 527917
rect 185535 527865 185547 527917
rect 185547 527865 185561 527917
rect 185585 527865 185599 527917
rect 185599 527865 185611 527917
rect 185611 527865 185641 527917
rect 185665 527865 185675 527917
rect 185675 527865 185721 527917
rect 185425 527863 185481 527865
rect 185505 527863 185561 527865
rect 185585 527863 185641 527865
rect 185665 527863 185721 527865
rect 182267 527373 182323 527375
rect 182347 527373 182403 527375
rect 182427 527373 182483 527375
rect 182507 527373 182563 527375
rect 182267 527321 182313 527373
rect 182313 527321 182323 527373
rect 182347 527321 182377 527373
rect 182377 527321 182389 527373
rect 182389 527321 182403 527373
rect 182427 527321 182441 527373
rect 182441 527321 182453 527373
rect 182453 527321 182483 527373
rect 182507 527321 182517 527373
rect 182517 527321 182563 527373
rect 182267 527319 182323 527321
rect 182347 527319 182403 527321
rect 182427 527319 182483 527321
rect 182507 527319 182563 527321
rect 186085 527373 186141 527375
rect 186165 527373 186221 527375
rect 186245 527373 186301 527375
rect 186325 527373 186381 527375
rect 186085 527321 186131 527373
rect 186131 527321 186141 527373
rect 186165 527321 186195 527373
rect 186195 527321 186207 527373
rect 186207 527321 186221 527373
rect 186245 527321 186259 527373
rect 186259 527321 186271 527373
rect 186271 527321 186301 527373
rect 186325 527321 186335 527373
rect 186335 527321 186381 527373
rect 186085 527319 186141 527321
rect 186165 527319 186221 527321
rect 186245 527319 186301 527321
rect 186325 527319 186381 527321
rect 181607 526829 181663 526831
rect 181687 526829 181743 526831
rect 181767 526829 181823 526831
rect 181847 526829 181903 526831
rect 181607 526777 181653 526829
rect 181653 526777 181663 526829
rect 181687 526777 181717 526829
rect 181717 526777 181729 526829
rect 181729 526777 181743 526829
rect 181767 526777 181781 526829
rect 181781 526777 181793 526829
rect 181793 526777 181823 526829
rect 181847 526777 181857 526829
rect 181857 526777 181903 526829
rect 181607 526775 181663 526777
rect 181687 526775 181743 526777
rect 181767 526775 181823 526777
rect 181847 526775 181903 526777
rect 185425 526829 185481 526831
rect 185505 526829 185561 526831
rect 185585 526829 185641 526831
rect 185665 526829 185721 526831
rect 185425 526777 185471 526829
rect 185471 526777 185481 526829
rect 185505 526777 185535 526829
rect 185535 526777 185547 526829
rect 185547 526777 185561 526829
rect 185585 526777 185599 526829
rect 185599 526777 185611 526829
rect 185611 526777 185641 526829
rect 185665 526777 185675 526829
rect 185675 526777 185721 526829
rect 185425 526775 185481 526777
rect 185505 526775 185561 526777
rect 185585 526775 185641 526777
rect 185665 526775 185721 526777
rect 182267 526285 182323 526287
rect 182347 526285 182403 526287
rect 182427 526285 182483 526287
rect 182507 526285 182563 526287
rect 182267 526233 182313 526285
rect 182313 526233 182323 526285
rect 182347 526233 182377 526285
rect 182377 526233 182389 526285
rect 182389 526233 182403 526285
rect 182427 526233 182441 526285
rect 182441 526233 182453 526285
rect 182453 526233 182483 526285
rect 182507 526233 182517 526285
rect 182517 526233 182563 526285
rect 182267 526231 182323 526233
rect 182347 526231 182403 526233
rect 182427 526231 182483 526233
rect 182507 526231 182563 526233
rect 186085 526285 186141 526287
rect 186165 526285 186221 526287
rect 186245 526285 186301 526287
rect 186325 526285 186381 526287
rect 186085 526233 186131 526285
rect 186131 526233 186141 526285
rect 186165 526233 186195 526285
rect 186195 526233 186207 526285
rect 186207 526233 186221 526285
rect 186245 526233 186259 526285
rect 186259 526233 186271 526285
rect 186271 526233 186301 526285
rect 186325 526233 186335 526285
rect 186335 526233 186381 526285
rect 186085 526231 186141 526233
rect 186165 526231 186221 526233
rect 186245 526231 186301 526233
rect 186325 526231 186381 526233
rect 181607 525741 181663 525743
rect 181687 525741 181743 525743
rect 181767 525741 181823 525743
rect 181847 525741 181903 525743
rect 181607 525689 181653 525741
rect 181653 525689 181663 525741
rect 181687 525689 181717 525741
rect 181717 525689 181729 525741
rect 181729 525689 181743 525741
rect 181767 525689 181781 525741
rect 181781 525689 181793 525741
rect 181793 525689 181823 525741
rect 181847 525689 181857 525741
rect 181857 525689 181903 525741
rect 181607 525687 181663 525689
rect 181687 525687 181743 525689
rect 181767 525687 181823 525689
rect 181847 525687 181903 525689
rect 185425 525741 185481 525743
rect 185505 525741 185561 525743
rect 185585 525741 185641 525743
rect 185665 525741 185721 525743
rect 185425 525689 185471 525741
rect 185471 525689 185481 525741
rect 185505 525689 185535 525741
rect 185535 525689 185547 525741
rect 185547 525689 185561 525741
rect 185585 525689 185599 525741
rect 185599 525689 185611 525741
rect 185611 525689 185641 525741
rect 185665 525689 185675 525741
rect 185675 525689 185721 525741
rect 185425 525687 185481 525689
rect 185505 525687 185561 525689
rect 185585 525687 185641 525689
rect 185665 525687 185721 525689
rect 182267 525197 182323 525199
rect 182347 525197 182403 525199
rect 182427 525197 182483 525199
rect 182507 525197 182563 525199
rect 182267 525145 182313 525197
rect 182313 525145 182323 525197
rect 182347 525145 182377 525197
rect 182377 525145 182389 525197
rect 182389 525145 182403 525197
rect 182427 525145 182441 525197
rect 182441 525145 182453 525197
rect 182453 525145 182483 525197
rect 182507 525145 182517 525197
rect 182517 525145 182563 525197
rect 182267 525143 182323 525145
rect 182347 525143 182403 525145
rect 182427 525143 182483 525145
rect 182507 525143 182563 525145
rect 186085 525197 186141 525199
rect 186165 525197 186221 525199
rect 186245 525197 186301 525199
rect 186325 525197 186381 525199
rect 186085 525145 186131 525197
rect 186131 525145 186141 525197
rect 186165 525145 186195 525197
rect 186195 525145 186207 525197
rect 186207 525145 186221 525197
rect 186245 525145 186259 525197
rect 186259 525145 186271 525197
rect 186271 525145 186301 525197
rect 186325 525145 186335 525197
rect 186335 525145 186381 525197
rect 186085 525143 186141 525145
rect 186165 525143 186221 525145
rect 186245 525143 186301 525145
rect 186325 525143 186381 525145
rect 181607 524653 181663 524655
rect 181687 524653 181743 524655
rect 181767 524653 181823 524655
rect 181847 524653 181903 524655
rect 181607 524601 181653 524653
rect 181653 524601 181663 524653
rect 181687 524601 181717 524653
rect 181717 524601 181729 524653
rect 181729 524601 181743 524653
rect 181767 524601 181781 524653
rect 181781 524601 181793 524653
rect 181793 524601 181823 524653
rect 181847 524601 181857 524653
rect 181857 524601 181903 524653
rect 181607 524599 181663 524601
rect 181687 524599 181743 524601
rect 181767 524599 181823 524601
rect 181847 524599 181903 524601
rect 185425 524653 185481 524655
rect 185505 524653 185561 524655
rect 185585 524653 185641 524655
rect 185665 524653 185721 524655
rect 185425 524601 185471 524653
rect 185471 524601 185481 524653
rect 185505 524601 185535 524653
rect 185535 524601 185547 524653
rect 185547 524601 185561 524653
rect 185585 524601 185599 524653
rect 185599 524601 185611 524653
rect 185611 524601 185641 524653
rect 185665 524601 185675 524653
rect 185675 524601 185721 524653
rect 185425 524599 185481 524601
rect 185505 524599 185561 524601
rect 185585 524599 185641 524601
rect 185665 524599 185721 524601
rect 182267 524109 182323 524111
rect 182347 524109 182403 524111
rect 182427 524109 182483 524111
rect 182507 524109 182563 524111
rect 182267 524057 182313 524109
rect 182313 524057 182323 524109
rect 182347 524057 182377 524109
rect 182377 524057 182389 524109
rect 182389 524057 182403 524109
rect 182427 524057 182441 524109
rect 182441 524057 182453 524109
rect 182453 524057 182483 524109
rect 182507 524057 182517 524109
rect 182517 524057 182563 524109
rect 182267 524055 182323 524057
rect 182347 524055 182403 524057
rect 182427 524055 182483 524057
rect 182507 524055 182563 524057
rect 186085 524109 186141 524111
rect 186165 524109 186221 524111
rect 186245 524109 186301 524111
rect 186325 524109 186381 524111
rect 186085 524057 186131 524109
rect 186131 524057 186141 524109
rect 186165 524057 186195 524109
rect 186195 524057 186207 524109
rect 186207 524057 186221 524109
rect 186245 524057 186259 524109
rect 186259 524057 186271 524109
rect 186271 524057 186301 524109
rect 186325 524057 186335 524109
rect 186335 524057 186381 524109
rect 186085 524055 186141 524057
rect 186165 524055 186221 524057
rect 186245 524055 186301 524057
rect 186325 524055 186381 524057
rect 181607 523565 181663 523567
rect 181687 523565 181743 523567
rect 181767 523565 181823 523567
rect 181847 523565 181903 523567
rect 181607 523513 181653 523565
rect 181653 523513 181663 523565
rect 181687 523513 181717 523565
rect 181717 523513 181729 523565
rect 181729 523513 181743 523565
rect 181767 523513 181781 523565
rect 181781 523513 181793 523565
rect 181793 523513 181823 523565
rect 181847 523513 181857 523565
rect 181857 523513 181903 523565
rect 181607 523511 181663 523513
rect 181687 523511 181743 523513
rect 181767 523511 181823 523513
rect 181847 523511 181903 523513
rect 185425 523565 185481 523567
rect 185505 523565 185561 523567
rect 185585 523565 185641 523567
rect 185665 523565 185721 523567
rect 185425 523513 185471 523565
rect 185471 523513 185481 523565
rect 185505 523513 185535 523565
rect 185535 523513 185547 523565
rect 185547 523513 185561 523565
rect 185585 523513 185599 523565
rect 185599 523513 185611 523565
rect 185611 523513 185641 523565
rect 185665 523513 185675 523565
rect 185675 523513 185721 523565
rect 185425 523511 185481 523513
rect 185505 523511 185561 523513
rect 185585 523511 185641 523513
rect 185665 523511 185721 523513
rect 182267 523021 182323 523023
rect 182347 523021 182403 523023
rect 182427 523021 182483 523023
rect 182507 523021 182563 523023
rect 182267 522969 182313 523021
rect 182313 522969 182323 523021
rect 182347 522969 182377 523021
rect 182377 522969 182389 523021
rect 182389 522969 182403 523021
rect 182427 522969 182441 523021
rect 182441 522969 182453 523021
rect 182453 522969 182483 523021
rect 182507 522969 182517 523021
rect 182517 522969 182563 523021
rect 182267 522967 182323 522969
rect 182347 522967 182403 522969
rect 182427 522967 182483 522969
rect 182507 522967 182563 522969
rect 186085 523021 186141 523023
rect 186165 523021 186221 523023
rect 186245 523021 186301 523023
rect 186325 523021 186381 523023
rect 186085 522969 186131 523021
rect 186131 522969 186141 523021
rect 186165 522969 186195 523021
rect 186195 522969 186207 523021
rect 186207 522969 186221 523021
rect 186245 522969 186259 523021
rect 186259 522969 186271 523021
rect 186271 522969 186301 523021
rect 186325 522969 186335 523021
rect 186335 522969 186381 523021
rect 186085 522967 186141 522969
rect 186165 522967 186221 522969
rect 186245 522967 186301 522969
rect 186325 522967 186381 522969
rect 181607 522477 181663 522479
rect 181687 522477 181743 522479
rect 181767 522477 181823 522479
rect 181847 522477 181903 522479
rect 181607 522425 181653 522477
rect 181653 522425 181663 522477
rect 181687 522425 181717 522477
rect 181717 522425 181729 522477
rect 181729 522425 181743 522477
rect 181767 522425 181781 522477
rect 181781 522425 181793 522477
rect 181793 522425 181823 522477
rect 181847 522425 181857 522477
rect 181857 522425 181903 522477
rect 181607 522423 181663 522425
rect 181687 522423 181743 522425
rect 181767 522423 181823 522425
rect 181847 522423 181903 522425
rect 185425 522477 185481 522479
rect 185505 522477 185561 522479
rect 185585 522477 185641 522479
rect 185665 522477 185721 522479
rect 185425 522425 185471 522477
rect 185471 522425 185481 522477
rect 185505 522425 185535 522477
rect 185535 522425 185547 522477
rect 185547 522425 185561 522477
rect 185585 522425 185599 522477
rect 185599 522425 185611 522477
rect 185611 522425 185641 522477
rect 185665 522425 185675 522477
rect 185675 522425 185721 522477
rect 185425 522423 185481 522425
rect 185505 522423 185561 522425
rect 185585 522423 185641 522425
rect 185665 522423 185721 522425
rect 182267 521933 182323 521935
rect 182347 521933 182403 521935
rect 182427 521933 182483 521935
rect 182507 521933 182563 521935
rect 182267 521881 182313 521933
rect 182313 521881 182323 521933
rect 182347 521881 182377 521933
rect 182377 521881 182389 521933
rect 182389 521881 182403 521933
rect 182427 521881 182441 521933
rect 182441 521881 182453 521933
rect 182453 521881 182483 521933
rect 182507 521881 182517 521933
rect 182517 521881 182563 521933
rect 182267 521879 182323 521881
rect 182347 521879 182403 521881
rect 182427 521879 182483 521881
rect 182507 521879 182563 521881
rect 186085 521933 186141 521935
rect 186165 521933 186221 521935
rect 186245 521933 186301 521935
rect 186325 521933 186381 521935
rect 186085 521881 186131 521933
rect 186131 521881 186141 521933
rect 186165 521881 186195 521933
rect 186195 521881 186207 521933
rect 186207 521881 186221 521933
rect 186245 521881 186259 521933
rect 186259 521881 186271 521933
rect 186271 521881 186301 521933
rect 186325 521881 186335 521933
rect 186335 521881 186381 521933
rect 186085 521879 186141 521881
rect 186165 521879 186221 521881
rect 186245 521879 186301 521881
rect 186325 521879 186381 521881
rect 181607 521389 181663 521391
rect 181687 521389 181743 521391
rect 181767 521389 181823 521391
rect 181847 521389 181903 521391
rect 181607 521337 181653 521389
rect 181653 521337 181663 521389
rect 181687 521337 181717 521389
rect 181717 521337 181729 521389
rect 181729 521337 181743 521389
rect 181767 521337 181781 521389
rect 181781 521337 181793 521389
rect 181793 521337 181823 521389
rect 181847 521337 181857 521389
rect 181857 521337 181903 521389
rect 181607 521335 181663 521337
rect 181687 521335 181743 521337
rect 181767 521335 181823 521337
rect 181847 521335 181903 521337
rect 185425 521389 185481 521391
rect 185505 521389 185561 521391
rect 185585 521389 185641 521391
rect 185665 521389 185721 521391
rect 185425 521337 185471 521389
rect 185471 521337 185481 521389
rect 185505 521337 185535 521389
rect 185535 521337 185547 521389
rect 185547 521337 185561 521389
rect 185585 521337 185599 521389
rect 185599 521337 185611 521389
rect 185611 521337 185641 521389
rect 185665 521337 185675 521389
rect 185675 521337 185721 521389
rect 185425 521335 185481 521337
rect 185505 521335 185561 521337
rect 185585 521335 185641 521337
rect 185665 521335 185721 521337
rect 182267 520845 182323 520847
rect 182347 520845 182403 520847
rect 182427 520845 182483 520847
rect 182507 520845 182563 520847
rect 182267 520793 182313 520845
rect 182313 520793 182323 520845
rect 182347 520793 182377 520845
rect 182377 520793 182389 520845
rect 182389 520793 182403 520845
rect 182427 520793 182441 520845
rect 182441 520793 182453 520845
rect 182453 520793 182483 520845
rect 182507 520793 182517 520845
rect 182517 520793 182563 520845
rect 182267 520791 182323 520793
rect 182347 520791 182403 520793
rect 182427 520791 182483 520793
rect 182507 520791 182563 520793
rect 186085 520845 186141 520847
rect 186165 520845 186221 520847
rect 186245 520845 186301 520847
rect 186325 520845 186381 520847
rect 186085 520793 186131 520845
rect 186131 520793 186141 520845
rect 186165 520793 186195 520845
rect 186195 520793 186207 520845
rect 186207 520793 186221 520845
rect 186245 520793 186259 520845
rect 186259 520793 186271 520845
rect 186271 520793 186301 520845
rect 186325 520793 186335 520845
rect 186335 520793 186381 520845
rect 186085 520791 186141 520793
rect 186165 520791 186221 520793
rect 186245 520791 186301 520793
rect 186325 520791 186381 520793
rect 181607 520301 181663 520303
rect 181687 520301 181743 520303
rect 181767 520301 181823 520303
rect 181847 520301 181903 520303
rect 181607 520249 181653 520301
rect 181653 520249 181663 520301
rect 181687 520249 181717 520301
rect 181717 520249 181729 520301
rect 181729 520249 181743 520301
rect 181767 520249 181781 520301
rect 181781 520249 181793 520301
rect 181793 520249 181823 520301
rect 181847 520249 181857 520301
rect 181857 520249 181903 520301
rect 181607 520247 181663 520249
rect 181687 520247 181743 520249
rect 181767 520247 181823 520249
rect 181847 520247 181903 520249
rect 185425 520301 185481 520303
rect 185505 520301 185561 520303
rect 185585 520301 185641 520303
rect 185665 520301 185721 520303
rect 185425 520249 185471 520301
rect 185471 520249 185481 520301
rect 185505 520249 185535 520301
rect 185535 520249 185547 520301
rect 185547 520249 185561 520301
rect 185585 520249 185599 520301
rect 185599 520249 185611 520301
rect 185611 520249 185641 520301
rect 185665 520249 185675 520301
rect 185675 520249 185721 520301
rect 185425 520247 185481 520249
rect 185505 520247 185561 520249
rect 185585 520247 185641 520249
rect 185665 520247 185721 520249
rect 182267 519757 182323 519759
rect 182347 519757 182403 519759
rect 182427 519757 182483 519759
rect 182507 519757 182563 519759
rect 182267 519705 182313 519757
rect 182313 519705 182323 519757
rect 182347 519705 182377 519757
rect 182377 519705 182389 519757
rect 182389 519705 182403 519757
rect 182427 519705 182441 519757
rect 182441 519705 182453 519757
rect 182453 519705 182483 519757
rect 182507 519705 182517 519757
rect 182517 519705 182563 519757
rect 182267 519703 182323 519705
rect 182347 519703 182403 519705
rect 182427 519703 182483 519705
rect 182507 519703 182563 519705
rect 186085 519757 186141 519759
rect 186165 519757 186221 519759
rect 186245 519757 186301 519759
rect 186325 519757 186381 519759
rect 186085 519705 186131 519757
rect 186131 519705 186141 519757
rect 186165 519705 186195 519757
rect 186195 519705 186207 519757
rect 186207 519705 186221 519757
rect 186245 519705 186259 519757
rect 186259 519705 186271 519757
rect 186271 519705 186301 519757
rect 186325 519705 186335 519757
rect 186335 519705 186381 519757
rect 186085 519703 186141 519705
rect 186165 519703 186221 519705
rect 186245 519703 186301 519705
rect 186325 519703 186381 519705
rect 181607 519213 181663 519215
rect 181687 519213 181743 519215
rect 181767 519213 181823 519215
rect 181847 519213 181903 519215
rect 181607 519161 181653 519213
rect 181653 519161 181663 519213
rect 181687 519161 181717 519213
rect 181717 519161 181729 519213
rect 181729 519161 181743 519213
rect 181767 519161 181781 519213
rect 181781 519161 181793 519213
rect 181793 519161 181823 519213
rect 181847 519161 181857 519213
rect 181857 519161 181903 519213
rect 181607 519159 181663 519161
rect 181687 519159 181743 519161
rect 181767 519159 181823 519161
rect 181847 519159 181903 519161
rect 185425 519213 185481 519215
rect 185505 519213 185561 519215
rect 185585 519213 185641 519215
rect 185665 519213 185721 519215
rect 185425 519161 185471 519213
rect 185471 519161 185481 519213
rect 185505 519161 185535 519213
rect 185535 519161 185547 519213
rect 185547 519161 185561 519213
rect 185585 519161 185599 519213
rect 185599 519161 185611 519213
rect 185611 519161 185641 519213
rect 185665 519161 185675 519213
rect 185675 519161 185721 519213
rect 185425 519159 185481 519161
rect 185505 519159 185561 519161
rect 185585 519159 185641 519161
rect 185665 519159 185721 519161
rect 182267 518669 182323 518671
rect 182347 518669 182403 518671
rect 182427 518669 182483 518671
rect 182507 518669 182563 518671
rect 182267 518617 182313 518669
rect 182313 518617 182323 518669
rect 182347 518617 182377 518669
rect 182377 518617 182389 518669
rect 182389 518617 182403 518669
rect 182427 518617 182441 518669
rect 182441 518617 182453 518669
rect 182453 518617 182483 518669
rect 182507 518617 182517 518669
rect 182517 518617 182563 518669
rect 182267 518615 182323 518617
rect 182347 518615 182403 518617
rect 182427 518615 182483 518617
rect 182507 518615 182563 518617
rect 186085 518669 186141 518671
rect 186165 518669 186221 518671
rect 186245 518669 186301 518671
rect 186325 518669 186381 518671
rect 186085 518617 186131 518669
rect 186131 518617 186141 518669
rect 186165 518617 186195 518669
rect 186195 518617 186207 518669
rect 186207 518617 186221 518669
rect 186245 518617 186259 518669
rect 186259 518617 186271 518669
rect 186271 518617 186301 518669
rect 186325 518617 186335 518669
rect 186335 518617 186381 518669
rect 186085 518615 186141 518617
rect 186165 518615 186221 518617
rect 186245 518615 186301 518617
rect 186325 518615 186381 518617
rect 181607 518125 181663 518127
rect 181687 518125 181743 518127
rect 181767 518125 181823 518127
rect 181847 518125 181903 518127
rect 181607 518073 181653 518125
rect 181653 518073 181663 518125
rect 181687 518073 181717 518125
rect 181717 518073 181729 518125
rect 181729 518073 181743 518125
rect 181767 518073 181781 518125
rect 181781 518073 181793 518125
rect 181793 518073 181823 518125
rect 181847 518073 181857 518125
rect 181857 518073 181903 518125
rect 181607 518071 181663 518073
rect 181687 518071 181743 518073
rect 181767 518071 181823 518073
rect 181847 518071 181903 518073
rect 185425 518125 185481 518127
rect 185505 518125 185561 518127
rect 185585 518125 185641 518127
rect 185665 518125 185721 518127
rect 185425 518073 185471 518125
rect 185471 518073 185481 518125
rect 185505 518073 185535 518125
rect 185535 518073 185547 518125
rect 185547 518073 185561 518125
rect 185585 518073 185599 518125
rect 185599 518073 185611 518125
rect 185611 518073 185641 518125
rect 185665 518073 185675 518125
rect 185675 518073 185721 518125
rect 185425 518071 185481 518073
rect 185505 518071 185561 518073
rect 185585 518071 185641 518073
rect 185665 518071 185721 518073
rect 182267 517581 182323 517583
rect 182347 517581 182403 517583
rect 182427 517581 182483 517583
rect 182507 517581 182563 517583
rect 182267 517529 182313 517581
rect 182313 517529 182323 517581
rect 182347 517529 182377 517581
rect 182377 517529 182389 517581
rect 182389 517529 182403 517581
rect 182427 517529 182441 517581
rect 182441 517529 182453 517581
rect 182453 517529 182483 517581
rect 182507 517529 182517 517581
rect 182517 517529 182563 517581
rect 182267 517527 182323 517529
rect 182347 517527 182403 517529
rect 182427 517527 182483 517529
rect 182507 517527 182563 517529
rect 186085 517581 186141 517583
rect 186165 517581 186221 517583
rect 186245 517581 186301 517583
rect 186325 517581 186381 517583
rect 186085 517529 186131 517581
rect 186131 517529 186141 517581
rect 186165 517529 186195 517581
rect 186195 517529 186207 517581
rect 186207 517529 186221 517581
rect 186245 517529 186259 517581
rect 186259 517529 186271 517581
rect 186271 517529 186301 517581
rect 186325 517529 186335 517581
rect 186335 517529 186381 517581
rect 186085 517527 186141 517529
rect 186165 517527 186221 517529
rect 186245 517527 186301 517529
rect 186325 517527 186381 517529
rect 181607 517037 181663 517039
rect 181687 517037 181743 517039
rect 181767 517037 181823 517039
rect 181847 517037 181903 517039
rect 181607 516985 181653 517037
rect 181653 516985 181663 517037
rect 181687 516985 181717 517037
rect 181717 516985 181729 517037
rect 181729 516985 181743 517037
rect 181767 516985 181781 517037
rect 181781 516985 181793 517037
rect 181793 516985 181823 517037
rect 181847 516985 181857 517037
rect 181857 516985 181903 517037
rect 181607 516983 181663 516985
rect 181687 516983 181743 516985
rect 181767 516983 181823 516985
rect 181847 516983 181903 516985
rect 185425 517037 185481 517039
rect 185505 517037 185561 517039
rect 185585 517037 185641 517039
rect 185665 517037 185721 517039
rect 185425 516985 185471 517037
rect 185471 516985 185481 517037
rect 185505 516985 185535 517037
rect 185535 516985 185547 517037
rect 185547 516985 185561 517037
rect 185585 516985 185599 517037
rect 185599 516985 185611 517037
rect 185611 516985 185641 517037
rect 185665 516985 185675 517037
rect 185675 516985 185721 517037
rect 185425 516983 185481 516985
rect 185505 516983 185561 516985
rect 185585 516983 185641 516985
rect 185665 516983 185721 516985
rect 182267 516493 182323 516495
rect 182347 516493 182403 516495
rect 182427 516493 182483 516495
rect 182507 516493 182563 516495
rect 182267 516441 182313 516493
rect 182313 516441 182323 516493
rect 182347 516441 182377 516493
rect 182377 516441 182389 516493
rect 182389 516441 182403 516493
rect 182427 516441 182441 516493
rect 182441 516441 182453 516493
rect 182453 516441 182483 516493
rect 182507 516441 182517 516493
rect 182517 516441 182563 516493
rect 182267 516439 182323 516441
rect 182347 516439 182403 516441
rect 182427 516439 182483 516441
rect 182507 516439 182563 516441
rect 186085 516493 186141 516495
rect 186165 516493 186221 516495
rect 186245 516493 186301 516495
rect 186325 516493 186381 516495
rect 186085 516441 186131 516493
rect 186131 516441 186141 516493
rect 186165 516441 186195 516493
rect 186195 516441 186207 516493
rect 186207 516441 186221 516493
rect 186245 516441 186259 516493
rect 186259 516441 186271 516493
rect 186271 516441 186301 516493
rect 186325 516441 186335 516493
rect 186335 516441 186381 516493
rect 186085 516439 186141 516441
rect 186165 516439 186221 516441
rect 186245 516439 186301 516441
rect 186325 516439 186381 516441
rect 181607 515949 181663 515951
rect 181687 515949 181743 515951
rect 181767 515949 181823 515951
rect 181847 515949 181903 515951
rect 181607 515897 181653 515949
rect 181653 515897 181663 515949
rect 181687 515897 181717 515949
rect 181717 515897 181729 515949
rect 181729 515897 181743 515949
rect 181767 515897 181781 515949
rect 181781 515897 181793 515949
rect 181793 515897 181823 515949
rect 181847 515897 181857 515949
rect 181857 515897 181903 515949
rect 181607 515895 181663 515897
rect 181687 515895 181743 515897
rect 181767 515895 181823 515897
rect 181847 515895 181903 515897
rect 185425 515949 185481 515951
rect 185505 515949 185561 515951
rect 185585 515949 185641 515951
rect 185665 515949 185721 515951
rect 185425 515897 185471 515949
rect 185471 515897 185481 515949
rect 185505 515897 185535 515949
rect 185535 515897 185547 515949
rect 185547 515897 185561 515949
rect 185585 515897 185599 515949
rect 185599 515897 185611 515949
rect 185611 515897 185641 515949
rect 185665 515897 185675 515949
rect 185675 515897 185721 515949
rect 185425 515895 185481 515897
rect 185505 515895 185561 515897
rect 185585 515895 185641 515897
rect 185665 515895 185721 515897
rect 178449 515405 178505 515407
rect 178529 515405 178585 515407
rect 178609 515405 178665 515407
rect 178689 515405 178745 515407
rect 178449 515353 178495 515405
rect 178495 515353 178505 515405
rect 178529 515353 178559 515405
rect 178559 515353 178571 515405
rect 178571 515353 178585 515405
rect 178609 515353 178623 515405
rect 178623 515353 178635 515405
rect 178635 515353 178665 515405
rect 178689 515353 178699 515405
rect 178699 515353 178745 515405
rect 178449 515351 178505 515353
rect 178529 515351 178585 515353
rect 178609 515351 178665 515353
rect 178689 515351 178745 515353
rect 182267 515405 182323 515407
rect 182347 515405 182403 515407
rect 182427 515405 182483 515407
rect 182507 515405 182563 515407
rect 182267 515353 182313 515405
rect 182313 515353 182323 515405
rect 182347 515353 182377 515405
rect 182377 515353 182389 515405
rect 182389 515353 182403 515405
rect 182427 515353 182441 515405
rect 182441 515353 182453 515405
rect 182453 515353 182483 515405
rect 182507 515353 182517 515405
rect 182517 515353 182563 515405
rect 182267 515351 182323 515353
rect 182347 515351 182403 515353
rect 182427 515351 182483 515353
rect 182507 515351 182563 515353
rect 186085 515405 186141 515407
rect 186165 515405 186221 515407
rect 186245 515405 186301 515407
rect 186325 515405 186381 515407
rect 186085 515353 186131 515405
rect 186131 515353 186141 515405
rect 186165 515353 186195 515405
rect 186195 515353 186207 515405
rect 186207 515353 186221 515405
rect 186245 515353 186259 515405
rect 186259 515353 186271 515405
rect 186271 515353 186301 515405
rect 186325 515353 186335 515405
rect 186335 515353 186381 515405
rect 186085 515351 186141 515353
rect 186165 515351 186221 515353
rect 186245 515351 186301 515353
rect 186325 515351 186381 515353
rect 2000 507000 4000 509000
rect 2000 464000 4000 466000
rect 2000 421000 4000 423000
rect 2000 378430 4000 380000
rect 2014 378318 4000 378430
rect 2000 378000 4000 378318
<< metal3 >>
rect 16194 701000 21194 703400
rect 16194 700900 18000 701000
rect 17990 699000 18000 700900
rect 20000 700900 21194 701000
rect 68194 701000 73194 703400
rect 68194 700900 70000 701000
rect 20000 699000 20010 700900
rect 17990 698995 20010 699000
rect 69990 699000 70000 700900
rect 72000 700900 73194 701000
rect 120194 701000 125194 703400
rect 120194 700900 122000 701000
rect 72000 699000 72010 700900
rect 69990 698995 72010 699000
rect 121990 699000 122000 700900
rect 124000 700900 125194 701000
rect 124000 699000 124010 700900
rect 121990 698995 124010 699000
rect 600 684005 3100 685242
rect 600 684000 5010 684005
rect 600 682000 3000 684000
rect 5000 682000 5010 684000
rect 600 681995 5010 682000
rect 600 680242 3100 681995
rect 157611 541869 162710 541897
rect 157611 538925 162626 541869
rect 162690 538925 162710 541869
rect 157611 538897 162710 538925
rect 163120 540287 192000 540297
rect 163120 540277 174190 540287
rect 163120 540097 166690 540277
rect 166870 540097 170490 540277
rect 170670 540107 174190 540277
rect 174370 540277 192000 540287
rect 174370 540107 177700 540277
rect 170670 540097 177700 540107
rect 177880 540097 181290 540277
rect 181470 540097 184590 540277
rect 184770 540097 187900 540277
rect 188080 540097 191190 540277
rect 191370 540097 191810 540277
rect 191990 540097 192000 540277
rect 163120 540077 192000 540097
rect 163120 538902 163340 540077
rect 163020 538897 163340 538902
rect 161380 538697 161530 538707
rect 159390 538687 159490 538697
rect 159390 538587 159400 538687
rect 159480 538587 159490 538687
rect 159390 538577 159490 538587
rect 161380 538577 161390 538697
rect 161510 538577 161530 538697
rect 163020 538697 163030 538897
rect 163330 538697 163340 538897
rect 163020 538692 163340 538697
rect 163120 538587 163340 538692
rect 163900 539347 192010 539357
rect 163900 539337 191200 539347
rect 163900 539157 166690 539337
rect 166870 539157 170490 539337
rect 170670 539157 174190 539337
rect 174370 539157 177690 539337
rect 177870 539157 181290 539337
rect 181470 539157 184590 539337
rect 184770 539157 187890 539337
rect 188070 539167 191200 539337
rect 191380 539337 192010 539347
rect 191380 539167 191820 539337
rect 188070 539157 191820 539167
rect 192000 539157 192010 539337
rect 163900 539137 192010 539157
rect 161380 538567 161530 538577
rect 163900 535657 164120 539137
rect 160200 535597 164120 535657
rect 160200 535457 160210 535597
rect 160360 535457 164120 535597
rect 160200 535437 164120 535457
rect 174621 530643 174937 530644
rect 174621 530579 174627 530643
rect 174691 530579 174707 530643
rect 174771 530579 174787 530643
rect 174851 530579 174867 530643
rect 174931 530579 174937 530643
rect 174621 530578 174937 530579
rect 178439 530643 178755 530644
rect 178439 530579 178445 530643
rect 178509 530579 178525 530643
rect 178589 530579 178605 530643
rect 178669 530579 178685 530643
rect 178749 530579 178755 530643
rect 178439 530578 178755 530579
rect 182257 530643 182573 530644
rect 182257 530579 182263 530643
rect 182327 530579 182343 530643
rect 182407 530579 182423 530643
rect 182487 530579 182503 530643
rect 182567 530579 182573 530643
rect 182257 530578 182573 530579
rect 186075 530643 186391 530644
rect 186075 530579 186081 530643
rect 186145 530579 186161 530643
rect 186225 530579 186241 530643
rect 186305 530579 186321 530643
rect 186385 530579 186391 530643
rect 186075 530578 186391 530579
rect 173961 530099 174277 530100
rect 173961 530035 173967 530099
rect 174031 530035 174047 530099
rect 174111 530035 174127 530099
rect 174191 530035 174207 530099
rect 174271 530035 174277 530099
rect 173961 530034 174277 530035
rect 177779 530099 178095 530100
rect 177779 530035 177785 530099
rect 177849 530035 177865 530099
rect 177929 530035 177945 530099
rect 178009 530035 178025 530099
rect 178089 530035 178095 530099
rect 177779 530034 178095 530035
rect 181597 530099 181913 530100
rect 181597 530035 181603 530099
rect 181667 530035 181683 530099
rect 181747 530035 181763 530099
rect 181827 530035 181843 530099
rect 181907 530035 181913 530099
rect 181597 530034 181913 530035
rect 185415 530099 185731 530100
rect 185415 530035 185421 530099
rect 185485 530035 185501 530099
rect 185565 530035 185581 530099
rect 185645 530035 185661 530099
rect 185725 530035 185731 530099
rect 185415 530034 185731 530035
rect 174621 529555 174937 529556
rect 174621 529491 174627 529555
rect 174691 529491 174707 529555
rect 174771 529491 174787 529555
rect 174851 529491 174867 529555
rect 174931 529491 174937 529555
rect 174621 529490 174937 529491
rect 178439 529555 178755 529556
rect 178439 529491 178445 529555
rect 178509 529491 178525 529555
rect 178589 529491 178605 529555
rect 178669 529491 178685 529555
rect 178749 529491 178755 529555
rect 178439 529490 178755 529491
rect 182257 529555 182573 529556
rect 182257 529491 182263 529555
rect 182327 529491 182343 529555
rect 182407 529491 182423 529555
rect 182487 529491 182503 529555
rect 182567 529491 182573 529555
rect 182257 529490 182573 529491
rect 186075 529555 186391 529556
rect 186075 529491 186081 529555
rect 186145 529491 186161 529555
rect 186225 529491 186241 529555
rect 186305 529491 186321 529555
rect 186385 529491 186391 529555
rect 186075 529490 186391 529491
rect 173961 529011 174277 529012
rect 173961 528947 173967 529011
rect 174031 528947 174047 529011
rect 174111 528947 174127 529011
rect 174191 528947 174207 529011
rect 174271 528947 174277 529011
rect 173961 528946 174277 528947
rect 177779 529011 178095 529012
rect 177779 528947 177785 529011
rect 177849 528947 177865 529011
rect 177929 528947 177945 529011
rect 178009 528947 178025 529011
rect 178089 528947 178095 529011
rect 177779 528946 178095 528947
rect 181597 529011 181913 529012
rect 181597 528947 181603 529011
rect 181667 528947 181683 529011
rect 181747 528947 181763 529011
rect 181827 528947 181843 529011
rect 181907 528947 181913 529011
rect 181597 528946 181913 528947
rect 185415 529011 185731 529012
rect 185415 528947 185421 529011
rect 185485 528947 185501 529011
rect 185565 528947 185581 529011
rect 185645 528947 185661 529011
rect 185725 528947 185731 529011
rect 185415 528946 185731 528947
rect 174621 528467 174937 528468
rect 174621 528403 174627 528467
rect 174691 528403 174707 528467
rect 174771 528403 174787 528467
rect 174851 528403 174867 528467
rect 174931 528403 174937 528467
rect 174621 528402 174937 528403
rect 178439 528467 178755 528468
rect 178439 528403 178445 528467
rect 178509 528403 178525 528467
rect 178589 528403 178605 528467
rect 178669 528403 178685 528467
rect 178749 528403 178755 528467
rect 178439 528402 178755 528403
rect 182257 528467 182573 528468
rect 182257 528403 182263 528467
rect 182327 528403 182343 528467
rect 182407 528403 182423 528467
rect 182487 528403 182503 528467
rect 182567 528403 182573 528467
rect 182257 528402 182573 528403
rect 186075 528467 186391 528468
rect 186075 528403 186081 528467
rect 186145 528403 186161 528467
rect 186225 528403 186241 528467
rect 186305 528403 186321 528467
rect 186385 528403 186391 528467
rect 186075 528402 186391 528403
rect 173961 527923 174277 527924
rect 173961 527859 173967 527923
rect 174031 527859 174047 527923
rect 174111 527859 174127 527923
rect 174191 527859 174207 527923
rect 174271 527859 174277 527923
rect 173961 527858 174277 527859
rect 177779 527923 178095 527924
rect 177779 527859 177785 527923
rect 177849 527859 177865 527923
rect 177929 527859 177945 527923
rect 178009 527859 178025 527923
rect 178089 527859 178095 527923
rect 177779 527858 178095 527859
rect 181597 527923 181913 527924
rect 181597 527859 181603 527923
rect 181667 527859 181683 527923
rect 181747 527859 181763 527923
rect 181827 527859 181843 527923
rect 181907 527859 181913 527923
rect 181597 527858 181913 527859
rect 185415 527923 185731 527924
rect 185415 527859 185421 527923
rect 185485 527859 185501 527923
rect 185565 527859 185581 527923
rect 185645 527859 185661 527923
rect 185725 527859 185731 527923
rect 185415 527858 185731 527859
rect 174621 527379 174937 527380
rect 174621 527315 174627 527379
rect 174691 527315 174707 527379
rect 174771 527315 174787 527379
rect 174851 527315 174867 527379
rect 174931 527315 174937 527379
rect 174621 527314 174937 527315
rect 178439 527379 178755 527380
rect 178439 527315 178445 527379
rect 178509 527315 178525 527379
rect 178589 527315 178605 527379
rect 178669 527315 178685 527379
rect 178749 527315 178755 527379
rect 178439 527314 178755 527315
rect 182257 527379 182573 527380
rect 182257 527315 182263 527379
rect 182327 527315 182343 527379
rect 182407 527315 182423 527379
rect 182487 527315 182503 527379
rect 182567 527315 182573 527379
rect 182257 527314 182573 527315
rect 186075 527379 186391 527380
rect 186075 527315 186081 527379
rect 186145 527315 186161 527379
rect 186225 527315 186241 527379
rect 186305 527315 186321 527379
rect 186385 527315 186391 527379
rect 186075 527314 186391 527315
rect 173961 526835 174277 526836
rect 173961 526771 173967 526835
rect 174031 526771 174047 526835
rect 174111 526771 174127 526835
rect 174191 526771 174207 526835
rect 174271 526771 174277 526835
rect 173961 526770 174277 526771
rect 177779 526835 178095 526836
rect 177779 526771 177785 526835
rect 177849 526771 177865 526835
rect 177929 526771 177945 526835
rect 178009 526771 178025 526835
rect 178089 526771 178095 526835
rect 177779 526770 178095 526771
rect 181597 526835 181913 526836
rect 181597 526771 181603 526835
rect 181667 526771 181683 526835
rect 181747 526771 181763 526835
rect 181827 526771 181843 526835
rect 181907 526771 181913 526835
rect 181597 526770 181913 526771
rect 185415 526835 185731 526836
rect 185415 526771 185421 526835
rect 185485 526771 185501 526835
rect 185565 526771 185581 526835
rect 185645 526771 185661 526835
rect 185725 526771 185731 526835
rect 185415 526770 185731 526771
rect 174621 526291 174937 526292
rect 174621 526227 174627 526291
rect 174691 526227 174707 526291
rect 174771 526227 174787 526291
rect 174851 526227 174867 526291
rect 174931 526227 174937 526291
rect 174621 526226 174937 526227
rect 178439 526291 178755 526292
rect 178439 526227 178445 526291
rect 178509 526227 178525 526291
rect 178589 526227 178605 526291
rect 178669 526227 178685 526291
rect 178749 526227 178755 526291
rect 178439 526226 178755 526227
rect 182257 526291 182573 526292
rect 182257 526227 182263 526291
rect 182327 526227 182343 526291
rect 182407 526227 182423 526291
rect 182487 526227 182503 526291
rect 182567 526227 182573 526291
rect 182257 526226 182573 526227
rect 186075 526291 186391 526292
rect 186075 526227 186081 526291
rect 186145 526227 186161 526291
rect 186225 526227 186241 526291
rect 186305 526227 186321 526291
rect 186385 526227 186391 526291
rect 186075 526226 186391 526227
rect 173961 525747 174277 525748
rect 173961 525683 173967 525747
rect 174031 525683 174047 525747
rect 174111 525683 174127 525747
rect 174191 525683 174207 525747
rect 174271 525683 174277 525747
rect 173961 525682 174277 525683
rect 177779 525747 178095 525748
rect 177779 525683 177785 525747
rect 177849 525683 177865 525747
rect 177929 525683 177945 525747
rect 178009 525683 178025 525747
rect 178089 525683 178095 525747
rect 177779 525682 178095 525683
rect 181597 525747 181913 525748
rect 181597 525683 181603 525747
rect 181667 525683 181683 525747
rect 181747 525683 181763 525747
rect 181827 525683 181843 525747
rect 181907 525683 181913 525747
rect 181597 525682 181913 525683
rect 185415 525747 185731 525748
rect 185415 525683 185421 525747
rect 185485 525683 185501 525747
rect 185565 525683 185581 525747
rect 185645 525683 185661 525747
rect 185725 525683 185731 525747
rect 185415 525682 185731 525683
rect 174621 525203 174937 525204
rect 174621 525139 174627 525203
rect 174691 525139 174707 525203
rect 174771 525139 174787 525203
rect 174851 525139 174867 525203
rect 174931 525139 174937 525203
rect 174621 525138 174937 525139
rect 178439 525203 178755 525204
rect 178439 525139 178445 525203
rect 178509 525139 178525 525203
rect 178589 525139 178605 525203
rect 178669 525139 178685 525203
rect 178749 525139 178755 525203
rect 178439 525138 178755 525139
rect 182257 525203 182573 525204
rect 182257 525139 182263 525203
rect 182327 525139 182343 525203
rect 182407 525139 182423 525203
rect 182487 525139 182503 525203
rect 182567 525139 182573 525203
rect 182257 525138 182573 525139
rect 186075 525203 186391 525204
rect 186075 525139 186081 525203
rect 186145 525139 186161 525203
rect 186225 525139 186241 525203
rect 186305 525139 186321 525203
rect 186385 525139 186391 525203
rect 186075 525138 186391 525139
rect 173961 524659 174277 524660
rect 173961 524595 173967 524659
rect 174031 524595 174047 524659
rect 174111 524595 174127 524659
rect 174191 524595 174207 524659
rect 174271 524595 174277 524659
rect 173961 524594 174277 524595
rect 177779 524659 178095 524660
rect 177779 524595 177785 524659
rect 177849 524595 177865 524659
rect 177929 524595 177945 524659
rect 178009 524595 178025 524659
rect 178089 524595 178095 524659
rect 177779 524594 178095 524595
rect 181597 524659 181913 524660
rect 181597 524595 181603 524659
rect 181667 524595 181683 524659
rect 181747 524595 181763 524659
rect 181827 524595 181843 524659
rect 181907 524595 181913 524659
rect 181597 524594 181913 524595
rect 185415 524659 185731 524660
rect 185415 524595 185421 524659
rect 185485 524595 185501 524659
rect 185565 524595 185581 524659
rect 185645 524595 185661 524659
rect 185725 524595 185731 524659
rect 185415 524594 185731 524595
rect 174621 524115 174937 524116
rect 174621 524051 174627 524115
rect 174691 524051 174707 524115
rect 174771 524051 174787 524115
rect 174851 524051 174867 524115
rect 174931 524051 174937 524115
rect 174621 524050 174937 524051
rect 178439 524115 178755 524116
rect 178439 524051 178445 524115
rect 178509 524051 178525 524115
rect 178589 524051 178605 524115
rect 178669 524051 178685 524115
rect 178749 524051 178755 524115
rect 178439 524050 178755 524051
rect 182257 524115 182573 524116
rect 182257 524051 182263 524115
rect 182327 524051 182343 524115
rect 182407 524051 182423 524115
rect 182487 524051 182503 524115
rect 182567 524051 182573 524115
rect 182257 524050 182573 524051
rect 186075 524115 186391 524116
rect 186075 524051 186081 524115
rect 186145 524051 186161 524115
rect 186225 524051 186241 524115
rect 186305 524051 186321 524115
rect 186385 524051 186391 524115
rect 186075 524050 186391 524051
rect 173961 523571 174277 523572
rect 173961 523507 173967 523571
rect 174031 523507 174047 523571
rect 174111 523507 174127 523571
rect 174191 523507 174207 523571
rect 174271 523507 174277 523571
rect 173961 523506 174277 523507
rect 177779 523571 178095 523572
rect 177779 523507 177785 523571
rect 177849 523507 177865 523571
rect 177929 523507 177945 523571
rect 178009 523507 178025 523571
rect 178089 523507 178095 523571
rect 177779 523506 178095 523507
rect 181597 523571 181913 523572
rect 181597 523507 181603 523571
rect 181667 523507 181683 523571
rect 181747 523507 181763 523571
rect 181827 523507 181843 523571
rect 181907 523507 181913 523571
rect 181597 523506 181913 523507
rect 185415 523571 185731 523572
rect 185415 523507 185421 523571
rect 185485 523507 185501 523571
rect 185565 523507 185581 523571
rect 185645 523507 185661 523571
rect 185725 523507 185731 523571
rect 185415 523506 185731 523507
rect 174621 523027 174937 523028
rect 174621 522963 174627 523027
rect 174691 522963 174707 523027
rect 174771 522963 174787 523027
rect 174851 522963 174867 523027
rect 174931 522963 174937 523027
rect 174621 522962 174937 522963
rect 178439 523027 178755 523028
rect 178439 522963 178445 523027
rect 178509 522963 178525 523027
rect 178589 522963 178605 523027
rect 178669 522963 178685 523027
rect 178749 522963 178755 523027
rect 178439 522962 178755 522963
rect 182257 523027 182573 523028
rect 182257 522963 182263 523027
rect 182327 522963 182343 523027
rect 182407 522963 182423 523027
rect 182487 522963 182503 523027
rect 182567 522963 182573 523027
rect 182257 522962 182573 522963
rect 186075 523027 186391 523028
rect 186075 522963 186081 523027
rect 186145 522963 186161 523027
rect 186225 522963 186241 523027
rect 186305 522963 186321 523027
rect 186385 522963 186391 523027
rect 186075 522962 186391 522963
rect 173961 522483 174277 522484
rect 173961 522419 173967 522483
rect 174031 522419 174047 522483
rect 174111 522419 174127 522483
rect 174191 522419 174207 522483
rect 174271 522419 174277 522483
rect 173961 522418 174277 522419
rect 177779 522483 178095 522484
rect 177779 522419 177785 522483
rect 177849 522419 177865 522483
rect 177929 522419 177945 522483
rect 178009 522419 178025 522483
rect 178089 522419 178095 522483
rect 177779 522418 178095 522419
rect 181597 522483 181913 522484
rect 181597 522419 181603 522483
rect 181667 522419 181683 522483
rect 181747 522419 181763 522483
rect 181827 522419 181843 522483
rect 181907 522419 181913 522483
rect 181597 522418 181913 522419
rect 185415 522483 185731 522484
rect 185415 522419 185421 522483
rect 185485 522419 185501 522483
rect 185565 522419 185581 522483
rect 185645 522419 185661 522483
rect 185725 522419 185731 522483
rect 185415 522418 185731 522419
rect 174621 521939 174937 521940
rect 174621 521875 174627 521939
rect 174691 521875 174707 521939
rect 174771 521875 174787 521939
rect 174851 521875 174867 521939
rect 174931 521875 174937 521939
rect 174621 521874 174937 521875
rect 178439 521939 178755 521940
rect 178439 521875 178445 521939
rect 178509 521875 178525 521939
rect 178589 521875 178605 521939
rect 178669 521875 178685 521939
rect 178749 521875 178755 521939
rect 178439 521874 178755 521875
rect 182257 521939 182573 521940
rect 182257 521875 182263 521939
rect 182327 521875 182343 521939
rect 182407 521875 182423 521939
rect 182487 521875 182503 521939
rect 182567 521875 182573 521939
rect 182257 521874 182573 521875
rect 186075 521939 186391 521940
rect 186075 521875 186081 521939
rect 186145 521875 186161 521939
rect 186225 521875 186241 521939
rect 186305 521875 186321 521939
rect 186385 521875 186391 521939
rect 186075 521874 186391 521875
rect 173961 521395 174277 521396
rect 173961 521331 173967 521395
rect 174031 521331 174047 521395
rect 174111 521331 174127 521395
rect 174191 521331 174207 521395
rect 174271 521331 174277 521395
rect 173961 521330 174277 521331
rect 177779 521395 178095 521396
rect 177779 521331 177785 521395
rect 177849 521331 177865 521395
rect 177929 521331 177945 521395
rect 178009 521331 178025 521395
rect 178089 521331 178095 521395
rect 177779 521330 178095 521331
rect 181597 521395 181913 521396
rect 181597 521331 181603 521395
rect 181667 521331 181683 521395
rect 181747 521331 181763 521395
rect 181827 521331 181843 521395
rect 181907 521331 181913 521395
rect 181597 521330 181913 521331
rect 185415 521395 185731 521396
rect 185415 521331 185421 521395
rect 185485 521331 185501 521395
rect 185565 521331 185581 521395
rect 185645 521331 185661 521395
rect 185725 521331 185731 521395
rect 185415 521330 185731 521331
rect 174621 520851 174937 520852
rect 174621 520787 174627 520851
rect 174691 520787 174707 520851
rect 174771 520787 174787 520851
rect 174851 520787 174867 520851
rect 174931 520787 174937 520851
rect 174621 520786 174937 520787
rect 178439 520851 178755 520852
rect 178439 520787 178445 520851
rect 178509 520787 178525 520851
rect 178589 520787 178605 520851
rect 178669 520787 178685 520851
rect 178749 520787 178755 520851
rect 178439 520786 178755 520787
rect 182257 520851 182573 520852
rect 182257 520787 182263 520851
rect 182327 520787 182343 520851
rect 182407 520787 182423 520851
rect 182487 520787 182503 520851
rect 182567 520787 182573 520851
rect 182257 520786 182573 520787
rect 186075 520851 186391 520852
rect 186075 520787 186081 520851
rect 186145 520787 186161 520851
rect 186225 520787 186241 520851
rect 186305 520787 186321 520851
rect 186385 520787 186391 520851
rect 186075 520786 186391 520787
rect 173961 520307 174277 520308
rect 173961 520243 173967 520307
rect 174031 520243 174047 520307
rect 174111 520243 174127 520307
rect 174191 520243 174207 520307
rect 174271 520243 174277 520307
rect 173961 520242 174277 520243
rect 177779 520307 178095 520308
rect 177779 520243 177785 520307
rect 177849 520243 177865 520307
rect 177929 520243 177945 520307
rect 178009 520243 178025 520307
rect 178089 520243 178095 520307
rect 177779 520242 178095 520243
rect 181597 520307 181913 520308
rect 181597 520243 181603 520307
rect 181667 520243 181683 520307
rect 181747 520243 181763 520307
rect 181827 520243 181843 520307
rect 181907 520243 181913 520307
rect 181597 520242 181913 520243
rect 185415 520307 185731 520308
rect 185415 520243 185421 520307
rect 185485 520243 185501 520307
rect 185565 520243 185581 520307
rect 185645 520243 185661 520307
rect 185725 520243 185731 520307
rect 185415 520242 185731 520243
rect 174621 519763 174937 519764
rect 174621 519699 174627 519763
rect 174691 519699 174707 519763
rect 174771 519699 174787 519763
rect 174851 519699 174867 519763
rect 174931 519699 174937 519763
rect 174621 519698 174937 519699
rect 178439 519763 178755 519764
rect 178439 519699 178445 519763
rect 178509 519699 178525 519763
rect 178589 519699 178605 519763
rect 178669 519699 178685 519763
rect 178749 519699 178755 519763
rect 178439 519698 178755 519699
rect 182257 519763 182573 519764
rect 182257 519699 182263 519763
rect 182327 519699 182343 519763
rect 182407 519699 182423 519763
rect 182487 519699 182503 519763
rect 182567 519699 182573 519763
rect 182257 519698 182573 519699
rect 186075 519763 186391 519764
rect 186075 519699 186081 519763
rect 186145 519699 186161 519763
rect 186225 519699 186241 519763
rect 186305 519699 186321 519763
rect 186385 519699 186391 519763
rect 186075 519698 186391 519699
rect 173961 519219 174277 519220
rect 173961 519155 173967 519219
rect 174031 519155 174047 519219
rect 174111 519155 174127 519219
rect 174191 519155 174207 519219
rect 174271 519155 174277 519219
rect 173961 519154 174277 519155
rect 177779 519219 178095 519220
rect 177779 519155 177785 519219
rect 177849 519155 177865 519219
rect 177929 519155 177945 519219
rect 178009 519155 178025 519219
rect 178089 519155 178095 519219
rect 177779 519154 178095 519155
rect 181597 519219 181913 519220
rect 181597 519155 181603 519219
rect 181667 519155 181683 519219
rect 181747 519155 181763 519219
rect 181827 519155 181843 519219
rect 181907 519155 181913 519219
rect 181597 519154 181913 519155
rect 185415 519219 185731 519220
rect 185415 519155 185421 519219
rect 185485 519155 185501 519219
rect 185565 519155 185581 519219
rect 185645 519155 185661 519219
rect 185725 519155 185731 519219
rect 185415 519154 185731 519155
rect 174621 518675 174937 518676
rect 174621 518611 174627 518675
rect 174691 518611 174707 518675
rect 174771 518611 174787 518675
rect 174851 518611 174867 518675
rect 174931 518611 174937 518675
rect 174621 518610 174937 518611
rect 178439 518675 178755 518676
rect 178439 518611 178445 518675
rect 178509 518611 178525 518675
rect 178589 518611 178605 518675
rect 178669 518611 178685 518675
rect 178749 518611 178755 518675
rect 178439 518610 178755 518611
rect 182257 518675 182573 518676
rect 182257 518611 182263 518675
rect 182327 518611 182343 518675
rect 182407 518611 182423 518675
rect 182487 518611 182503 518675
rect 182567 518611 182573 518675
rect 182257 518610 182573 518611
rect 186075 518675 186391 518676
rect 186075 518611 186081 518675
rect 186145 518611 186161 518675
rect 186225 518611 186241 518675
rect 186305 518611 186321 518675
rect 186385 518611 186391 518675
rect 186075 518610 186391 518611
rect 173961 518131 174277 518132
rect 173961 518067 173967 518131
rect 174031 518067 174047 518131
rect 174111 518067 174127 518131
rect 174191 518067 174207 518131
rect 174271 518067 174277 518131
rect 173961 518066 174277 518067
rect 177779 518131 178095 518132
rect 177779 518067 177785 518131
rect 177849 518067 177865 518131
rect 177929 518067 177945 518131
rect 178009 518067 178025 518131
rect 178089 518067 178095 518131
rect 177779 518066 178095 518067
rect 181597 518131 181913 518132
rect 181597 518067 181603 518131
rect 181667 518067 181683 518131
rect 181747 518067 181763 518131
rect 181827 518067 181843 518131
rect 181907 518067 181913 518131
rect 181597 518066 181913 518067
rect 185415 518131 185731 518132
rect 185415 518067 185421 518131
rect 185485 518067 185501 518131
rect 185565 518067 185581 518131
rect 185645 518067 185661 518131
rect 185725 518067 185731 518131
rect 185415 518066 185731 518067
rect 174621 517587 174937 517588
rect 174621 517523 174627 517587
rect 174691 517523 174707 517587
rect 174771 517523 174787 517587
rect 174851 517523 174867 517587
rect 174931 517523 174937 517587
rect 174621 517522 174937 517523
rect 178439 517587 178755 517588
rect 178439 517523 178445 517587
rect 178509 517523 178525 517587
rect 178589 517523 178605 517587
rect 178669 517523 178685 517587
rect 178749 517523 178755 517587
rect 178439 517522 178755 517523
rect 182257 517587 182573 517588
rect 182257 517523 182263 517587
rect 182327 517523 182343 517587
rect 182407 517523 182423 517587
rect 182487 517523 182503 517587
rect 182567 517523 182573 517587
rect 182257 517522 182573 517523
rect 186075 517587 186391 517588
rect 186075 517523 186081 517587
rect 186145 517523 186161 517587
rect 186225 517523 186241 517587
rect 186305 517523 186321 517587
rect 186385 517523 186391 517587
rect 186075 517522 186391 517523
rect 173961 517043 174277 517044
rect 173961 516979 173967 517043
rect 174031 516979 174047 517043
rect 174111 516979 174127 517043
rect 174191 516979 174207 517043
rect 174271 516979 174277 517043
rect 173961 516978 174277 516979
rect 177779 517043 178095 517044
rect 177779 516979 177785 517043
rect 177849 516979 177865 517043
rect 177929 516979 177945 517043
rect 178009 516979 178025 517043
rect 178089 516979 178095 517043
rect 177779 516978 178095 516979
rect 181597 517043 181913 517044
rect 181597 516979 181603 517043
rect 181667 516979 181683 517043
rect 181747 516979 181763 517043
rect 181827 516979 181843 517043
rect 181907 516979 181913 517043
rect 181597 516978 181913 516979
rect 185415 517043 185731 517044
rect 185415 516979 185421 517043
rect 185485 516979 185501 517043
rect 185565 516979 185581 517043
rect 185645 516979 185661 517043
rect 185725 516979 185731 517043
rect 185415 516978 185731 516979
rect 174621 516499 174937 516500
rect 174621 516435 174627 516499
rect 174691 516435 174707 516499
rect 174771 516435 174787 516499
rect 174851 516435 174867 516499
rect 174931 516435 174937 516499
rect 174621 516434 174937 516435
rect 178439 516499 178755 516500
rect 178439 516435 178445 516499
rect 178509 516435 178525 516499
rect 178589 516435 178605 516499
rect 178669 516435 178685 516499
rect 178749 516435 178755 516499
rect 178439 516434 178755 516435
rect 182257 516499 182573 516500
rect 182257 516435 182263 516499
rect 182327 516435 182343 516499
rect 182407 516435 182423 516499
rect 182487 516435 182503 516499
rect 182567 516435 182573 516499
rect 182257 516434 182573 516435
rect 186075 516499 186391 516500
rect 186075 516435 186081 516499
rect 186145 516435 186161 516499
rect 186225 516435 186241 516499
rect 186305 516435 186321 516499
rect 186385 516435 186391 516499
rect 186075 516434 186391 516435
rect 173961 515955 174277 515956
rect 173961 515891 173967 515955
rect 174031 515891 174047 515955
rect 174111 515891 174127 515955
rect 174191 515891 174207 515955
rect 174271 515891 174277 515955
rect 173961 515890 174277 515891
rect 177779 515955 178095 515956
rect 177779 515891 177785 515955
rect 177849 515891 177865 515955
rect 177929 515891 177945 515955
rect 178009 515891 178025 515955
rect 178089 515891 178095 515955
rect 177779 515890 178095 515891
rect 181597 515955 181913 515956
rect 181597 515891 181603 515955
rect 181667 515891 181683 515955
rect 181747 515891 181763 515955
rect 181827 515891 181843 515955
rect 181907 515891 181913 515955
rect 181597 515890 181913 515891
rect 185415 515955 185731 515956
rect 185415 515891 185421 515955
rect 185485 515891 185501 515955
rect 185565 515891 185581 515955
rect 185645 515891 185661 515955
rect 185725 515891 185731 515955
rect 185415 515890 185731 515891
rect 174621 515411 174937 515412
rect 174621 515347 174627 515411
rect 174691 515347 174707 515411
rect 174771 515347 174787 515411
rect 174851 515347 174867 515411
rect 174931 515347 174937 515411
rect 174621 515346 174937 515347
rect 178439 515411 178755 515412
rect 178439 515347 178445 515411
rect 178509 515347 178525 515411
rect 178589 515347 178605 515411
rect 178669 515347 178685 515411
rect 178749 515347 178755 515411
rect 178439 515346 178755 515347
rect 182257 515411 182573 515412
rect 182257 515347 182263 515411
rect 182327 515347 182343 515411
rect 182407 515347 182423 515411
rect 182487 515347 182503 515411
rect 182567 515347 182573 515411
rect 182257 515346 182573 515347
rect 186075 515411 186391 515412
rect 186075 515347 186081 515411
rect 186145 515347 186161 515411
rect 186225 515347 186241 515411
rect 186305 515347 186321 515411
rect 186385 515347 186391 515411
rect 186075 515346 186391 515347
rect 1990 509000 4010 509005
rect 1000 508200 2000 509000
rect 600 507800 2000 508200
rect 1000 507000 2000 507800
rect 4000 507000 4010 509000
rect 1990 506995 4010 507000
rect 1990 466000 4010 466005
rect 1000 465000 2000 466000
rect 600 464600 2000 465000
rect 1000 464000 2000 464600
rect 4000 464000 4010 466000
rect 1990 463995 4010 464000
rect 1990 423000 4010 423005
rect 1000 421700 2000 423000
rect 600 421000 2000 421700
rect 4000 421000 4010 423000
rect 1990 420995 4010 421000
rect 1990 380000 4010 380005
rect 1000 378700 2000 380000
rect 600 378430 2000 378700
rect 614 378318 2014 378430
rect 600 378000 2000 378318
rect 4000 378000 4010 380000
rect 1990 377995 4010 378000
<< via3 >>
rect 162626 538925 162690 541869
rect 159400 538587 159480 538687
rect 161390 538577 161510 538697
rect 174627 530639 174691 530643
rect 174627 530583 174631 530639
rect 174631 530583 174687 530639
rect 174687 530583 174691 530639
rect 174627 530579 174691 530583
rect 174707 530639 174771 530643
rect 174707 530583 174711 530639
rect 174711 530583 174767 530639
rect 174767 530583 174771 530639
rect 174707 530579 174771 530583
rect 174787 530639 174851 530643
rect 174787 530583 174791 530639
rect 174791 530583 174847 530639
rect 174847 530583 174851 530639
rect 174787 530579 174851 530583
rect 174867 530639 174931 530643
rect 174867 530583 174871 530639
rect 174871 530583 174927 530639
rect 174927 530583 174931 530639
rect 174867 530579 174931 530583
rect 178445 530639 178509 530643
rect 178445 530583 178449 530639
rect 178449 530583 178505 530639
rect 178505 530583 178509 530639
rect 178445 530579 178509 530583
rect 178525 530639 178589 530643
rect 178525 530583 178529 530639
rect 178529 530583 178585 530639
rect 178585 530583 178589 530639
rect 178525 530579 178589 530583
rect 178605 530639 178669 530643
rect 178605 530583 178609 530639
rect 178609 530583 178665 530639
rect 178665 530583 178669 530639
rect 178605 530579 178669 530583
rect 178685 530639 178749 530643
rect 178685 530583 178689 530639
rect 178689 530583 178745 530639
rect 178745 530583 178749 530639
rect 178685 530579 178749 530583
rect 182263 530639 182327 530643
rect 182263 530583 182267 530639
rect 182267 530583 182323 530639
rect 182323 530583 182327 530639
rect 182263 530579 182327 530583
rect 182343 530639 182407 530643
rect 182343 530583 182347 530639
rect 182347 530583 182403 530639
rect 182403 530583 182407 530639
rect 182343 530579 182407 530583
rect 182423 530639 182487 530643
rect 182423 530583 182427 530639
rect 182427 530583 182483 530639
rect 182483 530583 182487 530639
rect 182423 530579 182487 530583
rect 182503 530639 182567 530643
rect 182503 530583 182507 530639
rect 182507 530583 182563 530639
rect 182563 530583 182567 530639
rect 182503 530579 182567 530583
rect 186081 530639 186145 530643
rect 186081 530583 186085 530639
rect 186085 530583 186141 530639
rect 186141 530583 186145 530639
rect 186081 530579 186145 530583
rect 186161 530639 186225 530643
rect 186161 530583 186165 530639
rect 186165 530583 186221 530639
rect 186221 530583 186225 530639
rect 186161 530579 186225 530583
rect 186241 530639 186305 530643
rect 186241 530583 186245 530639
rect 186245 530583 186301 530639
rect 186301 530583 186305 530639
rect 186241 530579 186305 530583
rect 186321 530639 186385 530643
rect 186321 530583 186325 530639
rect 186325 530583 186381 530639
rect 186381 530583 186385 530639
rect 186321 530579 186385 530583
rect 173967 530095 174031 530099
rect 173967 530039 173971 530095
rect 173971 530039 174027 530095
rect 174027 530039 174031 530095
rect 173967 530035 174031 530039
rect 174047 530095 174111 530099
rect 174047 530039 174051 530095
rect 174051 530039 174107 530095
rect 174107 530039 174111 530095
rect 174047 530035 174111 530039
rect 174127 530095 174191 530099
rect 174127 530039 174131 530095
rect 174131 530039 174187 530095
rect 174187 530039 174191 530095
rect 174127 530035 174191 530039
rect 174207 530095 174271 530099
rect 174207 530039 174211 530095
rect 174211 530039 174267 530095
rect 174267 530039 174271 530095
rect 174207 530035 174271 530039
rect 177785 530095 177849 530099
rect 177785 530039 177789 530095
rect 177789 530039 177845 530095
rect 177845 530039 177849 530095
rect 177785 530035 177849 530039
rect 177865 530095 177929 530099
rect 177865 530039 177869 530095
rect 177869 530039 177925 530095
rect 177925 530039 177929 530095
rect 177865 530035 177929 530039
rect 177945 530095 178009 530099
rect 177945 530039 177949 530095
rect 177949 530039 178005 530095
rect 178005 530039 178009 530095
rect 177945 530035 178009 530039
rect 178025 530095 178089 530099
rect 178025 530039 178029 530095
rect 178029 530039 178085 530095
rect 178085 530039 178089 530095
rect 178025 530035 178089 530039
rect 181603 530095 181667 530099
rect 181603 530039 181607 530095
rect 181607 530039 181663 530095
rect 181663 530039 181667 530095
rect 181603 530035 181667 530039
rect 181683 530095 181747 530099
rect 181683 530039 181687 530095
rect 181687 530039 181743 530095
rect 181743 530039 181747 530095
rect 181683 530035 181747 530039
rect 181763 530095 181827 530099
rect 181763 530039 181767 530095
rect 181767 530039 181823 530095
rect 181823 530039 181827 530095
rect 181763 530035 181827 530039
rect 181843 530095 181907 530099
rect 181843 530039 181847 530095
rect 181847 530039 181903 530095
rect 181903 530039 181907 530095
rect 181843 530035 181907 530039
rect 185421 530095 185485 530099
rect 185421 530039 185425 530095
rect 185425 530039 185481 530095
rect 185481 530039 185485 530095
rect 185421 530035 185485 530039
rect 185501 530095 185565 530099
rect 185501 530039 185505 530095
rect 185505 530039 185561 530095
rect 185561 530039 185565 530095
rect 185501 530035 185565 530039
rect 185581 530095 185645 530099
rect 185581 530039 185585 530095
rect 185585 530039 185641 530095
rect 185641 530039 185645 530095
rect 185581 530035 185645 530039
rect 185661 530095 185725 530099
rect 185661 530039 185665 530095
rect 185665 530039 185721 530095
rect 185721 530039 185725 530095
rect 185661 530035 185725 530039
rect 174627 529551 174691 529555
rect 174627 529495 174631 529551
rect 174631 529495 174687 529551
rect 174687 529495 174691 529551
rect 174627 529491 174691 529495
rect 174707 529551 174771 529555
rect 174707 529495 174711 529551
rect 174711 529495 174767 529551
rect 174767 529495 174771 529551
rect 174707 529491 174771 529495
rect 174787 529551 174851 529555
rect 174787 529495 174791 529551
rect 174791 529495 174847 529551
rect 174847 529495 174851 529551
rect 174787 529491 174851 529495
rect 174867 529551 174931 529555
rect 174867 529495 174871 529551
rect 174871 529495 174927 529551
rect 174927 529495 174931 529551
rect 174867 529491 174931 529495
rect 178445 529551 178509 529555
rect 178445 529495 178449 529551
rect 178449 529495 178505 529551
rect 178505 529495 178509 529551
rect 178445 529491 178509 529495
rect 178525 529551 178589 529555
rect 178525 529495 178529 529551
rect 178529 529495 178585 529551
rect 178585 529495 178589 529551
rect 178525 529491 178589 529495
rect 178605 529551 178669 529555
rect 178605 529495 178609 529551
rect 178609 529495 178665 529551
rect 178665 529495 178669 529551
rect 178605 529491 178669 529495
rect 178685 529551 178749 529555
rect 178685 529495 178689 529551
rect 178689 529495 178745 529551
rect 178745 529495 178749 529551
rect 178685 529491 178749 529495
rect 182263 529551 182327 529555
rect 182263 529495 182267 529551
rect 182267 529495 182323 529551
rect 182323 529495 182327 529551
rect 182263 529491 182327 529495
rect 182343 529551 182407 529555
rect 182343 529495 182347 529551
rect 182347 529495 182403 529551
rect 182403 529495 182407 529551
rect 182343 529491 182407 529495
rect 182423 529551 182487 529555
rect 182423 529495 182427 529551
rect 182427 529495 182483 529551
rect 182483 529495 182487 529551
rect 182423 529491 182487 529495
rect 182503 529551 182567 529555
rect 182503 529495 182507 529551
rect 182507 529495 182563 529551
rect 182563 529495 182567 529551
rect 182503 529491 182567 529495
rect 186081 529551 186145 529555
rect 186081 529495 186085 529551
rect 186085 529495 186141 529551
rect 186141 529495 186145 529551
rect 186081 529491 186145 529495
rect 186161 529551 186225 529555
rect 186161 529495 186165 529551
rect 186165 529495 186221 529551
rect 186221 529495 186225 529551
rect 186161 529491 186225 529495
rect 186241 529551 186305 529555
rect 186241 529495 186245 529551
rect 186245 529495 186301 529551
rect 186301 529495 186305 529551
rect 186241 529491 186305 529495
rect 186321 529551 186385 529555
rect 186321 529495 186325 529551
rect 186325 529495 186381 529551
rect 186381 529495 186385 529551
rect 186321 529491 186385 529495
rect 173967 529007 174031 529011
rect 173967 528951 173971 529007
rect 173971 528951 174027 529007
rect 174027 528951 174031 529007
rect 173967 528947 174031 528951
rect 174047 529007 174111 529011
rect 174047 528951 174051 529007
rect 174051 528951 174107 529007
rect 174107 528951 174111 529007
rect 174047 528947 174111 528951
rect 174127 529007 174191 529011
rect 174127 528951 174131 529007
rect 174131 528951 174187 529007
rect 174187 528951 174191 529007
rect 174127 528947 174191 528951
rect 174207 529007 174271 529011
rect 174207 528951 174211 529007
rect 174211 528951 174267 529007
rect 174267 528951 174271 529007
rect 174207 528947 174271 528951
rect 177785 529007 177849 529011
rect 177785 528951 177789 529007
rect 177789 528951 177845 529007
rect 177845 528951 177849 529007
rect 177785 528947 177849 528951
rect 177865 529007 177929 529011
rect 177865 528951 177869 529007
rect 177869 528951 177925 529007
rect 177925 528951 177929 529007
rect 177865 528947 177929 528951
rect 177945 529007 178009 529011
rect 177945 528951 177949 529007
rect 177949 528951 178005 529007
rect 178005 528951 178009 529007
rect 177945 528947 178009 528951
rect 178025 529007 178089 529011
rect 178025 528951 178029 529007
rect 178029 528951 178085 529007
rect 178085 528951 178089 529007
rect 178025 528947 178089 528951
rect 181603 529007 181667 529011
rect 181603 528951 181607 529007
rect 181607 528951 181663 529007
rect 181663 528951 181667 529007
rect 181603 528947 181667 528951
rect 181683 529007 181747 529011
rect 181683 528951 181687 529007
rect 181687 528951 181743 529007
rect 181743 528951 181747 529007
rect 181683 528947 181747 528951
rect 181763 529007 181827 529011
rect 181763 528951 181767 529007
rect 181767 528951 181823 529007
rect 181823 528951 181827 529007
rect 181763 528947 181827 528951
rect 181843 529007 181907 529011
rect 181843 528951 181847 529007
rect 181847 528951 181903 529007
rect 181903 528951 181907 529007
rect 181843 528947 181907 528951
rect 185421 529007 185485 529011
rect 185421 528951 185425 529007
rect 185425 528951 185481 529007
rect 185481 528951 185485 529007
rect 185421 528947 185485 528951
rect 185501 529007 185565 529011
rect 185501 528951 185505 529007
rect 185505 528951 185561 529007
rect 185561 528951 185565 529007
rect 185501 528947 185565 528951
rect 185581 529007 185645 529011
rect 185581 528951 185585 529007
rect 185585 528951 185641 529007
rect 185641 528951 185645 529007
rect 185581 528947 185645 528951
rect 185661 529007 185725 529011
rect 185661 528951 185665 529007
rect 185665 528951 185721 529007
rect 185721 528951 185725 529007
rect 185661 528947 185725 528951
rect 174627 528463 174691 528467
rect 174627 528407 174631 528463
rect 174631 528407 174687 528463
rect 174687 528407 174691 528463
rect 174627 528403 174691 528407
rect 174707 528463 174771 528467
rect 174707 528407 174711 528463
rect 174711 528407 174767 528463
rect 174767 528407 174771 528463
rect 174707 528403 174771 528407
rect 174787 528463 174851 528467
rect 174787 528407 174791 528463
rect 174791 528407 174847 528463
rect 174847 528407 174851 528463
rect 174787 528403 174851 528407
rect 174867 528463 174931 528467
rect 174867 528407 174871 528463
rect 174871 528407 174927 528463
rect 174927 528407 174931 528463
rect 174867 528403 174931 528407
rect 178445 528463 178509 528467
rect 178445 528407 178449 528463
rect 178449 528407 178505 528463
rect 178505 528407 178509 528463
rect 178445 528403 178509 528407
rect 178525 528463 178589 528467
rect 178525 528407 178529 528463
rect 178529 528407 178585 528463
rect 178585 528407 178589 528463
rect 178525 528403 178589 528407
rect 178605 528463 178669 528467
rect 178605 528407 178609 528463
rect 178609 528407 178665 528463
rect 178665 528407 178669 528463
rect 178605 528403 178669 528407
rect 178685 528463 178749 528467
rect 178685 528407 178689 528463
rect 178689 528407 178745 528463
rect 178745 528407 178749 528463
rect 178685 528403 178749 528407
rect 182263 528463 182327 528467
rect 182263 528407 182267 528463
rect 182267 528407 182323 528463
rect 182323 528407 182327 528463
rect 182263 528403 182327 528407
rect 182343 528463 182407 528467
rect 182343 528407 182347 528463
rect 182347 528407 182403 528463
rect 182403 528407 182407 528463
rect 182343 528403 182407 528407
rect 182423 528463 182487 528467
rect 182423 528407 182427 528463
rect 182427 528407 182483 528463
rect 182483 528407 182487 528463
rect 182423 528403 182487 528407
rect 182503 528463 182567 528467
rect 182503 528407 182507 528463
rect 182507 528407 182563 528463
rect 182563 528407 182567 528463
rect 182503 528403 182567 528407
rect 186081 528463 186145 528467
rect 186081 528407 186085 528463
rect 186085 528407 186141 528463
rect 186141 528407 186145 528463
rect 186081 528403 186145 528407
rect 186161 528463 186225 528467
rect 186161 528407 186165 528463
rect 186165 528407 186221 528463
rect 186221 528407 186225 528463
rect 186161 528403 186225 528407
rect 186241 528463 186305 528467
rect 186241 528407 186245 528463
rect 186245 528407 186301 528463
rect 186301 528407 186305 528463
rect 186241 528403 186305 528407
rect 186321 528463 186385 528467
rect 186321 528407 186325 528463
rect 186325 528407 186381 528463
rect 186381 528407 186385 528463
rect 186321 528403 186385 528407
rect 173967 527919 174031 527923
rect 173967 527863 173971 527919
rect 173971 527863 174027 527919
rect 174027 527863 174031 527919
rect 173967 527859 174031 527863
rect 174047 527919 174111 527923
rect 174047 527863 174051 527919
rect 174051 527863 174107 527919
rect 174107 527863 174111 527919
rect 174047 527859 174111 527863
rect 174127 527919 174191 527923
rect 174127 527863 174131 527919
rect 174131 527863 174187 527919
rect 174187 527863 174191 527919
rect 174127 527859 174191 527863
rect 174207 527919 174271 527923
rect 174207 527863 174211 527919
rect 174211 527863 174267 527919
rect 174267 527863 174271 527919
rect 174207 527859 174271 527863
rect 177785 527919 177849 527923
rect 177785 527863 177789 527919
rect 177789 527863 177845 527919
rect 177845 527863 177849 527919
rect 177785 527859 177849 527863
rect 177865 527919 177929 527923
rect 177865 527863 177869 527919
rect 177869 527863 177925 527919
rect 177925 527863 177929 527919
rect 177865 527859 177929 527863
rect 177945 527919 178009 527923
rect 177945 527863 177949 527919
rect 177949 527863 178005 527919
rect 178005 527863 178009 527919
rect 177945 527859 178009 527863
rect 178025 527919 178089 527923
rect 178025 527863 178029 527919
rect 178029 527863 178085 527919
rect 178085 527863 178089 527919
rect 178025 527859 178089 527863
rect 181603 527919 181667 527923
rect 181603 527863 181607 527919
rect 181607 527863 181663 527919
rect 181663 527863 181667 527919
rect 181603 527859 181667 527863
rect 181683 527919 181747 527923
rect 181683 527863 181687 527919
rect 181687 527863 181743 527919
rect 181743 527863 181747 527919
rect 181683 527859 181747 527863
rect 181763 527919 181827 527923
rect 181763 527863 181767 527919
rect 181767 527863 181823 527919
rect 181823 527863 181827 527919
rect 181763 527859 181827 527863
rect 181843 527919 181907 527923
rect 181843 527863 181847 527919
rect 181847 527863 181903 527919
rect 181903 527863 181907 527919
rect 181843 527859 181907 527863
rect 185421 527919 185485 527923
rect 185421 527863 185425 527919
rect 185425 527863 185481 527919
rect 185481 527863 185485 527919
rect 185421 527859 185485 527863
rect 185501 527919 185565 527923
rect 185501 527863 185505 527919
rect 185505 527863 185561 527919
rect 185561 527863 185565 527919
rect 185501 527859 185565 527863
rect 185581 527919 185645 527923
rect 185581 527863 185585 527919
rect 185585 527863 185641 527919
rect 185641 527863 185645 527919
rect 185581 527859 185645 527863
rect 185661 527919 185725 527923
rect 185661 527863 185665 527919
rect 185665 527863 185721 527919
rect 185721 527863 185725 527919
rect 185661 527859 185725 527863
rect 174627 527375 174691 527379
rect 174627 527319 174631 527375
rect 174631 527319 174687 527375
rect 174687 527319 174691 527375
rect 174627 527315 174691 527319
rect 174707 527375 174771 527379
rect 174707 527319 174711 527375
rect 174711 527319 174767 527375
rect 174767 527319 174771 527375
rect 174707 527315 174771 527319
rect 174787 527375 174851 527379
rect 174787 527319 174791 527375
rect 174791 527319 174847 527375
rect 174847 527319 174851 527375
rect 174787 527315 174851 527319
rect 174867 527375 174931 527379
rect 174867 527319 174871 527375
rect 174871 527319 174927 527375
rect 174927 527319 174931 527375
rect 174867 527315 174931 527319
rect 178445 527375 178509 527379
rect 178445 527319 178449 527375
rect 178449 527319 178505 527375
rect 178505 527319 178509 527375
rect 178445 527315 178509 527319
rect 178525 527375 178589 527379
rect 178525 527319 178529 527375
rect 178529 527319 178585 527375
rect 178585 527319 178589 527375
rect 178525 527315 178589 527319
rect 178605 527375 178669 527379
rect 178605 527319 178609 527375
rect 178609 527319 178665 527375
rect 178665 527319 178669 527375
rect 178605 527315 178669 527319
rect 178685 527375 178749 527379
rect 178685 527319 178689 527375
rect 178689 527319 178745 527375
rect 178745 527319 178749 527375
rect 178685 527315 178749 527319
rect 182263 527375 182327 527379
rect 182263 527319 182267 527375
rect 182267 527319 182323 527375
rect 182323 527319 182327 527375
rect 182263 527315 182327 527319
rect 182343 527375 182407 527379
rect 182343 527319 182347 527375
rect 182347 527319 182403 527375
rect 182403 527319 182407 527375
rect 182343 527315 182407 527319
rect 182423 527375 182487 527379
rect 182423 527319 182427 527375
rect 182427 527319 182483 527375
rect 182483 527319 182487 527375
rect 182423 527315 182487 527319
rect 182503 527375 182567 527379
rect 182503 527319 182507 527375
rect 182507 527319 182563 527375
rect 182563 527319 182567 527375
rect 182503 527315 182567 527319
rect 186081 527375 186145 527379
rect 186081 527319 186085 527375
rect 186085 527319 186141 527375
rect 186141 527319 186145 527375
rect 186081 527315 186145 527319
rect 186161 527375 186225 527379
rect 186161 527319 186165 527375
rect 186165 527319 186221 527375
rect 186221 527319 186225 527375
rect 186161 527315 186225 527319
rect 186241 527375 186305 527379
rect 186241 527319 186245 527375
rect 186245 527319 186301 527375
rect 186301 527319 186305 527375
rect 186241 527315 186305 527319
rect 186321 527375 186385 527379
rect 186321 527319 186325 527375
rect 186325 527319 186381 527375
rect 186381 527319 186385 527375
rect 186321 527315 186385 527319
rect 173967 526831 174031 526835
rect 173967 526775 173971 526831
rect 173971 526775 174027 526831
rect 174027 526775 174031 526831
rect 173967 526771 174031 526775
rect 174047 526831 174111 526835
rect 174047 526775 174051 526831
rect 174051 526775 174107 526831
rect 174107 526775 174111 526831
rect 174047 526771 174111 526775
rect 174127 526831 174191 526835
rect 174127 526775 174131 526831
rect 174131 526775 174187 526831
rect 174187 526775 174191 526831
rect 174127 526771 174191 526775
rect 174207 526831 174271 526835
rect 174207 526775 174211 526831
rect 174211 526775 174267 526831
rect 174267 526775 174271 526831
rect 174207 526771 174271 526775
rect 177785 526831 177849 526835
rect 177785 526775 177789 526831
rect 177789 526775 177845 526831
rect 177845 526775 177849 526831
rect 177785 526771 177849 526775
rect 177865 526831 177929 526835
rect 177865 526775 177869 526831
rect 177869 526775 177925 526831
rect 177925 526775 177929 526831
rect 177865 526771 177929 526775
rect 177945 526831 178009 526835
rect 177945 526775 177949 526831
rect 177949 526775 178005 526831
rect 178005 526775 178009 526831
rect 177945 526771 178009 526775
rect 178025 526831 178089 526835
rect 178025 526775 178029 526831
rect 178029 526775 178085 526831
rect 178085 526775 178089 526831
rect 178025 526771 178089 526775
rect 181603 526831 181667 526835
rect 181603 526775 181607 526831
rect 181607 526775 181663 526831
rect 181663 526775 181667 526831
rect 181603 526771 181667 526775
rect 181683 526831 181747 526835
rect 181683 526775 181687 526831
rect 181687 526775 181743 526831
rect 181743 526775 181747 526831
rect 181683 526771 181747 526775
rect 181763 526831 181827 526835
rect 181763 526775 181767 526831
rect 181767 526775 181823 526831
rect 181823 526775 181827 526831
rect 181763 526771 181827 526775
rect 181843 526831 181907 526835
rect 181843 526775 181847 526831
rect 181847 526775 181903 526831
rect 181903 526775 181907 526831
rect 181843 526771 181907 526775
rect 185421 526831 185485 526835
rect 185421 526775 185425 526831
rect 185425 526775 185481 526831
rect 185481 526775 185485 526831
rect 185421 526771 185485 526775
rect 185501 526831 185565 526835
rect 185501 526775 185505 526831
rect 185505 526775 185561 526831
rect 185561 526775 185565 526831
rect 185501 526771 185565 526775
rect 185581 526831 185645 526835
rect 185581 526775 185585 526831
rect 185585 526775 185641 526831
rect 185641 526775 185645 526831
rect 185581 526771 185645 526775
rect 185661 526831 185725 526835
rect 185661 526775 185665 526831
rect 185665 526775 185721 526831
rect 185721 526775 185725 526831
rect 185661 526771 185725 526775
rect 174627 526287 174691 526291
rect 174627 526231 174631 526287
rect 174631 526231 174687 526287
rect 174687 526231 174691 526287
rect 174627 526227 174691 526231
rect 174707 526287 174771 526291
rect 174707 526231 174711 526287
rect 174711 526231 174767 526287
rect 174767 526231 174771 526287
rect 174707 526227 174771 526231
rect 174787 526287 174851 526291
rect 174787 526231 174791 526287
rect 174791 526231 174847 526287
rect 174847 526231 174851 526287
rect 174787 526227 174851 526231
rect 174867 526287 174931 526291
rect 174867 526231 174871 526287
rect 174871 526231 174927 526287
rect 174927 526231 174931 526287
rect 174867 526227 174931 526231
rect 178445 526287 178509 526291
rect 178445 526231 178449 526287
rect 178449 526231 178505 526287
rect 178505 526231 178509 526287
rect 178445 526227 178509 526231
rect 178525 526287 178589 526291
rect 178525 526231 178529 526287
rect 178529 526231 178585 526287
rect 178585 526231 178589 526287
rect 178525 526227 178589 526231
rect 178605 526287 178669 526291
rect 178605 526231 178609 526287
rect 178609 526231 178665 526287
rect 178665 526231 178669 526287
rect 178605 526227 178669 526231
rect 178685 526287 178749 526291
rect 178685 526231 178689 526287
rect 178689 526231 178745 526287
rect 178745 526231 178749 526287
rect 178685 526227 178749 526231
rect 182263 526287 182327 526291
rect 182263 526231 182267 526287
rect 182267 526231 182323 526287
rect 182323 526231 182327 526287
rect 182263 526227 182327 526231
rect 182343 526287 182407 526291
rect 182343 526231 182347 526287
rect 182347 526231 182403 526287
rect 182403 526231 182407 526287
rect 182343 526227 182407 526231
rect 182423 526287 182487 526291
rect 182423 526231 182427 526287
rect 182427 526231 182483 526287
rect 182483 526231 182487 526287
rect 182423 526227 182487 526231
rect 182503 526287 182567 526291
rect 182503 526231 182507 526287
rect 182507 526231 182563 526287
rect 182563 526231 182567 526287
rect 182503 526227 182567 526231
rect 186081 526287 186145 526291
rect 186081 526231 186085 526287
rect 186085 526231 186141 526287
rect 186141 526231 186145 526287
rect 186081 526227 186145 526231
rect 186161 526287 186225 526291
rect 186161 526231 186165 526287
rect 186165 526231 186221 526287
rect 186221 526231 186225 526287
rect 186161 526227 186225 526231
rect 186241 526287 186305 526291
rect 186241 526231 186245 526287
rect 186245 526231 186301 526287
rect 186301 526231 186305 526287
rect 186241 526227 186305 526231
rect 186321 526287 186385 526291
rect 186321 526231 186325 526287
rect 186325 526231 186381 526287
rect 186381 526231 186385 526287
rect 186321 526227 186385 526231
rect 173967 525743 174031 525747
rect 173967 525687 173971 525743
rect 173971 525687 174027 525743
rect 174027 525687 174031 525743
rect 173967 525683 174031 525687
rect 174047 525743 174111 525747
rect 174047 525687 174051 525743
rect 174051 525687 174107 525743
rect 174107 525687 174111 525743
rect 174047 525683 174111 525687
rect 174127 525743 174191 525747
rect 174127 525687 174131 525743
rect 174131 525687 174187 525743
rect 174187 525687 174191 525743
rect 174127 525683 174191 525687
rect 174207 525743 174271 525747
rect 174207 525687 174211 525743
rect 174211 525687 174267 525743
rect 174267 525687 174271 525743
rect 174207 525683 174271 525687
rect 177785 525743 177849 525747
rect 177785 525687 177789 525743
rect 177789 525687 177845 525743
rect 177845 525687 177849 525743
rect 177785 525683 177849 525687
rect 177865 525743 177929 525747
rect 177865 525687 177869 525743
rect 177869 525687 177925 525743
rect 177925 525687 177929 525743
rect 177865 525683 177929 525687
rect 177945 525743 178009 525747
rect 177945 525687 177949 525743
rect 177949 525687 178005 525743
rect 178005 525687 178009 525743
rect 177945 525683 178009 525687
rect 178025 525743 178089 525747
rect 178025 525687 178029 525743
rect 178029 525687 178085 525743
rect 178085 525687 178089 525743
rect 178025 525683 178089 525687
rect 181603 525743 181667 525747
rect 181603 525687 181607 525743
rect 181607 525687 181663 525743
rect 181663 525687 181667 525743
rect 181603 525683 181667 525687
rect 181683 525743 181747 525747
rect 181683 525687 181687 525743
rect 181687 525687 181743 525743
rect 181743 525687 181747 525743
rect 181683 525683 181747 525687
rect 181763 525743 181827 525747
rect 181763 525687 181767 525743
rect 181767 525687 181823 525743
rect 181823 525687 181827 525743
rect 181763 525683 181827 525687
rect 181843 525743 181907 525747
rect 181843 525687 181847 525743
rect 181847 525687 181903 525743
rect 181903 525687 181907 525743
rect 181843 525683 181907 525687
rect 185421 525743 185485 525747
rect 185421 525687 185425 525743
rect 185425 525687 185481 525743
rect 185481 525687 185485 525743
rect 185421 525683 185485 525687
rect 185501 525743 185565 525747
rect 185501 525687 185505 525743
rect 185505 525687 185561 525743
rect 185561 525687 185565 525743
rect 185501 525683 185565 525687
rect 185581 525743 185645 525747
rect 185581 525687 185585 525743
rect 185585 525687 185641 525743
rect 185641 525687 185645 525743
rect 185581 525683 185645 525687
rect 185661 525743 185725 525747
rect 185661 525687 185665 525743
rect 185665 525687 185721 525743
rect 185721 525687 185725 525743
rect 185661 525683 185725 525687
rect 174627 525199 174691 525203
rect 174627 525143 174631 525199
rect 174631 525143 174687 525199
rect 174687 525143 174691 525199
rect 174627 525139 174691 525143
rect 174707 525199 174771 525203
rect 174707 525143 174711 525199
rect 174711 525143 174767 525199
rect 174767 525143 174771 525199
rect 174707 525139 174771 525143
rect 174787 525199 174851 525203
rect 174787 525143 174791 525199
rect 174791 525143 174847 525199
rect 174847 525143 174851 525199
rect 174787 525139 174851 525143
rect 174867 525199 174931 525203
rect 174867 525143 174871 525199
rect 174871 525143 174927 525199
rect 174927 525143 174931 525199
rect 174867 525139 174931 525143
rect 178445 525199 178509 525203
rect 178445 525143 178449 525199
rect 178449 525143 178505 525199
rect 178505 525143 178509 525199
rect 178445 525139 178509 525143
rect 178525 525199 178589 525203
rect 178525 525143 178529 525199
rect 178529 525143 178585 525199
rect 178585 525143 178589 525199
rect 178525 525139 178589 525143
rect 178605 525199 178669 525203
rect 178605 525143 178609 525199
rect 178609 525143 178665 525199
rect 178665 525143 178669 525199
rect 178605 525139 178669 525143
rect 178685 525199 178749 525203
rect 178685 525143 178689 525199
rect 178689 525143 178745 525199
rect 178745 525143 178749 525199
rect 178685 525139 178749 525143
rect 182263 525199 182327 525203
rect 182263 525143 182267 525199
rect 182267 525143 182323 525199
rect 182323 525143 182327 525199
rect 182263 525139 182327 525143
rect 182343 525199 182407 525203
rect 182343 525143 182347 525199
rect 182347 525143 182403 525199
rect 182403 525143 182407 525199
rect 182343 525139 182407 525143
rect 182423 525199 182487 525203
rect 182423 525143 182427 525199
rect 182427 525143 182483 525199
rect 182483 525143 182487 525199
rect 182423 525139 182487 525143
rect 182503 525199 182567 525203
rect 182503 525143 182507 525199
rect 182507 525143 182563 525199
rect 182563 525143 182567 525199
rect 182503 525139 182567 525143
rect 186081 525199 186145 525203
rect 186081 525143 186085 525199
rect 186085 525143 186141 525199
rect 186141 525143 186145 525199
rect 186081 525139 186145 525143
rect 186161 525199 186225 525203
rect 186161 525143 186165 525199
rect 186165 525143 186221 525199
rect 186221 525143 186225 525199
rect 186161 525139 186225 525143
rect 186241 525199 186305 525203
rect 186241 525143 186245 525199
rect 186245 525143 186301 525199
rect 186301 525143 186305 525199
rect 186241 525139 186305 525143
rect 186321 525199 186385 525203
rect 186321 525143 186325 525199
rect 186325 525143 186381 525199
rect 186381 525143 186385 525199
rect 186321 525139 186385 525143
rect 173967 524655 174031 524659
rect 173967 524599 173971 524655
rect 173971 524599 174027 524655
rect 174027 524599 174031 524655
rect 173967 524595 174031 524599
rect 174047 524655 174111 524659
rect 174047 524599 174051 524655
rect 174051 524599 174107 524655
rect 174107 524599 174111 524655
rect 174047 524595 174111 524599
rect 174127 524655 174191 524659
rect 174127 524599 174131 524655
rect 174131 524599 174187 524655
rect 174187 524599 174191 524655
rect 174127 524595 174191 524599
rect 174207 524655 174271 524659
rect 174207 524599 174211 524655
rect 174211 524599 174267 524655
rect 174267 524599 174271 524655
rect 174207 524595 174271 524599
rect 177785 524655 177849 524659
rect 177785 524599 177789 524655
rect 177789 524599 177845 524655
rect 177845 524599 177849 524655
rect 177785 524595 177849 524599
rect 177865 524655 177929 524659
rect 177865 524599 177869 524655
rect 177869 524599 177925 524655
rect 177925 524599 177929 524655
rect 177865 524595 177929 524599
rect 177945 524655 178009 524659
rect 177945 524599 177949 524655
rect 177949 524599 178005 524655
rect 178005 524599 178009 524655
rect 177945 524595 178009 524599
rect 178025 524655 178089 524659
rect 178025 524599 178029 524655
rect 178029 524599 178085 524655
rect 178085 524599 178089 524655
rect 178025 524595 178089 524599
rect 181603 524655 181667 524659
rect 181603 524599 181607 524655
rect 181607 524599 181663 524655
rect 181663 524599 181667 524655
rect 181603 524595 181667 524599
rect 181683 524655 181747 524659
rect 181683 524599 181687 524655
rect 181687 524599 181743 524655
rect 181743 524599 181747 524655
rect 181683 524595 181747 524599
rect 181763 524655 181827 524659
rect 181763 524599 181767 524655
rect 181767 524599 181823 524655
rect 181823 524599 181827 524655
rect 181763 524595 181827 524599
rect 181843 524655 181907 524659
rect 181843 524599 181847 524655
rect 181847 524599 181903 524655
rect 181903 524599 181907 524655
rect 181843 524595 181907 524599
rect 185421 524655 185485 524659
rect 185421 524599 185425 524655
rect 185425 524599 185481 524655
rect 185481 524599 185485 524655
rect 185421 524595 185485 524599
rect 185501 524655 185565 524659
rect 185501 524599 185505 524655
rect 185505 524599 185561 524655
rect 185561 524599 185565 524655
rect 185501 524595 185565 524599
rect 185581 524655 185645 524659
rect 185581 524599 185585 524655
rect 185585 524599 185641 524655
rect 185641 524599 185645 524655
rect 185581 524595 185645 524599
rect 185661 524655 185725 524659
rect 185661 524599 185665 524655
rect 185665 524599 185721 524655
rect 185721 524599 185725 524655
rect 185661 524595 185725 524599
rect 174627 524111 174691 524115
rect 174627 524055 174631 524111
rect 174631 524055 174687 524111
rect 174687 524055 174691 524111
rect 174627 524051 174691 524055
rect 174707 524111 174771 524115
rect 174707 524055 174711 524111
rect 174711 524055 174767 524111
rect 174767 524055 174771 524111
rect 174707 524051 174771 524055
rect 174787 524111 174851 524115
rect 174787 524055 174791 524111
rect 174791 524055 174847 524111
rect 174847 524055 174851 524111
rect 174787 524051 174851 524055
rect 174867 524111 174931 524115
rect 174867 524055 174871 524111
rect 174871 524055 174927 524111
rect 174927 524055 174931 524111
rect 174867 524051 174931 524055
rect 178445 524111 178509 524115
rect 178445 524055 178449 524111
rect 178449 524055 178505 524111
rect 178505 524055 178509 524111
rect 178445 524051 178509 524055
rect 178525 524111 178589 524115
rect 178525 524055 178529 524111
rect 178529 524055 178585 524111
rect 178585 524055 178589 524111
rect 178525 524051 178589 524055
rect 178605 524111 178669 524115
rect 178605 524055 178609 524111
rect 178609 524055 178665 524111
rect 178665 524055 178669 524111
rect 178605 524051 178669 524055
rect 178685 524111 178749 524115
rect 178685 524055 178689 524111
rect 178689 524055 178745 524111
rect 178745 524055 178749 524111
rect 178685 524051 178749 524055
rect 182263 524111 182327 524115
rect 182263 524055 182267 524111
rect 182267 524055 182323 524111
rect 182323 524055 182327 524111
rect 182263 524051 182327 524055
rect 182343 524111 182407 524115
rect 182343 524055 182347 524111
rect 182347 524055 182403 524111
rect 182403 524055 182407 524111
rect 182343 524051 182407 524055
rect 182423 524111 182487 524115
rect 182423 524055 182427 524111
rect 182427 524055 182483 524111
rect 182483 524055 182487 524111
rect 182423 524051 182487 524055
rect 182503 524111 182567 524115
rect 182503 524055 182507 524111
rect 182507 524055 182563 524111
rect 182563 524055 182567 524111
rect 182503 524051 182567 524055
rect 186081 524111 186145 524115
rect 186081 524055 186085 524111
rect 186085 524055 186141 524111
rect 186141 524055 186145 524111
rect 186081 524051 186145 524055
rect 186161 524111 186225 524115
rect 186161 524055 186165 524111
rect 186165 524055 186221 524111
rect 186221 524055 186225 524111
rect 186161 524051 186225 524055
rect 186241 524111 186305 524115
rect 186241 524055 186245 524111
rect 186245 524055 186301 524111
rect 186301 524055 186305 524111
rect 186241 524051 186305 524055
rect 186321 524111 186385 524115
rect 186321 524055 186325 524111
rect 186325 524055 186381 524111
rect 186381 524055 186385 524111
rect 186321 524051 186385 524055
rect 173967 523567 174031 523571
rect 173967 523511 173971 523567
rect 173971 523511 174027 523567
rect 174027 523511 174031 523567
rect 173967 523507 174031 523511
rect 174047 523567 174111 523571
rect 174047 523511 174051 523567
rect 174051 523511 174107 523567
rect 174107 523511 174111 523567
rect 174047 523507 174111 523511
rect 174127 523567 174191 523571
rect 174127 523511 174131 523567
rect 174131 523511 174187 523567
rect 174187 523511 174191 523567
rect 174127 523507 174191 523511
rect 174207 523567 174271 523571
rect 174207 523511 174211 523567
rect 174211 523511 174267 523567
rect 174267 523511 174271 523567
rect 174207 523507 174271 523511
rect 177785 523567 177849 523571
rect 177785 523511 177789 523567
rect 177789 523511 177845 523567
rect 177845 523511 177849 523567
rect 177785 523507 177849 523511
rect 177865 523567 177929 523571
rect 177865 523511 177869 523567
rect 177869 523511 177925 523567
rect 177925 523511 177929 523567
rect 177865 523507 177929 523511
rect 177945 523567 178009 523571
rect 177945 523511 177949 523567
rect 177949 523511 178005 523567
rect 178005 523511 178009 523567
rect 177945 523507 178009 523511
rect 178025 523567 178089 523571
rect 178025 523511 178029 523567
rect 178029 523511 178085 523567
rect 178085 523511 178089 523567
rect 178025 523507 178089 523511
rect 181603 523567 181667 523571
rect 181603 523511 181607 523567
rect 181607 523511 181663 523567
rect 181663 523511 181667 523567
rect 181603 523507 181667 523511
rect 181683 523567 181747 523571
rect 181683 523511 181687 523567
rect 181687 523511 181743 523567
rect 181743 523511 181747 523567
rect 181683 523507 181747 523511
rect 181763 523567 181827 523571
rect 181763 523511 181767 523567
rect 181767 523511 181823 523567
rect 181823 523511 181827 523567
rect 181763 523507 181827 523511
rect 181843 523567 181907 523571
rect 181843 523511 181847 523567
rect 181847 523511 181903 523567
rect 181903 523511 181907 523567
rect 181843 523507 181907 523511
rect 185421 523567 185485 523571
rect 185421 523511 185425 523567
rect 185425 523511 185481 523567
rect 185481 523511 185485 523567
rect 185421 523507 185485 523511
rect 185501 523567 185565 523571
rect 185501 523511 185505 523567
rect 185505 523511 185561 523567
rect 185561 523511 185565 523567
rect 185501 523507 185565 523511
rect 185581 523567 185645 523571
rect 185581 523511 185585 523567
rect 185585 523511 185641 523567
rect 185641 523511 185645 523567
rect 185581 523507 185645 523511
rect 185661 523567 185725 523571
rect 185661 523511 185665 523567
rect 185665 523511 185721 523567
rect 185721 523511 185725 523567
rect 185661 523507 185725 523511
rect 174627 523023 174691 523027
rect 174627 522967 174631 523023
rect 174631 522967 174687 523023
rect 174687 522967 174691 523023
rect 174627 522963 174691 522967
rect 174707 523023 174771 523027
rect 174707 522967 174711 523023
rect 174711 522967 174767 523023
rect 174767 522967 174771 523023
rect 174707 522963 174771 522967
rect 174787 523023 174851 523027
rect 174787 522967 174791 523023
rect 174791 522967 174847 523023
rect 174847 522967 174851 523023
rect 174787 522963 174851 522967
rect 174867 523023 174931 523027
rect 174867 522967 174871 523023
rect 174871 522967 174927 523023
rect 174927 522967 174931 523023
rect 174867 522963 174931 522967
rect 178445 523023 178509 523027
rect 178445 522967 178449 523023
rect 178449 522967 178505 523023
rect 178505 522967 178509 523023
rect 178445 522963 178509 522967
rect 178525 523023 178589 523027
rect 178525 522967 178529 523023
rect 178529 522967 178585 523023
rect 178585 522967 178589 523023
rect 178525 522963 178589 522967
rect 178605 523023 178669 523027
rect 178605 522967 178609 523023
rect 178609 522967 178665 523023
rect 178665 522967 178669 523023
rect 178605 522963 178669 522967
rect 178685 523023 178749 523027
rect 178685 522967 178689 523023
rect 178689 522967 178745 523023
rect 178745 522967 178749 523023
rect 178685 522963 178749 522967
rect 182263 523023 182327 523027
rect 182263 522967 182267 523023
rect 182267 522967 182323 523023
rect 182323 522967 182327 523023
rect 182263 522963 182327 522967
rect 182343 523023 182407 523027
rect 182343 522967 182347 523023
rect 182347 522967 182403 523023
rect 182403 522967 182407 523023
rect 182343 522963 182407 522967
rect 182423 523023 182487 523027
rect 182423 522967 182427 523023
rect 182427 522967 182483 523023
rect 182483 522967 182487 523023
rect 182423 522963 182487 522967
rect 182503 523023 182567 523027
rect 182503 522967 182507 523023
rect 182507 522967 182563 523023
rect 182563 522967 182567 523023
rect 182503 522963 182567 522967
rect 186081 523023 186145 523027
rect 186081 522967 186085 523023
rect 186085 522967 186141 523023
rect 186141 522967 186145 523023
rect 186081 522963 186145 522967
rect 186161 523023 186225 523027
rect 186161 522967 186165 523023
rect 186165 522967 186221 523023
rect 186221 522967 186225 523023
rect 186161 522963 186225 522967
rect 186241 523023 186305 523027
rect 186241 522967 186245 523023
rect 186245 522967 186301 523023
rect 186301 522967 186305 523023
rect 186241 522963 186305 522967
rect 186321 523023 186385 523027
rect 186321 522967 186325 523023
rect 186325 522967 186381 523023
rect 186381 522967 186385 523023
rect 186321 522963 186385 522967
rect 173967 522479 174031 522483
rect 173967 522423 173971 522479
rect 173971 522423 174027 522479
rect 174027 522423 174031 522479
rect 173967 522419 174031 522423
rect 174047 522479 174111 522483
rect 174047 522423 174051 522479
rect 174051 522423 174107 522479
rect 174107 522423 174111 522479
rect 174047 522419 174111 522423
rect 174127 522479 174191 522483
rect 174127 522423 174131 522479
rect 174131 522423 174187 522479
rect 174187 522423 174191 522479
rect 174127 522419 174191 522423
rect 174207 522479 174271 522483
rect 174207 522423 174211 522479
rect 174211 522423 174267 522479
rect 174267 522423 174271 522479
rect 174207 522419 174271 522423
rect 177785 522479 177849 522483
rect 177785 522423 177789 522479
rect 177789 522423 177845 522479
rect 177845 522423 177849 522479
rect 177785 522419 177849 522423
rect 177865 522479 177929 522483
rect 177865 522423 177869 522479
rect 177869 522423 177925 522479
rect 177925 522423 177929 522479
rect 177865 522419 177929 522423
rect 177945 522479 178009 522483
rect 177945 522423 177949 522479
rect 177949 522423 178005 522479
rect 178005 522423 178009 522479
rect 177945 522419 178009 522423
rect 178025 522479 178089 522483
rect 178025 522423 178029 522479
rect 178029 522423 178085 522479
rect 178085 522423 178089 522479
rect 178025 522419 178089 522423
rect 181603 522479 181667 522483
rect 181603 522423 181607 522479
rect 181607 522423 181663 522479
rect 181663 522423 181667 522479
rect 181603 522419 181667 522423
rect 181683 522479 181747 522483
rect 181683 522423 181687 522479
rect 181687 522423 181743 522479
rect 181743 522423 181747 522479
rect 181683 522419 181747 522423
rect 181763 522479 181827 522483
rect 181763 522423 181767 522479
rect 181767 522423 181823 522479
rect 181823 522423 181827 522479
rect 181763 522419 181827 522423
rect 181843 522479 181907 522483
rect 181843 522423 181847 522479
rect 181847 522423 181903 522479
rect 181903 522423 181907 522479
rect 181843 522419 181907 522423
rect 185421 522479 185485 522483
rect 185421 522423 185425 522479
rect 185425 522423 185481 522479
rect 185481 522423 185485 522479
rect 185421 522419 185485 522423
rect 185501 522479 185565 522483
rect 185501 522423 185505 522479
rect 185505 522423 185561 522479
rect 185561 522423 185565 522479
rect 185501 522419 185565 522423
rect 185581 522479 185645 522483
rect 185581 522423 185585 522479
rect 185585 522423 185641 522479
rect 185641 522423 185645 522479
rect 185581 522419 185645 522423
rect 185661 522479 185725 522483
rect 185661 522423 185665 522479
rect 185665 522423 185721 522479
rect 185721 522423 185725 522479
rect 185661 522419 185725 522423
rect 174627 521935 174691 521939
rect 174627 521879 174631 521935
rect 174631 521879 174687 521935
rect 174687 521879 174691 521935
rect 174627 521875 174691 521879
rect 174707 521935 174771 521939
rect 174707 521879 174711 521935
rect 174711 521879 174767 521935
rect 174767 521879 174771 521935
rect 174707 521875 174771 521879
rect 174787 521935 174851 521939
rect 174787 521879 174791 521935
rect 174791 521879 174847 521935
rect 174847 521879 174851 521935
rect 174787 521875 174851 521879
rect 174867 521935 174931 521939
rect 174867 521879 174871 521935
rect 174871 521879 174927 521935
rect 174927 521879 174931 521935
rect 174867 521875 174931 521879
rect 178445 521935 178509 521939
rect 178445 521879 178449 521935
rect 178449 521879 178505 521935
rect 178505 521879 178509 521935
rect 178445 521875 178509 521879
rect 178525 521935 178589 521939
rect 178525 521879 178529 521935
rect 178529 521879 178585 521935
rect 178585 521879 178589 521935
rect 178525 521875 178589 521879
rect 178605 521935 178669 521939
rect 178605 521879 178609 521935
rect 178609 521879 178665 521935
rect 178665 521879 178669 521935
rect 178605 521875 178669 521879
rect 178685 521935 178749 521939
rect 178685 521879 178689 521935
rect 178689 521879 178745 521935
rect 178745 521879 178749 521935
rect 178685 521875 178749 521879
rect 182263 521935 182327 521939
rect 182263 521879 182267 521935
rect 182267 521879 182323 521935
rect 182323 521879 182327 521935
rect 182263 521875 182327 521879
rect 182343 521935 182407 521939
rect 182343 521879 182347 521935
rect 182347 521879 182403 521935
rect 182403 521879 182407 521935
rect 182343 521875 182407 521879
rect 182423 521935 182487 521939
rect 182423 521879 182427 521935
rect 182427 521879 182483 521935
rect 182483 521879 182487 521935
rect 182423 521875 182487 521879
rect 182503 521935 182567 521939
rect 182503 521879 182507 521935
rect 182507 521879 182563 521935
rect 182563 521879 182567 521935
rect 182503 521875 182567 521879
rect 186081 521935 186145 521939
rect 186081 521879 186085 521935
rect 186085 521879 186141 521935
rect 186141 521879 186145 521935
rect 186081 521875 186145 521879
rect 186161 521935 186225 521939
rect 186161 521879 186165 521935
rect 186165 521879 186221 521935
rect 186221 521879 186225 521935
rect 186161 521875 186225 521879
rect 186241 521935 186305 521939
rect 186241 521879 186245 521935
rect 186245 521879 186301 521935
rect 186301 521879 186305 521935
rect 186241 521875 186305 521879
rect 186321 521935 186385 521939
rect 186321 521879 186325 521935
rect 186325 521879 186381 521935
rect 186381 521879 186385 521935
rect 186321 521875 186385 521879
rect 173967 521391 174031 521395
rect 173967 521335 173971 521391
rect 173971 521335 174027 521391
rect 174027 521335 174031 521391
rect 173967 521331 174031 521335
rect 174047 521391 174111 521395
rect 174047 521335 174051 521391
rect 174051 521335 174107 521391
rect 174107 521335 174111 521391
rect 174047 521331 174111 521335
rect 174127 521391 174191 521395
rect 174127 521335 174131 521391
rect 174131 521335 174187 521391
rect 174187 521335 174191 521391
rect 174127 521331 174191 521335
rect 174207 521391 174271 521395
rect 174207 521335 174211 521391
rect 174211 521335 174267 521391
rect 174267 521335 174271 521391
rect 174207 521331 174271 521335
rect 177785 521391 177849 521395
rect 177785 521335 177789 521391
rect 177789 521335 177845 521391
rect 177845 521335 177849 521391
rect 177785 521331 177849 521335
rect 177865 521391 177929 521395
rect 177865 521335 177869 521391
rect 177869 521335 177925 521391
rect 177925 521335 177929 521391
rect 177865 521331 177929 521335
rect 177945 521391 178009 521395
rect 177945 521335 177949 521391
rect 177949 521335 178005 521391
rect 178005 521335 178009 521391
rect 177945 521331 178009 521335
rect 178025 521391 178089 521395
rect 178025 521335 178029 521391
rect 178029 521335 178085 521391
rect 178085 521335 178089 521391
rect 178025 521331 178089 521335
rect 181603 521391 181667 521395
rect 181603 521335 181607 521391
rect 181607 521335 181663 521391
rect 181663 521335 181667 521391
rect 181603 521331 181667 521335
rect 181683 521391 181747 521395
rect 181683 521335 181687 521391
rect 181687 521335 181743 521391
rect 181743 521335 181747 521391
rect 181683 521331 181747 521335
rect 181763 521391 181827 521395
rect 181763 521335 181767 521391
rect 181767 521335 181823 521391
rect 181823 521335 181827 521391
rect 181763 521331 181827 521335
rect 181843 521391 181907 521395
rect 181843 521335 181847 521391
rect 181847 521335 181903 521391
rect 181903 521335 181907 521391
rect 181843 521331 181907 521335
rect 185421 521391 185485 521395
rect 185421 521335 185425 521391
rect 185425 521335 185481 521391
rect 185481 521335 185485 521391
rect 185421 521331 185485 521335
rect 185501 521391 185565 521395
rect 185501 521335 185505 521391
rect 185505 521335 185561 521391
rect 185561 521335 185565 521391
rect 185501 521331 185565 521335
rect 185581 521391 185645 521395
rect 185581 521335 185585 521391
rect 185585 521335 185641 521391
rect 185641 521335 185645 521391
rect 185581 521331 185645 521335
rect 185661 521391 185725 521395
rect 185661 521335 185665 521391
rect 185665 521335 185721 521391
rect 185721 521335 185725 521391
rect 185661 521331 185725 521335
rect 174627 520847 174691 520851
rect 174627 520791 174631 520847
rect 174631 520791 174687 520847
rect 174687 520791 174691 520847
rect 174627 520787 174691 520791
rect 174707 520847 174771 520851
rect 174707 520791 174711 520847
rect 174711 520791 174767 520847
rect 174767 520791 174771 520847
rect 174707 520787 174771 520791
rect 174787 520847 174851 520851
rect 174787 520791 174791 520847
rect 174791 520791 174847 520847
rect 174847 520791 174851 520847
rect 174787 520787 174851 520791
rect 174867 520847 174931 520851
rect 174867 520791 174871 520847
rect 174871 520791 174927 520847
rect 174927 520791 174931 520847
rect 174867 520787 174931 520791
rect 178445 520847 178509 520851
rect 178445 520791 178449 520847
rect 178449 520791 178505 520847
rect 178505 520791 178509 520847
rect 178445 520787 178509 520791
rect 178525 520847 178589 520851
rect 178525 520791 178529 520847
rect 178529 520791 178585 520847
rect 178585 520791 178589 520847
rect 178525 520787 178589 520791
rect 178605 520847 178669 520851
rect 178605 520791 178609 520847
rect 178609 520791 178665 520847
rect 178665 520791 178669 520847
rect 178605 520787 178669 520791
rect 178685 520847 178749 520851
rect 178685 520791 178689 520847
rect 178689 520791 178745 520847
rect 178745 520791 178749 520847
rect 178685 520787 178749 520791
rect 182263 520847 182327 520851
rect 182263 520791 182267 520847
rect 182267 520791 182323 520847
rect 182323 520791 182327 520847
rect 182263 520787 182327 520791
rect 182343 520847 182407 520851
rect 182343 520791 182347 520847
rect 182347 520791 182403 520847
rect 182403 520791 182407 520847
rect 182343 520787 182407 520791
rect 182423 520847 182487 520851
rect 182423 520791 182427 520847
rect 182427 520791 182483 520847
rect 182483 520791 182487 520847
rect 182423 520787 182487 520791
rect 182503 520847 182567 520851
rect 182503 520791 182507 520847
rect 182507 520791 182563 520847
rect 182563 520791 182567 520847
rect 182503 520787 182567 520791
rect 186081 520847 186145 520851
rect 186081 520791 186085 520847
rect 186085 520791 186141 520847
rect 186141 520791 186145 520847
rect 186081 520787 186145 520791
rect 186161 520847 186225 520851
rect 186161 520791 186165 520847
rect 186165 520791 186221 520847
rect 186221 520791 186225 520847
rect 186161 520787 186225 520791
rect 186241 520847 186305 520851
rect 186241 520791 186245 520847
rect 186245 520791 186301 520847
rect 186301 520791 186305 520847
rect 186241 520787 186305 520791
rect 186321 520847 186385 520851
rect 186321 520791 186325 520847
rect 186325 520791 186381 520847
rect 186381 520791 186385 520847
rect 186321 520787 186385 520791
rect 173967 520303 174031 520307
rect 173967 520247 173971 520303
rect 173971 520247 174027 520303
rect 174027 520247 174031 520303
rect 173967 520243 174031 520247
rect 174047 520303 174111 520307
rect 174047 520247 174051 520303
rect 174051 520247 174107 520303
rect 174107 520247 174111 520303
rect 174047 520243 174111 520247
rect 174127 520303 174191 520307
rect 174127 520247 174131 520303
rect 174131 520247 174187 520303
rect 174187 520247 174191 520303
rect 174127 520243 174191 520247
rect 174207 520303 174271 520307
rect 174207 520247 174211 520303
rect 174211 520247 174267 520303
rect 174267 520247 174271 520303
rect 174207 520243 174271 520247
rect 177785 520303 177849 520307
rect 177785 520247 177789 520303
rect 177789 520247 177845 520303
rect 177845 520247 177849 520303
rect 177785 520243 177849 520247
rect 177865 520303 177929 520307
rect 177865 520247 177869 520303
rect 177869 520247 177925 520303
rect 177925 520247 177929 520303
rect 177865 520243 177929 520247
rect 177945 520303 178009 520307
rect 177945 520247 177949 520303
rect 177949 520247 178005 520303
rect 178005 520247 178009 520303
rect 177945 520243 178009 520247
rect 178025 520303 178089 520307
rect 178025 520247 178029 520303
rect 178029 520247 178085 520303
rect 178085 520247 178089 520303
rect 178025 520243 178089 520247
rect 181603 520303 181667 520307
rect 181603 520247 181607 520303
rect 181607 520247 181663 520303
rect 181663 520247 181667 520303
rect 181603 520243 181667 520247
rect 181683 520303 181747 520307
rect 181683 520247 181687 520303
rect 181687 520247 181743 520303
rect 181743 520247 181747 520303
rect 181683 520243 181747 520247
rect 181763 520303 181827 520307
rect 181763 520247 181767 520303
rect 181767 520247 181823 520303
rect 181823 520247 181827 520303
rect 181763 520243 181827 520247
rect 181843 520303 181907 520307
rect 181843 520247 181847 520303
rect 181847 520247 181903 520303
rect 181903 520247 181907 520303
rect 181843 520243 181907 520247
rect 185421 520303 185485 520307
rect 185421 520247 185425 520303
rect 185425 520247 185481 520303
rect 185481 520247 185485 520303
rect 185421 520243 185485 520247
rect 185501 520303 185565 520307
rect 185501 520247 185505 520303
rect 185505 520247 185561 520303
rect 185561 520247 185565 520303
rect 185501 520243 185565 520247
rect 185581 520303 185645 520307
rect 185581 520247 185585 520303
rect 185585 520247 185641 520303
rect 185641 520247 185645 520303
rect 185581 520243 185645 520247
rect 185661 520303 185725 520307
rect 185661 520247 185665 520303
rect 185665 520247 185721 520303
rect 185721 520247 185725 520303
rect 185661 520243 185725 520247
rect 174627 519759 174691 519763
rect 174627 519703 174631 519759
rect 174631 519703 174687 519759
rect 174687 519703 174691 519759
rect 174627 519699 174691 519703
rect 174707 519759 174771 519763
rect 174707 519703 174711 519759
rect 174711 519703 174767 519759
rect 174767 519703 174771 519759
rect 174707 519699 174771 519703
rect 174787 519759 174851 519763
rect 174787 519703 174791 519759
rect 174791 519703 174847 519759
rect 174847 519703 174851 519759
rect 174787 519699 174851 519703
rect 174867 519759 174931 519763
rect 174867 519703 174871 519759
rect 174871 519703 174927 519759
rect 174927 519703 174931 519759
rect 174867 519699 174931 519703
rect 178445 519759 178509 519763
rect 178445 519703 178449 519759
rect 178449 519703 178505 519759
rect 178505 519703 178509 519759
rect 178445 519699 178509 519703
rect 178525 519759 178589 519763
rect 178525 519703 178529 519759
rect 178529 519703 178585 519759
rect 178585 519703 178589 519759
rect 178525 519699 178589 519703
rect 178605 519759 178669 519763
rect 178605 519703 178609 519759
rect 178609 519703 178665 519759
rect 178665 519703 178669 519759
rect 178605 519699 178669 519703
rect 178685 519759 178749 519763
rect 178685 519703 178689 519759
rect 178689 519703 178745 519759
rect 178745 519703 178749 519759
rect 178685 519699 178749 519703
rect 182263 519759 182327 519763
rect 182263 519703 182267 519759
rect 182267 519703 182323 519759
rect 182323 519703 182327 519759
rect 182263 519699 182327 519703
rect 182343 519759 182407 519763
rect 182343 519703 182347 519759
rect 182347 519703 182403 519759
rect 182403 519703 182407 519759
rect 182343 519699 182407 519703
rect 182423 519759 182487 519763
rect 182423 519703 182427 519759
rect 182427 519703 182483 519759
rect 182483 519703 182487 519759
rect 182423 519699 182487 519703
rect 182503 519759 182567 519763
rect 182503 519703 182507 519759
rect 182507 519703 182563 519759
rect 182563 519703 182567 519759
rect 182503 519699 182567 519703
rect 186081 519759 186145 519763
rect 186081 519703 186085 519759
rect 186085 519703 186141 519759
rect 186141 519703 186145 519759
rect 186081 519699 186145 519703
rect 186161 519759 186225 519763
rect 186161 519703 186165 519759
rect 186165 519703 186221 519759
rect 186221 519703 186225 519759
rect 186161 519699 186225 519703
rect 186241 519759 186305 519763
rect 186241 519703 186245 519759
rect 186245 519703 186301 519759
rect 186301 519703 186305 519759
rect 186241 519699 186305 519703
rect 186321 519759 186385 519763
rect 186321 519703 186325 519759
rect 186325 519703 186381 519759
rect 186381 519703 186385 519759
rect 186321 519699 186385 519703
rect 173967 519215 174031 519219
rect 173967 519159 173971 519215
rect 173971 519159 174027 519215
rect 174027 519159 174031 519215
rect 173967 519155 174031 519159
rect 174047 519215 174111 519219
rect 174047 519159 174051 519215
rect 174051 519159 174107 519215
rect 174107 519159 174111 519215
rect 174047 519155 174111 519159
rect 174127 519215 174191 519219
rect 174127 519159 174131 519215
rect 174131 519159 174187 519215
rect 174187 519159 174191 519215
rect 174127 519155 174191 519159
rect 174207 519215 174271 519219
rect 174207 519159 174211 519215
rect 174211 519159 174267 519215
rect 174267 519159 174271 519215
rect 174207 519155 174271 519159
rect 177785 519215 177849 519219
rect 177785 519159 177789 519215
rect 177789 519159 177845 519215
rect 177845 519159 177849 519215
rect 177785 519155 177849 519159
rect 177865 519215 177929 519219
rect 177865 519159 177869 519215
rect 177869 519159 177925 519215
rect 177925 519159 177929 519215
rect 177865 519155 177929 519159
rect 177945 519215 178009 519219
rect 177945 519159 177949 519215
rect 177949 519159 178005 519215
rect 178005 519159 178009 519215
rect 177945 519155 178009 519159
rect 178025 519215 178089 519219
rect 178025 519159 178029 519215
rect 178029 519159 178085 519215
rect 178085 519159 178089 519215
rect 178025 519155 178089 519159
rect 181603 519215 181667 519219
rect 181603 519159 181607 519215
rect 181607 519159 181663 519215
rect 181663 519159 181667 519215
rect 181603 519155 181667 519159
rect 181683 519215 181747 519219
rect 181683 519159 181687 519215
rect 181687 519159 181743 519215
rect 181743 519159 181747 519215
rect 181683 519155 181747 519159
rect 181763 519215 181827 519219
rect 181763 519159 181767 519215
rect 181767 519159 181823 519215
rect 181823 519159 181827 519215
rect 181763 519155 181827 519159
rect 181843 519215 181907 519219
rect 181843 519159 181847 519215
rect 181847 519159 181903 519215
rect 181903 519159 181907 519215
rect 181843 519155 181907 519159
rect 185421 519215 185485 519219
rect 185421 519159 185425 519215
rect 185425 519159 185481 519215
rect 185481 519159 185485 519215
rect 185421 519155 185485 519159
rect 185501 519215 185565 519219
rect 185501 519159 185505 519215
rect 185505 519159 185561 519215
rect 185561 519159 185565 519215
rect 185501 519155 185565 519159
rect 185581 519215 185645 519219
rect 185581 519159 185585 519215
rect 185585 519159 185641 519215
rect 185641 519159 185645 519215
rect 185581 519155 185645 519159
rect 185661 519215 185725 519219
rect 185661 519159 185665 519215
rect 185665 519159 185721 519215
rect 185721 519159 185725 519215
rect 185661 519155 185725 519159
rect 174627 518671 174691 518675
rect 174627 518615 174631 518671
rect 174631 518615 174687 518671
rect 174687 518615 174691 518671
rect 174627 518611 174691 518615
rect 174707 518671 174771 518675
rect 174707 518615 174711 518671
rect 174711 518615 174767 518671
rect 174767 518615 174771 518671
rect 174707 518611 174771 518615
rect 174787 518671 174851 518675
rect 174787 518615 174791 518671
rect 174791 518615 174847 518671
rect 174847 518615 174851 518671
rect 174787 518611 174851 518615
rect 174867 518671 174931 518675
rect 174867 518615 174871 518671
rect 174871 518615 174927 518671
rect 174927 518615 174931 518671
rect 174867 518611 174931 518615
rect 178445 518671 178509 518675
rect 178445 518615 178449 518671
rect 178449 518615 178505 518671
rect 178505 518615 178509 518671
rect 178445 518611 178509 518615
rect 178525 518671 178589 518675
rect 178525 518615 178529 518671
rect 178529 518615 178585 518671
rect 178585 518615 178589 518671
rect 178525 518611 178589 518615
rect 178605 518671 178669 518675
rect 178605 518615 178609 518671
rect 178609 518615 178665 518671
rect 178665 518615 178669 518671
rect 178605 518611 178669 518615
rect 178685 518671 178749 518675
rect 178685 518615 178689 518671
rect 178689 518615 178745 518671
rect 178745 518615 178749 518671
rect 178685 518611 178749 518615
rect 182263 518671 182327 518675
rect 182263 518615 182267 518671
rect 182267 518615 182323 518671
rect 182323 518615 182327 518671
rect 182263 518611 182327 518615
rect 182343 518671 182407 518675
rect 182343 518615 182347 518671
rect 182347 518615 182403 518671
rect 182403 518615 182407 518671
rect 182343 518611 182407 518615
rect 182423 518671 182487 518675
rect 182423 518615 182427 518671
rect 182427 518615 182483 518671
rect 182483 518615 182487 518671
rect 182423 518611 182487 518615
rect 182503 518671 182567 518675
rect 182503 518615 182507 518671
rect 182507 518615 182563 518671
rect 182563 518615 182567 518671
rect 182503 518611 182567 518615
rect 186081 518671 186145 518675
rect 186081 518615 186085 518671
rect 186085 518615 186141 518671
rect 186141 518615 186145 518671
rect 186081 518611 186145 518615
rect 186161 518671 186225 518675
rect 186161 518615 186165 518671
rect 186165 518615 186221 518671
rect 186221 518615 186225 518671
rect 186161 518611 186225 518615
rect 186241 518671 186305 518675
rect 186241 518615 186245 518671
rect 186245 518615 186301 518671
rect 186301 518615 186305 518671
rect 186241 518611 186305 518615
rect 186321 518671 186385 518675
rect 186321 518615 186325 518671
rect 186325 518615 186381 518671
rect 186381 518615 186385 518671
rect 186321 518611 186385 518615
rect 173967 518127 174031 518131
rect 173967 518071 173971 518127
rect 173971 518071 174027 518127
rect 174027 518071 174031 518127
rect 173967 518067 174031 518071
rect 174047 518127 174111 518131
rect 174047 518071 174051 518127
rect 174051 518071 174107 518127
rect 174107 518071 174111 518127
rect 174047 518067 174111 518071
rect 174127 518127 174191 518131
rect 174127 518071 174131 518127
rect 174131 518071 174187 518127
rect 174187 518071 174191 518127
rect 174127 518067 174191 518071
rect 174207 518127 174271 518131
rect 174207 518071 174211 518127
rect 174211 518071 174267 518127
rect 174267 518071 174271 518127
rect 174207 518067 174271 518071
rect 177785 518127 177849 518131
rect 177785 518071 177789 518127
rect 177789 518071 177845 518127
rect 177845 518071 177849 518127
rect 177785 518067 177849 518071
rect 177865 518127 177929 518131
rect 177865 518071 177869 518127
rect 177869 518071 177925 518127
rect 177925 518071 177929 518127
rect 177865 518067 177929 518071
rect 177945 518127 178009 518131
rect 177945 518071 177949 518127
rect 177949 518071 178005 518127
rect 178005 518071 178009 518127
rect 177945 518067 178009 518071
rect 178025 518127 178089 518131
rect 178025 518071 178029 518127
rect 178029 518071 178085 518127
rect 178085 518071 178089 518127
rect 178025 518067 178089 518071
rect 181603 518127 181667 518131
rect 181603 518071 181607 518127
rect 181607 518071 181663 518127
rect 181663 518071 181667 518127
rect 181603 518067 181667 518071
rect 181683 518127 181747 518131
rect 181683 518071 181687 518127
rect 181687 518071 181743 518127
rect 181743 518071 181747 518127
rect 181683 518067 181747 518071
rect 181763 518127 181827 518131
rect 181763 518071 181767 518127
rect 181767 518071 181823 518127
rect 181823 518071 181827 518127
rect 181763 518067 181827 518071
rect 181843 518127 181907 518131
rect 181843 518071 181847 518127
rect 181847 518071 181903 518127
rect 181903 518071 181907 518127
rect 181843 518067 181907 518071
rect 185421 518127 185485 518131
rect 185421 518071 185425 518127
rect 185425 518071 185481 518127
rect 185481 518071 185485 518127
rect 185421 518067 185485 518071
rect 185501 518127 185565 518131
rect 185501 518071 185505 518127
rect 185505 518071 185561 518127
rect 185561 518071 185565 518127
rect 185501 518067 185565 518071
rect 185581 518127 185645 518131
rect 185581 518071 185585 518127
rect 185585 518071 185641 518127
rect 185641 518071 185645 518127
rect 185581 518067 185645 518071
rect 185661 518127 185725 518131
rect 185661 518071 185665 518127
rect 185665 518071 185721 518127
rect 185721 518071 185725 518127
rect 185661 518067 185725 518071
rect 174627 517583 174691 517587
rect 174627 517527 174631 517583
rect 174631 517527 174687 517583
rect 174687 517527 174691 517583
rect 174627 517523 174691 517527
rect 174707 517583 174771 517587
rect 174707 517527 174711 517583
rect 174711 517527 174767 517583
rect 174767 517527 174771 517583
rect 174707 517523 174771 517527
rect 174787 517583 174851 517587
rect 174787 517527 174791 517583
rect 174791 517527 174847 517583
rect 174847 517527 174851 517583
rect 174787 517523 174851 517527
rect 174867 517583 174931 517587
rect 174867 517527 174871 517583
rect 174871 517527 174927 517583
rect 174927 517527 174931 517583
rect 174867 517523 174931 517527
rect 178445 517583 178509 517587
rect 178445 517527 178449 517583
rect 178449 517527 178505 517583
rect 178505 517527 178509 517583
rect 178445 517523 178509 517527
rect 178525 517583 178589 517587
rect 178525 517527 178529 517583
rect 178529 517527 178585 517583
rect 178585 517527 178589 517583
rect 178525 517523 178589 517527
rect 178605 517583 178669 517587
rect 178605 517527 178609 517583
rect 178609 517527 178665 517583
rect 178665 517527 178669 517583
rect 178605 517523 178669 517527
rect 178685 517583 178749 517587
rect 178685 517527 178689 517583
rect 178689 517527 178745 517583
rect 178745 517527 178749 517583
rect 178685 517523 178749 517527
rect 182263 517583 182327 517587
rect 182263 517527 182267 517583
rect 182267 517527 182323 517583
rect 182323 517527 182327 517583
rect 182263 517523 182327 517527
rect 182343 517583 182407 517587
rect 182343 517527 182347 517583
rect 182347 517527 182403 517583
rect 182403 517527 182407 517583
rect 182343 517523 182407 517527
rect 182423 517583 182487 517587
rect 182423 517527 182427 517583
rect 182427 517527 182483 517583
rect 182483 517527 182487 517583
rect 182423 517523 182487 517527
rect 182503 517583 182567 517587
rect 182503 517527 182507 517583
rect 182507 517527 182563 517583
rect 182563 517527 182567 517583
rect 182503 517523 182567 517527
rect 186081 517583 186145 517587
rect 186081 517527 186085 517583
rect 186085 517527 186141 517583
rect 186141 517527 186145 517583
rect 186081 517523 186145 517527
rect 186161 517583 186225 517587
rect 186161 517527 186165 517583
rect 186165 517527 186221 517583
rect 186221 517527 186225 517583
rect 186161 517523 186225 517527
rect 186241 517583 186305 517587
rect 186241 517527 186245 517583
rect 186245 517527 186301 517583
rect 186301 517527 186305 517583
rect 186241 517523 186305 517527
rect 186321 517583 186385 517587
rect 186321 517527 186325 517583
rect 186325 517527 186381 517583
rect 186381 517527 186385 517583
rect 186321 517523 186385 517527
rect 173967 517039 174031 517043
rect 173967 516983 173971 517039
rect 173971 516983 174027 517039
rect 174027 516983 174031 517039
rect 173967 516979 174031 516983
rect 174047 517039 174111 517043
rect 174047 516983 174051 517039
rect 174051 516983 174107 517039
rect 174107 516983 174111 517039
rect 174047 516979 174111 516983
rect 174127 517039 174191 517043
rect 174127 516983 174131 517039
rect 174131 516983 174187 517039
rect 174187 516983 174191 517039
rect 174127 516979 174191 516983
rect 174207 517039 174271 517043
rect 174207 516983 174211 517039
rect 174211 516983 174267 517039
rect 174267 516983 174271 517039
rect 174207 516979 174271 516983
rect 177785 517039 177849 517043
rect 177785 516983 177789 517039
rect 177789 516983 177845 517039
rect 177845 516983 177849 517039
rect 177785 516979 177849 516983
rect 177865 517039 177929 517043
rect 177865 516983 177869 517039
rect 177869 516983 177925 517039
rect 177925 516983 177929 517039
rect 177865 516979 177929 516983
rect 177945 517039 178009 517043
rect 177945 516983 177949 517039
rect 177949 516983 178005 517039
rect 178005 516983 178009 517039
rect 177945 516979 178009 516983
rect 178025 517039 178089 517043
rect 178025 516983 178029 517039
rect 178029 516983 178085 517039
rect 178085 516983 178089 517039
rect 178025 516979 178089 516983
rect 181603 517039 181667 517043
rect 181603 516983 181607 517039
rect 181607 516983 181663 517039
rect 181663 516983 181667 517039
rect 181603 516979 181667 516983
rect 181683 517039 181747 517043
rect 181683 516983 181687 517039
rect 181687 516983 181743 517039
rect 181743 516983 181747 517039
rect 181683 516979 181747 516983
rect 181763 517039 181827 517043
rect 181763 516983 181767 517039
rect 181767 516983 181823 517039
rect 181823 516983 181827 517039
rect 181763 516979 181827 516983
rect 181843 517039 181907 517043
rect 181843 516983 181847 517039
rect 181847 516983 181903 517039
rect 181903 516983 181907 517039
rect 181843 516979 181907 516983
rect 185421 517039 185485 517043
rect 185421 516983 185425 517039
rect 185425 516983 185481 517039
rect 185481 516983 185485 517039
rect 185421 516979 185485 516983
rect 185501 517039 185565 517043
rect 185501 516983 185505 517039
rect 185505 516983 185561 517039
rect 185561 516983 185565 517039
rect 185501 516979 185565 516983
rect 185581 517039 185645 517043
rect 185581 516983 185585 517039
rect 185585 516983 185641 517039
rect 185641 516983 185645 517039
rect 185581 516979 185645 516983
rect 185661 517039 185725 517043
rect 185661 516983 185665 517039
rect 185665 516983 185721 517039
rect 185721 516983 185725 517039
rect 185661 516979 185725 516983
rect 174627 516495 174691 516499
rect 174627 516439 174631 516495
rect 174631 516439 174687 516495
rect 174687 516439 174691 516495
rect 174627 516435 174691 516439
rect 174707 516495 174771 516499
rect 174707 516439 174711 516495
rect 174711 516439 174767 516495
rect 174767 516439 174771 516495
rect 174707 516435 174771 516439
rect 174787 516495 174851 516499
rect 174787 516439 174791 516495
rect 174791 516439 174847 516495
rect 174847 516439 174851 516495
rect 174787 516435 174851 516439
rect 174867 516495 174931 516499
rect 174867 516439 174871 516495
rect 174871 516439 174927 516495
rect 174927 516439 174931 516495
rect 174867 516435 174931 516439
rect 178445 516495 178509 516499
rect 178445 516439 178449 516495
rect 178449 516439 178505 516495
rect 178505 516439 178509 516495
rect 178445 516435 178509 516439
rect 178525 516495 178589 516499
rect 178525 516439 178529 516495
rect 178529 516439 178585 516495
rect 178585 516439 178589 516495
rect 178525 516435 178589 516439
rect 178605 516495 178669 516499
rect 178605 516439 178609 516495
rect 178609 516439 178665 516495
rect 178665 516439 178669 516495
rect 178605 516435 178669 516439
rect 178685 516495 178749 516499
rect 178685 516439 178689 516495
rect 178689 516439 178745 516495
rect 178745 516439 178749 516495
rect 178685 516435 178749 516439
rect 182263 516495 182327 516499
rect 182263 516439 182267 516495
rect 182267 516439 182323 516495
rect 182323 516439 182327 516495
rect 182263 516435 182327 516439
rect 182343 516495 182407 516499
rect 182343 516439 182347 516495
rect 182347 516439 182403 516495
rect 182403 516439 182407 516495
rect 182343 516435 182407 516439
rect 182423 516495 182487 516499
rect 182423 516439 182427 516495
rect 182427 516439 182483 516495
rect 182483 516439 182487 516495
rect 182423 516435 182487 516439
rect 182503 516495 182567 516499
rect 182503 516439 182507 516495
rect 182507 516439 182563 516495
rect 182563 516439 182567 516495
rect 182503 516435 182567 516439
rect 186081 516495 186145 516499
rect 186081 516439 186085 516495
rect 186085 516439 186141 516495
rect 186141 516439 186145 516495
rect 186081 516435 186145 516439
rect 186161 516495 186225 516499
rect 186161 516439 186165 516495
rect 186165 516439 186221 516495
rect 186221 516439 186225 516495
rect 186161 516435 186225 516439
rect 186241 516495 186305 516499
rect 186241 516439 186245 516495
rect 186245 516439 186301 516495
rect 186301 516439 186305 516495
rect 186241 516435 186305 516439
rect 186321 516495 186385 516499
rect 186321 516439 186325 516495
rect 186325 516439 186381 516495
rect 186381 516439 186385 516495
rect 186321 516435 186385 516439
rect 173967 515951 174031 515955
rect 173967 515895 173971 515951
rect 173971 515895 174027 515951
rect 174027 515895 174031 515951
rect 173967 515891 174031 515895
rect 174047 515951 174111 515955
rect 174047 515895 174051 515951
rect 174051 515895 174107 515951
rect 174107 515895 174111 515951
rect 174047 515891 174111 515895
rect 174127 515951 174191 515955
rect 174127 515895 174131 515951
rect 174131 515895 174187 515951
rect 174187 515895 174191 515951
rect 174127 515891 174191 515895
rect 174207 515951 174271 515955
rect 174207 515895 174211 515951
rect 174211 515895 174267 515951
rect 174267 515895 174271 515951
rect 174207 515891 174271 515895
rect 177785 515951 177849 515955
rect 177785 515895 177789 515951
rect 177789 515895 177845 515951
rect 177845 515895 177849 515951
rect 177785 515891 177849 515895
rect 177865 515951 177929 515955
rect 177865 515895 177869 515951
rect 177869 515895 177925 515951
rect 177925 515895 177929 515951
rect 177865 515891 177929 515895
rect 177945 515951 178009 515955
rect 177945 515895 177949 515951
rect 177949 515895 178005 515951
rect 178005 515895 178009 515951
rect 177945 515891 178009 515895
rect 178025 515951 178089 515955
rect 178025 515895 178029 515951
rect 178029 515895 178085 515951
rect 178085 515895 178089 515951
rect 178025 515891 178089 515895
rect 181603 515951 181667 515955
rect 181603 515895 181607 515951
rect 181607 515895 181663 515951
rect 181663 515895 181667 515951
rect 181603 515891 181667 515895
rect 181683 515951 181747 515955
rect 181683 515895 181687 515951
rect 181687 515895 181743 515951
rect 181743 515895 181747 515951
rect 181683 515891 181747 515895
rect 181763 515951 181827 515955
rect 181763 515895 181767 515951
rect 181767 515895 181823 515951
rect 181823 515895 181827 515951
rect 181763 515891 181827 515895
rect 181843 515951 181907 515955
rect 181843 515895 181847 515951
rect 181847 515895 181903 515951
rect 181903 515895 181907 515951
rect 181843 515891 181907 515895
rect 185421 515951 185485 515955
rect 185421 515895 185425 515951
rect 185425 515895 185481 515951
rect 185481 515895 185485 515951
rect 185421 515891 185485 515895
rect 185501 515951 185565 515955
rect 185501 515895 185505 515951
rect 185505 515895 185561 515951
rect 185561 515895 185565 515951
rect 185501 515891 185565 515895
rect 185581 515951 185645 515955
rect 185581 515895 185585 515951
rect 185585 515895 185641 515951
rect 185641 515895 185645 515951
rect 185581 515891 185645 515895
rect 185661 515951 185725 515955
rect 185661 515895 185665 515951
rect 185665 515895 185721 515951
rect 185721 515895 185725 515951
rect 185661 515891 185725 515895
rect 174627 515407 174691 515411
rect 174627 515351 174631 515407
rect 174631 515351 174687 515407
rect 174687 515351 174691 515407
rect 174627 515347 174691 515351
rect 174707 515407 174771 515411
rect 174707 515351 174711 515407
rect 174711 515351 174767 515407
rect 174767 515351 174771 515407
rect 174707 515347 174771 515351
rect 174787 515407 174851 515411
rect 174787 515351 174791 515407
rect 174791 515351 174847 515407
rect 174847 515351 174851 515407
rect 174787 515347 174851 515351
rect 174867 515407 174931 515411
rect 174867 515351 174871 515407
rect 174871 515351 174927 515407
rect 174927 515351 174931 515407
rect 174867 515347 174931 515351
rect 178445 515407 178509 515411
rect 178445 515351 178449 515407
rect 178449 515351 178505 515407
rect 178505 515351 178509 515407
rect 178445 515347 178509 515351
rect 178525 515407 178589 515411
rect 178525 515351 178529 515407
rect 178529 515351 178585 515407
rect 178585 515351 178589 515407
rect 178525 515347 178589 515351
rect 178605 515407 178669 515411
rect 178605 515351 178609 515407
rect 178609 515351 178665 515407
rect 178665 515351 178669 515407
rect 178605 515347 178669 515351
rect 178685 515407 178749 515411
rect 178685 515351 178689 515407
rect 178689 515351 178745 515407
rect 178745 515351 178749 515407
rect 178685 515347 178749 515351
rect 182263 515407 182327 515411
rect 182263 515351 182267 515407
rect 182267 515351 182323 515407
rect 182323 515351 182327 515407
rect 182263 515347 182327 515351
rect 182343 515407 182407 515411
rect 182343 515351 182347 515407
rect 182347 515351 182403 515407
rect 182403 515351 182407 515407
rect 182343 515347 182407 515351
rect 182423 515407 182487 515411
rect 182423 515351 182427 515407
rect 182427 515351 182483 515407
rect 182483 515351 182487 515407
rect 182423 515347 182487 515351
rect 182503 515407 182567 515411
rect 182503 515351 182507 515407
rect 182507 515351 182563 515407
rect 182563 515351 182567 515407
rect 182503 515347 182567 515351
rect 186081 515407 186145 515411
rect 186081 515351 186085 515407
rect 186085 515351 186141 515407
rect 186141 515351 186145 515407
rect 186081 515347 186145 515351
rect 186161 515407 186225 515411
rect 186161 515351 186165 515407
rect 186165 515351 186221 515407
rect 186221 515351 186225 515407
rect 186161 515347 186225 515351
rect 186241 515407 186305 515411
rect 186241 515351 186245 515407
rect 186245 515351 186301 515407
rect 186301 515351 186305 515407
rect 186241 515347 186305 515351
rect 186321 515407 186385 515411
rect 186321 515351 186325 515407
rect 186325 515351 186381 515407
rect 186381 515351 186385 515407
rect 186321 515347 186385 515351
<< mimcap >>
rect 157711 541757 162511 541797
rect 157711 539037 157751 541757
rect 162471 539037 162511 541757
rect 157711 538997 162511 539037
<< mimcapcontact >>
rect 157751 539037 162471 541757
<< metal4 >>
rect 162610 541869 162706 541885
rect 157750 541757 162472 541758
rect 157750 539037 157751 541757
rect 162471 539037 162472 541757
rect 157750 539036 162472 539037
rect 159390 538687 159490 539036
rect 162610 538925 162626 541869
rect 162690 539112 162706 541869
rect 162690 538925 162765 539112
rect 162610 538909 162765 538925
rect 162630 538837 162765 538909
rect 159390 538587 159400 538687
rect 159480 538587 159490 538687
rect 159390 538577 159490 538587
rect 161380 538747 162765 538837
rect 161380 538697 161530 538747
rect 161380 538577 161390 538697
rect 161510 538577 161530 538697
rect 161380 538567 161530 538577
rect 173959 530099 174279 530659
rect 173959 530035 173967 530099
rect 174031 530035 174047 530099
rect 174111 530035 174127 530099
rect 174191 530035 174207 530099
rect 174271 530035 174279 530099
rect 173959 529011 174279 530035
rect 173959 528947 173967 529011
rect 174031 528947 174047 529011
rect 174111 528947 174127 529011
rect 174191 528947 174207 529011
rect 174271 528947 174279 529011
rect 173959 528825 174279 528947
rect 173959 528589 174001 528825
rect 174237 528589 174279 528825
rect 173959 527923 174279 528589
rect 173959 527859 173967 527923
rect 174031 527859 174047 527923
rect 174111 527859 174127 527923
rect 174191 527859 174207 527923
rect 174271 527859 174279 527923
rect 173959 526835 174279 527859
rect 173959 526771 173967 526835
rect 174031 526771 174047 526835
rect 174111 526771 174127 526835
rect 174191 526771 174207 526835
rect 174271 526771 174279 526835
rect 173959 525747 174279 526771
rect 173959 525683 173967 525747
rect 174031 525683 174047 525747
rect 174111 525683 174127 525747
rect 174191 525683 174207 525747
rect 174271 525683 174279 525747
rect 173959 525017 174279 525683
rect 173959 524781 174001 525017
rect 174237 524781 174279 525017
rect 173959 524659 174279 524781
rect 173959 524595 173967 524659
rect 174031 524595 174047 524659
rect 174111 524595 174127 524659
rect 174191 524595 174207 524659
rect 174271 524595 174279 524659
rect 173959 523571 174279 524595
rect 173959 523507 173967 523571
rect 174031 523507 174047 523571
rect 174111 523507 174127 523571
rect 174191 523507 174207 523571
rect 174271 523507 174279 523571
rect 173959 522483 174279 523507
rect 173959 522419 173967 522483
rect 174031 522419 174047 522483
rect 174111 522419 174127 522483
rect 174191 522419 174207 522483
rect 174271 522419 174279 522483
rect 173959 521395 174279 522419
rect 173959 521331 173967 521395
rect 174031 521331 174047 521395
rect 174111 521331 174127 521395
rect 174191 521331 174207 521395
rect 174271 521331 174279 521395
rect 173959 521209 174279 521331
rect 173959 520973 174001 521209
rect 174237 520973 174279 521209
rect 173959 520307 174279 520973
rect 173959 520243 173967 520307
rect 174031 520243 174047 520307
rect 174111 520243 174127 520307
rect 174191 520243 174207 520307
rect 174271 520243 174279 520307
rect 173959 519219 174279 520243
rect 173959 519155 173967 519219
rect 174031 519155 174047 519219
rect 174111 519155 174127 519219
rect 174191 519155 174207 519219
rect 174271 519155 174279 519219
rect 173959 518131 174279 519155
rect 173959 518067 173967 518131
rect 174031 518067 174047 518131
rect 174111 518067 174127 518131
rect 174191 518067 174207 518131
rect 174271 518067 174279 518131
rect 173959 517401 174279 518067
rect 173959 517165 174001 517401
rect 174237 517165 174279 517401
rect 173959 517043 174279 517165
rect 173959 516979 173967 517043
rect 174031 516979 174047 517043
rect 174111 516979 174127 517043
rect 174191 516979 174207 517043
rect 174271 516979 174279 517043
rect 173959 515955 174279 516979
rect 173959 515891 173967 515955
rect 174031 515891 174047 515955
rect 174111 515891 174127 515955
rect 174191 515891 174207 515955
rect 174271 515891 174279 515955
rect 173959 515331 174279 515891
rect 174619 530643 174939 530659
rect 174619 530579 174627 530643
rect 174691 530579 174707 530643
rect 174771 530579 174787 530643
rect 174851 530579 174867 530643
rect 174931 530579 174939 530643
rect 174619 529555 174939 530579
rect 174619 529491 174627 529555
rect 174691 529491 174707 529555
rect 174771 529491 174787 529555
rect 174851 529491 174867 529555
rect 174931 529491 174939 529555
rect 174619 528467 174939 529491
rect 174619 528403 174627 528467
rect 174691 528403 174707 528467
rect 174771 528403 174787 528467
rect 174851 528403 174867 528467
rect 174931 528403 174939 528467
rect 174619 528165 174939 528403
rect 174619 527929 174661 528165
rect 174897 527929 174939 528165
rect 174619 527379 174939 527929
rect 174619 527315 174627 527379
rect 174691 527315 174707 527379
rect 174771 527315 174787 527379
rect 174851 527315 174867 527379
rect 174931 527315 174939 527379
rect 174619 526291 174939 527315
rect 174619 526227 174627 526291
rect 174691 526227 174707 526291
rect 174771 526227 174787 526291
rect 174851 526227 174867 526291
rect 174931 526227 174939 526291
rect 174619 525203 174939 526227
rect 174619 525139 174627 525203
rect 174691 525139 174707 525203
rect 174771 525139 174787 525203
rect 174851 525139 174867 525203
rect 174931 525139 174939 525203
rect 174619 524357 174939 525139
rect 174619 524121 174661 524357
rect 174897 524121 174939 524357
rect 174619 524115 174939 524121
rect 174619 524051 174627 524115
rect 174691 524051 174707 524115
rect 174771 524051 174787 524115
rect 174851 524051 174867 524115
rect 174931 524051 174939 524115
rect 174619 523027 174939 524051
rect 174619 522963 174627 523027
rect 174691 522963 174707 523027
rect 174771 522963 174787 523027
rect 174851 522963 174867 523027
rect 174931 522963 174939 523027
rect 174619 521939 174939 522963
rect 174619 521875 174627 521939
rect 174691 521875 174707 521939
rect 174771 521875 174787 521939
rect 174851 521875 174867 521939
rect 174931 521875 174939 521939
rect 174619 520851 174939 521875
rect 174619 520787 174627 520851
rect 174691 520787 174707 520851
rect 174771 520787 174787 520851
rect 174851 520787 174867 520851
rect 174931 520787 174939 520851
rect 174619 520549 174939 520787
rect 174619 520313 174661 520549
rect 174897 520313 174939 520549
rect 174619 519763 174939 520313
rect 174619 519699 174627 519763
rect 174691 519699 174707 519763
rect 174771 519699 174787 519763
rect 174851 519699 174867 519763
rect 174931 519699 174939 519763
rect 174619 518675 174939 519699
rect 174619 518611 174627 518675
rect 174691 518611 174707 518675
rect 174771 518611 174787 518675
rect 174851 518611 174867 518675
rect 174931 518611 174939 518675
rect 174619 517587 174939 518611
rect 174619 517523 174627 517587
rect 174691 517523 174707 517587
rect 174771 517523 174787 517587
rect 174851 517523 174867 517587
rect 174931 517523 174939 517587
rect 174619 516741 174939 517523
rect 174619 516505 174661 516741
rect 174897 516505 174939 516741
rect 174619 516499 174939 516505
rect 174619 516435 174627 516499
rect 174691 516435 174707 516499
rect 174771 516435 174787 516499
rect 174851 516435 174867 516499
rect 174931 516435 174939 516499
rect 174619 515411 174939 516435
rect 174619 515347 174627 515411
rect 174691 515347 174707 515411
rect 174771 515347 174787 515411
rect 174851 515347 174867 515411
rect 174931 515347 174939 515411
rect 174619 515331 174939 515347
rect 177777 530099 178097 530659
rect 177777 530035 177785 530099
rect 177849 530035 177865 530099
rect 177929 530035 177945 530099
rect 178009 530035 178025 530099
rect 178089 530035 178097 530099
rect 177777 529011 178097 530035
rect 177777 528947 177785 529011
rect 177849 528947 177865 529011
rect 177929 528947 177945 529011
rect 178009 528947 178025 529011
rect 178089 528947 178097 529011
rect 177777 528825 178097 528947
rect 177777 528589 177819 528825
rect 178055 528589 178097 528825
rect 177777 527923 178097 528589
rect 177777 527859 177785 527923
rect 177849 527859 177865 527923
rect 177929 527859 177945 527923
rect 178009 527859 178025 527923
rect 178089 527859 178097 527923
rect 177777 526835 178097 527859
rect 177777 526771 177785 526835
rect 177849 526771 177865 526835
rect 177929 526771 177945 526835
rect 178009 526771 178025 526835
rect 178089 526771 178097 526835
rect 177777 525747 178097 526771
rect 177777 525683 177785 525747
rect 177849 525683 177865 525747
rect 177929 525683 177945 525747
rect 178009 525683 178025 525747
rect 178089 525683 178097 525747
rect 177777 525017 178097 525683
rect 177777 524781 177819 525017
rect 178055 524781 178097 525017
rect 177777 524659 178097 524781
rect 177777 524595 177785 524659
rect 177849 524595 177865 524659
rect 177929 524595 177945 524659
rect 178009 524595 178025 524659
rect 178089 524595 178097 524659
rect 177777 523571 178097 524595
rect 177777 523507 177785 523571
rect 177849 523507 177865 523571
rect 177929 523507 177945 523571
rect 178009 523507 178025 523571
rect 178089 523507 178097 523571
rect 177777 522483 178097 523507
rect 177777 522419 177785 522483
rect 177849 522419 177865 522483
rect 177929 522419 177945 522483
rect 178009 522419 178025 522483
rect 178089 522419 178097 522483
rect 177777 521395 178097 522419
rect 177777 521331 177785 521395
rect 177849 521331 177865 521395
rect 177929 521331 177945 521395
rect 178009 521331 178025 521395
rect 178089 521331 178097 521395
rect 177777 521209 178097 521331
rect 177777 520973 177819 521209
rect 178055 520973 178097 521209
rect 177777 520307 178097 520973
rect 177777 520243 177785 520307
rect 177849 520243 177865 520307
rect 177929 520243 177945 520307
rect 178009 520243 178025 520307
rect 178089 520243 178097 520307
rect 177777 519219 178097 520243
rect 177777 519155 177785 519219
rect 177849 519155 177865 519219
rect 177929 519155 177945 519219
rect 178009 519155 178025 519219
rect 178089 519155 178097 519219
rect 177777 518131 178097 519155
rect 177777 518067 177785 518131
rect 177849 518067 177865 518131
rect 177929 518067 177945 518131
rect 178009 518067 178025 518131
rect 178089 518067 178097 518131
rect 177777 517401 178097 518067
rect 177777 517165 177819 517401
rect 178055 517165 178097 517401
rect 177777 517043 178097 517165
rect 177777 516979 177785 517043
rect 177849 516979 177865 517043
rect 177929 516979 177945 517043
rect 178009 516979 178025 517043
rect 178089 516979 178097 517043
rect 177777 515955 178097 516979
rect 177777 515891 177785 515955
rect 177849 515891 177865 515955
rect 177929 515891 177945 515955
rect 178009 515891 178025 515955
rect 178089 515891 178097 515955
rect 177777 515331 178097 515891
rect 178437 530643 178757 530659
rect 178437 530579 178445 530643
rect 178509 530579 178525 530643
rect 178589 530579 178605 530643
rect 178669 530579 178685 530643
rect 178749 530579 178757 530643
rect 178437 529555 178757 530579
rect 178437 529491 178445 529555
rect 178509 529491 178525 529555
rect 178589 529491 178605 529555
rect 178669 529491 178685 529555
rect 178749 529491 178757 529555
rect 178437 528467 178757 529491
rect 178437 528403 178445 528467
rect 178509 528403 178525 528467
rect 178589 528403 178605 528467
rect 178669 528403 178685 528467
rect 178749 528403 178757 528467
rect 178437 528165 178757 528403
rect 178437 527929 178479 528165
rect 178715 527929 178757 528165
rect 178437 527379 178757 527929
rect 178437 527315 178445 527379
rect 178509 527315 178525 527379
rect 178589 527315 178605 527379
rect 178669 527315 178685 527379
rect 178749 527315 178757 527379
rect 178437 526291 178757 527315
rect 178437 526227 178445 526291
rect 178509 526227 178525 526291
rect 178589 526227 178605 526291
rect 178669 526227 178685 526291
rect 178749 526227 178757 526291
rect 178437 525203 178757 526227
rect 178437 525139 178445 525203
rect 178509 525139 178525 525203
rect 178589 525139 178605 525203
rect 178669 525139 178685 525203
rect 178749 525139 178757 525203
rect 178437 524357 178757 525139
rect 178437 524121 178479 524357
rect 178715 524121 178757 524357
rect 178437 524115 178757 524121
rect 178437 524051 178445 524115
rect 178509 524051 178525 524115
rect 178589 524051 178605 524115
rect 178669 524051 178685 524115
rect 178749 524051 178757 524115
rect 178437 523027 178757 524051
rect 178437 522963 178445 523027
rect 178509 522963 178525 523027
rect 178589 522963 178605 523027
rect 178669 522963 178685 523027
rect 178749 522963 178757 523027
rect 178437 521939 178757 522963
rect 178437 521875 178445 521939
rect 178509 521875 178525 521939
rect 178589 521875 178605 521939
rect 178669 521875 178685 521939
rect 178749 521875 178757 521939
rect 178437 520851 178757 521875
rect 178437 520787 178445 520851
rect 178509 520787 178525 520851
rect 178589 520787 178605 520851
rect 178669 520787 178685 520851
rect 178749 520787 178757 520851
rect 178437 520549 178757 520787
rect 178437 520313 178479 520549
rect 178715 520313 178757 520549
rect 178437 519763 178757 520313
rect 178437 519699 178445 519763
rect 178509 519699 178525 519763
rect 178589 519699 178605 519763
rect 178669 519699 178685 519763
rect 178749 519699 178757 519763
rect 178437 518675 178757 519699
rect 178437 518611 178445 518675
rect 178509 518611 178525 518675
rect 178589 518611 178605 518675
rect 178669 518611 178685 518675
rect 178749 518611 178757 518675
rect 178437 517587 178757 518611
rect 178437 517523 178445 517587
rect 178509 517523 178525 517587
rect 178589 517523 178605 517587
rect 178669 517523 178685 517587
rect 178749 517523 178757 517587
rect 178437 516741 178757 517523
rect 178437 516505 178479 516741
rect 178715 516505 178757 516741
rect 178437 516499 178757 516505
rect 178437 516435 178445 516499
rect 178509 516435 178525 516499
rect 178589 516435 178605 516499
rect 178669 516435 178685 516499
rect 178749 516435 178757 516499
rect 178437 515411 178757 516435
rect 178437 515347 178445 515411
rect 178509 515347 178525 515411
rect 178589 515347 178605 515411
rect 178669 515347 178685 515411
rect 178749 515347 178757 515411
rect 178437 515331 178757 515347
rect 181595 530099 181915 530659
rect 181595 530035 181603 530099
rect 181667 530035 181683 530099
rect 181747 530035 181763 530099
rect 181827 530035 181843 530099
rect 181907 530035 181915 530099
rect 181595 529011 181915 530035
rect 181595 528947 181603 529011
rect 181667 528947 181683 529011
rect 181747 528947 181763 529011
rect 181827 528947 181843 529011
rect 181907 528947 181915 529011
rect 181595 528825 181915 528947
rect 181595 528589 181637 528825
rect 181873 528589 181915 528825
rect 181595 527923 181915 528589
rect 181595 527859 181603 527923
rect 181667 527859 181683 527923
rect 181747 527859 181763 527923
rect 181827 527859 181843 527923
rect 181907 527859 181915 527923
rect 181595 526835 181915 527859
rect 181595 526771 181603 526835
rect 181667 526771 181683 526835
rect 181747 526771 181763 526835
rect 181827 526771 181843 526835
rect 181907 526771 181915 526835
rect 181595 525747 181915 526771
rect 181595 525683 181603 525747
rect 181667 525683 181683 525747
rect 181747 525683 181763 525747
rect 181827 525683 181843 525747
rect 181907 525683 181915 525747
rect 181595 525017 181915 525683
rect 181595 524781 181637 525017
rect 181873 524781 181915 525017
rect 181595 524659 181915 524781
rect 181595 524595 181603 524659
rect 181667 524595 181683 524659
rect 181747 524595 181763 524659
rect 181827 524595 181843 524659
rect 181907 524595 181915 524659
rect 181595 523571 181915 524595
rect 181595 523507 181603 523571
rect 181667 523507 181683 523571
rect 181747 523507 181763 523571
rect 181827 523507 181843 523571
rect 181907 523507 181915 523571
rect 181595 522483 181915 523507
rect 181595 522419 181603 522483
rect 181667 522419 181683 522483
rect 181747 522419 181763 522483
rect 181827 522419 181843 522483
rect 181907 522419 181915 522483
rect 181595 521395 181915 522419
rect 181595 521331 181603 521395
rect 181667 521331 181683 521395
rect 181747 521331 181763 521395
rect 181827 521331 181843 521395
rect 181907 521331 181915 521395
rect 181595 521209 181915 521331
rect 181595 520973 181637 521209
rect 181873 520973 181915 521209
rect 181595 520307 181915 520973
rect 181595 520243 181603 520307
rect 181667 520243 181683 520307
rect 181747 520243 181763 520307
rect 181827 520243 181843 520307
rect 181907 520243 181915 520307
rect 181595 519219 181915 520243
rect 181595 519155 181603 519219
rect 181667 519155 181683 519219
rect 181747 519155 181763 519219
rect 181827 519155 181843 519219
rect 181907 519155 181915 519219
rect 181595 518131 181915 519155
rect 181595 518067 181603 518131
rect 181667 518067 181683 518131
rect 181747 518067 181763 518131
rect 181827 518067 181843 518131
rect 181907 518067 181915 518131
rect 181595 517401 181915 518067
rect 181595 517165 181637 517401
rect 181873 517165 181915 517401
rect 181595 517043 181915 517165
rect 181595 516979 181603 517043
rect 181667 516979 181683 517043
rect 181747 516979 181763 517043
rect 181827 516979 181843 517043
rect 181907 516979 181915 517043
rect 181595 515955 181915 516979
rect 181595 515891 181603 515955
rect 181667 515891 181683 515955
rect 181747 515891 181763 515955
rect 181827 515891 181843 515955
rect 181907 515891 181915 515955
rect 181595 515331 181915 515891
rect 182255 530643 182575 530659
rect 182255 530579 182263 530643
rect 182327 530579 182343 530643
rect 182407 530579 182423 530643
rect 182487 530579 182503 530643
rect 182567 530579 182575 530643
rect 182255 529555 182575 530579
rect 182255 529491 182263 529555
rect 182327 529491 182343 529555
rect 182407 529491 182423 529555
rect 182487 529491 182503 529555
rect 182567 529491 182575 529555
rect 182255 528467 182575 529491
rect 182255 528403 182263 528467
rect 182327 528403 182343 528467
rect 182407 528403 182423 528467
rect 182487 528403 182503 528467
rect 182567 528403 182575 528467
rect 182255 528165 182575 528403
rect 182255 527929 182297 528165
rect 182533 527929 182575 528165
rect 182255 527379 182575 527929
rect 182255 527315 182263 527379
rect 182327 527315 182343 527379
rect 182407 527315 182423 527379
rect 182487 527315 182503 527379
rect 182567 527315 182575 527379
rect 182255 526291 182575 527315
rect 182255 526227 182263 526291
rect 182327 526227 182343 526291
rect 182407 526227 182423 526291
rect 182487 526227 182503 526291
rect 182567 526227 182575 526291
rect 182255 525203 182575 526227
rect 182255 525139 182263 525203
rect 182327 525139 182343 525203
rect 182407 525139 182423 525203
rect 182487 525139 182503 525203
rect 182567 525139 182575 525203
rect 182255 524357 182575 525139
rect 182255 524121 182297 524357
rect 182533 524121 182575 524357
rect 182255 524115 182575 524121
rect 182255 524051 182263 524115
rect 182327 524051 182343 524115
rect 182407 524051 182423 524115
rect 182487 524051 182503 524115
rect 182567 524051 182575 524115
rect 182255 523027 182575 524051
rect 182255 522963 182263 523027
rect 182327 522963 182343 523027
rect 182407 522963 182423 523027
rect 182487 522963 182503 523027
rect 182567 522963 182575 523027
rect 182255 521939 182575 522963
rect 182255 521875 182263 521939
rect 182327 521875 182343 521939
rect 182407 521875 182423 521939
rect 182487 521875 182503 521939
rect 182567 521875 182575 521939
rect 182255 520851 182575 521875
rect 182255 520787 182263 520851
rect 182327 520787 182343 520851
rect 182407 520787 182423 520851
rect 182487 520787 182503 520851
rect 182567 520787 182575 520851
rect 182255 520549 182575 520787
rect 182255 520313 182297 520549
rect 182533 520313 182575 520549
rect 182255 519763 182575 520313
rect 182255 519699 182263 519763
rect 182327 519699 182343 519763
rect 182407 519699 182423 519763
rect 182487 519699 182503 519763
rect 182567 519699 182575 519763
rect 182255 518675 182575 519699
rect 182255 518611 182263 518675
rect 182327 518611 182343 518675
rect 182407 518611 182423 518675
rect 182487 518611 182503 518675
rect 182567 518611 182575 518675
rect 182255 517587 182575 518611
rect 182255 517523 182263 517587
rect 182327 517523 182343 517587
rect 182407 517523 182423 517587
rect 182487 517523 182503 517587
rect 182567 517523 182575 517587
rect 182255 516741 182575 517523
rect 182255 516505 182297 516741
rect 182533 516505 182575 516741
rect 182255 516499 182575 516505
rect 182255 516435 182263 516499
rect 182327 516435 182343 516499
rect 182407 516435 182423 516499
rect 182487 516435 182503 516499
rect 182567 516435 182575 516499
rect 182255 515411 182575 516435
rect 182255 515347 182263 515411
rect 182327 515347 182343 515411
rect 182407 515347 182423 515411
rect 182487 515347 182503 515411
rect 182567 515347 182575 515411
rect 182255 515331 182575 515347
rect 185413 530099 185733 530659
rect 185413 530035 185421 530099
rect 185485 530035 185501 530099
rect 185565 530035 185581 530099
rect 185645 530035 185661 530099
rect 185725 530035 185733 530099
rect 185413 529011 185733 530035
rect 185413 528947 185421 529011
rect 185485 528947 185501 529011
rect 185565 528947 185581 529011
rect 185645 528947 185661 529011
rect 185725 528947 185733 529011
rect 185413 528825 185733 528947
rect 185413 528589 185455 528825
rect 185691 528589 185733 528825
rect 185413 527923 185733 528589
rect 185413 527859 185421 527923
rect 185485 527859 185501 527923
rect 185565 527859 185581 527923
rect 185645 527859 185661 527923
rect 185725 527859 185733 527923
rect 185413 526835 185733 527859
rect 185413 526771 185421 526835
rect 185485 526771 185501 526835
rect 185565 526771 185581 526835
rect 185645 526771 185661 526835
rect 185725 526771 185733 526835
rect 185413 525747 185733 526771
rect 185413 525683 185421 525747
rect 185485 525683 185501 525747
rect 185565 525683 185581 525747
rect 185645 525683 185661 525747
rect 185725 525683 185733 525747
rect 185413 525017 185733 525683
rect 185413 524781 185455 525017
rect 185691 524781 185733 525017
rect 185413 524659 185733 524781
rect 185413 524595 185421 524659
rect 185485 524595 185501 524659
rect 185565 524595 185581 524659
rect 185645 524595 185661 524659
rect 185725 524595 185733 524659
rect 185413 523571 185733 524595
rect 185413 523507 185421 523571
rect 185485 523507 185501 523571
rect 185565 523507 185581 523571
rect 185645 523507 185661 523571
rect 185725 523507 185733 523571
rect 185413 522483 185733 523507
rect 185413 522419 185421 522483
rect 185485 522419 185501 522483
rect 185565 522419 185581 522483
rect 185645 522419 185661 522483
rect 185725 522419 185733 522483
rect 185413 521395 185733 522419
rect 185413 521331 185421 521395
rect 185485 521331 185501 521395
rect 185565 521331 185581 521395
rect 185645 521331 185661 521395
rect 185725 521331 185733 521395
rect 185413 521209 185733 521331
rect 185413 520973 185455 521209
rect 185691 520973 185733 521209
rect 185413 520307 185733 520973
rect 185413 520243 185421 520307
rect 185485 520243 185501 520307
rect 185565 520243 185581 520307
rect 185645 520243 185661 520307
rect 185725 520243 185733 520307
rect 185413 519219 185733 520243
rect 185413 519155 185421 519219
rect 185485 519155 185501 519219
rect 185565 519155 185581 519219
rect 185645 519155 185661 519219
rect 185725 519155 185733 519219
rect 185413 518131 185733 519155
rect 185413 518067 185421 518131
rect 185485 518067 185501 518131
rect 185565 518067 185581 518131
rect 185645 518067 185661 518131
rect 185725 518067 185733 518131
rect 185413 517401 185733 518067
rect 185413 517165 185455 517401
rect 185691 517165 185733 517401
rect 185413 517043 185733 517165
rect 185413 516979 185421 517043
rect 185485 516979 185501 517043
rect 185565 516979 185581 517043
rect 185645 516979 185661 517043
rect 185725 516979 185733 517043
rect 185413 515955 185733 516979
rect 185413 515891 185421 515955
rect 185485 515891 185501 515955
rect 185565 515891 185581 515955
rect 185645 515891 185661 515955
rect 185725 515891 185733 515955
rect 185413 515331 185733 515891
rect 186073 530643 186393 530659
rect 186073 530579 186081 530643
rect 186145 530579 186161 530643
rect 186225 530579 186241 530643
rect 186305 530579 186321 530643
rect 186385 530579 186393 530643
rect 186073 529555 186393 530579
rect 186073 529491 186081 529555
rect 186145 529491 186161 529555
rect 186225 529491 186241 529555
rect 186305 529491 186321 529555
rect 186385 529491 186393 529555
rect 186073 528467 186393 529491
rect 186073 528403 186081 528467
rect 186145 528403 186161 528467
rect 186225 528403 186241 528467
rect 186305 528403 186321 528467
rect 186385 528403 186393 528467
rect 186073 528165 186393 528403
rect 186073 527929 186115 528165
rect 186351 527929 186393 528165
rect 186073 527379 186393 527929
rect 186073 527315 186081 527379
rect 186145 527315 186161 527379
rect 186225 527315 186241 527379
rect 186305 527315 186321 527379
rect 186385 527315 186393 527379
rect 186073 526291 186393 527315
rect 186073 526227 186081 526291
rect 186145 526227 186161 526291
rect 186225 526227 186241 526291
rect 186305 526227 186321 526291
rect 186385 526227 186393 526291
rect 186073 525203 186393 526227
rect 186073 525139 186081 525203
rect 186145 525139 186161 525203
rect 186225 525139 186241 525203
rect 186305 525139 186321 525203
rect 186385 525139 186393 525203
rect 186073 524357 186393 525139
rect 186073 524121 186115 524357
rect 186351 524121 186393 524357
rect 186073 524115 186393 524121
rect 186073 524051 186081 524115
rect 186145 524051 186161 524115
rect 186225 524051 186241 524115
rect 186305 524051 186321 524115
rect 186385 524051 186393 524115
rect 186073 523027 186393 524051
rect 186073 522963 186081 523027
rect 186145 522963 186161 523027
rect 186225 522963 186241 523027
rect 186305 522963 186321 523027
rect 186385 522963 186393 523027
rect 186073 521939 186393 522963
rect 186073 521875 186081 521939
rect 186145 521875 186161 521939
rect 186225 521875 186241 521939
rect 186305 521875 186321 521939
rect 186385 521875 186393 521939
rect 186073 520851 186393 521875
rect 186073 520787 186081 520851
rect 186145 520787 186161 520851
rect 186225 520787 186241 520851
rect 186305 520787 186321 520851
rect 186385 520787 186393 520851
rect 186073 520549 186393 520787
rect 186073 520313 186115 520549
rect 186351 520313 186393 520549
rect 186073 519763 186393 520313
rect 186073 519699 186081 519763
rect 186145 519699 186161 519763
rect 186225 519699 186241 519763
rect 186305 519699 186321 519763
rect 186385 519699 186393 519763
rect 186073 518675 186393 519699
rect 186073 518611 186081 518675
rect 186145 518611 186161 518675
rect 186225 518611 186241 518675
rect 186305 518611 186321 518675
rect 186385 518611 186393 518675
rect 186073 517587 186393 518611
rect 186073 517523 186081 517587
rect 186145 517523 186161 517587
rect 186225 517523 186241 517587
rect 186305 517523 186321 517587
rect 186385 517523 186393 517587
rect 186073 516741 186393 517523
rect 186073 516505 186115 516741
rect 186351 516505 186393 516741
rect 186073 516499 186393 516505
rect 186073 516435 186081 516499
rect 186145 516435 186161 516499
rect 186225 516435 186241 516499
rect 186305 516435 186321 516499
rect 186385 516435 186393 516499
rect 186073 515411 186393 516435
rect 186073 515347 186081 515411
rect 186145 515347 186161 515411
rect 186225 515347 186241 515411
rect 186305 515347 186321 515411
rect 186385 515347 186393 515411
rect 186073 515331 186393 515347
<< via4 >>
rect 174001 528589 174237 528825
rect 174001 524781 174237 525017
rect 174001 520973 174237 521209
rect 174001 517165 174237 517401
rect 174661 527929 174897 528165
rect 174661 524121 174897 524357
rect 174661 520313 174897 520549
rect 174661 516505 174897 516741
rect 177819 528589 178055 528825
rect 177819 524781 178055 525017
rect 177819 520973 178055 521209
rect 177819 517165 178055 517401
rect 178479 527929 178715 528165
rect 178479 524121 178715 524357
rect 178479 520313 178715 520549
rect 178479 516505 178715 516741
rect 181637 528589 181873 528825
rect 181637 524781 181873 525017
rect 181637 520973 181873 521209
rect 181637 517165 181873 517401
rect 182297 527929 182533 528165
rect 182297 524121 182533 524357
rect 182297 520313 182533 520549
rect 182297 516505 182533 516741
rect 185455 528589 185691 528825
rect 185455 524781 185691 525017
rect 185455 520973 185691 521209
rect 185455 517165 185691 517401
rect 186115 527929 186351 528165
rect 186115 524121 186351 524357
rect 186115 520313 186351 520549
rect 186115 516505 186351 516741
<< metal5 >>
rect 172162 528825 187530 528867
rect 172162 528589 174001 528825
rect 174237 528589 177819 528825
rect 178055 528589 181637 528825
rect 181873 528589 185455 528825
rect 185691 528589 187530 528825
rect 172162 528547 187530 528589
rect 172162 528165 187530 528207
rect 172162 527929 174661 528165
rect 174897 527929 178479 528165
rect 178715 527929 182297 528165
rect 182533 527929 186115 528165
rect 186351 527929 187530 528165
rect 172162 527887 187530 527929
rect 172162 525017 187530 525059
rect 172162 524781 174001 525017
rect 174237 524781 177819 525017
rect 178055 524781 181637 525017
rect 181873 524781 185455 525017
rect 185691 524781 187530 525017
rect 172162 524739 187530 524781
rect 172162 524357 187530 524399
rect 172162 524121 174661 524357
rect 174897 524121 178479 524357
rect 178715 524121 182297 524357
rect 182533 524121 186115 524357
rect 186351 524121 187530 524357
rect 172162 524079 187530 524121
rect 172162 521209 187530 521251
rect 172162 520973 174001 521209
rect 174237 520973 177819 521209
rect 178055 520973 181637 521209
rect 181873 520973 185455 521209
rect 185691 520973 187530 521209
rect 172162 520931 187530 520973
rect 172162 520549 187530 520591
rect 172162 520313 174661 520549
rect 174897 520313 178479 520549
rect 178715 520313 182297 520549
rect 182533 520313 186115 520549
rect 186351 520313 187530 520549
rect 172162 520271 187530 520313
rect 172162 517401 187530 517443
rect 172162 517165 174001 517401
rect 174237 517165 177819 517401
rect 178055 517165 181637 517401
rect 181873 517165 185455 517401
rect 185691 517165 187530 517401
rect 172162 517123 187530 517165
rect 172162 516741 187530 516783
rect 172162 516505 174661 516741
rect 174897 516505 178479 516741
rect 178715 516505 182297 516741
rect 182533 516505 186115 516741
rect 186351 516505 187530 516741
rect 172162 516463 187530 516505
<< res0p35 >>
rect 164316 536463 164390 537551
rect 164634 536463 164708 537551
rect 164952 536463 165026 537551
rect 165270 536463 165344 537551
rect 165588 536463 165662 537551
rect 165906 536463 165980 537551
rect 166224 536463 166298 537551
rect 166542 536463 166616 537551
rect 168088 536463 168162 537551
rect 168406 536463 168480 537551
rect 168724 536463 168798 537551
rect 169042 536463 169116 537551
rect 171824 536463 171898 537551
rect 172142 536463 172216 537551
rect 175342 536463 175416 537551
rect 178942 537023 179016 537551
rect 182242 537303 182316 537551
rect 185542 537443 185616 537551
rect 188842 537347 188916 537551
rect 164286 534123 164360 535211
rect 164604 534123 164678 535211
rect 164922 534123 164996 535211
rect 165240 534123 165314 535211
rect 165558 534123 165632 535211
rect 165876 534123 165950 535211
rect 166194 534123 166268 535211
rect 166512 534123 166586 535211
<< labels >>
flabel metal1 193000 521000 195000 523000 0 FreeSans 1600 0 0 0 gnd_spi
port 71 nsew
flabel metal1 193000 524000 195000 526000 0 FreeSans 1600 0 0 0 vd_spi
port 73 nsew
flabel metal3 s 614 378318 1894 378430 0 FreeSans 1120 0 0 0 reset
port 64 nsew signal input
flabel metal3 s 600 421540 1880 421652 0 FreeSans 1120 0 0 0 sdi
port 63 nsew signal input
flabel metal3 s 600 464762 1880 464874 0 FreeSans 1120 0 0 0 sclk
port 62 nsew signal input
flabel metal3 s 600 507984 1880 508096 0 FreeSans 1120 0 0 0 ss
port 61 nsew signal input
flabel metal3 s 1400 680242 3100 685242 0 FreeSans 1120 0 0 0 ib
port 37 nsew signal bidirectional
flabel metal3 s 16194 700900 21194 703400 0 FreeSans 1920 180 0 0 inp
port 46 nsew signal bidirectional
flabel metal3 s 68194 700900 73194 703400 0 FreeSans 1920 180 0 0 inn
port 45 nsew signal bidirectional
flabel metal3 s 120194 700900 125194 703400 0 FreeSans 1920 180 0 0 out
port 44 nsew signal bidirectional
flabel metal1 193000 540036 195000 542036 0 FreeSans 1600 0 0 0 gnd_ota
port 70 nsew
flabel metal1 193000 537356 195000 539356 0 FreeSans 1600 0 0 0 vd_ota
port 68 nsew
flabel space 163530 542597 163730 542787 0 FreeSans 1600 0 0 0 dpga_flat_0.inp
flabel metal2 186230 513087 186430 513277 0 FreeSans 1600 0 0 0 dpga_flat_0.reset
flabel metal2 181910 513127 182110 513317 0 FreeSans 1600 0 0 0 dpga_flat_0.sdi
flabel metal1 192430 539147 192630 539347 0 FreeSans 1600 0 0 0 dpga_flat_0.vd
flabel metal1 192430 540087 192630 540287 0 FreeSans 1600 0 0 0 dpga_flat_0.gnd
flabel metal1 178180 542747 178380 542947 0 FreeSans 1600 0 0 0 dpga_flat_0.inn
flabel metal1 163530 542787 163730 542987 0 FreeSans 1600 0 0 0 dpga_flat_0.inp
flabel metal1 156800 536797 157000 536997 0 FreeSans 1600 0 0 0 dpga_flat_0.out
flabel metal1 163030 533147 163230 533347 0 FreeSans 1600 0 0 0 dpga_flat_0.ib
flabel metal1 192430 522907 192630 523097 0 FreeSans 1600 0 0 0 dpga_flat_0.gndd
flabel metal2 177580 513127 177780 513317 0 FreeSans 1600 0 0 0 dpga_flat_0.sclk
flabel metal2 173250 513127 173450 513317 0 FreeSans 1600 0 0 0 dpga_flat_0.ss
flabel metal1 192430 523427 192630 523617 0 FreeSans 1600 0 0 0 dpga_flat_0.vpwr
flabel metal1 190922 522999 191012 523017 0 FreeSans 1600 0 0 0 dpga_flat_0.vgnd
flabel metal4 174619 515331 174939 530659 0 FreeSans 1920 90 0 0 dpga_flat_0.sr_0.VGND
flabel metal4 178437 515331 178757 530659 0 FreeSans 1920 90 0 0 dpga_flat_0.sr_0.VGND
flabel metal4 182255 515331 182575 530659 0 FreeSans 1920 90 0 0 dpga_flat_0.sr_0.VGND
flabel metal4 186073 515331 186393 530659 0 FreeSans 1920 90 0 0 dpga_flat_0.sr_0.VGND
flabel metal5 172162 527887 187530 528207 0 FreeSans 2560 0 0 0 dpga_flat_0.sr_0.VGND
flabel metal5 172162 524079 187530 524399 0 FreeSans 2560 0 0 0 dpga_flat_0.sr_0.VGND
flabel metal5 172162 520271 187530 520591 0 FreeSans 2560 0 0 0 dpga_flat_0.sr_0.VGND
flabel metal5 172162 516463 187530 516783 0 FreeSans 2560 0 0 0 dpga_flat_0.sr_0.VGND
flabel metal4 173959 515331 174279 530659 0 FreeSans 1920 90 0 0 dpga_flat_0.sr_0.VPWR
flabel metal4 177777 515331 178097 530659 0 FreeSans 1920 90 0 0 dpga_flat_0.sr_0.VPWR
flabel metal4 181595 515331 181915 530659 0 FreeSans 1920 90 0 0 dpga_flat_0.sr_0.VPWR
flabel metal4 185413 515331 185733 530659 0 FreeSans 1920 90 0 0 dpga_flat_0.sr_0.VPWR
flabel metal5 172162 528547 187530 528867 0 FreeSans 2560 0 0 0 dpga_flat_0.sr_0.VPWR
flabel metal5 172162 524739 187530 525059 0 FreeSans 2560 0 0 0 dpga_flat_0.sr_0.VPWR
flabel metal5 172162 520931 187530 521251 0 FreeSans 2560 0 0 0 dpga_flat_0.sr_0.VPWR
flabel metal5 172162 517123 187530 517443 0 FreeSans 2560 0 0 0 dpga_flat_0.sr_0.VPWR
flabel metal2 172412 531987 172468 532787 0 FreeSans 224 90 0 0 dpga_flat_0.sr_0.data[0]
flabel metal2 174528 531987 174584 532787 0 FreeSans 224 90 0 0 dpga_flat_0.sr_0.data[1]
flabel metal2 176644 531987 176700 532787 0 FreeSans 224 90 0 0 dpga_flat_0.sr_0.data[2]
flabel metal2 178760 531987 178816 532787 0 FreeSans 224 90 0 0 dpga_flat_0.sr_0.data[3]
flabel metal2 180876 531987 180932 532787 0 FreeSans 224 90 0 0 dpga_flat_0.sr_0.data[4]
flabel metal2 182992 531987 183048 532787 0 FreeSans 224 90 0 0 dpga_flat_0.sr_0.data[5]
flabel metal2 185108 531987 185164 532787 0 FreeSans 224 90 0 0 dpga_flat_0.sr_0.data[6]
flabel metal2 187224 531987 187280 532787 0 FreeSans 224 90 0 0 dpga_flat_0.sr_0.data[7]
flabel metal2 186304 513131 186360 513931 0 FreeSans 224 90 0 0 dpga_flat_0.sr_0.reset
flabel metal2 177656 513131 177712 513931 0 FreeSans 224 90 0 0 dpga_flat_0.sr_0.sclk
flabel metal2 181980 513131 182036 513931 0 FreeSans 224 90 0 0 dpga_flat_0.sr_0.sdi
flabel metal2 173332 513131 173388 513931 0 FreeSans 224 90 0 0 dpga_flat_0.sr_0.ss
rlabel metal1 179846 515379 179846 515379 0 dpga_flat_0.sr_0.VGND
rlabel metal1 179846 515923 179846 515923 0 dpga_flat_0.sr_0.VPWR
rlabel metal1 176626 529829 176626 529829 0 dpga_flat_0.sr_0._00_
rlabel metal1 178374 530169 178374 530169 0 dpga_flat_0.sr_0._01_
rlabel metal2 179892 529625 179892 529625 0 dpga_flat_0.sr_0._02_
rlabel metal1 181180 529829 181180 529829 0 dpga_flat_0.sr_0._03_
rlabel metal1 180720 528741 180720 528741 0 dpga_flat_0.sr_0._04_
rlabel metal1 176856 530305 176856 530305 0 dpga_flat_0.sr_0._05_
rlabel metal2 176396 528401 176396 528401 0 dpga_flat_0.sr_0._06_
rlabel metal1 175890 529081 175890 529081 0 dpga_flat_0.sr_0._07_
rlabel metal1 177132 528537 177132 528537 0 dpga_flat_0.sr_0._08_
rlabel metal1 178236 529897 178236 529897 0 dpga_flat_0.sr_0._09_
rlabel metal1 178788 530373 178788 530373 0 dpga_flat_0.sr_0._10_
rlabel metal1 179984 530169 179984 530169 0 dpga_flat_0.sr_0._11_
rlabel metal1 182330 530237 182330 530237 0 dpga_flat_0.sr_0._12_
rlabel metal1 180398 528673 180398 528673 0 dpga_flat_0.sr_0._13_
rlabel metal2 177684 529081 177684 529081 0 dpga_flat_0.sr_0.clknet_0_sclk
rlabel metal1 176166 529081 176166 529081 0 dpga_flat_0.sr_0.clknet_1_0__leaf_sclk
rlabel metal2 180536 528911 180536 528911 0 dpga_flat_0.sr_0.clknet_1_1__leaf_sclk
rlabel metal2 172440 531233 172440 531233 0 dpga_flat_0.sr_0.data[0]
rlabel metal2 174556 531233 174556 531233 0 dpga_flat_0.sr_0.data[1]
rlabel metal2 176672 531828 176672 531828 0 dpga_flat_0.sr_0.data[2]
rlabel metal2 178788 531828 178788 531828 0 dpga_flat_0.sr_0.data[3]
rlabel metal2 180904 530995 180904 530995 0 dpga_flat_0.sr_0.data[4]
rlabel metal2 183020 531267 183020 531267 0 dpga_flat_0.sr_0.data[5]
rlabel metal2 185136 531267 185136 531267 0 dpga_flat_0.sr_0.data[6]
rlabel metal1 176895 529761 176895 529761 0 dpga_flat_0.sr_0.net1
rlabel metal1 182100 530373 182100 530373 0 dpga_flat_0.sr_0.net10
rlabel metal2 187252 531760 187252 531760 0 dpga_flat_0.sr_0.net11
rlabel metal1 175430 529625 175430 529625 0 dpga_flat_0.sr_0.net12
rlabel metal1 177178 528673 177178 528673 0 dpga_flat_0.sr_0.net13
rlabel metal1 176258 528673 176258 528673 0 dpga_flat_0.sr_0.net14
rlabel metal1 179340 528095 179340 528095 0 dpga_flat_0.sr_0.net15
rlabel metal1 182054 530305 182054 530305 0 dpga_flat_0.sr_0.net16
rlabel metal2 177684 529931 177684 529931 0 dpga_flat_0.sr_0.net17
rlabel metal1 181732 515821 181732 515821 0 dpga_flat_0.sr_0.net2
rlabel metal1 174464 529217 174464 529217 0 dpga_flat_0.sr_0.net3
rlabel metal2 174832 530101 174832 530101 0 dpga_flat_0.sr_0.net4
rlabel metal2 176764 528435 176764 528435 0 dpga_flat_0.sr_0.net5
rlabel metal2 178236 529353 178236 529353 0 dpga_flat_0.sr_0.net6
rlabel metal1 177960 529795 177960 529795 0 dpga_flat_0.sr_0.net7
rlabel metal1 178972 529965 178972 529965 0 dpga_flat_0.sr_0.net8
rlabel metal1 182606 529829 182606 529829 0 dpga_flat_0.sr_0.net9
rlabel metal2 186516 514682 186516 514682 0 dpga_flat_0.sr_0.reset
rlabel metal2 177684 515641 177684 515641 0 dpga_flat_0.sr_0.sclk
rlabel metal1 182238 515617 182238 515617 0 dpga_flat_0.sr_0.sdi
rlabel metal1 173452 515549 173452 515549 0 dpga_flat_0.sr_0.ss
flabel metal1 173067 530594 173101 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_9.VGND
flabel metal1 173067 530050 173101 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_9.VPWR
flabel nwell 173067 530050 173101 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_9.VPB
flabel pwell 173067 530594 173101 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_9.VNB
rlabel comment 173038 530611 173038 530611 2 dpga_flat_0.sr_0.FILLER_0_0_9.decap_12
flabel metal1 172515 529506 172549 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_3.VGND
flabel metal1 172515 530050 172549 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_3.VPWR
flabel nwell 172515 530050 172549 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_3.VPB
flabel pwell 172515 529506 172549 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_3.VNB
rlabel comment 172486 529523 172486 529523 4 dpga_flat_0.sr_0.FILLER_0_1_3.decap_12
flabel metal1 173619 529506 173653 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_15.VGND
flabel metal1 173619 530050 173653 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_15.VPWR
flabel nwell 173619 530050 173653 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_15.VPB
flabel pwell 173619 529506 173653 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_15.VNB
rlabel comment 173590 529523 173590 529523 4 dpga_flat_0.sr_0.FILLER_0_1_15.decap_12
flabel metal1 172239 530050 172273 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_0_Left_28.VPWR
flabel metal1 172239 530594 172273 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_0_Left_28.VGND
flabel nwell 172239 530050 172273 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_0_Left_28.VPB
flabel pwell 172239 530594 172273 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_0_Left_28.VNB
rlabel comment 172210 530611 172210 530611 2 dpga_flat_0.sr_0.PHY_EDGE_ROW_0_Left_28.decap_3
rlabel metal1 172210 530563 172486 530659 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_0_Left_28.VGND
rlabel metal1 172210 530019 172486 530115 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_0_Left_28.VPWR
flabel metal1 172239 530050 172273 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_1_Left_29.VPWR
flabel metal1 172239 529506 172273 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_1_Left_29.VGND
flabel nwell 172239 530050 172273 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_1_Left_29.VPB
flabel pwell 172239 529506 172273 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_1_Left_29.VNB
rlabel comment 172210 529523 172210 529523 4 dpga_flat_0.sr_0.PHY_EDGE_ROW_1_Left_29.decap_3
rlabel metal1 172210 529475 172486 529571 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_1_Left_29.VGND
rlabel metal1 172210 530019 172486 530115 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_1_Left_29.VPWR
flabel locali 172607 530288 172641 530322 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output4.X
flabel locali 172883 530424 172917 530458 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output4.A
flabel locali 172515 530424 172549 530458 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output4.X
flabel locali 172883 530356 172917 530390 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output4.A
flabel locali 172515 530356 172549 530390 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output4.X
flabel metal1 172975 530594 173009 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output4.VGND
flabel metal1 172975 530050 173009 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output4.VPWR
flabel nwell 172975 530050 173009 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output4.VPB
flabel pwell 172975 530594 173009 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output4.VNB
rlabel comment 173038 530611 173038 530611 8 dpga_flat_0.sr_0.output4.clkbuf_4
rlabel metal1 172486 530563 173038 530659 5 dpga_flat_0.sr_0.output4.VGND
rlabel metal1 172486 530019 173038 530115 5 dpga_flat_0.sr_0.output4.VPWR
flabel metal1 174171 530050 174205 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_21.VPWR
flabel metal1 174171 530594 174205 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_21.VGND
flabel nwell 174171 530050 174205 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_21.VPB
flabel pwell 174171 530594 174205 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_21.VNB
rlabel comment 174142 530611 174142 530611 2 dpga_flat_0.sr_0.FILLER_0_0_21.decap_6
rlabel metal1 174142 530563 174694 530659 5 dpga_flat_0.sr_0.FILLER_0_0_21.VGND
rlabel metal1 174142 530019 174694 530115 5 dpga_flat_0.sr_0.FILLER_0_0_21.VPWR
flabel metal1 174716 530054 174752 530084 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_27.VPWR
flabel metal1 174716 530595 174752 530624 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_27.VGND
flabel nwell 174725 530060 174745 530077 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_27.VPB
flabel pwell 174722 530600 174746 530622 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_27.VNB
rlabel comment 174694 530611 174694 530611 2 dpga_flat_0.sr_0.FILLER_0_0_27.fill_1
rlabel metal1 174694 530563 174786 530659 5 dpga_flat_0.sr_0.FILLER_0_0_27.VGND
rlabel metal1 174694 530019 174786 530115 5 dpga_flat_0.sr_0.FILLER_0_0_27.VPWR
flabel metal1 175452 530054 175488 530084 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_35.VPWR
flabel metal1 175452 530595 175488 530624 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_35.VGND
flabel nwell 175461 530060 175481 530077 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_35.VPB
flabel pwell 175458 530600 175482 530622 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_35.VNB
rlabel comment 175430 530611 175430 530611 2 dpga_flat_0.sr_0.FILLER_0_0_35.fill_1
rlabel metal1 175430 530563 175522 530659 5 dpga_flat_0.sr_0.FILLER_0_0_35.VGND
rlabel metal1 175430 530019 175522 530115 5 dpga_flat_0.sr_0.FILLER_0_0_35.VPWR
flabel metal1 174716 530050 174752 530080 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_27.VPWR
flabel metal1 174716 529510 174752 529539 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_27.VGND
flabel nwell 174725 530057 174745 530074 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_27.VPB
flabel pwell 174722 529512 174746 529534 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_27.VNB
rlabel comment 174694 529523 174694 529523 4 dpga_flat_0.sr_0.FILLER_0_1_27.fill_1
rlabel metal1 174694 529475 174786 529571 1 dpga_flat_0.sr_0.FILLER_0_1_27.VGND
rlabel metal1 174694 530019 174786 530115 1 dpga_flat_0.sr_0.FILLER_0_1_27.VPWR
flabel metal1 174808 530058 174861 530087 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_56.VPWR
flabel metal1 174807 530591 174858 530629 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_56.VGND
rlabel comment 174786 530611 174786 530611 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_56.tapvpwrvgnd_1
rlabel metal1 174786 530563 174878 530659 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_56.VGND
rlabel metal1 174786 530019 174878 530115 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_56.VPWR
flabel locali 175552 530152 175586 530186 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._28_.Q
flabel locali 175552 530220 175586 530254 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._28_.Q
flabel locali 175552 530288 175586 530322 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._28_.Q
flabel locali 175552 530492 175586 530526 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._28_.Q
flabel locali 175847 530424 175881 530458 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._28_.RESET_B
flabel locali 177023 530288 177057 530322 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._28_.D
flabel locali 177298 530288 177332 530322 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._28_.CLK
flabel locali 177298 530356 177332 530390 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._28_.CLK
flabel locali 175847 530356 175881 530390 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._28_.RESET_B
flabel metal1 177299 530594 177333 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._28_.VGND
flabel metal1 177299 530050 177333 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._28_.VPWR
flabel nwell 177299 530050 177333 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._28_.VPB
flabel pwell 177299 530594 177333 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._28_.VNB
rlabel comment 177362 530611 177362 530611 8 dpga_flat_0.sr_0._28_.dfrtp_1
rlabel locali 175833 530404 175881 530484 5 dpga_flat_0.sr_0._28_.RESET_B
rlabel locali 175833 530330 175941 530404 5 dpga_flat_0.sr_0._28_.RESET_B
rlabel metal1 175835 530455 175893 530464 5 dpga_flat_0.sr_0._28_.RESET_B
rlabel metal1 175895 530355 175953 530418 5 dpga_flat_0.sr_0._28_.RESET_B
rlabel metal1 175835 530418 175953 530427 5 dpga_flat_0.sr_0._28_.RESET_B
rlabel metal1 176483 530418 176613 530427 5 dpga_flat_0.sr_0._28_.RESET_B
rlabel metal1 175835 530427 176613 530455 5 dpga_flat_0.sr_0._28_.RESET_B
rlabel metal1 176483 530455 176613 530464 5 dpga_flat_0.sr_0._28_.RESET_B
rlabel metal1 175522 530563 177362 530659 5 dpga_flat_0.sr_0._28_.VGND
rlabel metal1 175522 530019 177362 530115 5 dpga_flat_0.sr_0._28_.VPWR
flabel locali 177298 529948 177332 529982 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._30_.Q
flabel locali 177298 529880 177332 529914 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._30_.Q
flabel locali 177298 529812 177332 529846 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._30_.Q
flabel locali 177298 529608 177332 529642 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._30_.Q
flabel locali 177003 529676 177037 529710 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._30_.RESET_B
flabel locali 175827 529812 175861 529846 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._30_.D
flabel locali 175552 529812 175586 529846 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._30_.CLK
flabel locali 175552 529744 175586 529778 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._30_.CLK
flabel locali 177003 529744 177037 529778 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._30_.RESET_B
flabel metal1 175551 529506 175585 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._30_.VGND
flabel metal1 175551 530050 175585 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._30_.VPWR
flabel nwell 175551 530050 175585 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._30_.VPB
flabel pwell 175551 529506 175585 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._30_.VNB
rlabel comment 175522 529523 175522 529523 4 dpga_flat_0.sr_0._30_.dfrtp_1
rlabel locali 177003 529650 177051 529730 1 dpga_flat_0.sr_0._30_.RESET_B
rlabel locali 176943 529730 177051 529804 1 dpga_flat_0.sr_0._30_.RESET_B
rlabel metal1 176991 529670 177049 529679 1 dpga_flat_0.sr_0._30_.RESET_B
rlabel metal1 176931 529716 176989 529779 1 dpga_flat_0.sr_0._30_.RESET_B
rlabel metal1 176931 529707 177049 529716 1 dpga_flat_0.sr_0._30_.RESET_B
rlabel metal1 176271 529707 176401 529716 1 dpga_flat_0.sr_0._30_.RESET_B
rlabel metal1 176271 529679 177049 529707 1 dpga_flat_0.sr_0._30_.RESET_B
rlabel metal1 176271 529670 176401 529679 1 dpga_flat_0.sr_0._30_.RESET_B
rlabel metal1 175522 529475 177362 529571 1 dpga_flat_0.sr_0._30_.VGND
rlabel metal1 175522 530019 177362 530115 1 dpga_flat_0.sr_0._30_.VPWR
flabel locali 174815 529744 174849 529778 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold1.A
flabel locali 175463 529676 175497 529710 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold1.X
flabel locali 174815 529812 174849 529846 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold1.A
flabel locali 175463 529608 175497 529642 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold1.X
flabel locali 174907 529744 174941 529778 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold1.A
flabel locali 174907 529812 174941 529846 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold1.A
flabel locali 175463 529948 175497 529982 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold1.X
flabel locali 175463 529812 175497 529846 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold1.X
flabel locali 175463 529880 175497 529914 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold1.X
flabel locali 175463 529744 175497 529778 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold1.X
flabel nwell 174815 530050 174849 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold1.VPB
flabel pwell 174815 529506 174849 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold1.VNB
flabel metal1 174815 529506 174849 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold1.VGND
flabel metal1 174815 530050 174849 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold1.VPWR
rlabel comment 174786 529523 174786 529523 4 dpga_flat_0.sr_0.hold1.dlygate4sd3_1
rlabel metal1 174786 529475 175522 529571 1 dpga_flat_0.sr_0.hold1.VGND
rlabel metal1 174786 530019 175522 530115 1 dpga_flat_0.sr_0.hold1.VPWR
flabel locali 174999 530288 175033 530322 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output5.X
flabel locali 175275 530424 175309 530458 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output5.A
flabel locali 174907 530424 174941 530458 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output5.X
flabel locali 175275 530356 175309 530390 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output5.A
flabel locali 174907 530356 174941 530390 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output5.X
flabel metal1 175367 530594 175401 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output5.VGND
flabel metal1 175367 530050 175401 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output5.VPWR
flabel nwell 175367 530050 175401 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output5.VPB
flabel pwell 175367 530594 175401 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output5.VNB
rlabel comment 175430 530611 175430 530611 8 dpga_flat_0.sr_0.output5.clkbuf_4
rlabel metal1 174878 530563 175430 530659 5 dpga_flat_0.sr_0.output5.VGND
rlabel metal1 174878 530019 175430 530115 5 dpga_flat_0.sr_0.output5.VPWR
flabel metal1 177474 530593 177527 530625 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_57.VGND
flabel metal1 177475 530050 177527 530081 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_57.VPWR
flabel nwell 177482 530058 177516 530076 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_57.VPB
flabel pwell 177485 530599 177517 530621 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_57.VNB
rlabel comment 177454 530611 177454 530611 2 dpga_flat_0.sr_0.FILLER_0_0_57.fill_2
rlabel metal1 177454 530563 177638 530659 5 dpga_flat_0.sr_0.FILLER_0_0_57.VGND
rlabel metal1 177454 530019 177638 530115 5 dpga_flat_0.sr_0.FILLER_0_0_57.VPWR
flabel metal1 177476 530050 177512 530080 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_57.VPWR
flabel metal1 177476 529510 177512 529539 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_57.VGND
flabel nwell 177485 530057 177505 530074 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_57.VPB
flabel pwell 177482 529512 177506 529534 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_57.VNB
rlabel comment 177454 529523 177454 529523 4 dpga_flat_0.sr_0.FILLER_0_1_57.fill_1
rlabel metal1 177454 529475 177546 529571 1 dpga_flat_0.sr_0.FILLER_0_1_57.VGND
rlabel metal1 177454 530019 177546 530115 1 dpga_flat_0.sr_0.FILLER_0_1_57.VPWR
flabel metal1 177384 530058 177437 530087 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_57.VPWR
flabel metal1 177383 530591 177434 530629 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_57.VGND
rlabel comment 177362 530611 177362 530611 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_57.tapvpwrvgnd_1
rlabel metal1 177362 530563 177454 530659 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_57.VGND
rlabel metal1 177362 530019 177454 530115 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_57.VPWR
flabel metal1 177384 530047 177437 530076 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_1_61.VPWR
flabel metal1 177383 529505 177434 529543 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_1_61.VGND
rlabel comment 177362 529523 177362 529523 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_1_61.tapvpwrvgnd_1
rlabel metal1 177362 529475 177454 529571 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_1_61.VGND
rlabel metal1 177362 530019 177454 530115 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_1_61.VPWR
flabel metal1 178310 529506 178344 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._18_.VGND
flabel metal1 178310 530050 178344 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._18_.VPWR
flabel locali 177666 529812 177700 529846 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._18_.S
flabel locali 177758 529812 177792 529846 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._18_.S
flabel locali 177850 529676 177884 529710 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._18_.A1
flabel locali 177850 529744 177884 529778 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._18_.A1
flabel locali 177942 529744 177976 529778 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._18_.A0
flabel locali 178310 529608 178344 529642 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._18_.X
flabel locali 178310 529880 178344 529914 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._18_.X
flabel locali 178310 529948 178344 529982 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._18_.X
flabel nwell 178266 530050 178300 530084 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._18_.VPB
flabel pwell 178256 529506 178290 529540 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._18_.VNB
rlabel comment 178374 529523 178374 529523 6 dpga_flat_0.sr_0._18_.mux2_1
rlabel metal1 177546 529475 178374 529571 1 dpga_flat_0.sr_0._18_.VGND
rlabel metal1 177546 530019 178374 530115 1 dpga_flat_0.sr_0._18_.VPWR
flabel locali 178311 530356 178345 530390 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold6.A
flabel locali 177663 530424 177697 530458 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold6.X
flabel locali 178311 530288 178345 530322 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold6.A
flabel locali 177663 530492 177697 530526 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold6.X
flabel locali 178219 530356 178253 530390 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold6.A
flabel locali 178219 530288 178253 530322 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold6.A
flabel locali 177663 530152 177697 530186 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold6.X
flabel locali 177663 530288 177697 530322 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold6.X
flabel locali 177663 530220 177697 530254 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold6.X
flabel locali 177663 530356 177697 530390 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold6.X
flabel nwell 178311 530050 178345 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold6.VPB
flabel pwell 178311 530594 178345 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold6.VNB
flabel metal1 178311 530594 178345 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold6.VGND
flabel metal1 178311 530050 178345 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold6.VPWR
rlabel comment 178374 530611 178374 530611 8 dpga_flat_0.sr_0.hold6.dlygate4sd3_1
rlabel metal1 177638 530563 178374 530659 5 dpga_flat_0.sr_0.hold6.VGND
rlabel metal1 177638 530019 178374 530115 5 dpga_flat_0.sr_0.hold6.VPWR
flabel metal1 179774 530593 179827 530625 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_82.VGND
flabel metal1 179775 530050 179827 530081 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_82.VPWR
flabel nwell 179782 530058 179816 530076 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_82.VPB
flabel pwell 179785 530599 179817 530621 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_82.VNB
rlabel comment 179754 530611 179754 530611 2 dpga_flat_0.sr_0.FILLER_0_0_82.fill_2
rlabel metal1 179754 530563 179938 530659 5 dpga_flat_0.sr_0.FILLER_0_0_82.VGND
rlabel metal1 179754 530019 179938 530115 5 dpga_flat_0.sr_0.FILLER_0_0_82.VPWR
flabel metal1 178587 530594 178621 530628 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._21_.VGND
flabel metal1 178587 530050 178621 530084 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._21_.VPWR
flabel locali 178403 530492 178437 530526 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._21_.X
flabel locali 178403 530220 178437 530254 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._21_.X
flabel locali 178403 530152 178437 530186 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._21_.X
flabel locali 178587 530356 178621 530390 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._21_.A
flabel nwell 178587 530050 178621 530084 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._21_.VPB
flabel pwell 178587 530594 178621 530628 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._21_.VNB
rlabel comment 178374 530611 178374 530611 2 dpga_flat_0.sr_0._21_.clkbuf_1
rlabel metal1 178374 530563 178650 530659 5 dpga_flat_0.sr_0._21_.VGND
rlabel metal1 178374 530019 178650 530115 5 dpga_flat_0.sr_0._21_.VPWR
flabel locali 178404 529948 178438 529982 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._32_.Q
flabel locali 178404 529880 178438 529914 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._32_.Q
flabel locali 178404 529812 178438 529846 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._32_.Q
flabel locali 178404 529608 178438 529642 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._32_.Q
flabel locali 178699 529676 178733 529710 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._32_.RESET_B
flabel locali 179875 529812 179909 529846 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._32_.D
flabel locali 180150 529812 180184 529846 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._32_.CLK
flabel locali 180150 529744 180184 529778 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._32_.CLK
flabel locali 178699 529744 178733 529778 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._32_.RESET_B
flabel metal1 180151 529506 180185 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._32_.VGND
flabel metal1 180151 530050 180185 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._32_.VPWR
flabel nwell 180151 530050 180185 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._32_.VPB
flabel pwell 180151 529506 180185 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._32_.VNB
rlabel comment 180214 529523 180214 529523 6 dpga_flat_0.sr_0._32_.dfrtp_1
rlabel locali 178685 529650 178733 529730 1 dpga_flat_0.sr_0._32_.RESET_B
rlabel locali 178685 529730 178793 529804 1 dpga_flat_0.sr_0._32_.RESET_B
rlabel metal1 178687 529670 178745 529679 1 dpga_flat_0.sr_0._32_.RESET_B
rlabel metal1 178747 529716 178805 529779 1 dpga_flat_0.sr_0._32_.RESET_B
rlabel metal1 178687 529707 178805 529716 1 dpga_flat_0.sr_0._32_.RESET_B
rlabel metal1 179335 529707 179465 529716 1 dpga_flat_0.sr_0._32_.RESET_B
rlabel metal1 178687 529679 179465 529707 1 dpga_flat_0.sr_0._32_.RESET_B
rlabel metal1 179335 529670 179465 529679 1 dpga_flat_0.sr_0._32_.RESET_B
rlabel metal1 178374 529475 180214 529571 1 dpga_flat_0.sr_0._32_.VGND
rlabel metal1 178374 530019 180214 530115 1 dpga_flat_0.sr_0._32_.VPWR
flabel locali 179599 530288 179633 530322 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output6.X
flabel locali 179323 530424 179357 530458 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output6.A
flabel locali 179691 530424 179725 530458 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output6.X
flabel locali 179323 530356 179357 530390 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output6.A
flabel locali 179691 530356 179725 530390 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output6.X
flabel metal1 179231 530594 179265 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output6.VGND
flabel metal1 179231 530050 179265 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output6.VPWR
flabel nwell 179231 530050 179265 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output6.VPB
flabel pwell 179231 530594 179265 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output6.VNB
rlabel comment 179202 530611 179202 530611 2 dpga_flat_0.sr_0.output6.clkbuf_4
rlabel metal1 179202 530563 179754 530659 5 dpga_flat_0.sr_0.output6.VGND
rlabel metal1 179202 530019 179754 530115 5 dpga_flat_0.sr_0.output6.VPWR
flabel locali 178771 530288 178805 530322 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output7.X
flabel locali 179047 530424 179081 530458 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output7.A
flabel locali 178679 530424 178713 530458 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output7.X
flabel locali 179047 530356 179081 530390 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output7.A
flabel locali 178679 530356 178713 530390 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output7.X
flabel metal1 179139 530594 179173 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output7.VGND
flabel metal1 179139 530050 179173 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output7.VPWR
flabel nwell 179139 530050 179173 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output7.VPB
flabel pwell 179139 530594 179173 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output7.VNB
rlabel comment 179202 530611 179202 530611 8 dpga_flat_0.sr_0.output7.clkbuf_4
rlabel metal1 178650 530563 179202 530659 5 dpga_flat_0.sr_0.output7.VGND
rlabel metal1 178650 530019 179202 530115 5 dpga_flat_0.sr_0.output7.VPWR
flabel metal1 180050 530593 180103 530625 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_85.VGND
flabel metal1 180051 530050 180103 530081 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_85.VPWR
flabel nwell 180058 530058 180092 530076 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_85.VPB
flabel pwell 180061 530599 180093 530621 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_85.VNB
rlabel comment 180030 530611 180030 530611 2 dpga_flat_0.sr_0.FILLER_0_0_85.fill_2
rlabel metal1 180030 530563 180214 530659 5 dpga_flat_0.sr_0.FILLER_0_0_85.VGND
rlabel metal1 180030 530019 180214 530115 5 dpga_flat_0.sr_0.FILLER_0_0_85.VPWR
flabel metal1 181064 530054 181100 530084 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_96.VPWR
flabel metal1 181064 530595 181100 530624 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_96.VGND
flabel nwell 181073 530060 181093 530077 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_96.VPB
flabel pwell 181070 530600 181094 530622 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_96.VNB
rlabel comment 181042 530611 181042 530611 2 dpga_flat_0.sr_0.FILLER_0_0_96.fill_1
rlabel metal1 181042 530563 181134 530659 5 dpga_flat_0.sr_0.FILLER_0_0_96.VGND
rlabel metal1 181042 530019 181134 530115 5 dpga_flat_0.sr_0.FILLER_0_0_96.VPWR
flabel metal1 179960 530058 180013 530087 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_58.VPWR
flabel metal1 179959 530591 180010 530629 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_58.VGND
rlabel comment 179938 530611 179938 530611 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_58.tapvpwrvgnd_1
rlabel metal1 179938 530563 180030 530659 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_58.VGND
rlabel metal1 179938 530019 180030 530115 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_58.VPWR
flabel metal1 180244 530594 180278 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._22_.VGND
flabel metal1 180244 530050 180278 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._22_.VPWR
flabel locali 180888 530288 180922 530322 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._22_.S
flabel locali 180796 530288 180830 530322 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._22_.S
flabel locali 180704 530424 180738 530458 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._22_.A1
flabel locali 180704 530356 180738 530390 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._22_.A1
flabel locali 180612 530356 180646 530390 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._22_.A0
flabel locali 180244 530492 180278 530526 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._22_.X
flabel locali 180244 530220 180278 530254 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._22_.X
flabel locali 180244 530152 180278 530186 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._22_.X
flabel nwell 180288 530050 180322 530084 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._22_.VPB
flabel pwell 180298 530594 180332 530628 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._22_.VNB
rlabel comment 180214 530611 180214 530611 2 dpga_flat_0.sr_0._22_.mux2_1
rlabel metal1 180214 530563 181042 530659 5 dpga_flat_0.sr_0._22_.VGND
rlabel metal1 180214 530019 181042 530115 5 dpga_flat_0.sr_0._22_.VPWR
flabel metal1 181898 530594 181932 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._24_.VGND
flabel metal1 181898 530050 181932 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._24_.VPWR
flabel locali 181254 530288 181288 530322 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._24_.S
flabel locali 181346 530288 181380 530322 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._24_.S
flabel locali 181438 530424 181472 530458 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._24_.A1
flabel locali 181438 530356 181472 530390 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._24_.A1
flabel locali 181530 530356 181564 530390 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._24_.A0
flabel locali 181898 530492 181932 530526 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._24_.X
flabel locali 181898 530220 181932 530254 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._24_.X
flabel locali 181898 530152 181932 530186 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._24_.X
flabel nwell 181854 530050 181888 530084 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._24_.VPB
flabel pwell 181844 530594 181878 530628 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._24_.VNB
rlabel comment 181962 530611 181962 530611 8 dpga_flat_0.sr_0._24_.mux2_1
rlabel metal1 181134 530563 181962 530659 5 dpga_flat_0.sr_0._24_.VGND
rlabel metal1 181134 530019 181962 530115 5 dpga_flat_0.sr_0._24_.VPWR
flabel locali 181990 529948 182024 529982 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._33_.Q
flabel locali 181990 529880 182024 529914 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._33_.Q
flabel locali 181990 529812 182024 529846 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._33_.Q
flabel locali 181990 529608 182024 529642 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._33_.Q
flabel locali 181695 529676 181729 529710 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._33_.RESET_B
flabel locali 180519 529812 180553 529846 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._33_.D
flabel locali 180244 529812 180278 529846 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._33_.CLK
flabel locali 180244 529744 180278 529778 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._33_.CLK
flabel locali 181695 529744 181729 529778 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._33_.RESET_B
flabel metal1 180243 529506 180277 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._33_.VGND
flabel metal1 180243 530050 180277 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._33_.VPWR
flabel nwell 180243 530050 180277 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._33_.VPB
flabel pwell 180243 529506 180277 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._33_.VNB
rlabel comment 180214 529523 180214 529523 4 dpga_flat_0.sr_0._33_.dfrtp_1
rlabel locali 181695 529650 181743 529730 1 dpga_flat_0.sr_0._33_.RESET_B
rlabel locali 181635 529730 181743 529804 1 dpga_flat_0.sr_0._33_.RESET_B
rlabel metal1 181683 529670 181741 529679 1 dpga_flat_0.sr_0._33_.RESET_B
rlabel metal1 181623 529716 181681 529779 1 dpga_flat_0.sr_0._33_.RESET_B
rlabel metal1 181623 529707 181741 529716 1 dpga_flat_0.sr_0._33_.RESET_B
rlabel metal1 180963 529707 181093 529716 1 dpga_flat_0.sr_0._33_.RESET_B
rlabel metal1 180963 529679 181741 529707 1 dpga_flat_0.sr_0._33_.RESET_B
rlabel metal1 180963 529670 181093 529679 1 dpga_flat_0.sr_0._33_.RESET_B
rlabel metal1 180214 529475 182054 529571 1 dpga_flat_0.sr_0._33_.VGND
rlabel metal1 180214 530019 182054 530115 1 dpga_flat_0.sr_0._33_.VPWR
flabel locali 182359 530288 182393 530322 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output8.X
flabel locali 182083 530424 182117 530458 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output8.A
flabel locali 182451 530424 182485 530458 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output8.X
flabel locali 182083 530356 182117 530390 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output8.A
flabel locali 182451 530356 182485 530390 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output8.X
flabel metal1 181991 530594 182025 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output8.VGND
flabel metal1 181991 530050 182025 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output8.VPWR
flabel nwell 181991 530050 182025 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output8.VPB
flabel pwell 181991 530594 182025 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output8.VNB
rlabel comment 181962 530611 181962 530611 2 dpga_flat_0.sr_0.output8.clkbuf_4
rlabel metal1 181962 530563 182514 530659 5 dpga_flat_0.sr_0.output8.VGND
rlabel metal1 181962 530019 182514 530115 5 dpga_flat_0.sr_0.output8.VPWR
flabel locali 183279 529744 183313 529778 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold5.A
flabel locali 182631 529676 182665 529710 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold5.X
flabel locali 183279 529812 183313 529846 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold5.A
flabel locali 182631 529608 182665 529642 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold5.X
flabel locali 183187 529744 183221 529778 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold5.A
flabel locali 183187 529812 183221 529846 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold5.A
flabel locali 182631 529948 182665 529982 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold5.X
flabel locali 182631 529812 182665 529846 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold5.X
flabel locali 182631 529880 182665 529914 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold5.X
flabel locali 182631 529744 182665 529778 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold5.X
flabel nwell 183279 530050 183313 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold5.VPB
flabel pwell 183279 529506 183313 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold5.VNB
flabel metal1 183279 529506 183313 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold5.VGND
flabel metal1 183279 530050 183313 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold5.VPWR
rlabel comment 183342 529523 183342 529523 6 dpga_flat_0.sr_0.hold5.dlygate4sd3_1
rlabel metal1 182606 529475 183342 529571 1 dpga_flat_0.sr_0.hold5.VGND
rlabel metal1 182606 530019 183342 530115 1 dpga_flat_0.sr_0.hold5.VPWR
flabel metal1 182536 530047 182589 530076 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_1_62.VPWR
flabel metal1 182535 529505 182586 529543 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_1_62.VGND
rlabel comment 182514 529523 182514 529523 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_1_62.tapvpwrvgnd_1
rlabel metal1 182514 529475 182606 529571 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_1_62.VGND
rlabel metal1 182514 530019 182606 530115 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_1_62.VPWR
flabel metal1 182536 530058 182589 530087 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_59.VPWR
flabel metal1 182535 530591 182586 530629 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_59.VGND
rlabel comment 182514 530611 182514 530611 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_59.tapvpwrvgnd_1
rlabel metal1 182514 530563 182606 530659 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_59.VGND
rlabel metal1 182514 530019 182606 530115 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_59.VPWR
flabel metal1 182444 530050 182480 530080 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_111.VPWR
flabel metal1 182444 529510 182480 529539 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_111.VGND
flabel nwell 182453 530057 182473 530074 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_111.VPB
flabel pwell 182450 529512 182474 529534 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_111.VNB
rlabel comment 182422 529523 182422 529523 4 dpga_flat_0.sr_0.FILLER_0_1_111.fill_1
rlabel metal1 182422 529475 182514 529571 1 dpga_flat_0.sr_0.FILLER_0_1_111.VGND
rlabel metal1 182422 530019 182514 530115 1 dpga_flat_0.sr_0.FILLER_0_1_111.VPWR
flabel metal1 182083 529506 182117 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_107.VGND
flabel metal1 182083 530050 182117 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_107.VPWR
flabel nwell 182083 530050 182117 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_107.VPB
flabel pwell 182083 529506 182117 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_107.VNB
rlabel comment 182054 529523 182054 529523 4 dpga_flat_0.sr_0.FILLER_0_1_107.decap_4
rlabel metal1 182054 529475 182422 529571 1 dpga_flat_0.sr_0.FILLER_0_1_107.VGND
rlabel metal1 182054 530019 182422 530115 1 dpga_flat_0.sr_0.FILLER_0_1_107.VPWR
flabel metal1 182635 530594 182669 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_113.VGND
flabel metal1 182635 530050 182669 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_113.VPWR
flabel nwell 182635 530050 182669 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_113.VPB
flabel pwell 182635 530594 182669 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_113.VNB
rlabel comment 182606 530611 182606 530611 2 dpga_flat_0.sr_0.FILLER_0_0_113.decap_4
rlabel metal1 182606 530563 182974 530659 5 dpga_flat_0.sr_0.FILLER_0_0_113.VGND
rlabel metal1 182606 530019 182974 530115 5 dpga_flat_0.sr_0.FILLER_0_0_113.VPWR
flabel locali 183463 530288 183497 530322 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output9.X
flabel locali 183187 530424 183221 530458 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output9.A
flabel locali 183555 530424 183589 530458 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output9.X
flabel locali 183187 530356 183221 530390 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output9.A
flabel locali 183555 530356 183589 530390 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output9.X
flabel metal1 183095 530594 183129 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output9.VGND
flabel metal1 183095 530050 183129 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output9.VPWR
flabel nwell 183095 530050 183129 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output9.VPB
flabel pwell 183095 530594 183129 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output9.VNB
rlabel comment 183066 530611 183066 530611 2 dpga_flat_0.sr_0.output9.clkbuf_4
rlabel metal1 183066 530563 183618 530659 5 dpga_flat_0.sr_0.output9.VGND
rlabel metal1 183066 530019 183618 530115 5 dpga_flat_0.sr_0.output9.VPWR
flabel metal1 182996 530054 183032 530084 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_117.VPWR
flabel metal1 182996 530595 183032 530624 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_117.VGND
flabel nwell 183005 530060 183025 530077 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_117.VPB
flabel pwell 183002 530600 183026 530622 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_117.VNB
rlabel comment 182974 530611 182974 530611 2 dpga_flat_0.sr_0.FILLER_0_0_117.fill_1
rlabel metal1 182974 530563 183066 530659 5 dpga_flat_0.sr_0.FILLER_0_0_117.VGND
rlabel metal1 182974 530019 183066 530115 5 dpga_flat_0.sr_0.FILLER_0_0_117.VPWR
flabel metal1 183371 529506 183405 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_121.VGND
flabel metal1 183371 530050 183405 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_121.VPWR
flabel nwell 183371 530050 183405 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_121.VPB
flabel pwell 183371 529506 183405 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_121.VNB
rlabel comment 183342 529523 183342 529523 4 dpga_flat_0.sr_0.FILLER_0_1_121.decap_12
flabel metal1 183647 530594 183681 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_124.VGND
flabel metal1 183647 530050 183681 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_124.VPWR
flabel nwell 183647 530050 183681 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_124.VPB
flabel pwell 183647 530594 183681 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_124.VNB
rlabel comment 183618 530611 183618 530611 2 dpga_flat_0.sr_0.FILLER_0_0_124.decap_12
flabel metal1 184751 530594 184785 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_136.VGND
flabel metal1 184751 530050 184785 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_136.VPWR
flabel nwell 184751 530050 184785 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_136.VPB
flabel pwell 184751 530594 184785 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_136.VNB
rlabel comment 184722 530611 184722 530611 2 dpga_flat_0.sr_0.FILLER_0_0_136.decap_4
rlabel metal1 184722 530563 185090 530659 5 dpga_flat_0.sr_0.FILLER_0_0_136.VGND
rlabel metal1 184722 530019 185090 530115 5 dpga_flat_0.sr_0.FILLER_0_0_136.VPWR
flabel metal1 184475 529506 184509 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_133.VGND
flabel metal1 184475 530050 184509 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_133.VPWR
flabel nwell 184475 530050 184509 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_133.VPB
flabel pwell 184475 529506 184509 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_133.VNB
rlabel comment 184446 529523 184446 529523 4 dpga_flat_0.sr_0.FILLER_0_1_133.decap_12
flabel metal1 185579 529506 185613 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_145.VGND
flabel metal1 185579 530050 185613 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_145.VPWR
flabel nwell 185579 530050 185613 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_145.VPB
flabel pwell 185579 529506 185613 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_145.VNB
rlabel comment 185550 529523 185550 529523 4 dpga_flat_0.sr_0.FILLER_0_1_145.decap_12
flabel metal1 185112 530058 185165 530087 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_60.VPWR
flabel metal1 185111 530591 185162 530629 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_60.VGND
rlabel comment 185090 530611 185090 530611 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_60.tapvpwrvgnd_1
rlabel metal1 185090 530563 185182 530659 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_60.VGND
rlabel metal1 185090 530019 185182 530115 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_0_60.VPWR
flabel locali 185579 530288 185613 530322 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output10.X
flabel locali 185303 530424 185337 530458 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output10.A
flabel locali 185671 530424 185705 530458 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output10.X
flabel locali 185303 530356 185337 530390 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output10.A
flabel locali 185671 530356 185705 530390 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output10.X
flabel metal1 185211 530594 185245 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output10.VGND
flabel metal1 185211 530050 185245 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output10.VPWR
flabel nwell 185211 530050 185245 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output10.VPB
flabel pwell 185211 530594 185245 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.output10.VNB
rlabel comment 185182 530611 185182 530611 2 dpga_flat_0.sr_0.output10.clkbuf_4
rlabel metal1 185182 530563 185734 530659 5 dpga_flat_0.sr_0.output10.VGND
rlabel metal1 185182 530019 185734 530115 5 dpga_flat_0.sr_0.output10.VPWR
flabel metal1 185763 530594 185797 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_147.VGND
flabel metal1 185763 530050 185797 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_147.VPWR
flabel nwell 185763 530050 185797 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_147.VPB
flabel pwell 185763 530594 185797 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_147.VNB
rlabel comment 185734 530611 185734 530611 2 dpga_flat_0.sr_0.FILLER_0_0_147.decap_12
flabel metal1 186860 530054 186896 530084 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_159.VPWR
flabel metal1 186860 530595 186896 530624 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_159.VGND
flabel nwell 186869 530060 186889 530077 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_159.VPB
flabel pwell 186866 530600 186890 530622 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_0_159.VNB
rlabel comment 186838 530611 186838 530611 2 dpga_flat_0.sr_0.FILLER_0_0_159.fill_1
rlabel metal1 186838 530563 186930 530659 5 dpga_flat_0.sr_0.FILLER_0_0_159.VGND
rlabel metal1 186838 530019 186930 530115 5 dpga_flat_0.sr_0.FILLER_0_0_159.VPWR
flabel metal1 186683 530050 186717 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_157.VPWR
flabel metal1 186683 529506 186717 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_157.VGND
flabel nwell 186683 530050 186717 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_157.VPB
flabel pwell 186683 529506 186717 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_1_157.VNB
rlabel comment 186654 529523 186654 529523 4 dpga_flat_0.sr_0.FILLER_0_1_157.decap_6
rlabel metal1 186654 529475 187206 529571 1 dpga_flat_0.sr_0.FILLER_0_1_157.VGND
rlabel metal1 186654 530019 187206 530115 1 dpga_flat_0.sr_0.FILLER_0_1_157.VPWR
flabel metal1 187419 530050 187453 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_0_Right_0.VPWR
flabel metal1 187419 530594 187453 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_0_Right_0.VGND
flabel nwell 187419 530050 187453 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_0_Right_0.VPB
flabel pwell 187419 530594 187453 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_0_Right_0.VNB
rlabel comment 187482 530611 187482 530611 8 dpga_flat_0.sr_0.PHY_EDGE_ROW_0_Right_0.decap_3
rlabel metal1 187206 530563 187482 530659 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_0_Right_0.VGND
rlabel metal1 187206 530019 187482 530115 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_0_Right_0.VPWR
flabel metal1 187419 530050 187453 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_1_Right_1.VPWR
flabel metal1 187419 529506 187453 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_1_Right_1.VGND
flabel nwell 187419 530050 187453 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_1_Right_1.VPB
flabel pwell 187419 529506 187453 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_1_Right_1.VNB
rlabel comment 187482 529523 187482 529523 6 dpga_flat_0.sr_0.PHY_EDGE_ROW_1_Right_1.decap_3
rlabel metal1 187206 529475 187482 529571 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_1_Right_1.VGND
rlabel metal1 187206 530019 187482 530115 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_1_Right_1.VPWR
flabel locali 187124 530288 187158 530322 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.sr_11.LO
flabel locali 186997 530352 187031 530386 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.sr_11.HI
flabel nwell 186959 530050 186993 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.sr_11.VPB
flabel pwell 186959 530594 186993 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.sr_11.VNB
flabel metal1 186959 530594 186993 530628 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.sr_11.VGND
flabel metal1 186959 530050 186993 530084 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.sr_11.VPWR
rlabel comment 186930 530611 186930 530611 2 dpga_flat_0.sr_0.sr_11.conb_1
flabel comment 186975 530338 186975 530338 0 FreeSans 200 90 0 0 dpga_flat_0.sr_0.sr_11.resistive_li1_ok
flabel comment 187163 530338 187163 530338 0 FreeSans 200 90 0 0 dpga_flat_0.sr_0.sr_11.resistive_li1_ok
flabel comment 187116 530353 187116 530353 0 FreeSans 200 90 0 0 dpga_flat_0.sr_0.sr_11.no_jumper_check
flabel comment 187013 530353 187013 530353 0 FreeSans 200 90 0 0 dpga_flat_0.sr_0.sr_11.no_jumper_check
rlabel metal1 186930 530563 187206 530659 5 dpga_flat_0.sr_0.sr_11.VGND
rlabel metal1 186930 530019 187206 530115 5 dpga_flat_0.sr_0.sr_11.VPWR
flabel metal1 172515 529506 172549 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_3.VGND
flabel metal1 172515 528962 172549 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_3.VPWR
flabel nwell 172515 528962 172549 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_3.VPB
flabel pwell 172515 529506 172549 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_3.VNB
rlabel comment 172486 529523 172486 529523 2 dpga_flat_0.sr_0.FILLER_0_2_3.decap_12
flabel metal1 173619 529506 173653 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_15.VGND
flabel metal1 173619 528962 173653 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_15.VPWR
flabel nwell 173619 528962 173653 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_15.VPB
flabel pwell 173619 529506 173653 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_15.VNB
rlabel comment 173590 529523 173590 529523 2 dpga_flat_0.sr_0.FILLER_0_2_15.decap_12
flabel metal1 172239 528962 172273 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_2_Left_30.VPWR
flabel metal1 172239 529506 172273 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_2_Left_30.VGND
flabel nwell 172239 528962 172273 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_2_Left_30.VPB
flabel pwell 172239 529506 172273 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_2_Left_30.VNB
rlabel comment 172210 529523 172210 529523 2 dpga_flat_0.sr_0.PHY_EDGE_ROW_2_Left_30.decap_3
rlabel metal1 172210 529475 172486 529571 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_2_Left_30.VGND
rlabel metal1 172210 528931 172486 529027 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_2_Left_30.VPWR
flabel metal1 174716 528966 174752 528996 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_27.VPWR
flabel metal1 174716 529507 174752 529536 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_27.VGND
flabel nwell 174725 528972 174745 528989 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_27.VPB
flabel pwell 174722 529512 174746 529534 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_27.VNB
rlabel comment 174694 529523 174694 529523 2 dpga_flat_0.sr_0.FILLER_0_2_27.fill_1
rlabel metal1 174694 529475 174786 529571 5 dpga_flat_0.sr_0.FILLER_0_2_27.VGND
rlabel metal1 174694 528931 174786 529027 5 dpga_flat_0.sr_0.FILLER_0_2_27.VPWR
flabel metal1 174898 529505 174951 529537 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_29.VGND
flabel metal1 174899 528962 174951 528993 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_29.VPWR
flabel nwell 174906 528970 174940 528988 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_29.VPB
flabel pwell 174909 529511 174941 529533 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_29.VNB
rlabel comment 174878 529523 174878 529523 2 dpga_flat_0.sr_0.FILLER_0_2_29.fill_2
rlabel metal1 174878 529475 175062 529571 5 dpga_flat_0.sr_0.FILLER_0_2_29.VGND
rlabel metal1 174878 528931 175062 529027 5 dpga_flat_0.sr_0.FILLER_0_2_29.VPWR
flabel metal1 174808 528970 174861 528999 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_2_63.VPWR
flabel metal1 174807 529503 174858 529541 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_2_63.VGND
rlabel comment 174786 529523 174786 529523 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_2_63.tapvpwrvgnd_1
rlabel metal1 174786 529475 174878 529571 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_2_63.VGND
rlabel metal1 174786 528931 174878 529027 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_2_63.VPWR
flabel metal1 175826 529506 175860 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._14_.VGND
flabel metal1 175826 528962 175860 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._14_.VPWR
flabel locali 175182 529200 175216 529234 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._14_.S
flabel locali 175274 529200 175308 529234 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._14_.S
flabel locali 175366 529336 175400 529370 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._14_.A1
flabel locali 175366 529268 175400 529302 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._14_.A1
flabel locali 175458 529268 175492 529302 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._14_.A0
flabel locali 175826 529404 175860 529438 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._14_.X
flabel locali 175826 529132 175860 529166 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._14_.X
flabel locali 175826 529064 175860 529098 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._14_.X
flabel nwell 175782 528962 175816 528996 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._14_.VPB
flabel pwell 175772 529506 175806 529540 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._14_.VNB
rlabel comment 175890 529523 175890 529523 8 dpga_flat_0.sr_0._14_.mux2_1
rlabel metal1 175062 529475 175890 529571 5 dpga_flat_0.sr_0._14_.VGND
rlabel metal1 175062 528931 175890 529027 5 dpga_flat_0.sr_0._14_.VPWR
flabel locali 176103 529200 176137 529234 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_0__f_sclk.X
flabel locali 176011 529200 176045 529234 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_0__f_sclk.X
flabel locali 176011 529268 176045 529302 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_0__f_sclk.X
flabel locali 176103 529268 176137 529302 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_0__f_sclk.X
flabel locali 176103 529336 176137 529370 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_0__f_sclk.X
flabel locali 176011 529336 176045 529370 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_0__f_sclk.X
flabel locali 177667 529336 177701 529370 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_0__f_sclk.A
flabel locali 177667 529268 177701 529302 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_0__f_sclk.A
flabel pwell 177667 529506 177701 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_0__f_sclk.VNB
flabel pwell 177684 529523 177684 529523 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_0__f_sclk.VNB
flabel nwell 177667 528962 177701 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_0__f_sclk.VPB
flabel nwell 177684 528979 177684 528979 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_0__f_sclk.VPB
flabel metal1 177667 529506 177701 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_0__f_sclk.VGND
flabel metal1 177667 528962 177701 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_0__f_sclk.VPWR
rlabel comment 177730 529523 177730 529523 8 dpga_flat_0.sr_0.clkbuf_1_0__f_sclk.clkbuf_16
rlabel metal1 175890 529475 177730 529571 5 dpga_flat_0.sr_0.clkbuf_1_0__f_sclk.VGND
rlabel metal1 175890 528931 177730 529027 5 dpga_flat_0.sr_0.clkbuf_1_0__f_sclk.VPWR
flabel locali 179506 529064 179540 529098 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._31_.Q
flabel locali 179506 529132 179540 529166 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._31_.Q
flabel locali 179506 529200 179540 529234 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._31_.Q
flabel locali 179506 529404 179540 529438 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._31_.Q
flabel locali 179211 529336 179245 529370 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._31_.RESET_B
flabel locali 178035 529200 178069 529234 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._31_.D
flabel locali 177760 529200 177794 529234 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._31_.CLK
flabel locali 177760 529268 177794 529302 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._31_.CLK
flabel locali 179211 529268 179245 529302 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._31_.RESET_B
flabel metal1 177759 529506 177793 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._31_.VGND
flabel metal1 177759 528962 177793 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._31_.VPWR
flabel nwell 177759 528962 177793 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._31_.VPB
flabel pwell 177759 529506 177793 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._31_.VNB
rlabel comment 177730 529523 177730 529523 2 dpga_flat_0.sr_0._31_.dfrtp_1
rlabel locali 179211 529316 179259 529396 5 dpga_flat_0.sr_0._31_.RESET_B
rlabel locali 179151 529242 179259 529316 5 dpga_flat_0.sr_0._31_.RESET_B
rlabel metal1 179199 529367 179257 529376 5 dpga_flat_0.sr_0._31_.RESET_B
rlabel metal1 179139 529267 179197 529330 5 dpga_flat_0.sr_0._31_.RESET_B
rlabel metal1 179139 529330 179257 529339 5 dpga_flat_0.sr_0._31_.RESET_B
rlabel metal1 178479 529330 178609 529339 5 dpga_flat_0.sr_0._31_.RESET_B
rlabel metal1 178479 529339 179257 529367 5 dpga_flat_0.sr_0._31_.RESET_B
rlabel metal1 178479 529367 178609 529376 5 dpga_flat_0.sr_0._31_.RESET_B
rlabel metal1 177730 529475 179570 529571 5 dpga_flat_0.sr_0._31_.VGND
rlabel metal1 177730 528931 179570 529027 5 dpga_flat_0.sr_0._31_.VPWR
flabel metal1 179592 528966 179628 528996 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_80.VPWR
flabel metal1 179592 529507 179628 529536 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_80.VGND
flabel nwell 179601 528972 179621 528989 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_80.VPB
flabel pwell 179598 529512 179622 529534 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_80.VNB
rlabel comment 179570 529523 179570 529523 2 dpga_flat_0.sr_0.FILLER_0_2_80.fill_1
rlabel metal1 179570 529475 179662 529571 5 dpga_flat_0.sr_0.FILLER_0_2_80.VGND
rlabel metal1 179570 528931 179662 529027 5 dpga_flat_0.sr_0.FILLER_0_2_80.VPWR
flabel metal1 179691 529506 179725 529540 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._23_.VGND
flabel metal1 179691 528962 179725 528996 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._23_.VPWR
flabel locali 179875 529404 179909 529438 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._23_.X
flabel locali 179875 529132 179909 529166 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._23_.X
flabel locali 179875 529064 179909 529098 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._23_.X
flabel locali 179691 529268 179725 529302 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._23_.A
flabel nwell 179691 528962 179725 528996 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._23_.VPB
flabel pwell 179691 529506 179725 529540 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._23_.VNB
rlabel comment 179938 529523 179938 529523 8 dpga_flat_0.sr_0._23_.clkbuf_1
rlabel metal1 179662 529475 179938 529571 5 dpga_flat_0.sr_0._23_.VGND
rlabel metal1 179662 528931 179938 529027 5 dpga_flat_0.sr_0._23_.VPWR
flabel metal1 180059 528962 180093 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_85.VPWR
flabel metal1 180059 529506 180093 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_85.VGND
flabel nwell 180059 528962 180093 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_85.VPB
flabel pwell 180059 529506 180093 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_85.VNB
rlabel comment 180030 529523 180030 529523 2 dpga_flat_0.sr_0.FILLER_0_2_85.decap_6
rlabel metal1 180030 529475 180582 529571 5 dpga_flat_0.sr_0.FILLER_0_2_85.VGND
rlabel metal1 180030 528931 180582 529027 5 dpga_flat_0.sr_0.FILLER_0_2_85.VPWR
flabel metal1 180604 528966 180640 528996 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_91.VPWR
flabel metal1 180604 529507 180640 529536 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_91.VGND
flabel nwell 180613 528972 180633 528989 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_91.VPB
flabel pwell 180610 529512 180634 529534 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_91.VNB
rlabel comment 180582 529523 180582 529523 2 dpga_flat_0.sr_0.FILLER_0_2_91.fill_1
rlabel metal1 180582 529475 180674 529571 5 dpga_flat_0.sr_0.FILLER_0_2_91.VGND
rlabel metal1 180582 528931 180674 529027 5 dpga_flat_0.sr_0.FILLER_0_2_91.VPWR
flabel metal1 179960 528970 180013 528999 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_2_64.VPWR
flabel metal1 179959 529503 180010 529541 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_2_64.VGND
rlabel comment 179938 529523 179938 529523 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_2_64.tapvpwrvgnd_1
rlabel metal1 179938 529475 180030 529571 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_2_64.VGND
rlabel metal1 179938 528931 180030 529027 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_2_64.VPWR
flabel locali 182267 529200 182301 529234 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_1__f_sclk.X
flabel locali 182359 529200 182393 529234 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_1__f_sclk.X
flabel locali 182359 529268 182393 529302 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_1__f_sclk.X
flabel locali 182267 529268 182301 529302 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_1__f_sclk.X
flabel locali 182267 529336 182301 529370 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_1__f_sclk.X
flabel locali 182359 529336 182393 529370 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_1__f_sclk.X
flabel locali 180703 529336 180737 529370 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_1__f_sclk.A
flabel locali 180703 529268 180737 529302 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_1__f_sclk.A
flabel pwell 180703 529506 180737 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_1__f_sclk.VNB
flabel pwell 180720 529523 180720 529523 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_1__f_sclk.VNB
flabel nwell 180703 528962 180737 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_1__f_sclk.VPB
flabel nwell 180720 528979 180720 528979 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_1__f_sclk.VPB
flabel metal1 180703 529506 180737 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_1__f_sclk.VGND
flabel metal1 180703 528962 180737 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_1_1__f_sclk.VPWR
rlabel comment 180674 529523 180674 529523 2 dpga_flat_0.sr_0.clkbuf_1_1__f_sclk.clkbuf_16
rlabel metal1 180674 529475 182514 529571 5 dpga_flat_0.sr_0.clkbuf_1_1__f_sclk.VGND
rlabel metal1 180674 528931 182514 529027 5 dpga_flat_0.sr_0.clkbuf_1_1__f_sclk.VPWR
flabel metal1 182819 529506 182853 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_115.VGND
flabel metal1 182819 528962 182853 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_115.VPWR
flabel nwell 182819 528962 182853 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_115.VPB
flabel pwell 182819 529506 182853 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_115.VNB
rlabel comment 182790 529523 182790 529523 2 dpga_flat_0.sr_0.FILLER_0_2_115.decap_12
flabel metal1 182727 529506 182761 529540 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._25_.VGND
flabel metal1 182727 528962 182761 528996 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._25_.VPWR
flabel locali 182543 529404 182577 529438 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._25_.X
flabel locali 182543 529132 182577 529166 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._25_.X
flabel locali 182543 529064 182577 529098 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._25_.X
flabel locali 182727 529268 182761 529302 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._25_.A
flabel nwell 182727 528962 182761 528996 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._25_.VPB
flabel pwell 182727 529506 182761 529540 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._25_.VNB
rlabel comment 182514 529523 182514 529523 2 dpga_flat_0.sr_0._25_.clkbuf_1
rlabel metal1 182514 529475 182790 529571 5 dpga_flat_0.sr_0._25_.VGND
rlabel metal1 182514 528931 182790 529027 5 dpga_flat_0.sr_0._25_.VPWR
flabel metal1 183923 529506 183957 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_127.VGND
flabel metal1 183923 528962 183957 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_127.VPWR
flabel nwell 183923 528962 183957 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_127.VPB
flabel pwell 183923 529506 183957 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_127.VNB
rlabel comment 183894 529523 183894 529523 2 dpga_flat_0.sr_0.FILLER_0_2_127.decap_12
flabel metal1 185020 528966 185056 528996 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_139.VPWR
flabel metal1 185020 529507 185056 529536 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_139.VGND
flabel nwell 185029 528972 185049 528989 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_139.VPB
flabel pwell 185026 529512 185050 529534 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_139.VNB
rlabel comment 184998 529523 184998 529523 2 dpga_flat_0.sr_0.FILLER_0_2_139.fill_1
rlabel metal1 184998 529475 185090 529571 5 dpga_flat_0.sr_0.FILLER_0_2_139.VGND
rlabel metal1 184998 528931 185090 529027 5 dpga_flat_0.sr_0.FILLER_0_2_139.VPWR
flabel metal1 185211 529506 185245 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_141.VGND
flabel metal1 185211 528962 185245 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_141.VPWR
flabel nwell 185211 528962 185245 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_141.VPB
flabel pwell 185211 529506 185245 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_141.VNB
rlabel comment 185182 529523 185182 529523 2 dpga_flat_0.sr_0.FILLER_0_2_141.decap_12
flabel metal1 185112 528970 185165 528999 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_2_65.VPWR
flabel metal1 185111 529503 185162 529541 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_2_65.VGND
rlabel comment 185090 529523 185090 529523 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_2_65.tapvpwrvgnd_1
rlabel metal1 185090 529475 185182 529571 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_2_65.VGND
rlabel metal1 185090 528931 185182 529027 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_2_65.VPWR
flabel metal1 186315 528962 186349 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_153.VPWR
flabel metal1 186315 529506 186349 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_153.VGND
flabel nwell 186315 528962 186349 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_153.VPB
flabel pwell 186315 529506 186349 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_153.VNB
rlabel comment 186286 529523 186286 529523 2 dpga_flat_0.sr_0.FILLER_0_2_153.decap_8
rlabel metal1 186286 529475 187022 529571 5 dpga_flat_0.sr_0.FILLER_0_2_153.VGND
rlabel metal1 186286 528931 187022 529027 5 dpga_flat_0.sr_0.FILLER_0_2_153.VPWR
flabel metal1 187042 529505 187095 529537 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_161.VGND
flabel metal1 187043 528962 187095 528993 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_161.VPWR
flabel nwell 187050 528970 187084 528988 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_161.VPB
flabel pwell 187053 529511 187085 529533 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_2_161.VNB
rlabel comment 187022 529523 187022 529523 2 dpga_flat_0.sr_0.FILLER_0_2_161.fill_2
rlabel metal1 187022 529475 187206 529571 5 dpga_flat_0.sr_0.FILLER_0_2_161.VGND
rlabel metal1 187022 528931 187206 529027 5 dpga_flat_0.sr_0.FILLER_0_2_161.VPWR
flabel metal1 187419 528962 187453 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_2_Right_2.VPWR
flabel metal1 187419 529506 187453 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_2_Right_2.VGND
flabel nwell 187419 528962 187453 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_2_Right_2.VPB
flabel pwell 187419 529506 187453 529540 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_2_Right_2.VNB
rlabel comment 187482 529523 187482 529523 8 dpga_flat_0.sr_0.PHY_EDGE_ROW_2_Right_2.decap_3
rlabel metal1 187206 529475 187482 529571 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_2_Right_2.VGND
rlabel metal1 187206 528931 187482 529027 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_2_Right_2.VPWR
flabel metal1 172515 528418 172549 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_3.VGND
flabel metal1 172515 528962 172549 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_3.VPWR
flabel nwell 172515 528962 172549 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_3.VPB
flabel pwell 172515 528418 172549 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_3.VNB
rlabel comment 172486 528435 172486 528435 4 dpga_flat_0.sr_0.FILLER_0_3_3.decap_12
flabel metal1 173619 528418 173653 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_15.VGND
flabel metal1 173619 528962 173653 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_15.VPWR
flabel nwell 173619 528962 173653 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_15.VPB
flabel pwell 173619 528418 173653 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_15.VNB
rlabel comment 173590 528435 173590 528435 4 dpga_flat_0.sr_0.FILLER_0_3_15.decap_12
flabel metal1 172239 528962 172273 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_3_Left_31.VPWR
flabel metal1 172239 528418 172273 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_3_Left_31.VGND
flabel nwell 172239 528962 172273 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_3_Left_31.VPB
flabel pwell 172239 528418 172273 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_3_Left_31.VNB
rlabel comment 172210 528435 172210 528435 4 dpga_flat_0.sr_0.PHY_EDGE_ROW_3_Left_31.decap_3
rlabel metal1 172210 528387 172486 528483 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_3_Left_31.VGND
rlabel metal1 172210 528931 172486 529027 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_3_Left_31.VPWR
flabel metal1 174723 528418 174757 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_27.VGND
flabel metal1 174723 528962 174757 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_27.VPWR
flabel nwell 174723 528962 174757 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_27.VPB
flabel pwell 174723 528418 174757 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_27.VNB
rlabel comment 174694 528435 174694 528435 4 dpga_flat_0.sr_0.FILLER_0_3_27.decap_12
flabel metal1 175820 528962 175856 528992 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_39.VPWR
flabel metal1 175820 528422 175856 528451 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_39.VGND
flabel nwell 175829 528969 175849 528986 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_39.VPB
flabel pwell 175826 528424 175850 528446 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_39.VNB
rlabel comment 175798 528435 175798 528435 4 dpga_flat_0.sr_0.FILLER_0_3_39.fill_1
rlabel metal1 175798 528387 175890 528483 1 dpga_flat_0.sr_0.FILLER_0_3_39.VGND
rlabel metal1 175798 528931 175890 529027 1 dpga_flat_0.sr_0.FILLER_0_3_39.VPWR
flabel metal1 175919 528418 175953 528452 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._15_.VGND
flabel metal1 175919 528962 175953 528996 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._15_.VPWR
flabel locali 176103 528520 176137 528554 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._15_.X
flabel locali 176103 528792 176137 528826 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._15_.X
flabel locali 176103 528860 176137 528894 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._15_.X
flabel locali 175919 528656 175953 528690 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._15_.A
flabel nwell 175919 528962 175953 528996 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._15_.VPB
flabel pwell 175919 528418 175953 528452 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._15_.VNB
rlabel comment 176166 528435 176166 528435 6 dpga_flat_0.sr_0._15_.clkbuf_1
rlabel metal1 175890 528387 176166 528483 1 dpga_flat_0.sr_0._15_.VGND
rlabel metal1 175890 528931 176166 529027 1 dpga_flat_0.sr_0._15_.VPWR
flabel metal1 177292 528962 177328 528992 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_55.VPWR
flabel metal1 177292 528422 177328 528451 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_55.VGND
flabel nwell 177301 528969 177321 528986 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_55.VPB
flabel pwell 177298 528424 177322 528446 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_55.VNB
rlabel comment 177270 528435 177270 528435 4 dpga_flat_0.sr_0.FILLER_0_3_55.fill_1
rlabel metal1 177270 528387 177362 528483 1 dpga_flat_0.sr_0.FILLER_0_3_55.VGND
rlabel metal1 177270 528931 177362 529027 1 dpga_flat_0.sr_0.FILLER_0_3_55.VPWR
flabel metal1 177384 528959 177437 528988 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_3_66.VPWR
flabel metal1 177383 528417 177434 528455 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_3_66.VGND
rlabel comment 177362 528435 177362 528435 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_3_66.tapvpwrvgnd_1
rlabel metal1 177362 528387 177454 528483 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_3_66.VGND
rlabel metal1 177362 528931 177454 529027 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_3_66.VPWR
flabel metal1 177206 528418 177240 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._16_.VGND
flabel metal1 177206 528962 177240 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._16_.VPWR
flabel locali 176562 528724 176596 528758 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._16_.S
flabel locali 176654 528724 176688 528758 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._16_.S
flabel locali 176746 528588 176780 528622 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._16_.A1
flabel locali 176746 528656 176780 528690 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._16_.A1
flabel locali 176838 528656 176872 528690 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._16_.A0
flabel locali 177206 528520 177240 528554 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._16_.X
flabel locali 177206 528792 177240 528826 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._16_.X
flabel locali 177206 528860 177240 528894 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._16_.X
flabel nwell 177162 528962 177196 528996 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._16_.VPB
flabel pwell 177152 528418 177186 528452 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._16_.VNB
rlabel comment 177270 528435 177270 528435 6 dpga_flat_0.sr_0._16_.mux2_1
rlabel metal1 176442 528387 177270 528483 1 dpga_flat_0.sr_0._16_.VGND
rlabel metal1 176442 528931 177270 529027 1 dpga_flat_0.sr_0._16_.VPWR
flabel metal1 176195 528418 176229 528452 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._17_.VGND
flabel metal1 176195 528962 176229 528996 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._17_.VPWR
flabel locali 176379 528520 176413 528554 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._17_.X
flabel locali 176379 528792 176413 528826 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._17_.X
flabel locali 176379 528860 176413 528894 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._17_.X
flabel locali 176195 528656 176229 528690 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._17_.A
flabel nwell 176195 528962 176229 528996 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._17_.VPB
flabel pwell 176195 528418 176229 528452 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._17_.VNB
rlabel comment 176442 528435 176442 528435 6 dpga_flat_0.sr_0._17_.clkbuf_1
rlabel metal1 176166 528387 176442 528483 1 dpga_flat_0.sr_0._17_.VGND
rlabel metal1 176166 528931 176442 529027 1 dpga_flat_0.sr_0._17_.VPWR
flabel locali 178127 528656 178161 528690 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold2.A
flabel locali 177479 528588 177513 528622 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold2.X
flabel locali 178127 528724 178161 528758 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold2.A
flabel locali 177479 528520 177513 528554 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold2.X
flabel locali 178035 528656 178069 528690 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold2.A
flabel locali 178035 528724 178069 528758 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold2.A
flabel locali 177479 528860 177513 528894 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold2.X
flabel locali 177479 528724 177513 528758 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold2.X
flabel locali 177479 528792 177513 528826 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold2.X
flabel locali 177479 528656 177513 528690 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold2.X
flabel nwell 178127 528962 178161 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold2.VPB
flabel pwell 178127 528418 178161 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold2.VNB
flabel metal1 178127 528418 178161 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold2.VGND
flabel metal1 178127 528962 178161 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold2.VPWR
rlabel comment 178190 528435 178190 528435 6 dpga_flat_0.sr_0.hold2.dlygate4sd3_1
rlabel metal1 177454 528387 178190 528483 1 dpga_flat_0.sr_0.hold2.VGND
rlabel metal1 177454 528931 178190 529027 1 dpga_flat_0.sr_0.hold2.VPWR
flabel metal1 178210 528421 178263 528453 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_65.VGND
flabel metal1 178211 528965 178263 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_65.VPWR
flabel nwell 178218 528970 178252 528988 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_65.VPB
flabel pwell 178221 528425 178253 528447 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_65.VNB
rlabel comment 178190 528435 178190 528435 4 dpga_flat_0.sr_0.FILLER_0_3_65.fill_2
rlabel metal1 178190 528387 178374 528483 1 dpga_flat_0.sr_0.FILLER_0_3_65.VGND
rlabel metal1 178190 528931 178374 529027 1 dpga_flat_0.sr_0.FILLER_0_3_65.VPWR
flabel locali 179967 528724 180001 528758 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_0_sclk.X
flabel locali 180059 528724 180093 528758 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_0_sclk.X
flabel locali 180059 528656 180093 528690 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_0_sclk.X
flabel locali 179967 528656 180001 528690 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_0_sclk.X
flabel locali 179967 528588 180001 528622 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_0_sclk.X
flabel locali 180059 528588 180093 528622 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_0_sclk.X
flabel locali 178403 528588 178437 528622 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_0_sclk.A
flabel locali 178403 528656 178437 528690 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_0_sclk.A
flabel pwell 178403 528418 178437 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_0_sclk.VNB
flabel pwell 178420 528435 178420 528435 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_0_sclk.VNB
flabel nwell 178403 528962 178437 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_0_sclk.VPB
flabel nwell 178420 528979 178420 528979 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_0_sclk.VPB
flabel metal1 178403 528418 178437 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_0_sclk.VGND
flabel metal1 178403 528962 178437 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.clkbuf_0_sclk.VPWR
rlabel comment 178374 528435 178374 528435 4 dpga_flat_0.sr_0.clkbuf_0_sclk.clkbuf_16
rlabel metal1 178374 528387 180214 528483 1 dpga_flat_0.sr_0.clkbuf_0_sclk.VGND
rlabel metal1 178374 528931 180214 529027 1 dpga_flat_0.sr_0.clkbuf_0_sclk.VPWR
flabel metal1 180243 528418 180277 528452 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._27_.VGND
flabel metal1 180243 528962 180277 528996 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._27_.VPWR
flabel locali 180427 528520 180461 528554 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._27_.X
flabel locali 180427 528792 180461 528826 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._27_.X
flabel locali 180427 528860 180461 528894 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._27_.X
flabel locali 180243 528656 180277 528690 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._27_.A
flabel nwell 180243 528962 180277 528996 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._27_.VPB
flabel pwell 180243 528418 180277 528452 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._27_.VNB
rlabel comment 180490 528435 180490 528435 6 dpga_flat_0.sr_0._27_.clkbuf_1
rlabel metal1 180214 528387 180490 528483 1 dpga_flat_0.sr_0._27_.VGND
rlabel metal1 180214 528931 180490 529027 1 dpga_flat_0.sr_0._27_.VPWR
flabel locali 182266 528860 182300 528894 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._34_.Q
flabel locali 182266 528792 182300 528826 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._34_.Q
flabel locali 182266 528724 182300 528758 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._34_.Q
flabel locali 182266 528520 182300 528554 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._34_.Q
flabel locali 181971 528588 182005 528622 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._34_.RESET_B
flabel locali 180795 528724 180829 528758 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._34_.D
flabel locali 180520 528724 180554 528758 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._34_.CLK
flabel locali 180520 528656 180554 528690 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._34_.CLK
flabel locali 181971 528656 182005 528690 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._34_.RESET_B
flabel metal1 180519 528418 180553 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._34_.VGND
flabel metal1 180519 528962 180553 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._34_.VPWR
flabel nwell 180519 528962 180553 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._34_.VPB
flabel pwell 180519 528418 180553 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._34_.VNB
rlabel comment 180490 528435 180490 528435 4 dpga_flat_0.sr_0._34_.dfrtp_1
rlabel locali 181971 528562 182019 528642 1 dpga_flat_0.sr_0._34_.RESET_B
rlabel locali 181911 528642 182019 528716 1 dpga_flat_0.sr_0._34_.RESET_B
rlabel metal1 181959 528582 182017 528591 1 dpga_flat_0.sr_0._34_.RESET_B
rlabel metal1 181899 528628 181957 528691 1 dpga_flat_0.sr_0._34_.RESET_B
rlabel metal1 181899 528619 182017 528628 1 dpga_flat_0.sr_0._34_.RESET_B
rlabel metal1 181239 528619 181369 528628 1 dpga_flat_0.sr_0._34_.RESET_B
rlabel metal1 181239 528591 182017 528619 1 dpga_flat_0.sr_0._34_.RESET_B
rlabel metal1 181239 528582 181369 528591 1 dpga_flat_0.sr_0._34_.RESET_B
rlabel metal1 180490 528387 182330 528483 1 dpga_flat_0.sr_0._34_.VGND
rlabel metal1 180490 528931 182330 529027 1 dpga_flat_0.sr_0._34_.VPWR
flabel metal1 182350 528421 182403 528453 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_110.VGND
flabel metal1 182351 528965 182403 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_110.VPWR
flabel nwell 182358 528970 182392 528988 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_110.VPB
flabel pwell 182361 528425 182393 528447 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_110.VNB
rlabel comment 182330 528435 182330 528435 4 dpga_flat_0.sr_0.FILLER_0_3_110.fill_2
rlabel metal1 182330 528387 182514 528483 1 dpga_flat_0.sr_0.FILLER_0_3_110.VGND
rlabel metal1 182330 528931 182514 529027 1 dpga_flat_0.sr_0.FILLER_0_3_110.VPWR
flabel metal1 182635 528418 182669 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_113.VGND
flabel metal1 182635 528962 182669 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_113.VPWR
flabel nwell 182635 528962 182669 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_113.VPB
flabel pwell 182635 528418 182669 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_113.VNB
rlabel comment 182606 528435 182606 528435 4 dpga_flat_0.sr_0.FILLER_0_3_113.decap_12
flabel metal1 183739 528418 183773 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_125.VGND
flabel metal1 183739 528962 183773 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_125.VPWR
flabel nwell 183739 528962 183773 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_125.VPB
flabel pwell 183739 528418 183773 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_125.VNB
rlabel comment 183710 528435 183710 528435 4 dpga_flat_0.sr_0.FILLER_0_3_125.decap_12
flabel metal1 182536 528959 182589 528988 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_3_67.VPWR
flabel metal1 182535 528417 182586 528455 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_3_67.VGND
rlabel comment 182514 528435 182514 528435 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_3_67.tapvpwrvgnd_1
rlabel metal1 182514 528387 182606 528483 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_3_67.VGND
rlabel metal1 182514 528931 182606 529027 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_3_67.VPWR
flabel metal1 184843 528418 184877 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_137.VGND
flabel metal1 184843 528962 184877 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_137.VPWR
flabel nwell 184843 528962 184877 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_137.VPB
flabel pwell 184843 528418 184877 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_137.VNB
rlabel comment 184814 528435 184814 528435 4 dpga_flat_0.sr_0.FILLER_0_3_137.decap_12
flabel metal1 185947 528418 185981 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_149.VGND
flabel metal1 185947 528962 185981 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_149.VPWR
flabel nwell 185947 528962 185981 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_149.VPB
flabel pwell 185947 528418 185981 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_149.VNB
rlabel comment 185918 528435 185918 528435 4 dpga_flat_0.sr_0.FILLER_0_3_149.decap_12
flabel metal1 187042 528421 187095 528453 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_161.VGND
flabel metal1 187043 528965 187095 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_161.VPWR
flabel nwell 187050 528970 187084 528988 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_161.VPB
flabel pwell 187053 528425 187085 528447 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_3_161.VNB
rlabel comment 187022 528435 187022 528435 4 dpga_flat_0.sr_0.FILLER_0_3_161.fill_2
rlabel metal1 187022 528387 187206 528483 1 dpga_flat_0.sr_0.FILLER_0_3_161.VGND
rlabel metal1 187022 528931 187206 529027 1 dpga_flat_0.sr_0.FILLER_0_3_161.VPWR
flabel metal1 187419 528962 187453 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_3_Right_3.VPWR
flabel metal1 187419 528418 187453 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_3_Right_3.VGND
flabel nwell 187419 528962 187453 528996 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_3_Right_3.VPB
flabel pwell 187419 528418 187453 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_3_Right_3.VNB
rlabel comment 187482 528435 187482 528435 6 dpga_flat_0.sr_0.PHY_EDGE_ROW_3_Right_3.decap_3
rlabel metal1 187206 528387 187482 528483 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_3_Right_3.VGND
rlabel metal1 187206 528931 187482 529027 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_3_Right_3.VPWR
flabel metal1 172515 528418 172549 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_3.VGND
flabel metal1 172515 527874 172549 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_3.VPWR
flabel nwell 172515 527874 172549 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_3.VPB
flabel pwell 172515 528418 172549 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_3.VNB
rlabel comment 172486 528435 172486 528435 2 dpga_flat_0.sr_0.FILLER_0_4_3.decap_12
flabel metal1 173619 528418 173653 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_15.VGND
flabel metal1 173619 527874 173653 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_15.VPWR
flabel nwell 173619 527874 173653 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_15.VPB
flabel pwell 173619 528418 173653 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_15.VNB
rlabel comment 173590 528435 173590 528435 2 dpga_flat_0.sr_0.FILLER_0_4_15.decap_12
flabel metal1 172239 527874 172273 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_4_Left_32.VPWR
flabel metal1 172239 528418 172273 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_4_Left_32.VGND
flabel nwell 172239 527874 172273 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_4_Left_32.VPB
flabel pwell 172239 528418 172273 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_4_Left_32.VNB
rlabel comment 172210 528435 172210 528435 2 dpga_flat_0.sr_0.PHY_EDGE_ROW_4_Left_32.decap_3
rlabel metal1 172210 528387 172486 528483 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_4_Left_32.VGND
rlabel metal1 172210 527843 172486 527939 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_4_Left_32.VPWR
flabel metal1 174716 527878 174752 527908 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_27.VPWR
flabel metal1 174716 528419 174752 528448 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_27.VGND
flabel nwell 174725 527884 174745 527901 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_27.VPB
flabel pwell 174722 528424 174746 528446 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_27.VNB
rlabel comment 174694 528435 174694 528435 2 dpga_flat_0.sr_0.FILLER_0_4_27.fill_1
rlabel metal1 174694 528387 174786 528483 5 dpga_flat_0.sr_0.FILLER_0_4_27.VGND
rlabel metal1 174694 527843 174786 527939 5 dpga_flat_0.sr_0.FILLER_0_4_27.VPWR
flabel metal1 174907 528418 174941 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_29.VGND
flabel metal1 174907 527874 174941 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_29.VPWR
flabel nwell 174907 527874 174941 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_29.VPB
flabel pwell 174907 528418 174941 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_29.VNB
rlabel comment 174878 528435 174878 528435 2 dpga_flat_0.sr_0.FILLER_0_4_29.decap_12
flabel metal1 176004 527878 176040 527908 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_41.VPWR
flabel metal1 176004 528419 176040 528448 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_41.VGND
flabel nwell 176013 527884 176033 527901 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_41.VPB
flabel pwell 176010 528424 176034 528446 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_41.VNB
rlabel comment 175982 528435 175982 528435 2 dpga_flat_0.sr_0.FILLER_0_4_41.fill_1
rlabel metal1 175982 528387 176074 528483 5 dpga_flat_0.sr_0.FILLER_0_4_41.VGND
rlabel metal1 175982 527843 176074 527939 5 dpga_flat_0.sr_0.FILLER_0_4_41.VPWR
flabel metal1 174808 527882 174861 527911 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_4_68.VPWR
flabel metal1 174807 528415 174858 528453 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_4_68.VGND
rlabel comment 174786 528435 174786 528435 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_4_68.tapvpwrvgnd_1
rlabel metal1 174786 528387 174878 528483 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_4_68.VGND
rlabel metal1 174786 527843 174878 527939 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_4_68.VPWR
flabel metal1 178127 528418 178161 528452 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._19_.VGND
flabel metal1 178127 527874 178161 527908 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._19_.VPWR
flabel locali 177943 528316 177977 528350 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._19_.X
flabel locali 177943 528044 177977 528078 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._19_.X
flabel locali 177943 527976 177977 528010 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._19_.X
flabel locali 178127 528180 178161 528214 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._19_.A
flabel nwell 178127 527874 178161 527908 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._19_.VPB
flabel pwell 178127 528418 178161 528452 0 FreeSans 200 180 0 0 dpga_flat_0.sr_0._19_.VNB
rlabel comment 177914 528435 177914 528435 2 dpga_flat_0.sr_0._19_.clkbuf_1
rlabel metal1 177914 528387 178190 528483 5 dpga_flat_0.sr_0._19_.VGND
rlabel metal1 177914 527843 178190 527939 5 dpga_flat_0.sr_0._19_.VPWR
flabel locali 177850 527976 177884 528010 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._29_.Q
flabel locali 177850 528044 177884 528078 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._29_.Q
flabel locali 177850 528112 177884 528146 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._29_.Q
flabel locali 177850 528316 177884 528350 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._29_.Q
flabel locali 177555 528248 177589 528282 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._29_.RESET_B
flabel locali 176379 528112 176413 528146 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._29_.D
flabel locali 176104 528112 176138 528146 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._29_.CLK
flabel locali 176104 528180 176138 528214 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._29_.CLK
flabel locali 177555 528180 177589 528214 0 FreeSans 400 0 0 0 dpga_flat_0.sr_0._29_.RESET_B
flabel metal1 176103 528418 176137 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._29_.VGND
flabel metal1 176103 527874 176137 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._29_.VPWR
flabel nwell 176103 527874 176137 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._29_.VPB
flabel pwell 176103 528418 176137 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._29_.VNB
rlabel comment 176074 528435 176074 528435 2 dpga_flat_0.sr_0._29_.dfrtp_1
rlabel locali 177555 528228 177603 528308 5 dpga_flat_0.sr_0._29_.RESET_B
rlabel locali 177495 528154 177603 528228 5 dpga_flat_0.sr_0._29_.RESET_B
rlabel metal1 177543 528279 177601 528288 5 dpga_flat_0.sr_0._29_.RESET_B
rlabel metal1 177483 528179 177541 528242 5 dpga_flat_0.sr_0._29_.RESET_B
rlabel metal1 177483 528242 177601 528251 5 dpga_flat_0.sr_0._29_.RESET_B
rlabel metal1 176823 528242 176953 528251 5 dpga_flat_0.sr_0._29_.RESET_B
rlabel metal1 176823 528251 177601 528279 5 dpga_flat_0.sr_0._29_.RESET_B
rlabel metal1 176823 528279 176953 528288 5 dpga_flat_0.sr_0._29_.RESET_B
rlabel metal1 176074 528387 177914 528483 5 dpga_flat_0.sr_0._29_.VGND
rlabel metal1 176074 527843 177914 527939 5 dpga_flat_0.sr_0._29_.VPWR
flabel metal1 178219 527874 178253 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_65.VPWR
flabel metal1 178219 528418 178253 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_65.VGND
flabel nwell 178219 527874 178253 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_65.VPB
flabel pwell 178219 528418 178253 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_65.VNB
rlabel comment 178190 528435 178190 528435 2 dpga_flat_0.sr_0.FILLER_0_4_65.decap_8
rlabel metal1 178190 528387 178926 528483 5 dpga_flat_0.sr_0.FILLER_0_4_65.VGND
rlabel metal1 178190 527843 178926 527939 5 dpga_flat_0.sr_0.FILLER_0_4_65.VPWR
flabel metal1 179774 528417 179827 528449 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_82.VGND
flabel metal1 179775 527874 179827 527905 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_82.VPWR
flabel nwell 179782 527882 179816 527900 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_82.VPB
flabel pwell 179785 528423 179817 528445 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_82.VNB
rlabel comment 179754 528435 179754 528435 2 dpga_flat_0.sr_0.FILLER_0_4_82.fill_2
rlabel metal1 179754 528387 179938 528483 5 dpga_flat_0.sr_0.FILLER_0_4_82.VGND
rlabel metal1 179754 527843 179938 527939 5 dpga_flat_0.sr_0.FILLER_0_4_82.VPWR
flabel metal1 178956 528418 178990 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._20_.VGND
flabel metal1 178956 527874 178990 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._20_.VPWR
flabel locali 179600 528112 179634 528146 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._20_.S
flabel locali 179508 528112 179542 528146 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._20_.S
flabel locali 179416 528248 179450 528282 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._20_.A1
flabel locali 179416 528180 179450 528214 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._20_.A1
flabel locali 179324 528180 179358 528214 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._20_.A0
flabel locali 178956 528316 178990 528350 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._20_.X
flabel locali 178956 528044 178990 528078 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._20_.X
flabel locali 178956 527976 178990 528010 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._20_.X
flabel nwell 179000 527874 179034 527908 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._20_.VPB
flabel pwell 179010 528418 179044 528452 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._20_.VNB
rlabel comment 178926 528435 178926 528435 2 dpga_flat_0.sr_0._20_.mux2_1
rlabel metal1 178926 528387 179754 528483 5 dpga_flat_0.sr_0._20_.VGND
rlabel metal1 178926 527843 179754 527939 5 dpga_flat_0.sr_0._20_.VPWR
flabel metal1 180059 527874 180093 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_85.VPWR
flabel metal1 180059 528418 180093 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_85.VGND
flabel nwell 180059 527874 180093 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_85.VPB
flabel pwell 180059 528418 180093 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_85.VNB
rlabel comment 180030 528435 180030 528435 2 dpga_flat_0.sr_0.FILLER_0_4_85.decap_8
rlabel metal1 180030 528387 180766 528483 5 dpga_flat_0.sr_0.FILLER_0_4_85.VGND
rlabel metal1 180030 527843 180766 527939 5 dpga_flat_0.sr_0.FILLER_0_4_85.VPWR
flabel metal1 180786 528417 180839 528449 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_93.VGND
flabel metal1 180787 527874 180839 527905 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_93.VPWR
flabel nwell 180794 527882 180828 527900 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_93.VPB
flabel pwell 180797 528423 180829 528445 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_93.VNB
rlabel comment 180766 528435 180766 528435 2 dpga_flat_0.sr_0.FILLER_0_4_93.fill_2
rlabel metal1 180766 528387 180950 528483 5 dpga_flat_0.sr_0.FILLER_0_4_93.VGND
rlabel metal1 180766 527843 180950 527939 5 dpga_flat_0.sr_0.FILLER_0_4_93.VPWR
flabel metal1 181807 528418 181841 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_104.VGND
flabel metal1 181807 527874 181841 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_104.VPWR
flabel nwell 181807 527874 181841 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_104.VPB
flabel pwell 181807 528418 181841 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_104.VNB
rlabel comment 181778 528435 181778 528435 2 dpga_flat_0.sr_0.FILLER_0_4_104.decap_12
flabel metal1 179960 527882 180013 527911 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_4_69.VPWR
flabel metal1 179959 528415 180010 528453 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_4_69.VGND
rlabel comment 179938 528435 179938 528435 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_4_69.tapvpwrvgnd_1
rlabel metal1 179938 528387 180030 528483 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_4_69.VGND
rlabel metal1 179938 527843 180030 527939 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_4_69.VPWR
flabel metal1 180980 528418 181014 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._26_.VGND
flabel metal1 180980 527874 181014 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0._26_.VPWR
flabel locali 181624 528112 181658 528146 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._26_.S
flabel locali 181532 528112 181566 528146 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._26_.S
flabel locali 181440 528248 181474 528282 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._26_.A1
flabel locali 181440 528180 181474 528214 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._26_.A1
flabel locali 181348 528180 181382 528214 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._26_.A0
flabel locali 180980 528316 181014 528350 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._26_.X
flabel locali 180980 528044 181014 528078 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._26_.X
flabel locali 180980 527976 181014 528010 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._26_.X
flabel nwell 181024 527874 181058 527908 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._26_.VPB
flabel pwell 181034 528418 181068 528452 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0._26_.VNB
rlabel comment 180950 528435 180950 528435 2 dpga_flat_0.sr_0._26_.mux2_1
rlabel metal1 180950 528387 181778 528483 5 dpga_flat_0.sr_0._26_.VGND
rlabel metal1 180950 527843 181778 527939 5 dpga_flat_0.sr_0._26_.VPWR
flabel metal1 182911 528418 182945 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_116.VGND
flabel metal1 182911 527874 182945 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_116.VPWR
flabel nwell 182911 527874 182945 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_116.VPB
flabel pwell 182911 528418 182945 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_116.VNB
rlabel comment 182882 528435 182882 528435 2 dpga_flat_0.sr_0.FILLER_0_4_116.decap_12
flabel metal1 184015 528418 184049 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_128.VGND
flabel metal1 184015 527874 184049 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_128.VPWR
flabel nwell 184015 527874 184049 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_128.VPB
flabel pwell 184015 528418 184049 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_128.VNB
rlabel comment 183986 528435 183986 528435 2 dpga_flat_0.sr_0.FILLER_0_4_128.decap_12
flabel metal1 185211 528418 185245 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_141.VGND
flabel metal1 185211 527874 185245 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_141.VPWR
flabel nwell 185211 527874 185245 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_141.VPB
flabel pwell 185211 528418 185245 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_141.VNB
rlabel comment 185182 528435 185182 528435 2 dpga_flat_0.sr_0.FILLER_0_4_141.decap_12
flabel metal1 185112 527882 185165 527911 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_4_70.VPWR
flabel metal1 185111 528415 185162 528453 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_4_70.VGND
rlabel comment 185090 528435 185090 528435 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_4_70.tapvpwrvgnd_1
rlabel metal1 185090 528387 185182 528483 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_4_70.VGND
rlabel metal1 185090 527843 185182 527939 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_4_70.VPWR
flabel metal1 186315 527874 186349 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_153.VPWR
flabel metal1 186315 528418 186349 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_153.VGND
flabel nwell 186315 527874 186349 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_153.VPB
flabel pwell 186315 528418 186349 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_153.VNB
rlabel comment 186286 528435 186286 528435 2 dpga_flat_0.sr_0.FILLER_0_4_153.decap_8
rlabel metal1 186286 528387 187022 528483 5 dpga_flat_0.sr_0.FILLER_0_4_153.VGND
rlabel metal1 186286 527843 187022 527939 5 dpga_flat_0.sr_0.FILLER_0_4_153.VPWR
flabel metal1 187042 528417 187095 528449 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_161.VGND
flabel metal1 187043 527874 187095 527905 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_161.VPWR
flabel nwell 187050 527882 187084 527900 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_161.VPB
flabel pwell 187053 528423 187085 528445 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_4_161.VNB
rlabel comment 187022 528435 187022 528435 2 dpga_flat_0.sr_0.FILLER_0_4_161.fill_2
rlabel metal1 187022 528387 187206 528483 5 dpga_flat_0.sr_0.FILLER_0_4_161.VGND
rlabel metal1 187022 527843 187206 527939 5 dpga_flat_0.sr_0.FILLER_0_4_161.VPWR
flabel metal1 187419 527874 187453 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_4_Right_4.VPWR
flabel metal1 187419 528418 187453 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_4_Right_4.VGND
flabel nwell 187419 527874 187453 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_4_Right_4.VPB
flabel pwell 187419 528418 187453 528452 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_4_Right_4.VNB
rlabel comment 187482 528435 187482 528435 8 dpga_flat_0.sr_0.PHY_EDGE_ROW_4_Right_4.decap_3
rlabel metal1 187206 528387 187482 528483 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_4_Right_4.VGND
rlabel metal1 187206 527843 187482 527939 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_4_Right_4.VPWR
flabel metal1 172515 527330 172549 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_3.VGND
flabel metal1 172515 527874 172549 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_3.VPWR
flabel nwell 172515 527874 172549 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_3.VPB
flabel pwell 172515 527330 172549 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_3.VNB
rlabel comment 172486 527347 172486 527347 4 dpga_flat_0.sr_0.FILLER_0_5_3.decap_12
flabel metal1 173619 527330 173653 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_15.VGND
flabel metal1 173619 527874 173653 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_15.VPWR
flabel nwell 173619 527874 173653 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_15.VPB
flabel pwell 173619 527330 173653 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_15.VNB
rlabel comment 173590 527347 173590 527347 4 dpga_flat_0.sr_0.FILLER_0_5_15.decap_12
flabel metal1 172239 527874 172273 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_5_Left_33.VPWR
flabel metal1 172239 527330 172273 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_5_Left_33.VGND
flabel nwell 172239 527874 172273 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_5_Left_33.VPB
flabel pwell 172239 527330 172273 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_5_Left_33.VNB
rlabel comment 172210 527347 172210 527347 4 dpga_flat_0.sr_0.PHY_EDGE_ROW_5_Left_33.decap_3
rlabel metal1 172210 527299 172486 527395 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_5_Left_33.VGND
rlabel metal1 172210 527843 172486 527939 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_5_Left_33.VPWR
flabel metal1 174723 527330 174757 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_27.VGND
flabel metal1 174723 527874 174757 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_27.VPWR
flabel nwell 174723 527874 174757 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_27.VPB
flabel pwell 174723 527330 174757 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_27.VNB
rlabel comment 174694 527347 174694 527347 4 dpga_flat_0.sr_0.FILLER_0_5_27.decap_12
flabel metal1 175827 527874 175861 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_39.VPWR
flabel metal1 175827 527330 175861 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_39.VGND
flabel nwell 175827 527874 175861 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_39.VPB
flabel pwell 175827 527330 175861 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_39.VNB
rlabel comment 175798 527347 175798 527347 4 dpga_flat_0.sr_0.FILLER_0_5_39.decap_6
rlabel metal1 175798 527299 176350 527395 1 dpga_flat_0.sr_0.FILLER_0_5_39.VGND
rlabel metal1 175798 527843 176350 527939 1 dpga_flat_0.sr_0.FILLER_0_5_39.VPWR
flabel metal1 177115 527874 177149 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_53.VPWR
flabel metal1 177115 527330 177149 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_53.VGND
flabel nwell 177115 527874 177149 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_53.VPB
flabel pwell 177115 527330 177149 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_53.VNB
rlabel comment 177086 527347 177086 527347 4 dpga_flat_0.sr_0.FILLER_0_5_53.decap_3
rlabel metal1 177086 527299 177362 527395 1 dpga_flat_0.sr_0.FILLER_0_5_53.VGND
rlabel metal1 177086 527843 177362 527939 1 dpga_flat_0.sr_0.FILLER_0_5_53.VPWR
flabel metal1 177483 527330 177517 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_57.VGND
flabel metal1 177483 527874 177517 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_57.VPWR
flabel nwell 177483 527874 177517 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_57.VPB
flabel pwell 177483 527330 177517 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_57.VNB
rlabel comment 177454 527347 177454 527347 4 dpga_flat_0.sr_0.FILLER_0_5_57.decap_12
flabel metal1 177384 527871 177437 527900 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_5_71.VPWR
flabel metal1 177383 527329 177434 527367 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_5_71.VGND
rlabel comment 177362 527347 177362 527347 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_5_71.tapvpwrvgnd_1
rlabel metal1 177362 527299 177454 527395 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_5_71.VGND
rlabel metal1 177362 527843 177454 527939 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_5_71.VPWR
flabel locali 177023 527568 177057 527602 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold3.A
flabel locali 176375 527500 176409 527534 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold3.X
flabel locali 177023 527636 177057 527670 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold3.A
flabel locali 176375 527432 176409 527466 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold3.X
flabel locali 176931 527568 176965 527602 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold3.A
flabel locali 176931 527636 176965 527670 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold3.A
flabel locali 176375 527772 176409 527806 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold3.X
flabel locali 176375 527636 176409 527670 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold3.X
flabel locali 176375 527704 176409 527738 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold3.X
flabel locali 176375 527568 176409 527602 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold3.X
flabel nwell 177023 527874 177057 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold3.VPB
flabel pwell 177023 527330 177057 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold3.VNB
flabel metal1 177023 527330 177057 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold3.VGND
flabel metal1 177023 527874 177057 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold3.VPWR
rlabel comment 177086 527347 177086 527347 6 dpga_flat_0.sr_0.hold3.dlygate4sd3_1
rlabel metal1 176350 527299 177086 527395 1 dpga_flat_0.sr_0.hold3.VGND
rlabel metal1 176350 527843 177086 527939 1 dpga_flat_0.sr_0.hold3.VPWR
flabel metal1 178587 527330 178621 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_69.VGND
flabel metal1 178587 527874 178621 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_69.VPWR
flabel nwell 178587 527874 178621 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_69.VPB
flabel pwell 178587 527330 178621 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_69.VNB
rlabel comment 178558 527347 178558 527347 4 dpga_flat_0.sr_0.FILLER_0_5_69.decap_4
rlabel metal1 178558 527299 178926 527395 1 dpga_flat_0.sr_0.FILLER_0_5_69.VGND
rlabel metal1 178558 527843 178926 527939 1 dpga_flat_0.sr_0.FILLER_0_5_69.VPWR
flabel metal1 179691 527330 179725 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_81.VGND
flabel metal1 179691 527874 179725 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_81.VPWR
flabel nwell 179691 527874 179725 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_81.VPB
flabel pwell 179691 527330 179725 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_81.VNB
rlabel comment 179662 527347 179662 527347 4 dpga_flat_0.sr_0.FILLER_0_5_81.decap_12
flabel locali 179599 527568 179633 527602 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold4.A
flabel locali 178951 527500 178985 527534 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold4.X
flabel locali 179599 527636 179633 527670 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold4.A
flabel locali 178951 527432 178985 527466 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold4.X
flabel locali 179507 527568 179541 527602 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold4.A
flabel locali 179507 527636 179541 527670 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold4.A
flabel locali 178951 527772 178985 527806 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold4.X
flabel locali 178951 527636 178985 527670 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold4.X
flabel locali 178951 527704 178985 527738 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold4.X
flabel locali 178951 527568 178985 527602 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold4.X
flabel nwell 179599 527874 179633 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold4.VPB
flabel pwell 179599 527330 179633 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold4.VNB
flabel metal1 179599 527330 179633 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold4.VGND
flabel metal1 179599 527874 179633 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.hold4.VPWR
rlabel comment 179662 527347 179662 527347 6 dpga_flat_0.sr_0.hold4.dlygate4sd3_1
rlabel metal1 178926 527299 179662 527395 1 dpga_flat_0.sr_0.hold4.VGND
rlabel metal1 178926 527843 179662 527939 1 dpga_flat_0.sr_0.hold4.VPWR
flabel metal1 180795 527330 180829 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_93.VGND
flabel metal1 180795 527874 180829 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_93.VPWR
flabel nwell 180795 527874 180829 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_93.VPB
flabel pwell 180795 527330 180829 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_93.VNB
rlabel comment 180766 527347 180766 527347 4 dpga_flat_0.sr_0.FILLER_0_5_93.decap_12
flabel metal1 181899 527874 181933 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_105.VPWR
flabel metal1 181899 527330 181933 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_105.VGND
flabel nwell 181899 527874 181933 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_105.VPB
flabel pwell 181899 527330 181933 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_105.VNB
rlabel comment 181870 527347 181870 527347 4 dpga_flat_0.sr_0.FILLER_0_5_105.decap_6
rlabel metal1 181870 527299 182422 527395 1 dpga_flat_0.sr_0.FILLER_0_5_105.VGND
rlabel metal1 181870 527843 182422 527939 1 dpga_flat_0.sr_0.FILLER_0_5_105.VPWR
flabel metal1 182444 527874 182480 527904 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_111.VPWR
flabel metal1 182444 527334 182480 527363 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_111.VGND
flabel nwell 182453 527881 182473 527898 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_111.VPB
flabel pwell 182450 527336 182474 527358 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_111.VNB
rlabel comment 182422 527347 182422 527347 4 dpga_flat_0.sr_0.FILLER_0_5_111.fill_1
rlabel metal1 182422 527299 182514 527395 1 dpga_flat_0.sr_0.FILLER_0_5_111.VGND
rlabel metal1 182422 527843 182514 527939 1 dpga_flat_0.sr_0.FILLER_0_5_111.VPWR
flabel metal1 182635 527330 182669 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_113.VGND
flabel metal1 182635 527874 182669 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_113.VPWR
flabel nwell 182635 527874 182669 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_113.VPB
flabel pwell 182635 527330 182669 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_113.VNB
rlabel comment 182606 527347 182606 527347 4 dpga_flat_0.sr_0.FILLER_0_5_113.decap_12
flabel metal1 183739 527330 183773 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_125.VGND
flabel metal1 183739 527874 183773 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_125.VPWR
flabel nwell 183739 527874 183773 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_125.VPB
flabel pwell 183739 527330 183773 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_125.VNB
rlabel comment 183710 527347 183710 527347 4 dpga_flat_0.sr_0.FILLER_0_5_125.decap_12
flabel metal1 182536 527871 182589 527900 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_5_72.VPWR
flabel metal1 182535 527329 182586 527367 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_5_72.VGND
rlabel comment 182514 527347 182514 527347 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_5_72.tapvpwrvgnd_1
rlabel metal1 182514 527299 182606 527395 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_5_72.VGND
rlabel metal1 182514 527843 182606 527939 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_5_72.VPWR
flabel metal1 184843 527330 184877 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_137.VGND
flabel metal1 184843 527874 184877 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_137.VPWR
flabel nwell 184843 527874 184877 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_137.VPB
flabel pwell 184843 527330 184877 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_137.VNB
rlabel comment 184814 527347 184814 527347 4 dpga_flat_0.sr_0.FILLER_0_5_137.decap_12
flabel metal1 185947 527330 185981 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_149.VGND
flabel metal1 185947 527874 185981 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_149.VPWR
flabel nwell 185947 527874 185981 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_149.VPB
flabel pwell 185947 527330 185981 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_149.VNB
rlabel comment 185918 527347 185918 527347 4 dpga_flat_0.sr_0.FILLER_0_5_149.decap_12
flabel metal1 187042 527333 187095 527365 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_161.VGND
flabel metal1 187043 527877 187095 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_161.VPWR
flabel nwell 187050 527882 187084 527900 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_161.VPB
flabel pwell 187053 527337 187085 527359 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_5_161.VNB
rlabel comment 187022 527347 187022 527347 4 dpga_flat_0.sr_0.FILLER_0_5_161.fill_2
rlabel metal1 187022 527299 187206 527395 1 dpga_flat_0.sr_0.FILLER_0_5_161.VGND
rlabel metal1 187022 527843 187206 527939 1 dpga_flat_0.sr_0.FILLER_0_5_161.VPWR
flabel metal1 187419 527874 187453 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_5_Right_5.VPWR
flabel metal1 187419 527330 187453 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_5_Right_5.VGND
flabel nwell 187419 527874 187453 527908 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_5_Right_5.VPB
flabel pwell 187419 527330 187453 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_5_Right_5.VNB
rlabel comment 187482 527347 187482 527347 6 dpga_flat_0.sr_0.PHY_EDGE_ROW_5_Right_5.decap_3
rlabel metal1 187206 527299 187482 527395 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_5_Right_5.VGND
rlabel metal1 187206 527843 187482 527939 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_5_Right_5.VPWR
flabel metal1 172515 527330 172549 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_3.VGND
flabel metal1 172515 526786 172549 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_3.VPWR
flabel nwell 172515 526786 172549 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_3.VPB
flabel pwell 172515 527330 172549 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_3.VNB
rlabel comment 172486 527347 172486 527347 2 dpga_flat_0.sr_0.FILLER_0_6_3.decap_12
flabel metal1 173619 527330 173653 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_15.VGND
flabel metal1 173619 526786 173653 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_15.VPWR
flabel nwell 173619 526786 173653 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_15.VPB
flabel pwell 173619 527330 173653 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_15.VNB
rlabel comment 173590 527347 173590 527347 2 dpga_flat_0.sr_0.FILLER_0_6_15.decap_12
flabel metal1 172515 526242 172549 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_3.VGND
flabel metal1 172515 526786 172549 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_3.VPWR
flabel nwell 172515 526786 172549 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_3.VPB
flabel pwell 172515 526242 172549 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_3.VNB
rlabel comment 172486 526259 172486 526259 4 dpga_flat_0.sr_0.FILLER_0_7_3.decap_12
flabel metal1 173619 526242 173653 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_15.VGND
flabel metal1 173619 526786 173653 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_15.VPWR
flabel nwell 173619 526786 173653 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_15.VPB
flabel pwell 173619 526242 173653 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_15.VNB
rlabel comment 173590 526259 173590 526259 4 dpga_flat_0.sr_0.FILLER_0_7_15.decap_12
flabel metal1 172239 526786 172273 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_6_Left_34.VPWR
flabel metal1 172239 527330 172273 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_6_Left_34.VGND
flabel nwell 172239 526786 172273 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_6_Left_34.VPB
flabel pwell 172239 527330 172273 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_6_Left_34.VNB
rlabel comment 172210 527347 172210 527347 2 dpga_flat_0.sr_0.PHY_EDGE_ROW_6_Left_34.decap_3
rlabel metal1 172210 527299 172486 527395 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_6_Left_34.VGND
rlabel metal1 172210 526755 172486 526851 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_6_Left_34.VPWR
flabel metal1 172239 526786 172273 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_7_Left_35.VPWR
flabel metal1 172239 526242 172273 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_7_Left_35.VGND
flabel nwell 172239 526786 172273 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_7_Left_35.VPB
flabel pwell 172239 526242 172273 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_7_Left_35.VNB
rlabel comment 172210 526259 172210 526259 4 dpga_flat_0.sr_0.PHY_EDGE_ROW_7_Left_35.decap_3
rlabel metal1 172210 526211 172486 526307 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_7_Left_35.VGND
rlabel metal1 172210 526755 172486 526851 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_7_Left_35.VPWR
flabel metal1 174716 526790 174752 526820 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_27.VPWR
flabel metal1 174716 527331 174752 527360 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_27.VGND
flabel nwell 174725 526796 174745 526813 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_27.VPB
flabel pwell 174722 527336 174746 527358 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_27.VNB
rlabel comment 174694 527347 174694 527347 2 dpga_flat_0.sr_0.FILLER_0_6_27.fill_1
rlabel metal1 174694 527299 174786 527395 5 dpga_flat_0.sr_0.FILLER_0_6_27.VGND
rlabel metal1 174694 526755 174786 526851 5 dpga_flat_0.sr_0.FILLER_0_6_27.VPWR
flabel metal1 174907 527330 174941 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_29.VGND
flabel metal1 174907 526786 174941 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_29.VPWR
flabel nwell 174907 526786 174941 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_29.VPB
flabel pwell 174907 527330 174941 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_29.VNB
rlabel comment 174878 527347 174878 527347 2 dpga_flat_0.sr_0.FILLER_0_6_29.decap_12
flabel metal1 176011 527330 176045 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_41.VGND
flabel metal1 176011 526786 176045 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_41.VPWR
flabel nwell 176011 526786 176045 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_41.VPB
flabel pwell 176011 527330 176045 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_41.VNB
rlabel comment 175982 527347 175982 527347 2 dpga_flat_0.sr_0.FILLER_0_6_41.decap_12
flabel metal1 174723 526242 174757 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_27.VGND
flabel metal1 174723 526786 174757 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_27.VPWR
flabel nwell 174723 526786 174757 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_27.VPB
flabel pwell 174723 526242 174757 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_27.VNB
rlabel comment 174694 526259 174694 526259 4 dpga_flat_0.sr_0.FILLER_0_7_27.decap_12
flabel metal1 175827 526242 175861 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_39.VGND
flabel metal1 175827 526786 175861 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_39.VPWR
flabel nwell 175827 526786 175861 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_39.VPB
flabel pwell 175827 526242 175861 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_39.VNB
rlabel comment 175798 526259 175798 526259 4 dpga_flat_0.sr_0.FILLER_0_7_39.decap_12
flabel metal1 174808 526794 174861 526823 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_6_73.VPWR
flabel metal1 174807 527327 174858 527365 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_6_73.VGND
rlabel comment 174786 527347 174786 527347 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_6_73.tapvpwrvgnd_1
rlabel metal1 174786 527299 174878 527395 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_6_73.VGND
rlabel metal1 174786 526755 174878 526851 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_6_73.VPWR
flabel metal1 177115 527330 177149 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_53.VGND
flabel metal1 177115 526786 177149 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_53.VPWR
flabel nwell 177115 526786 177149 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_53.VPB
flabel pwell 177115 527330 177149 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_53.VNB
rlabel comment 177086 527347 177086 527347 2 dpga_flat_0.sr_0.FILLER_0_6_53.decap_12
flabel metal1 176931 526242 176965 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_51.VGND
flabel metal1 176931 526786 176965 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_51.VPWR
flabel nwell 176931 526786 176965 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_51.VPB
flabel pwell 176931 526242 176965 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_51.VNB
rlabel comment 176902 526259 176902 526259 4 dpga_flat_0.sr_0.FILLER_0_7_51.decap_4
rlabel metal1 176902 526211 177270 526307 1 dpga_flat_0.sr_0.FILLER_0_7_51.VGND
rlabel metal1 176902 526755 177270 526851 1 dpga_flat_0.sr_0.FILLER_0_7_51.VPWR
flabel metal1 177292 526786 177328 526816 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_55.VPWR
flabel metal1 177292 526246 177328 526275 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_55.VGND
flabel nwell 177301 526793 177321 526810 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_55.VPB
flabel pwell 177298 526248 177322 526270 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_55.VNB
rlabel comment 177270 526259 177270 526259 4 dpga_flat_0.sr_0.FILLER_0_7_55.fill_1
rlabel metal1 177270 526211 177362 526307 1 dpga_flat_0.sr_0.FILLER_0_7_55.VGND
rlabel metal1 177270 526755 177362 526851 1 dpga_flat_0.sr_0.FILLER_0_7_55.VPWR
flabel metal1 177483 526242 177517 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_57.VGND
flabel metal1 177483 526786 177517 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_57.VPWR
flabel nwell 177483 526786 177517 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_57.VPB
flabel pwell 177483 526242 177517 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_57.VNB
rlabel comment 177454 526259 177454 526259 4 dpga_flat_0.sr_0.FILLER_0_7_57.decap_12
flabel metal1 177384 526783 177437 526812 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_7_76.VPWR
flabel metal1 177383 526241 177434 526279 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_7_76.VGND
rlabel comment 177362 526259 177362 526259 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_7_76.tapvpwrvgnd_1
rlabel metal1 177362 526211 177454 526307 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_7_76.VGND
rlabel metal1 177362 526755 177454 526851 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_7_76.VPWR
flabel metal1 178219 527330 178253 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_65.VGND
flabel metal1 178219 526786 178253 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_65.VPWR
flabel nwell 178219 526786 178253 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_65.VPB
flabel pwell 178219 527330 178253 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_65.VNB
rlabel comment 178190 527347 178190 527347 2 dpga_flat_0.sr_0.FILLER_0_6_65.decap_12
flabel metal1 179323 526786 179357 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_77.VPWR
flabel metal1 179323 527330 179357 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_77.VGND
flabel nwell 179323 526786 179357 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_77.VPB
flabel pwell 179323 527330 179357 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_77.VNB
rlabel comment 179294 527347 179294 527347 2 dpga_flat_0.sr_0.FILLER_0_6_77.decap_6
rlabel metal1 179294 527299 179846 527395 5 dpga_flat_0.sr_0.FILLER_0_6_77.VGND
rlabel metal1 179294 526755 179846 526851 5 dpga_flat_0.sr_0.FILLER_0_6_77.VPWR
flabel metal1 179868 526790 179904 526820 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_83.VPWR
flabel metal1 179868 527331 179904 527360 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_83.VGND
flabel nwell 179877 526796 179897 526813 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_83.VPB
flabel pwell 179874 527336 179898 527358 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_83.VNB
rlabel comment 179846 527347 179846 527347 2 dpga_flat_0.sr_0.FILLER_0_6_83.fill_1
rlabel metal1 179846 527299 179938 527395 5 dpga_flat_0.sr_0.FILLER_0_6_83.VGND
rlabel metal1 179846 526755 179938 526851 5 dpga_flat_0.sr_0.FILLER_0_6_83.VPWR
flabel metal1 178587 526242 178621 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_69.VGND
flabel metal1 178587 526786 178621 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_69.VPWR
flabel nwell 178587 526786 178621 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_69.VPB
flabel pwell 178587 526242 178621 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_69.VNB
rlabel comment 178558 526259 178558 526259 4 dpga_flat_0.sr_0.FILLER_0_7_69.decap_12
flabel metal1 179691 526242 179725 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_81.VGND
flabel metal1 179691 526786 179725 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_81.VPWR
flabel nwell 179691 526786 179725 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_81.VPB
flabel pwell 179691 526242 179725 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_81.VNB
rlabel comment 179662 526259 179662 526259 4 dpga_flat_0.sr_0.FILLER_0_7_81.decap_12
flabel metal1 180059 527330 180093 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_85.VGND
flabel metal1 180059 526786 180093 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_85.VPWR
flabel nwell 180059 526786 180093 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_85.VPB
flabel pwell 180059 527330 180093 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_85.VNB
rlabel comment 180030 527347 180030 527347 2 dpga_flat_0.sr_0.FILLER_0_6_85.decap_12
flabel metal1 181163 527330 181197 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_97.VGND
flabel metal1 181163 526786 181197 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_97.VPWR
flabel nwell 181163 526786 181197 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_97.VPB
flabel pwell 181163 527330 181197 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_97.VNB
rlabel comment 181134 527347 181134 527347 2 dpga_flat_0.sr_0.FILLER_0_6_97.decap_12
flabel metal1 180795 526242 180829 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_93.VGND
flabel metal1 180795 526786 180829 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_93.VPWR
flabel nwell 180795 526786 180829 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_93.VPB
flabel pwell 180795 526242 180829 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_93.VNB
rlabel comment 180766 526259 180766 526259 4 dpga_flat_0.sr_0.FILLER_0_7_93.decap_12
flabel metal1 179960 526794 180013 526823 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_6_74.VPWR
flabel metal1 179959 527327 180010 527365 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_6_74.VGND
rlabel comment 179938 527347 179938 527347 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_6_74.tapvpwrvgnd_1
rlabel metal1 179938 527299 180030 527395 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_6_74.VGND
rlabel metal1 179938 526755 180030 526851 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_6_74.VPWR
flabel metal1 182267 527330 182301 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_109.VGND
flabel metal1 182267 526786 182301 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_109.VPWR
flabel nwell 182267 526786 182301 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_109.VPB
flabel pwell 182267 527330 182301 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_109.VNB
rlabel comment 182238 527347 182238 527347 2 dpga_flat_0.sr_0.FILLER_0_6_109.decap_12
flabel metal1 183371 527330 183405 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_121.VGND
flabel metal1 183371 526786 183405 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_121.VPWR
flabel nwell 183371 526786 183405 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_121.VPB
flabel pwell 183371 527330 183405 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_121.VNB
rlabel comment 183342 527347 183342 527347 2 dpga_flat_0.sr_0.FILLER_0_6_121.decap_12
flabel metal1 181899 526786 181933 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_105.VPWR
flabel metal1 181899 526242 181933 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_105.VGND
flabel nwell 181899 526786 181933 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_105.VPB
flabel pwell 181899 526242 181933 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_105.VNB
rlabel comment 181870 526259 181870 526259 4 dpga_flat_0.sr_0.FILLER_0_7_105.decap_6
rlabel metal1 181870 526211 182422 526307 1 dpga_flat_0.sr_0.FILLER_0_7_105.VGND
rlabel metal1 181870 526755 182422 526851 1 dpga_flat_0.sr_0.FILLER_0_7_105.VPWR
flabel metal1 182444 526786 182480 526816 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_111.VPWR
flabel metal1 182444 526246 182480 526275 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_111.VGND
flabel nwell 182453 526793 182473 526810 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_111.VPB
flabel pwell 182450 526248 182474 526270 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_111.VNB
rlabel comment 182422 526259 182422 526259 4 dpga_flat_0.sr_0.FILLER_0_7_111.fill_1
rlabel metal1 182422 526211 182514 526307 1 dpga_flat_0.sr_0.FILLER_0_7_111.VGND
rlabel metal1 182422 526755 182514 526851 1 dpga_flat_0.sr_0.FILLER_0_7_111.VPWR
flabel metal1 182635 526242 182669 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_113.VGND
flabel metal1 182635 526786 182669 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_113.VPWR
flabel nwell 182635 526786 182669 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_113.VPB
flabel pwell 182635 526242 182669 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_113.VNB
rlabel comment 182606 526259 182606 526259 4 dpga_flat_0.sr_0.FILLER_0_7_113.decap_12
flabel metal1 183739 526242 183773 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_125.VGND
flabel metal1 183739 526786 183773 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_125.VPWR
flabel nwell 183739 526786 183773 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_125.VPB
flabel pwell 183739 526242 183773 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_125.VNB
rlabel comment 183710 526259 183710 526259 4 dpga_flat_0.sr_0.FILLER_0_7_125.decap_12
flabel metal1 182536 526783 182589 526812 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_7_77.VPWR
flabel metal1 182535 526241 182586 526279 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_7_77.VGND
rlabel comment 182514 526259 182514 526259 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_7_77.tapvpwrvgnd_1
rlabel metal1 182514 526211 182606 526307 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_7_77.VGND
rlabel metal1 182514 526755 182606 526851 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_7_77.VPWR
flabel metal1 184475 526786 184509 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_133.VPWR
flabel metal1 184475 527330 184509 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_133.VGND
flabel nwell 184475 526786 184509 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_133.VPB
flabel pwell 184475 527330 184509 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_133.VNB
rlabel comment 184446 527347 184446 527347 2 dpga_flat_0.sr_0.FILLER_0_6_133.decap_6
rlabel metal1 184446 527299 184998 527395 5 dpga_flat_0.sr_0.FILLER_0_6_133.VGND
rlabel metal1 184446 526755 184998 526851 5 dpga_flat_0.sr_0.FILLER_0_6_133.VPWR
flabel metal1 185020 526790 185056 526820 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_139.VPWR
flabel metal1 185020 527331 185056 527360 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_139.VGND
flabel nwell 185029 526796 185049 526813 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_139.VPB
flabel pwell 185026 527336 185050 527358 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_139.VNB
rlabel comment 184998 527347 184998 527347 2 dpga_flat_0.sr_0.FILLER_0_6_139.fill_1
rlabel metal1 184998 527299 185090 527395 5 dpga_flat_0.sr_0.FILLER_0_6_139.VGND
rlabel metal1 184998 526755 185090 526851 5 dpga_flat_0.sr_0.FILLER_0_6_139.VPWR
flabel metal1 185211 527330 185245 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_141.VGND
flabel metal1 185211 526786 185245 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_141.VPWR
flabel nwell 185211 526786 185245 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_141.VPB
flabel pwell 185211 527330 185245 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_141.VNB
rlabel comment 185182 527347 185182 527347 2 dpga_flat_0.sr_0.FILLER_0_6_141.decap_12
flabel metal1 184843 526242 184877 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_137.VGND
flabel metal1 184843 526786 184877 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_137.VPWR
flabel nwell 184843 526786 184877 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_137.VPB
flabel pwell 184843 526242 184877 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_137.VNB
rlabel comment 184814 526259 184814 526259 4 dpga_flat_0.sr_0.FILLER_0_7_137.decap_12
flabel metal1 185112 526794 185165 526823 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_6_75.VPWR
flabel metal1 185111 527327 185162 527365 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_6_75.VGND
rlabel comment 185090 527347 185090 527347 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_6_75.tapvpwrvgnd_1
rlabel metal1 185090 527299 185182 527395 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_6_75.VGND
rlabel metal1 185090 526755 185182 526851 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_6_75.VPWR
flabel metal1 186315 526786 186349 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_153.VPWR
flabel metal1 186315 527330 186349 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_153.VGND
flabel nwell 186315 526786 186349 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_153.VPB
flabel pwell 186315 527330 186349 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_153.VNB
rlabel comment 186286 527347 186286 527347 2 dpga_flat_0.sr_0.FILLER_0_6_153.decap_8
rlabel metal1 186286 527299 187022 527395 5 dpga_flat_0.sr_0.FILLER_0_6_153.VGND
rlabel metal1 186286 526755 187022 526851 5 dpga_flat_0.sr_0.FILLER_0_6_153.VPWR
flabel metal1 187042 527329 187095 527361 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_161.VGND
flabel metal1 187043 526786 187095 526817 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_161.VPWR
flabel nwell 187050 526794 187084 526812 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_161.VPB
flabel pwell 187053 527335 187085 527357 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_6_161.VNB
rlabel comment 187022 527347 187022 527347 2 dpga_flat_0.sr_0.FILLER_0_6_161.fill_2
rlabel metal1 187022 527299 187206 527395 5 dpga_flat_0.sr_0.FILLER_0_6_161.VGND
rlabel metal1 187022 526755 187206 526851 5 dpga_flat_0.sr_0.FILLER_0_6_161.VPWR
flabel metal1 185947 526242 185981 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_149.VGND
flabel metal1 185947 526786 185981 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_149.VPWR
flabel nwell 185947 526786 185981 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_149.VPB
flabel pwell 185947 526242 185981 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_149.VNB
rlabel comment 185918 526259 185918 526259 4 dpga_flat_0.sr_0.FILLER_0_7_149.decap_12
flabel metal1 187042 526245 187095 526277 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_161.VGND
flabel metal1 187043 526789 187095 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_161.VPWR
flabel nwell 187050 526794 187084 526812 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_161.VPB
flabel pwell 187053 526249 187085 526271 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_7_161.VNB
rlabel comment 187022 526259 187022 526259 4 dpga_flat_0.sr_0.FILLER_0_7_161.fill_2
rlabel metal1 187022 526211 187206 526307 1 dpga_flat_0.sr_0.FILLER_0_7_161.VGND
rlabel metal1 187022 526755 187206 526851 1 dpga_flat_0.sr_0.FILLER_0_7_161.VPWR
flabel metal1 187419 526786 187453 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_6_Right_6.VPWR
flabel metal1 187419 527330 187453 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_6_Right_6.VGND
flabel nwell 187419 526786 187453 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_6_Right_6.VPB
flabel pwell 187419 527330 187453 527364 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_6_Right_6.VNB
rlabel comment 187482 527347 187482 527347 8 dpga_flat_0.sr_0.PHY_EDGE_ROW_6_Right_6.decap_3
rlabel metal1 187206 527299 187482 527395 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_6_Right_6.VGND
rlabel metal1 187206 526755 187482 526851 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_6_Right_6.VPWR
flabel metal1 187419 526786 187453 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_7_Right_7.VPWR
flabel metal1 187419 526242 187453 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_7_Right_7.VGND
flabel nwell 187419 526786 187453 526820 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_7_Right_7.VPB
flabel pwell 187419 526242 187453 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_7_Right_7.VNB
rlabel comment 187482 526259 187482 526259 6 dpga_flat_0.sr_0.PHY_EDGE_ROW_7_Right_7.decap_3
rlabel metal1 187206 526211 187482 526307 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_7_Right_7.VGND
rlabel metal1 187206 526755 187482 526851 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_7_Right_7.VPWR
flabel metal1 172515 526242 172549 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_3.VGND
flabel metal1 172515 525698 172549 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_3.VPWR
flabel nwell 172515 525698 172549 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_3.VPB
flabel pwell 172515 526242 172549 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_3.VNB
rlabel comment 172486 526259 172486 526259 2 dpga_flat_0.sr_0.FILLER_0_8_3.decap_12
flabel metal1 173619 526242 173653 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_15.VGND
flabel metal1 173619 525698 173653 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_15.VPWR
flabel nwell 173619 525698 173653 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_15.VPB
flabel pwell 173619 526242 173653 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_15.VNB
rlabel comment 173590 526259 173590 526259 2 dpga_flat_0.sr_0.FILLER_0_8_15.decap_12
flabel metal1 172239 525698 172273 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_8_Left_36.VPWR
flabel metal1 172239 526242 172273 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_8_Left_36.VGND
flabel nwell 172239 525698 172273 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_8_Left_36.VPB
flabel pwell 172239 526242 172273 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_8_Left_36.VNB
rlabel comment 172210 526259 172210 526259 2 dpga_flat_0.sr_0.PHY_EDGE_ROW_8_Left_36.decap_3
rlabel metal1 172210 526211 172486 526307 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_8_Left_36.VGND
rlabel metal1 172210 525667 172486 525763 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_8_Left_36.VPWR
flabel metal1 174716 525702 174752 525732 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_27.VPWR
flabel metal1 174716 526243 174752 526272 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_27.VGND
flabel nwell 174725 525708 174745 525725 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_27.VPB
flabel pwell 174722 526248 174746 526270 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_27.VNB
rlabel comment 174694 526259 174694 526259 2 dpga_flat_0.sr_0.FILLER_0_8_27.fill_1
rlabel metal1 174694 526211 174786 526307 5 dpga_flat_0.sr_0.FILLER_0_8_27.VGND
rlabel metal1 174694 525667 174786 525763 5 dpga_flat_0.sr_0.FILLER_0_8_27.VPWR
flabel metal1 174907 526242 174941 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_29.VGND
flabel metal1 174907 525698 174941 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_29.VPWR
flabel nwell 174907 525698 174941 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_29.VPB
flabel pwell 174907 526242 174941 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_29.VNB
rlabel comment 174878 526259 174878 526259 2 dpga_flat_0.sr_0.FILLER_0_8_29.decap_12
flabel metal1 176011 526242 176045 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_41.VGND
flabel metal1 176011 525698 176045 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_41.VPWR
flabel nwell 176011 525698 176045 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_41.VPB
flabel pwell 176011 526242 176045 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_41.VNB
rlabel comment 175982 526259 175982 526259 2 dpga_flat_0.sr_0.FILLER_0_8_41.decap_12
flabel metal1 174808 525706 174861 525735 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_8_78.VPWR
flabel metal1 174807 526239 174858 526277 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_8_78.VGND
rlabel comment 174786 526259 174786 526259 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_8_78.tapvpwrvgnd_1
rlabel metal1 174786 526211 174878 526307 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_8_78.VGND
rlabel metal1 174786 525667 174878 525763 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_8_78.VPWR
flabel metal1 177115 526242 177149 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_53.VGND
flabel metal1 177115 525698 177149 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_53.VPWR
flabel nwell 177115 525698 177149 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_53.VPB
flabel pwell 177115 526242 177149 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_53.VNB
rlabel comment 177086 526259 177086 526259 2 dpga_flat_0.sr_0.FILLER_0_8_53.decap_12
flabel metal1 178219 526242 178253 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_65.VGND
flabel metal1 178219 525698 178253 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_65.VPWR
flabel nwell 178219 525698 178253 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_65.VPB
flabel pwell 178219 526242 178253 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_65.VNB
rlabel comment 178190 526259 178190 526259 2 dpga_flat_0.sr_0.FILLER_0_8_65.decap_12
flabel metal1 179323 525698 179357 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_77.VPWR
flabel metal1 179323 526242 179357 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_77.VGND
flabel nwell 179323 525698 179357 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_77.VPB
flabel pwell 179323 526242 179357 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_77.VNB
rlabel comment 179294 526259 179294 526259 2 dpga_flat_0.sr_0.FILLER_0_8_77.decap_6
rlabel metal1 179294 526211 179846 526307 5 dpga_flat_0.sr_0.FILLER_0_8_77.VGND
rlabel metal1 179294 525667 179846 525763 5 dpga_flat_0.sr_0.FILLER_0_8_77.VPWR
flabel metal1 179868 525702 179904 525732 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_83.VPWR
flabel metal1 179868 526243 179904 526272 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_83.VGND
flabel nwell 179877 525708 179897 525725 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_83.VPB
flabel pwell 179874 526248 179898 526270 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_83.VNB
rlabel comment 179846 526259 179846 526259 2 dpga_flat_0.sr_0.FILLER_0_8_83.fill_1
rlabel metal1 179846 526211 179938 526307 5 dpga_flat_0.sr_0.FILLER_0_8_83.VGND
rlabel metal1 179846 525667 179938 525763 5 dpga_flat_0.sr_0.FILLER_0_8_83.VPWR
flabel metal1 180059 526242 180093 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_85.VGND
flabel metal1 180059 525698 180093 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_85.VPWR
flabel nwell 180059 525698 180093 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_85.VPB
flabel pwell 180059 526242 180093 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_85.VNB
rlabel comment 180030 526259 180030 526259 2 dpga_flat_0.sr_0.FILLER_0_8_85.decap_12
flabel metal1 181163 526242 181197 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_97.VGND
flabel metal1 181163 525698 181197 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_97.VPWR
flabel nwell 181163 525698 181197 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_97.VPB
flabel pwell 181163 526242 181197 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_97.VNB
rlabel comment 181134 526259 181134 526259 2 dpga_flat_0.sr_0.FILLER_0_8_97.decap_12
flabel metal1 179960 525706 180013 525735 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_8_79.VPWR
flabel metal1 179959 526239 180010 526277 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_8_79.VGND
rlabel comment 179938 526259 179938 526259 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_8_79.tapvpwrvgnd_1
rlabel metal1 179938 526211 180030 526307 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_8_79.VGND
rlabel metal1 179938 525667 180030 525763 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_8_79.VPWR
flabel metal1 182267 526242 182301 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_109.VGND
flabel metal1 182267 525698 182301 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_109.VPWR
flabel nwell 182267 525698 182301 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_109.VPB
flabel pwell 182267 526242 182301 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_109.VNB
rlabel comment 182238 526259 182238 526259 2 dpga_flat_0.sr_0.FILLER_0_8_109.decap_12
flabel metal1 183371 526242 183405 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_121.VGND
flabel metal1 183371 525698 183405 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_121.VPWR
flabel nwell 183371 525698 183405 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_121.VPB
flabel pwell 183371 526242 183405 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_121.VNB
rlabel comment 183342 526259 183342 526259 2 dpga_flat_0.sr_0.FILLER_0_8_121.decap_12
flabel metal1 184475 525698 184509 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_133.VPWR
flabel metal1 184475 526242 184509 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_133.VGND
flabel nwell 184475 525698 184509 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_133.VPB
flabel pwell 184475 526242 184509 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_133.VNB
rlabel comment 184446 526259 184446 526259 2 dpga_flat_0.sr_0.FILLER_0_8_133.decap_6
rlabel metal1 184446 526211 184998 526307 5 dpga_flat_0.sr_0.FILLER_0_8_133.VGND
rlabel metal1 184446 525667 184998 525763 5 dpga_flat_0.sr_0.FILLER_0_8_133.VPWR
flabel metal1 185020 525702 185056 525732 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_139.VPWR
flabel metal1 185020 526243 185056 526272 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_139.VGND
flabel nwell 185029 525708 185049 525725 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_139.VPB
flabel pwell 185026 526248 185050 526270 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_139.VNB
rlabel comment 184998 526259 184998 526259 2 dpga_flat_0.sr_0.FILLER_0_8_139.fill_1
rlabel metal1 184998 526211 185090 526307 5 dpga_flat_0.sr_0.FILLER_0_8_139.VGND
rlabel metal1 184998 525667 185090 525763 5 dpga_flat_0.sr_0.FILLER_0_8_139.VPWR
flabel metal1 185211 526242 185245 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_141.VGND
flabel metal1 185211 525698 185245 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_141.VPWR
flabel nwell 185211 525698 185245 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_141.VPB
flabel pwell 185211 526242 185245 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_141.VNB
rlabel comment 185182 526259 185182 526259 2 dpga_flat_0.sr_0.FILLER_0_8_141.decap_12
flabel metal1 185112 525706 185165 525735 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_8_80.VPWR
flabel metal1 185111 526239 185162 526277 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_8_80.VGND
rlabel comment 185090 526259 185090 526259 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_8_80.tapvpwrvgnd_1
rlabel metal1 185090 526211 185182 526307 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_8_80.VGND
rlabel metal1 185090 525667 185182 525763 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_8_80.VPWR
flabel metal1 186315 525698 186349 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_153.VPWR
flabel metal1 186315 526242 186349 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_153.VGND
flabel nwell 186315 525698 186349 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_153.VPB
flabel pwell 186315 526242 186349 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_153.VNB
rlabel comment 186286 526259 186286 526259 2 dpga_flat_0.sr_0.FILLER_0_8_153.decap_8
rlabel metal1 186286 526211 187022 526307 5 dpga_flat_0.sr_0.FILLER_0_8_153.VGND
rlabel metal1 186286 525667 187022 525763 5 dpga_flat_0.sr_0.FILLER_0_8_153.VPWR
flabel metal1 187042 526241 187095 526273 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_161.VGND
flabel metal1 187043 525698 187095 525729 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_161.VPWR
flabel nwell 187050 525706 187084 525724 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_161.VPB
flabel pwell 187053 526247 187085 526269 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_8_161.VNB
rlabel comment 187022 526259 187022 526259 2 dpga_flat_0.sr_0.FILLER_0_8_161.fill_2
rlabel metal1 187022 526211 187206 526307 5 dpga_flat_0.sr_0.FILLER_0_8_161.VGND
rlabel metal1 187022 525667 187206 525763 5 dpga_flat_0.sr_0.FILLER_0_8_161.VPWR
flabel metal1 187419 525698 187453 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_8_Right_8.VPWR
flabel metal1 187419 526242 187453 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_8_Right_8.VGND
flabel nwell 187419 525698 187453 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_8_Right_8.VPB
flabel pwell 187419 526242 187453 526276 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_8_Right_8.VNB
rlabel comment 187482 526259 187482 526259 8 dpga_flat_0.sr_0.PHY_EDGE_ROW_8_Right_8.decap_3
rlabel metal1 187206 526211 187482 526307 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_8_Right_8.VGND
rlabel metal1 187206 525667 187482 525763 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_8_Right_8.VPWR
flabel metal1 172515 525154 172549 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_3.VGND
flabel metal1 172515 525698 172549 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_3.VPWR
flabel nwell 172515 525698 172549 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_3.VPB
flabel pwell 172515 525154 172549 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_3.VNB
rlabel comment 172486 525171 172486 525171 4 dpga_flat_0.sr_0.FILLER_0_9_3.decap_12
flabel metal1 173619 525154 173653 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_15.VGND
flabel metal1 173619 525698 173653 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_15.VPWR
flabel nwell 173619 525698 173653 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_15.VPB
flabel pwell 173619 525154 173653 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_15.VNB
rlabel comment 173590 525171 173590 525171 4 dpga_flat_0.sr_0.FILLER_0_9_15.decap_12
flabel metal1 172239 525698 172273 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_9_Left_37.VPWR
flabel metal1 172239 525154 172273 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_9_Left_37.VGND
flabel nwell 172239 525698 172273 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_9_Left_37.VPB
flabel pwell 172239 525154 172273 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_9_Left_37.VNB
rlabel comment 172210 525171 172210 525171 4 dpga_flat_0.sr_0.PHY_EDGE_ROW_9_Left_37.decap_3
rlabel metal1 172210 525123 172486 525219 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_9_Left_37.VGND
rlabel metal1 172210 525667 172486 525763 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_9_Left_37.VPWR
flabel metal1 174723 525154 174757 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_27.VGND
flabel metal1 174723 525698 174757 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_27.VPWR
flabel nwell 174723 525698 174757 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_27.VPB
flabel pwell 174723 525154 174757 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_27.VNB
rlabel comment 174694 525171 174694 525171 4 dpga_flat_0.sr_0.FILLER_0_9_27.decap_12
flabel metal1 175827 525154 175861 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_39.VGND
flabel metal1 175827 525698 175861 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_39.VPWR
flabel nwell 175827 525698 175861 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_39.VPB
flabel pwell 175827 525154 175861 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_39.VNB
rlabel comment 175798 525171 175798 525171 4 dpga_flat_0.sr_0.FILLER_0_9_39.decap_12
flabel metal1 176931 525154 176965 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_51.VGND
flabel metal1 176931 525698 176965 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_51.VPWR
flabel nwell 176931 525698 176965 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_51.VPB
flabel pwell 176931 525154 176965 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_51.VNB
rlabel comment 176902 525171 176902 525171 4 dpga_flat_0.sr_0.FILLER_0_9_51.decap_4
rlabel metal1 176902 525123 177270 525219 1 dpga_flat_0.sr_0.FILLER_0_9_51.VGND
rlabel metal1 176902 525667 177270 525763 1 dpga_flat_0.sr_0.FILLER_0_9_51.VPWR
flabel metal1 177292 525698 177328 525728 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_55.VPWR
flabel metal1 177292 525158 177328 525187 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_55.VGND
flabel nwell 177301 525705 177321 525722 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_55.VPB
flabel pwell 177298 525160 177322 525182 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_55.VNB
rlabel comment 177270 525171 177270 525171 4 dpga_flat_0.sr_0.FILLER_0_9_55.fill_1
rlabel metal1 177270 525123 177362 525219 1 dpga_flat_0.sr_0.FILLER_0_9_55.VGND
rlabel metal1 177270 525667 177362 525763 1 dpga_flat_0.sr_0.FILLER_0_9_55.VPWR
flabel metal1 177483 525154 177517 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_57.VGND
flabel metal1 177483 525698 177517 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_57.VPWR
flabel nwell 177483 525698 177517 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_57.VPB
flabel pwell 177483 525154 177517 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_57.VNB
rlabel comment 177454 525171 177454 525171 4 dpga_flat_0.sr_0.FILLER_0_9_57.decap_12
flabel metal1 177384 525695 177437 525724 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_9_81.VPWR
flabel metal1 177383 525153 177434 525191 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_9_81.VGND
rlabel comment 177362 525171 177362 525171 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_9_81.tapvpwrvgnd_1
rlabel metal1 177362 525123 177454 525219 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_9_81.VGND
rlabel metal1 177362 525667 177454 525763 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_9_81.VPWR
flabel metal1 178587 525154 178621 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_69.VGND
flabel metal1 178587 525698 178621 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_69.VPWR
flabel nwell 178587 525698 178621 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_69.VPB
flabel pwell 178587 525154 178621 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_69.VNB
rlabel comment 178558 525171 178558 525171 4 dpga_flat_0.sr_0.FILLER_0_9_69.decap_12
flabel metal1 179691 525154 179725 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_81.VGND
flabel metal1 179691 525698 179725 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_81.VPWR
flabel nwell 179691 525698 179725 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_81.VPB
flabel pwell 179691 525154 179725 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_81.VNB
rlabel comment 179662 525171 179662 525171 4 dpga_flat_0.sr_0.FILLER_0_9_81.decap_12
flabel metal1 180795 525154 180829 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_93.VGND
flabel metal1 180795 525698 180829 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_93.VPWR
flabel nwell 180795 525698 180829 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_93.VPB
flabel pwell 180795 525154 180829 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_93.VNB
rlabel comment 180766 525171 180766 525171 4 dpga_flat_0.sr_0.FILLER_0_9_93.decap_12
flabel metal1 181899 525698 181933 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_105.VPWR
flabel metal1 181899 525154 181933 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_105.VGND
flabel nwell 181899 525698 181933 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_105.VPB
flabel pwell 181899 525154 181933 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_105.VNB
rlabel comment 181870 525171 181870 525171 4 dpga_flat_0.sr_0.FILLER_0_9_105.decap_6
rlabel metal1 181870 525123 182422 525219 1 dpga_flat_0.sr_0.FILLER_0_9_105.VGND
rlabel metal1 181870 525667 182422 525763 1 dpga_flat_0.sr_0.FILLER_0_9_105.VPWR
flabel metal1 182444 525698 182480 525728 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_111.VPWR
flabel metal1 182444 525158 182480 525187 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_111.VGND
flabel nwell 182453 525705 182473 525722 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_111.VPB
flabel pwell 182450 525160 182474 525182 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_111.VNB
rlabel comment 182422 525171 182422 525171 4 dpga_flat_0.sr_0.FILLER_0_9_111.fill_1
rlabel metal1 182422 525123 182514 525219 1 dpga_flat_0.sr_0.FILLER_0_9_111.VGND
rlabel metal1 182422 525667 182514 525763 1 dpga_flat_0.sr_0.FILLER_0_9_111.VPWR
flabel metal1 182635 525154 182669 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_113.VGND
flabel metal1 182635 525698 182669 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_113.VPWR
flabel nwell 182635 525698 182669 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_113.VPB
flabel pwell 182635 525154 182669 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_113.VNB
rlabel comment 182606 525171 182606 525171 4 dpga_flat_0.sr_0.FILLER_0_9_113.decap_12
flabel metal1 183739 525154 183773 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_125.VGND
flabel metal1 183739 525698 183773 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_125.VPWR
flabel nwell 183739 525698 183773 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_125.VPB
flabel pwell 183739 525154 183773 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_125.VNB
rlabel comment 183710 525171 183710 525171 4 dpga_flat_0.sr_0.FILLER_0_9_125.decap_12
flabel metal1 182536 525695 182589 525724 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_9_82.VPWR
flabel metal1 182535 525153 182586 525191 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_9_82.VGND
rlabel comment 182514 525171 182514 525171 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_9_82.tapvpwrvgnd_1
rlabel metal1 182514 525123 182606 525219 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_9_82.VGND
rlabel metal1 182514 525667 182606 525763 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_9_82.VPWR
flabel metal1 184843 525154 184877 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_137.VGND
flabel metal1 184843 525698 184877 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_137.VPWR
flabel nwell 184843 525698 184877 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_137.VPB
flabel pwell 184843 525154 184877 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_137.VNB
rlabel comment 184814 525171 184814 525171 4 dpga_flat_0.sr_0.FILLER_0_9_137.decap_12
flabel metal1 185947 525154 185981 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_149.VGND
flabel metal1 185947 525698 185981 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_149.VPWR
flabel nwell 185947 525698 185981 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_149.VPB
flabel pwell 185947 525154 185981 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_149.VNB
rlabel comment 185918 525171 185918 525171 4 dpga_flat_0.sr_0.FILLER_0_9_149.decap_12
flabel metal1 187042 525157 187095 525189 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_161.VGND
flabel metal1 187043 525701 187095 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_161.VPWR
flabel nwell 187050 525706 187084 525724 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_161.VPB
flabel pwell 187053 525161 187085 525183 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_9_161.VNB
rlabel comment 187022 525171 187022 525171 4 dpga_flat_0.sr_0.FILLER_0_9_161.fill_2
rlabel metal1 187022 525123 187206 525219 1 dpga_flat_0.sr_0.FILLER_0_9_161.VGND
rlabel metal1 187022 525667 187206 525763 1 dpga_flat_0.sr_0.FILLER_0_9_161.VPWR
flabel metal1 187419 525698 187453 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_9_Right_9.VPWR
flabel metal1 187419 525154 187453 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_9_Right_9.VGND
flabel nwell 187419 525698 187453 525732 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_9_Right_9.VPB
flabel pwell 187419 525154 187453 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_9_Right_9.VNB
rlabel comment 187482 525171 187482 525171 6 dpga_flat_0.sr_0.PHY_EDGE_ROW_9_Right_9.decap_3
rlabel metal1 187206 525123 187482 525219 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_9_Right_9.VGND
rlabel metal1 187206 525667 187482 525763 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_9_Right_9.VPWR
flabel metal1 172515 525154 172549 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_3.VGND
flabel metal1 172515 524610 172549 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_3.VPWR
flabel nwell 172515 524610 172549 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_3.VPB
flabel pwell 172515 525154 172549 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_3.VNB
rlabel comment 172486 525171 172486 525171 2 dpga_flat_0.sr_0.FILLER_0_10_3.decap_12
flabel metal1 173619 525154 173653 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_15.VGND
flabel metal1 173619 524610 173653 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_15.VPWR
flabel nwell 173619 524610 173653 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_15.VPB
flabel pwell 173619 525154 173653 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_15.VNB
rlabel comment 173590 525171 173590 525171 2 dpga_flat_0.sr_0.FILLER_0_10_15.decap_12
flabel metal1 172239 524610 172273 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_10_Left_38.VPWR
flabel metal1 172239 525154 172273 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_10_Left_38.VGND
flabel nwell 172239 524610 172273 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_10_Left_38.VPB
flabel pwell 172239 525154 172273 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_10_Left_38.VNB
rlabel comment 172210 525171 172210 525171 2 dpga_flat_0.sr_0.PHY_EDGE_ROW_10_Left_38.decap_3
rlabel metal1 172210 525123 172486 525219 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_10_Left_38.VGND
rlabel metal1 172210 524579 172486 524675 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_10_Left_38.VPWR
flabel metal1 174716 524614 174752 524644 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_27.VPWR
flabel metal1 174716 525155 174752 525184 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_27.VGND
flabel nwell 174725 524620 174745 524637 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_27.VPB
flabel pwell 174722 525160 174746 525182 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_27.VNB
rlabel comment 174694 525171 174694 525171 2 dpga_flat_0.sr_0.FILLER_0_10_27.fill_1
rlabel metal1 174694 525123 174786 525219 5 dpga_flat_0.sr_0.FILLER_0_10_27.VGND
rlabel metal1 174694 524579 174786 524675 5 dpga_flat_0.sr_0.FILLER_0_10_27.VPWR
flabel metal1 174907 525154 174941 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_29.VGND
flabel metal1 174907 524610 174941 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_29.VPWR
flabel nwell 174907 524610 174941 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_29.VPB
flabel pwell 174907 525154 174941 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_29.VNB
rlabel comment 174878 525171 174878 525171 2 dpga_flat_0.sr_0.FILLER_0_10_29.decap_12
flabel metal1 176011 525154 176045 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_41.VGND
flabel metal1 176011 524610 176045 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_41.VPWR
flabel nwell 176011 524610 176045 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_41.VPB
flabel pwell 176011 525154 176045 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_41.VNB
rlabel comment 175982 525171 175982 525171 2 dpga_flat_0.sr_0.FILLER_0_10_41.decap_12
flabel metal1 174808 524618 174861 524647 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_10_83.VPWR
flabel metal1 174807 525151 174858 525189 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_10_83.VGND
rlabel comment 174786 525171 174786 525171 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_10_83.tapvpwrvgnd_1
rlabel metal1 174786 525123 174878 525219 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_10_83.VGND
rlabel metal1 174786 524579 174878 524675 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_10_83.VPWR
flabel metal1 177115 525154 177149 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_53.VGND
flabel metal1 177115 524610 177149 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_53.VPWR
flabel nwell 177115 524610 177149 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_53.VPB
flabel pwell 177115 525154 177149 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_53.VNB
rlabel comment 177086 525171 177086 525171 2 dpga_flat_0.sr_0.FILLER_0_10_53.decap_12
flabel metal1 178219 525154 178253 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_65.VGND
flabel metal1 178219 524610 178253 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_65.VPWR
flabel nwell 178219 524610 178253 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_65.VPB
flabel pwell 178219 525154 178253 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_65.VNB
rlabel comment 178190 525171 178190 525171 2 dpga_flat_0.sr_0.FILLER_0_10_65.decap_12
flabel metal1 179323 524610 179357 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_77.VPWR
flabel metal1 179323 525154 179357 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_77.VGND
flabel nwell 179323 524610 179357 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_77.VPB
flabel pwell 179323 525154 179357 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_77.VNB
rlabel comment 179294 525171 179294 525171 2 dpga_flat_0.sr_0.FILLER_0_10_77.decap_6
rlabel metal1 179294 525123 179846 525219 5 dpga_flat_0.sr_0.FILLER_0_10_77.VGND
rlabel metal1 179294 524579 179846 524675 5 dpga_flat_0.sr_0.FILLER_0_10_77.VPWR
flabel metal1 179868 524614 179904 524644 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_83.VPWR
flabel metal1 179868 525155 179904 525184 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_83.VGND
flabel nwell 179877 524620 179897 524637 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_83.VPB
flabel pwell 179874 525160 179898 525182 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_83.VNB
rlabel comment 179846 525171 179846 525171 2 dpga_flat_0.sr_0.FILLER_0_10_83.fill_1
rlabel metal1 179846 525123 179938 525219 5 dpga_flat_0.sr_0.FILLER_0_10_83.VGND
rlabel metal1 179846 524579 179938 524675 5 dpga_flat_0.sr_0.FILLER_0_10_83.VPWR
flabel metal1 180059 525154 180093 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_85.VGND
flabel metal1 180059 524610 180093 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_85.VPWR
flabel nwell 180059 524610 180093 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_85.VPB
flabel pwell 180059 525154 180093 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_85.VNB
rlabel comment 180030 525171 180030 525171 2 dpga_flat_0.sr_0.FILLER_0_10_85.decap_12
flabel metal1 181163 525154 181197 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_97.VGND
flabel metal1 181163 524610 181197 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_97.VPWR
flabel nwell 181163 524610 181197 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_97.VPB
flabel pwell 181163 525154 181197 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_97.VNB
rlabel comment 181134 525171 181134 525171 2 dpga_flat_0.sr_0.FILLER_0_10_97.decap_12
flabel metal1 179960 524618 180013 524647 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_10_84.VPWR
flabel metal1 179959 525151 180010 525189 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_10_84.VGND
rlabel comment 179938 525171 179938 525171 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_10_84.tapvpwrvgnd_1
rlabel metal1 179938 525123 180030 525219 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_10_84.VGND
rlabel metal1 179938 524579 180030 524675 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_10_84.VPWR
flabel metal1 182267 525154 182301 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_109.VGND
flabel metal1 182267 524610 182301 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_109.VPWR
flabel nwell 182267 524610 182301 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_109.VPB
flabel pwell 182267 525154 182301 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_109.VNB
rlabel comment 182238 525171 182238 525171 2 dpga_flat_0.sr_0.FILLER_0_10_109.decap_12
flabel metal1 183371 525154 183405 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_121.VGND
flabel metal1 183371 524610 183405 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_121.VPWR
flabel nwell 183371 524610 183405 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_121.VPB
flabel pwell 183371 525154 183405 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_121.VNB
rlabel comment 183342 525171 183342 525171 2 dpga_flat_0.sr_0.FILLER_0_10_121.decap_12
flabel metal1 184475 524610 184509 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_133.VPWR
flabel metal1 184475 525154 184509 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_133.VGND
flabel nwell 184475 524610 184509 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_133.VPB
flabel pwell 184475 525154 184509 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_133.VNB
rlabel comment 184446 525171 184446 525171 2 dpga_flat_0.sr_0.FILLER_0_10_133.decap_6
rlabel metal1 184446 525123 184998 525219 5 dpga_flat_0.sr_0.FILLER_0_10_133.VGND
rlabel metal1 184446 524579 184998 524675 5 dpga_flat_0.sr_0.FILLER_0_10_133.VPWR
flabel metal1 185020 524614 185056 524644 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_139.VPWR
flabel metal1 185020 525155 185056 525184 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_139.VGND
flabel nwell 185029 524620 185049 524637 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_139.VPB
flabel pwell 185026 525160 185050 525182 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_139.VNB
rlabel comment 184998 525171 184998 525171 2 dpga_flat_0.sr_0.FILLER_0_10_139.fill_1
rlabel metal1 184998 525123 185090 525219 5 dpga_flat_0.sr_0.FILLER_0_10_139.VGND
rlabel metal1 184998 524579 185090 524675 5 dpga_flat_0.sr_0.FILLER_0_10_139.VPWR
flabel metal1 185211 525154 185245 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_141.VGND
flabel metal1 185211 524610 185245 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_141.VPWR
flabel nwell 185211 524610 185245 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_141.VPB
flabel pwell 185211 525154 185245 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_141.VNB
rlabel comment 185182 525171 185182 525171 2 dpga_flat_0.sr_0.FILLER_0_10_141.decap_12
flabel metal1 185112 524618 185165 524647 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_10_85.VPWR
flabel metal1 185111 525151 185162 525189 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_10_85.VGND
rlabel comment 185090 525171 185090 525171 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_10_85.tapvpwrvgnd_1
rlabel metal1 185090 525123 185182 525219 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_10_85.VGND
rlabel metal1 185090 524579 185182 524675 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_10_85.VPWR
flabel metal1 186315 524610 186349 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_153.VPWR
flabel metal1 186315 525154 186349 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_153.VGND
flabel nwell 186315 524610 186349 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_153.VPB
flabel pwell 186315 525154 186349 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_153.VNB
rlabel comment 186286 525171 186286 525171 2 dpga_flat_0.sr_0.FILLER_0_10_153.decap_8
rlabel metal1 186286 525123 187022 525219 5 dpga_flat_0.sr_0.FILLER_0_10_153.VGND
rlabel metal1 186286 524579 187022 524675 5 dpga_flat_0.sr_0.FILLER_0_10_153.VPWR
flabel metal1 187042 525153 187095 525185 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_161.VGND
flabel metal1 187043 524610 187095 524641 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_161.VPWR
flabel nwell 187050 524618 187084 524636 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_161.VPB
flabel pwell 187053 525159 187085 525181 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_10_161.VNB
rlabel comment 187022 525171 187022 525171 2 dpga_flat_0.sr_0.FILLER_0_10_161.fill_2
rlabel metal1 187022 525123 187206 525219 5 dpga_flat_0.sr_0.FILLER_0_10_161.VGND
rlabel metal1 187022 524579 187206 524675 5 dpga_flat_0.sr_0.FILLER_0_10_161.VPWR
flabel metal1 187419 524610 187453 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_10_Right_10.VPWR
flabel metal1 187419 525154 187453 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_10_Right_10.VGND
flabel nwell 187419 524610 187453 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_10_Right_10.VPB
flabel pwell 187419 525154 187453 525188 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_10_Right_10.VNB
rlabel comment 187482 525171 187482 525171 8 dpga_flat_0.sr_0.PHY_EDGE_ROW_10_Right_10.decap_3
rlabel metal1 187206 525123 187482 525219 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_10_Right_10.VGND
rlabel metal1 187206 524579 187482 524675 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_10_Right_10.VPWR
flabel metal1 172515 524066 172549 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_3.VGND
flabel metal1 172515 524610 172549 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_3.VPWR
flabel nwell 172515 524610 172549 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_3.VPB
flabel pwell 172515 524066 172549 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_3.VNB
rlabel comment 172486 524083 172486 524083 4 dpga_flat_0.sr_0.FILLER_0_11_3.decap_12
flabel metal1 173619 524066 173653 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_15.VGND
flabel metal1 173619 524610 173653 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_15.VPWR
flabel nwell 173619 524610 173653 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_15.VPB
flabel pwell 173619 524066 173653 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_15.VNB
rlabel comment 173590 524083 173590 524083 4 dpga_flat_0.sr_0.FILLER_0_11_15.decap_12
flabel metal1 172239 524610 172273 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_11_Left_39.VPWR
flabel metal1 172239 524066 172273 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_11_Left_39.VGND
flabel nwell 172239 524610 172273 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_11_Left_39.VPB
flabel pwell 172239 524066 172273 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_11_Left_39.VNB
rlabel comment 172210 524083 172210 524083 4 dpga_flat_0.sr_0.PHY_EDGE_ROW_11_Left_39.decap_3
rlabel metal1 172210 524035 172486 524131 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_11_Left_39.VGND
rlabel metal1 172210 524579 172486 524675 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_11_Left_39.VPWR
flabel metal1 174723 524066 174757 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_27.VGND
flabel metal1 174723 524610 174757 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_27.VPWR
flabel nwell 174723 524610 174757 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_27.VPB
flabel pwell 174723 524066 174757 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_27.VNB
rlabel comment 174694 524083 174694 524083 4 dpga_flat_0.sr_0.FILLER_0_11_27.decap_12
flabel metal1 175827 524066 175861 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_39.VGND
flabel metal1 175827 524610 175861 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_39.VPWR
flabel nwell 175827 524610 175861 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_39.VPB
flabel pwell 175827 524066 175861 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_39.VNB
rlabel comment 175798 524083 175798 524083 4 dpga_flat_0.sr_0.FILLER_0_11_39.decap_12
flabel metal1 176931 524066 176965 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_51.VGND
flabel metal1 176931 524610 176965 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_51.VPWR
flabel nwell 176931 524610 176965 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_51.VPB
flabel pwell 176931 524066 176965 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_51.VNB
rlabel comment 176902 524083 176902 524083 4 dpga_flat_0.sr_0.FILLER_0_11_51.decap_4
rlabel metal1 176902 524035 177270 524131 1 dpga_flat_0.sr_0.FILLER_0_11_51.VGND
rlabel metal1 176902 524579 177270 524675 1 dpga_flat_0.sr_0.FILLER_0_11_51.VPWR
flabel metal1 177292 524610 177328 524640 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_55.VPWR
flabel metal1 177292 524070 177328 524099 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_55.VGND
flabel nwell 177301 524617 177321 524634 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_55.VPB
flabel pwell 177298 524072 177322 524094 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_55.VNB
rlabel comment 177270 524083 177270 524083 4 dpga_flat_0.sr_0.FILLER_0_11_55.fill_1
rlabel metal1 177270 524035 177362 524131 1 dpga_flat_0.sr_0.FILLER_0_11_55.VGND
rlabel metal1 177270 524579 177362 524675 1 dpga_flat_0.sr_0.FILLER_0_11_55.VPWR
flabel metal1 177483 524066 177517 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_57.VGND
flabel metal1 177483 524610 177517 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_57.VPWR
flabel nwell 177483 524610 177517 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_57.VPB
flabel pwell 177483 524066 177517 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_57.VNB
rlabel comment 177454 524083 177454 524083 4 dpga_flat_0.sr_0.FILLER_0_11_57.decap_12
flabel metal1 177384 524607 177437 524636 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_11_86.VPWR
flabel metal1 177383 524065 177434 524103 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_11_86.VGND
rlabel comment 177362 524083 177362 524083 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_11_86.tapvpwrvgnd_1
rlabel metal1 177362 524035 177454 524131 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_11_86.VGND
rlabel metal1 177362 524579 177454 524675 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_11_86.VPWR
flabel metal1 178587 524066 178621 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_69.VGND
flabel metal1 178587 524610 178621 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_69.VPWR
flabel nwell 178587 524610 178621 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_69.VPB
flabel pwell 178587 524066 178621 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_69.VNB
rlabel comment 178558 524083 178558 524083 4 dpga_flat_0.sr_0.FILLER_0_11_69.decap_12
flabel metal1 179691 524066 179725 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_81.VGND
flabel metal1 179691 524610 179725 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_81.VPWR
flabel nwell 179691 524610 179725 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_81.VPB
flabel pwell 179691 524066 179725 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_81.VNB
rlabel comment 179662 524083 179662 524083 4 dpga_flat_0.sr_0.FILLER_0_11_81.decap_12
flabel metal1 180795 524066 180829 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_93.VGND
flabel metal1 180795 524610 180829 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_93.VPWR
flabel nwell 180795 524610 180829 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_93.VPB
flabel pwell 180795 524066 180829 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_93.VNB
rlabel comment 180766 524083 180766 524083 4 dpga_flat_0.sr_0.FILLER_0_11_93.decap_12
flabel metal1 181899 524610 181933 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_105.VPWR
flabel metal1 181899 524066 181933 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_105.VGND
flabel nwell 181899 524610 181933 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_105.VPB
flabel pwell 181899 524066 181933 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_105.VNB
rlabel comment 181870 524083 181870 524083 4 dpga_flat_0.sr_0.FILLER_0_11_105.decap_6
rlabel metal1 181870 524035 182422 524131 1 dpga_flat_0.sr_0.FILLER_0_11_105.VGND
rlabel metal1 181870 524579 182422 524675 1 dpga_flat_0.sr_0.FILLER_0_11_105.VPWR
flabel metal1 182444 524610 182480 524640 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_111.VPWR
flabel metal1 182444 524070 182480 524099 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_111.VGND
flabel nwell 182453 524617 182473 524634 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_111.VPB
flabel pwell 182450 524072 182474 524094 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_111.VNB
rlabel comment 182422 524083 182422 524083 4 dpga_flat_0.sr_0.FILLER_0_11_111.fill_1
rlabel metal1 182422 524035 182514 524131 1 dpga_flat_0.sr_0.FILLER_0_11_111.VGND
rlabel metal1 182422 524579 182514 524675 1 dpga_flat_0.sr_0.FILLER_0_11_111.VPWR
flabel metal1 182635 524066 182669 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_113.VGND
flabel metal1 182635 524610 182669 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_113.VPWR
flabel nwell 182635 524610 182669 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_113.VPB
flabel pwell 182635 524066 182669 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_113.VNB
rlabel comment 182606 524083 182606 524083 4 dpga_flat_0.sr_0.FILLER_0_11_113.decap_12
flabel metal1 183739 524066 183773 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_125.VGND
flabel metal1 183739 524610 183773 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_125.VPWR
flabel nwell 183739 524610 183773 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_125.VPB
flabel pwell 183739 524066 183773 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_125.VNB
rlabel comment 183710 524083 183710 524083 4 dpga_flat_0.sr_0.FILLER_0_11_125.decap_12
flabel metal1 182536 524607 182589 524636 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_11_87.VPWR
flabel metal1 182535 524065 182586 524103 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_11_87.VGND
rlabel comment 182514 524083 182514 524083 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_11_87.tapvpwrvgnd_1
rlabel metal1 182514 524035 182606 524131 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_11_87.VGND
rlabel metal1 182514 524579 182606 524675 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_11_87.VPWR
flabel metal1 184843 524066 184877 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_137.VGND
flabel metal1 184843 524610 184877 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_137.VPWR
flabel nwell 184843 524610 184877 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_137.VPB
flabel pwell 184843 524066 184877 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_137.VNB
rlabel comment 184814 524083 184814 524083 4 dpga_flat_0.sr_0.FILLER_0_11_137.decap_12
flabel metal1 185947 524066 185981 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_149.VGND
flabel metal1 185947 524610 185981 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_149.VPWR
flabel nwell 185947 524610 185981 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_149.VPB
flabel pwell 185947 524066 185981 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_149.VNB
rlabel comment 185918 524083 185918 524083 4 dpga_flat_0.sr_0.FILLER_0_11_149.decap_12
flabel metal1 187042 524069 187095 524101 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_161.VGND
flabel metal1 187043 524613 187095 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_161.VPWR
flabel nwell 187050 524618 187084 524636 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_161.VPB
flabel pwell 187053 524073 187085 524095 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_11_161.VNB
rlabel comment 187022 524083 187022 524083 4 dpga_flat_0.sr_0.FILLER_0_11_161.fill_2
rlabel metal1 187022 524035 187206 524131 1 dpga_flat_0.sr_0.FILLER_0_11_161.VGND
rlabel metal1 187022 524579 187206 524675 1 dpga_flat_0.sr_0.FILLER_0_11_161.VPWR
flabel metal1 187419 524610 187453 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_11_Right_11.VPWR
flabel metal1 187419 524066 187453 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_11_Right_11.VGND
flabel nwell 187419 524610 187453 524644 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_11_Right_11.VPB
flabel pwell 187419 524066 187453 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_11_Right_11.VNB
rlabel comment 187482 524083 187482 524083 6 dpga_flat_0.sr_0.PHY_EDGE_ROW_11_Right_11.decap_3
rlabel metal1 187206 524035 187482 524131 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_11_Right_11.VGND
rlabel metal1 187206 524579 187482 524675 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_11_Right_11.VPWR
flabel metal1 172515 524066 172549 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_3.VGND
flabel metal1 172515 523522 172549 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_3.VPWR
flabel nwell 172515 523522 172549 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_3.VPB
flabel pwell 172515 524066 172549 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_3.VNB
rlabel comment 172486 524083 172486 524083 2 dpga_flat_0.sr_0.FILLER_0_12_3.decap_12
flabel metal1 173619 524066 173653 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_15.VGND
flabel metal1 173619 523522 173653 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_15.VPWR
flabel nwell 173619 523522 173653 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_15.VPB
flabel pwell 173619 524066 173653 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_15.VNB
rlabel comment 173590 524083 173590 524083 2 dpga_flat_0.sr_0.FILLER_0_12_15.decap_12
flabel metal1 172239 523522 172273 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_12_Left_40.VPWR
flabel metal1 172239 524066 172273 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_12_Left_40.VGND
flabel nwell 172239 523522 172273 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_12_Left_40.VPB
flabel pwell 172239 524066 172273 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_12_Left_40.VNB
rlabel comment 172210 524083 172210 524083 2 dpga_flat_0.sr_0.PHY_EDGE_ROW_12_Left_40.decap_3
rlabel metal1 172210 524035 172486 524131 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_12_Left_40.VGND
rlabel metal1 172210 523491 172486 523587 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_12_Left_40.VPWR
flabel metal1 174716 523526 174752 523556 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_27.VPWR
flabel metal1 174716 524067 174752 524096 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_27.VGND
flabel nwell 174725 523532 174745 523549 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_27.VPB
flabel pwell 174722 524072 174746 524094 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_27.VNB
rlabel comment 174694 524083 174694 524083 2 dpga_flat_0.sr_0.FILLER_0_12_27.fill_1
rlabel metal1 174694 524035 174786 524131 5 dpga_flat_0.sr_0.FILLER_0_12_27.VGND
rlabel metal1 174694 523491 174786 523587 5 dpga_flat_0.sr_0.FILLER_0_12_27.VPWR
flabel metal1 174907 524066 174941 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_29.VGND
flabel metal1 174907 523522 174941 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_29.VPWR
flabel nwell 174907 523522 174941 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_29.VPB
flabel pwell 174907 524066 174941 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_29.VNB
rlabel comment 174878 524083 174878 524083 2 dpga_flat_0.sr_0.FILLER_0_12_29.decap_12
flabel metal1 176011 524066 176045 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_41.VGND
flabel metal1 176011 523522 176045 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_41.VPWR
flabel nwell 176011 523522 176045 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_41.VPB
flabel pwell 176011 524066 176045 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_41.VNB
rlabel comment 175982 524083 175982 524083 2 dpga_flat_0.sr_0.FILLER_0_12_41.decap_12
flabel metal1 174808 523530 174861 523559 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_12_88.VPWR
flabel metal1 174807 524063 174858 524101 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_12_88.VGND
rlabel comment 174786 524083 174786 524083 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_12_88.tapvpwrvgnd_1
rlabel metal1 174786 524035 174878 524131 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_12_88.VGND
rlabel metal1 174786 523491 174878 523587 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_12_88.VPWR
flabel metal1 177115 524066 177149 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_53.VGND
flabel metal1 177115 523522 177149 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_53.VPWR
flabel nwell 177115 523522 177149 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_53.VPB
flabel pwell 177115 524066 177149 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_53.VNB
rlabel comment 177086 524083 177086 524083 2 dpga_flat_0.sr_0.FILLER_0_12_53.decap_12
flabel metal1 178219 524066 178253 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_65.VGND
flabel metal1 178219 523522 178253 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_65.VPWR
flabel nwell 178219 523522 178253 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_65.VPB
flabel pwell 178219 524066 178253 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_65.VNB
rlabel comment 178190 524083 178190 524083 2 dpga_flat_0.sr_0.FILLER_0_12_65.decap_12
flabel metal1 179323 523522 179357 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_77.VPWR
flabel metal1 179323 524066 179357 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_77.VGND
flabel nwell 179323 523522 179357 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_77.VPB
flabel pwell 179323 524066 179357 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_77.VNB
rlabel comment 179294 524083 179294 524083 2 dpga_flat_0.sr_0.FILLER_0_12_77.decap_6
rlabel metal1 179294 524035 179846 524131 5 dpga_flat_0.sr_0.FILLER_0_12_77.VGND
rlabel metal1 179294 523491 179846 523587 5 dpga_flat_0.sr_0.FILLER_0_12_77.VPWR
flabel metal1 179868 523526 179904 523556 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_83.VPWR
flabel metal1 179868 524067 179904 524096 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_83.VGND
flabel nwell 179877 523532 179897 523549 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_83.VPB
flabel pwell 179874 524072 179898 524094 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_83.VNB
rlabel comment 179846 524083 179846 524083 2 dpga_flat_0.sr_0.FILLER_0_12_83.fill_1
rlabel metal1 179846 524035 179938 524131 5 dpga_flat_0.sr_0.FILLER_0_12_83.VGND
rlabel metal1 179846 523491 179938 523587 5 dpga_flat_0.sr_0.FILLER_0_12_83.VPWR
flabel metal1 180059 524066 180093 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_85.VGND
flabel metal1 180059 523522 180093 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_85.VPWR
flabel nwell 180059 523522 180093 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_85.VPB
flabel pwell 180059 524066 180093 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_85.VNB
rlabel comment 180030 524083 180030 524083 2 dpga_flat_0.sr_0.FILLER_0_12_85.decap_12
flabel metal1 181163 524066 181197 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_97.VGND
flabel metal1 181163 523522 181197 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_97.VPWR
flabel nwell 181163 523522 181197 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_97.VPB
flabel pwell 181163 524066 181197 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_97.VNB
rlabel comment 181134 524083 181134 524083 2 dpga_flat_0.sr_0.FILLER_0_12_97.decap_12
flabel metal1 179960 523530 180013 523559 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_12_89.VPWR
flabel metal1 179959 524063 180010 524101 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_12_89.VGND
rlabel comment 179938 524083 179938 524083 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_12_89.tapvpwrvgnd_1
rlabel metal1 179938 524035 180030 524131 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_12_89.VGND
rlabel metal1 179938 523491 180030 523587 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_12_89.VPWR
flabel metal1 182267 524066 182301 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_109.VGND
flabel metal1 182267 523522 182301 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_109.VPWR
flabel nwell 182267 523522 182301 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_109.VPB
flabel pwell 182267 524066 182301 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_109.VNB
rlabel comment 182238 524083 182238 524083 2 dpga_flat_0.sr_0.FILLER_0_12_109.decap_12
flabel metal1 183371 524066 183405 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_121.VGND
flabel metal1 183371 523522 183405 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_121.VPWR
flabel nwell 183371 523522 183405 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_121.VPB
flabel pwell 183371 524066 183405 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_121.VNB
rlabel comment 183342 524083 183342 524083 2 dpga_flat_0.sr_0.FILLER_0_12_121.decap_12
flabel metal1 184475 523522 184509 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_133.VPWR
flabel metal1 184475 524066 184509 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_133.VGND
flabel nwell 184475 523522 184509 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_133.VPB
flabel pwell 184475 524066 184509 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_133.VNB
rlabel comment 184446 524083 184446 524083 2 dpga_flat_0.sr_0.FILLER_0_12_133.decap_6
rlabel metal1 184446 524035 184998 524131 5 dpga_flat_0.sr_0.FILLER_0_12_133.VGND
rlabel metal1 184446 523491 184998 523587 5 dpga_flat_0.sr_0.FILLER_0_12_133.VPWR
flabel metal1 185020 523526 185056 523556 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_139.VPWR
flabel metal1 185020 524067 185056 524096 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_139.VGND
flabel nwell 185029 523532 185049 523549 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_139.VPB
flabel pwell 185026 524072 185050 524094 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_139.VNB
rlabel comment 184998 524083 184998 524083 2 dpga_flat_0.sr_0.FILLER_0_12_139.fill_1
rlabel metal1 184998 524035 185090 524131 5 dpga_flat_0.sr_0.FILLER_0_12_139.VGND
rlabel metal1 184998 523491 185090 523587 5 dpga_flat_0.sr_0.FILLER_0_12_139.VPWR
flabel metal1 185211 524066 185245 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_141.VGND
flabel metal1 185211 523522 185245 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_141.VPWR
flabel nwell 185211 523522 185245 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_141.VPB
flabel pwell 185211 524066 185245 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_141.VNB
rlabel comment 185182 524083 185182 524083 2 dpga_flat_0.sr_0.FILLER_0_12_141.decap_12
flabel metal1 185112 523530 185165 523559 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_12_90.VPWR
flabel metal1 185111 524063 185162 524101 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_12_90.VGND
rlabel comment 185090 524083 185090 524083 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_12_90.tapvpwrvgnd_1
rlabel metal1 185090 524035 185182 524131 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_12_90.VGND
rlabel metal1 185090 523491 185182 523587 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_12_90.VPWR
flabel metal1 186315 523522 186349 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_153.VPWR
flabel metal1 186315 524066 186349 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_153.VGND
flabel nwell 186315 523522 186349 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_153.VPB
flabel pwell 186315 524066 186349 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_153.VNB
rlabel comment 186286 524083 186286 524083 2 dpga_flat_0.sr_0.FILLER_0_12_153.decap_8
rlabel metal1 186286 524035 187022 524131 5 dpga_flat_0.sr_0.FILLER_0_12_153.VGND
rlabel metal1 186286 523491 187022 523587 5 dpga_flat_0.sr_0.FILLER_0_12_153.VPWR
flabel metal1 187042 524065 187095 524097 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_161.VGND
flabel metal1 187043 523522 187095 523553 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_161.VPWR
flabel nwell 187050 523530 187084 523548 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_161.VPB
flabel pwell 187053 524071 187085 524093 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_12_161.VNB
rlabel comment 187022 524083 187022 524083 2 dpga_flat_0.sr_0.FILLER_0_12_161.fill_2
rlabel metal1 187022 524035 187206 524131 5 dpga_flat_0.sr_0.FILLER_0_12_161.VGND
rlabel metal1 187022 523491 187206 523587 5 dpga_flat_0.sr_0.FILLER_0_12_161.VPWR
flabel metal1 187419 523522 187453 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_12_Right_12.VPWR
flabel metal1 187419 524066 187453 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_12_Right_12.VGND
flabel nwell 187419 523522 187453 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_12_Right_12.VPB
flabel pwell 187419 524066 187453 524100 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_12_Right_12.VNB
rlabel comment 187482 524083 187482 524083 8 dpga_flat_0.sr_0.PHY_EDGE_ROW_12_Right_12.decap_3
rlabel metal1 187206 524035 187482 524131 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_12_Right_12.VGND
rlabel metal1 187206 523491 187482 523587 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_12_Right_12.VPWR
flabel metal1 172515 522978 172549 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_3.VGND
flabel metal1 172515 523522 172549 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_3.VPWR
flabel nwell 172515 523522 172549 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_3.VPB
flabel pwell 172515 522978 172549 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_3.VNB
rlabel comment 172486 522995 172486 522995 4 dpga_flat_0.sr_0.FILLER_0_13_3.decap_12
flabel metal1 173619 522978 173653 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_15.VGND
flabel metal1 173619 523522 173653 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_15.VPWR
flabel nwell 173619 523522 173653 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_15.VPB
flabel pwell 173619 522978 173653 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_15.VNB
rlabel comment 173590 522995 173590 522995 4 dpga_flat_0.sr_0.FILLER_0_13_15.decap_12
flabel metal1 172515 522978 172549 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_3.VGND
flabel metal1 172515 522434 172549 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_3.VPWR
flabel nwell 172515 522434 172549 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_3.VPB
flabel pwell 172515 522978 172549 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_3.VNB
rlabel comment 172486 522995 172486 522995 2 dpga_flat_0.sr_0.FILLER_0_14_3.decap_12
flabel metal1 173619 522978 173653 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_15.VGND
flabel metal1 173619 522434 173653 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_15.VPWR
flabel nwell 173619 522434 173653 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_15.VPB
flabel pwell 173619 522978 173653 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_15.VNB
rlabel comment 173590 522995 173590 522995 2 dpga_flat_0.sr_0.FILLER_0_14_15.decap_12
flabel metal1 172239 523522 172273 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_13_Left_41.VPWR
flabel metal1 172239 522978 172273 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_13_Left_41.VGND
flabel nwell 172239 523522 172273 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_13_Left_41.VPB
flabel pwell 172239 522978 172273 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_13_Left_41.VNB
rlabel comment 172210 522995 172210 522995 4 dpga_flat_0.sr_0.PHY_EDGE_ROW_13_Left_41.decap_3
rlabel metal1 172210 522947 172486 523043 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_13_Left_41.VGND
rlabel metal1 172210 523491 172486 523587 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_13_Left_41.VPWR
flabel metal1 172239 522434 172273 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_14_Left_42.VPWR
flabel metal1 172239 522978 172273 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_14_Left_42.VGND
flabel nwell 172239 522434 172273 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_14_Left_42.VPB
flabel pwell 172239 522978 172273 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_14_Left_42.VNB
rlabel comment 172210 522995 172210 522995 2 dpga_flat_0.sr_0.PHY_EDGE_ROW_14_Left_42.decap_3
rlabel metal1 172210 522947 172486 523043 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_14_Left_42.VGND
rlabel metal1 172210 522403 172486 522499 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_14_Left_42.VPWR
flabel metal1 174723 522978 174757 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_27.VGND
flabel metal1 174723 523522 174757 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_27.VPWR
flabel nwell 174723 523522 174757 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_27.VPB
flabel pwell 174723 522978 174757 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_27.VNB
rlabel comment 174694 522995 174694 522995 4 dpga_flat_0.sr_0.FILLER_0_13_27.decap_12
flabel metal1 175827 522978 175861 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_39.VGND
flabel metal1 175827 523522 175861 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_39.VPWR
flabel nwell 175827 523522 175861 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_39.VPB
flabel pwell 175827 522978 175861 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_39.VNB
rlabel comment 175798 522995 175798 522995 4 dpga_flat_0.sr_0.FILLER_0_13_39.decap_12
flabel metal1 174716 522438 174752 522468 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_27.VPWR
flabel metal1 174716 522979 174752 523008 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_27.VGND
flabel nwell 174725 522444 174745 522461 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_27.VPB
flabel pwell 174722 522984 174746 523006 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_27.VNB
rlabel comment 174694 522995 174694 522995 2 dpga_flat_0.sr_0.FILLER_0_14_27.fill_1
rlabel metal1 174694 522947 174786 523043 5 dpga_flat_0.sr_0.FILLER_0_14_27.VGND
rlabel metal1 174694 522403 174786 522499 5 dpga_flat_0.sr_0.FILLER_0_14_27.VPWR
flabel metal1 174907 522978 174941 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_29.VGND
flabel metal1 174907 522434 174941 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_29.VPWR
flabel nwell 174907 522434 174941 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_29.VPB
flabel pwell 174907 522978 174941 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_29.VNB
rlabel comment 174878 522995 174878 522995 2 dpga_flat_0.sr_0.FILLER_0_14_29.decap_12
flabel metal1 176011 522978 176045 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_41.VGND
flabel metal1 176011 522434 176045 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_41.VPWR
flabel nwell 176011 522434 176045 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_41.VPB
flabel pwell 176011 522978 176045 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_41.VNB
rlabel comment 175982 522995 175982 522995 2 dpga_flat_0.sr_0.FILLER_0_14_41.decap_12
flabel metal1 174808 522442 174861 522471 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_14_93.VPWR
flabel metal1 174807 522975 174858 523013 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_14_93.VGND
rlabel comment 174786 522995 174786 522995 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_14_93.tapvpwrvgnd_1
rlabel metal1 174786 522947 174878 523043 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_14_93.VGND
rlabel metal1 174786 522403 174878 522499 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_14_93.VPWR
flabel metal1 176931 522978 176965 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_51.VGND
flabel metal1 176931 523522 176965 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_51.VPWR
flabel nwell 176931 523522 176965 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_51.VPB
flabel pwell 176931 522978 176965 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_51.VNB
rlabel comment 176902 522995 176902 522995 4 dpga_flat_0.sr_0.FILLER_0_13_51.decap_4
rlabel metal1 176902 522947 177270 523043 1 dpga_flat_0.sr_0.FILLER_0_13_51.VGND
rlabel metal1 176902 523491 177270 523587 1 dpga_flat_0.sr_0.FILLER_0_13_51.VPWR
flabel metal1 177292 523522 177328 523552 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_55.VPWR
flabel metal1 177292 522982 177328 523011 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_55.VGND
flabel nwell 177301 523529 177321 523546 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_55.VPB
flabel pwell 177298 522984 177322 523006 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_55.VNB
rlabel comment 177270 522995 177270 522995 4 dpga_flat_0.sr_0.FILLER_0_13_55.fill_1
rlabel metal1 177270 522947 177362 523043 1 dpga_flat_0.sr_0.FILLER_0_13_55.VGND
rlabel metal1 177270 523491 177362 523587 1 dpga_flat_0.sr_0.FILLER_0_13_55.VPWR
flabel metal1 177483 522978 177517 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_57.VGND
flabel metal1 177483 523522 177517 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_57.VPWR
flabel nwell 177483 523522 177517 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_57.VPB
flabel pwell 177483 522978 177517 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_57.VNB
rlabel comment 177454 522995 177454 522995 4 dpga_flat_0.sr_0.FILLER_0_13_57.decap_12
flabel metal1 177115 522978 177149 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_53.VGND
flabel metal1 177115 522434 177149 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_53.VPWR
flabel nwell 177115 522434 177149 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_53.VPB
flabel pwell 177115 522978 177149 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_53.VNB
rlabel comment 177086 522995 177086 522995 2 dpga_flat_0.sr_0.FILLER_0_14_53.decap_12
flabel metal1 177384 523519 177437 523548 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_13_91.VPWR
flabel metal1 177383 522977 177434 523015 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_13_91.VGND
rlabel comment 177362 522995 177362 522995 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_13_91.tapvpwrvgnd_1
rlabel metal1 177362 522947 177454 523043 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_13_91.VGND
rlabel metal1 177362 523491 177454 523587 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_13_91.VPWR
flabel metal1 178587 522978 178621 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_69.VGND
flabel metal1 178587 523522 178621 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_69.VPWR
flabel nwell 178587 523522 178621 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_69.VPB
flabel pwell 178587 522978 178621 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_69.VNB
rlabel comment 178558 522995 178558 522995 4 dpga_flat_0.sr_0.FILLER_0_13_69.decap_12
flabel metal1 179691 522978 179725 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_81.VGND
flabel metal1 179691 523522 179725 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_81.VPWR
flabel nwell 179691 523522 179725 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_81.VPB
flabel pwell 179691 522978 179725 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_81.VNB
rlabel comment 179662 522995 179662 522995 4 dpga_flat_0.sr_0.FILLER_0_13_81.decap_12
flabel metal1 178219 522978 178253 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_65.VGND
flabel metal1 178219 522434 178253 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_65.VPWR
flabel nwell 178219 522434 178253 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_65.VPB
flabel pwell 178219 522978 178253 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_65.VNB
rlabel comment 178190 522995 178190 522995 2 dpga_flat_0.sr_0.FILLER_0_14_65.decap_12
flabel metal1 179323 522434 179357 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_77.VPWR
flabel metal1 179323 522978 179357 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_77.VGND
flabel nwell 179323 522434 179357 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_77.VPB
flabel pwell 179323 522978 179357 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_77.VNB
rlabel comment 179294 522995 179294 522995 2 dpga_flat_0.sr_0.FILLER_0_14_77.decap_6
rlabel metal1 179294 522947 179846 523043 5 dpga_flat_0.sr_0.FILLER_0_14_77.VGND
rlabel metal1 179294 522403 179846 522499 5 dpga_flat_0.sr_0.FILLER_0_14_77.VPWR
flabel metal1 179868 522438 179904 522468 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_83.VPWR
flabel metal1 179868 522979 179904 523008 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_83.VGND
flabel nwell 179877 522444 179897 522461 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_83.VPB
flabel pwell 179874 522984 179898 523006 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_83.VNB
rlabel comment 179846 522995 179846 522995 2 dpga_flat_0.sr_0.FILLER_0_14_83.fill_1
rlabel metal1 179846 522947 179938 523043 5 dpga_flat_0.sr_0.FILLER_0_14_83.VGND
rlabel metal1 179846 522403 179938 522499 5 dpga_flat_0.sr_0.FILLER_0_14_83.VPWR
flabel metal1 180795 522978 180829 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_93.VGND
flabel metal1 180795 523522 180829 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_93.VPWR
flabel nwell 180795 523522 180829 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_93.VPB
flabel pwell 180795 522978 180829 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_93.VNB
rlabel comment 180766 522995 180766 522995 4 dpga_flat_0.sr_0.FILLER_0_13_93.decap_12
flabel metal1 180059 522978 180093 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_85.VGND
flabel metal1 180059 522434 180093 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_85.VPWR
flabel nwell 180059 522434 180093 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_85.VPB
flabel pwell 180059 522978 180093 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_85.VNB
rlabel comment 180030 522995 180030 522995 2 dpga_flat_0.sr_0.FILLER_0_14_85.decap_12
flabel metal1 181163 522978 181197 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_97.VGND
flabel metal1 181163 522434 181197 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_97.VPWR
flabel nwell 181163 522434 181197 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_97.VPB
flabel pwell 181163 522978 181197 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_97.VNB
rlabel comment 181134 522995 181134 522995 2 dpga_flat_0.sr_0.FILLER_0_14_97.decap_12
flabel metal1 179960 522442 180013 522471 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_14_94.VPWR
flabel metal1 179959 522975 180010 523013 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_14_94.VGND
rlabel comment 179938 522995 179938 522995 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_14_94.tapvpwrvgnd_1
rlabel metal1 179938 522947 180030 523043 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_14_94.VGND
rlabel metal1 179938 522403 180030 522499 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_14_94.VPWR
flabel metal1 181899 523522 181933 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_105.VPWR
flabel metal1 181899 522978 181933 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_105.VGND
flabel nwell 181899 523522 181933 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_105.VPB
flabel pwell 181899 522978 181933 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_105.VNB
rlabel comment 181870 522995 181870 522995 4 dpga_flat_0.sr_0.FILLER_0_13_105.decap_6
rlabel metal1 181870 522947 182422 523043 1 dpga_flat_0.sr_0.FILLER_0_13_105.VGND
rlabel metal1 181870 523491 182422 523587 1 dpga_flat_0.sr_0.FILLER_0_13_105.VPWR
flabel metal1 182444 523522 182480 523552 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_111.VPWR
flabel metal1 182444 522982 182480 523011 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_111.VGND
flabel nwell 182453 523529 182473 523546 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_111.VPB
flabel pwell 182450 522984 182474 523006 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_111.VNB
rlabel comment 182422 522995 182422 522995 4 dpga_flat_0.sr_0.FILLER_0_13_111.fill_1
rlabel metal1 182422 522947 182514 523043 1 dpga_flat_0.sr_0.FILLER_0_13_111.VGND
rlabel metal1 182422 523491 182514 523587 1 dpga_flat_0.sr_0.FILLER_0_13_111.VPWR
flabel metal1 182635 522978 182669 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_113.VGND
flabel metal1 182635 523522 182669 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_113.VPWR
flabel nwell 182635 523522 182669 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_113.VPB
flabel pwell 182635 522978 182669 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_113.VNB
rlabel comment 182606 522995 182606 522995 4 dpga_flat_0.sr_0.FILLER_0_13_113.decap_12
flabel metal1 183739 522978 183773 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_125.VGND
flabel metal1 183739 523522 183773 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_125.VPWR
flabel nwell 183739 523522 183773 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_125.VPB
flabel pwell 183739 522978 183773 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_125.VNB
rlabel comment 183710 522995 183710 522995 4 dpga_flat_0.sr_0.FILLER_0_13_125.decap_12
flabel metal1 182267 522978 182301 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_109.VGND
flabel metal1 182267 522434 182301 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_109.VPWR
flabel nwell 182267 522434 182301 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_109.VPB
flabel pwell 182267 522978 182301 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_109.VNB
rlabel comment 182238 522995 182238 522995 2 dpga_flat_0.sr_0.FILLER_0_14_109.decap_12
flabel metal1 183371 522978 183405 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_121.VGND
flabel metal1 183371 522434 183405 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_121.VPWR
flabel nwell 183371 522434 183405 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_121.VPB
flabel pwell 183371 522978 183405 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_121.VNB
rlabel comment 183342 522995 183342 522995 2 dpga_flat_0.sr_0.FILLER_0_14_121.decap_12
flabel metal1 182536 523519 182589 523548 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_13_92.VPWR
flabel metal1 182535 522977 182586 523015 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_13_92.VGND
rlabel comment 182514 522995 182514 522995 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_13_92.tapvpwrvgnd_1
rlabel metal1 182514 522947 182606 523043 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_13_92.VGND
rlabel metal1 182514 523491 182606 523587 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_13_92.VPWR
flabel metal1 184843 522978 184877 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_137.VGND
flabel metal1 184843 523522 184877 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_137.VPWR
flabel nwell 184843 523522 184877 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_137.VPB
flabel pwell 184843 522978 184877 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_137.VNB
rlabel comment 184814 522995 184814 522995 4 dpga_flat_0.sr_0.FILLER_0_13_137.decap_12
flabel metal1 184475 522434 184509 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_133.VPWR
flabel metal1 184475 522978 184509 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_133.VGND
flabel nwell 184475 522434 184509 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_133.VPB
flabel pwell 184475 522978 184509 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_133.VNB
rlabel comment 184446 522995 184446 522995 2 dpga_flat_0.sr_0.FILLER_0_14_133.decap_6
rlabel metal1 184446 522947 184998 523043 5 dpga_flat_0.sr_0.FILLER_0_14_133.VGND
rlabel metal1 184446 522403 184998 522499 5 dpga_flat_0.sr_0.FILLER_0_14_133.VPWR
flabel metal1 185020 522438 185056 522468 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_139.VPWR
flabel metal1 185020 522979 185056 523008 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_139.VGND
flabel nwell 185029 522444 185049 522461 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_139.VPB
flabel pwell 185026 522984 185050 523006 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_139.VNB
rlabel comment 184998 522995 184998 522995 2 dpga_flat_0.sr_0.FILLER_0_14_139.fill_1
rlabel metal1 184998 522947 185090 523043 5 dpga_flat_0.sr_0.FILLER_0_14_139.VGND
rlabel metal1 184998 522403 185090 522499 5 dpga_flat_0.sr_0.FILLER_0_14_139.VPWR
flabel metal1 185211 522978 185245 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_141.VGND
flabel metal1 185211 522434 185245 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_141.VPWR
flabel nwell 185211 522434 185245 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_141.VPB
flabel pwell 185211 522978 185245 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_141.VNB
rlabel comment 185182 522995 185182 522995 2 dpga_flat_0.sr_0.FILLER_0_14_141.decap_12
flabel metal1 185112 522442 185165 522471 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_14_95.VPWR
flabel metal1 185111 522975 185162 523013 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_14_95.VGND
rlabel comment 185090 522995 185090 522995 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_14_95.tapvpwrvgnd_1
rlabel metal1 185090 522947 185182 523043 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_14_95.VGND
rlabel metal1 185090 522403 185182 522499 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_14_95.VPWR
flabel metal1 185947 522978 185981 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_149.VGND
flabel metal1 185947 523522 185981 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_149.VPWR
flabel nwell 185947 523522 185981 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_149.VPB
flabel pwell 185947 522978 185981 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_149.VNB
rlabel comment 185918 522995 185918 522995 4 dpga_flat_0.sr_0.FILLER_0_13_149.decap_12
flabel metal1 187042 522981 187095 523013 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_161.VGND
flabel metal1 187043 523525 187095 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_161.VPWR
flabel nwell 187050 523530 187084 523548 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_161.VPB
flabel pwell 187053 522985 187085 523007 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_13_161.VNB
rlabel comment 187022 522995 187022 522995 4 dpga_flat_0.sr_0.FILLER_0_13_161.fill_2
rlabel metal1 187022 522947 187206 523043 1 dpga_flat_0.sr_0.FILLER_0_13_161.VGND
rlabel metal1 187022 523491 187206 523587 1 dpga_flat_0.sr_0.FILLER_0_13_161.VPWR
flabel metal1 186315 522434 186349 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_153.VPWR
flabel metal1 186315 522978 186349 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_153.VGND
flabel nwell 186315 522434 186349 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_153.VPB
flabel pwell 186315 522978 186349 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_153.VNB
rlabel comment 186286 522995 186286 522995 2 dpga_flat_0.sr_0.FILLER_0_14_153.decap_8
rlabel metal1 186286 522947 187022 523043 5 dpga_flat_0.sr_0.FILLER_0_14_153.VGND
rlabel metal1 186286 522403 187022 522499 5 dpga_flat_0.sr_0.FILLER_0_14_153.VPWR
flabel metal1 187042 522977 187095 523009 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_161.VGND
flabel metal1 187043 522434 187095 522465 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_161.VPWR
flabel nwell 187050 522442 187084 522460 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_161.VPB
flabel pwell 187053 522983 187085 523005 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_14_161.VNB
rlabel comment 187022 522995 187022 522995 2 dpga_flat_0.sr_0.FILLER_0_14_161.fill_2
rlabel metal1 187022 522947 187206 523043 5 dpga_flat_0.sr_0.FILLER_0_14_161.VGND
rlabel metal1 187022 522403 187206 522499 5 dpga_flat_0.sr_0.FILLER_0_14_161.VPWR
flabel metal1 187419 523522 187453 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_13_Right_13.VPWR
flabel metal1 187419 522978 187453 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_13_Right_13.VGND
flabel nwell 187419 523522 187453 523556 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_13_Right_13.VPB
flabel pwell 187419 522978 187453 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_13_Right_13.VNB
rlabel comment 187482 522995 187482 522995 6 dpga_flat_0.sr_0.PHY_EDGE_ROW_13_Right_13.decap_3
rlabel metal1 187206 522947 187482 523043 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_13_Right_13.VGND
rlabel metal1 187206 523491 187482 523587 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_13_Right_13.VPWR
flabel metal1 187419 522434 187453 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_14_Right_14.VPWR
flabel metal1 187419 522978 187453 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_14_Right_14.VGND
flabel nwell 187419 522434 187453 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_14_Right_14.VPB
flabel pwell 187419 522978 187453 523012 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_14_Right_14.VNB
rlabel comment 187482 522995 187482 522995 8 dpga_flat_0.sr_0.PHY_EDGE_ROW_14_Right_14.decap_3
rlabel metal1 187206 522947 187482 523043 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_14_Right_14.VGND
rlabel metal1 187206 522403 187482 522499 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_14_Right_14.VPWR
flabel metal1 172515 521890 172549 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_3.VGND
flabel metal1 172515 522434 172549 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_3.VPWR
flabel nwell 172515 522434 172549 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_3.VPB
flabel pwell 172515 521890 172549 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_3.VNB
rlabel comment 172486 521907 172486 521907 4 dpga_flat_0.sr_0.FILLER_0_15_3.decap_12
flabel metal1 173619 521890 173653 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_15.VGND
flabel metal1 173619 522434 173653 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_15.VPWR
flabel nwell 173619 522434 173653 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_15.VPB
flabel pwell 173619 521890 173653 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_15.VNB
rlabel comment 173590 521907 173590 521907 4 dpga_flat_0.sr_0.FILLER_0_15_15.decap_12
flabel metal1 172239 522434 172273 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_15_Left_43.VPWR
flabel metal1 172239 521890 172273 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_15_Left_43.VGND
flabel nwell 172239 522434 172273 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_15_Left_43.VPB
flabel pwell 172239 521890 172273 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_15_Left_43.VNB
rlabel comment 172210 521907 172210 521907 4 dpga_flat_0.sr_0.PHY_EDGE_ROW_15_Left_43.decap_3
rlabel metal1 172210 521859 172486 521955 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_15_Left_43.VGND
rlabel metal1 172210 522403 172486 522499 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_15_Left_43.VPWR
flabel metal1 174723 521890 174757 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_27.VGND
flabel metal1 174723 522434 174757 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_27.VPWR
flabel nwell 174723 522434 174757 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_27.VPB
flabel pwell 174723 521890 174757 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_27.VNB
rlabel comment 174694 521907 174694 521907 4 dpga_flat_0.sr_0.FILLER_0_15_27.decap_12
flabel metal1 175827 521890 175861 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_39.VGND
flabel metal1 175827 522434 175861 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_39.VPWR
flabel nwell 175827 522434 175861 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_39.VPB
flabel pwell 175827 521890 175861 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_39.VNB
rlabel comment 175798 521907 175798 521907 4 dpga_flat_0.sr_0.FILLER_0_15_39.decap_12
flabel metal1 176931 521890 176965 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_51.VGND
flabel metal1 176931 522434 176965 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_51.VPWR
flabel nwell 176931 522434 176965 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_51.VPB
flabel pwell 176931 521890 176965 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_51.VNB
rlabel comment 176902 521907 176902 521907 4 dpga_flat_0.sr_0.FILLER_0_15_51.decap_4
rlabel metal1 176902 521859 177270 521955 1 dpga_flat_0.sr_0.FILLER_0_15_51.VGND
rlabel metal1 176902 522403 177270 522499 1 dpga_flat_0.sr_0.FILLER_0_15_51.VPWR
flabel metal1 177292 522434 177328 522464 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_55.VPWR
flabel metal1 177292 521894 177328 521923 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_55.VGND
flabel nwell 177301 522441 177321 522458 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_55.VPB
flabel pwell 177298 521896 177322 521918 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_55.VNB
rlabel comment 177270 521907 177270 521907 4 dpga_flat_0.sr_0.FILLER_0_15_55.fill_1
rlabel metal1 177270 521859 177362 521955 1 dpga_flat_0.sr_0.FILLER_0_15_55.VGND
rlabel metal1 177270 522403 177362 522499 1 dpga_flat_0.sr_0.FILLER_0_15_55.VPWR
flabel metal1 177483 521890 177517 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_57.VGND
flabel metal1 177483 522434 177517 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_57.VPWR
flabel nwell 177483 522434 177517 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_57.VPB
flabel pwell 177483 521890 177517 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_57.VNB
rlabel comment 177454 521907 177454 521907 4 dpga_flat_0.sr_0.FILLER_0_15_57.decap_12
flabel metal1 177384 522431 177437 522460 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_15_96.VPWR
flabel metal1 177383 521889 177434 521927 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_15_96.VGND
rlabel comment 177362 521907 177362 521907 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_15_96.tapvpwrvgnd_1
rlabel metal1 177362 521859 177454 521955 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_15_96.VGND
rlabel metal1 177362 522403 177454 522499 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_15_96.VPWR
flabel metal1 178587 521890 178621 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_69.VGND
flabel metal1 178587 522434 178621 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_69.VPWR
flabel nwell 178587 522434 178621 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_69.VPB
flabel pwell 178587 521890 178621 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_69.VNB
rlabel comment 178558 521907 178558 521907 4 dpga_flat_0.sr_0.FILLER_0_15_69.decap_12
flabel metal1 179691 521890 179725 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_81.VGND
flabel metal1 179691 522434 179725 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_81.VPWR
flabel nwell 179691 522434 179725 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_81.VPB
flabel pwell 179691 521890 179725 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_81.VNB
rlabel comment 179662 521907 179662 521907 4 dpga_flat_0.sr_0.FILLER_0_15_81.decap_12
flabel metal1 180795 521890 180829 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_93.VGND
flabel metal1 180795 522434 180829 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_93.VPWR
flabel nwell 180795 522434 180829 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_93.VPB
flabel pwell 180795 521890 180829 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_93.VNB
rlabel comment 180766 521907 180766 521907 4 dpga_flat_0.sr_0.FILLER_0_15_93.decap_12
flabel metal1 181899 522434 181933 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_105.VPWR
flabel metal1 181899 521890 181933 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_105.VGND
flabel nwell 181899 522434 181933 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_105.VPB
flabel pwell 181899 521890 181933 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_105.VNB
rlabel comment 181870 521907 181870 521907 4 dpga_flat_0.sr_0.FILLER_0_15_105.decap_6
rlabel metal1 181870 521859 182422 521955 1 dpga_flat_0.sr_0.FILLER_0_15_105.VGND
rlabel metal1 181870 522403 182422 522499 1 dpga_flat_0.sr_0.FILLER_0_15_105.VPWR
flabel metal1 182444 522434 182480 522464 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_111.VPWR
flabel metal1 182444 521894 182480 521923 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_111.VGND
flabel nwell 182453 522441 182473 522458 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_111.VPB
flabel pwell 182450 521896 182474 521918 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_111.VNB
rlabel comment 182422 521907 182422 521907 4 dpga_flat_0.sr_0.FILLER_0_15_111.fill_1
rlabel metal1 182422 521859 182514 521955 1 dpga_flat_0.sr_0.FILLER_0_15_111.VGND
rlabel metal1 182422 522403 182514 522499 1 dpga_flat_0.sr_0.FILLER_0_15_111.VPWR
flabel metal1 182635 521890 182669 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_113.VGND
flabel metal1 182635 522434 182669 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_113.VPWR
flabel nwell 182635 522434 182669 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_113.VPB
flabel pwell 182635 521890 182669 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_113.VNB
rlabel comment 182606 521907 182606 521907 4 dpga_flat_0.sr_0.FILLER_0_15_113.decap_12
flabel metal1 183739 521890 183773 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_125.VGND
flabel metal1 183739 522434 183773 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_125.VPWR
flabel nwell 183739 522434 183773 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_125.VPB
flabel pwell 183739 521890 183773 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_125.VNB
rlabel comment 183710 521907 183710 521907 4 dpga_flat_0.sr_0.FILLER_0_15_125.decap_12
flabel metal1 182536 522431 182589 522460 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_15_97.VPWR
flabel metal1 182535 521889 182586 521927 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_15_97.VGND
rlabel comment 182514 521907 182514 521907 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_15_97.tapvpwrvgnd_1
rlabel metal1 182514 521859 182606 521955 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_15_97.VGND
rlabel metal1 182514 522403 182606 522499 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_15_97.VPWR
flabel metal1 184843 521890 184877 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_137.VGND
flabel metal1 184843 522434 184877 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_137.VPWR
flabel nwell 184843 522434 184877 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_137.VPB
flabel pwell 184843 521890 184877 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_137.VNB
rlabel comment 184814 521907 184814 521907 4 dpga_flat_0.sr_0.FILLER_0_15_137.decap_12
flabel metal1 185947 521890 185981 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_149.VGND
flabel metal1 185947 522434 185981 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_149.VPWR
flabel nwell 185947 522434 185981 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_149.VPB
flabel pwell 185947 521890 185981 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_149.VNB
rlabel comment 185918 521907 185918 521907 4 dpga_flat_0.sr_0.FILLER_0_15_149.decap_12
flabel metal1 187042 521893 187095 521925 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_161.VGND
flabel metal1 187043 522437 187095 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_161.VPWR
flabel nwell 187050 522442 187084 522460 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_161.VPB
flabel pwell 187053 521897 187085 521919 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_15_161.VNB
rlabel comment 187022 521907 187022 521907 4 dpga_flat_0.sr_0.FILLER_0_15_161.fill_2
rlabel metal1 187022 521859 187206 521955 1 dpga_flat_0.sr_0.FILLER_0_15_161.VGND
rlabel metal1 187022 522403 187206 522499 1 dpga_flat_0.sr_0.FILLER_0_15_161.VPWR
flabel metal1 187419 522434 187453 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_15_Right_15.VPWR
flabel metal1 187419 521890 187453 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_15_Right_15.VGND
flabel nwell 187419 522434 187453 522468 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_15_Right_15.VPB
flabel pwell 187419 521890 187453 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_15_Right_15.VNB
rlabel comment 187482 521907 187482 521907 6 dpga_flat_0.sr_0.PHY_EDGE_ROW_15_Right_15.decap_3
rlabel metal1 187206 521859 187482 521955 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_15_Right_15.VGND
rlabel metal1 187206 522403 187482 522499 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_15_Right_15.VPWR
flabel metal1 172515 521890 172549 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_3.VGND
flabel metal1 172515 521346 172549 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_3.VPWR
flabel nwell 172515 521346 172549 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_3.VPB
flabel pwell 172515 521890 172549 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_3.VNB
rlabel comment 172486 521907 172486 521907 2 dpga_flat_0.sr_0.FILLER_0_16_3.decap_12
flabel metal1 173619 521890 173653 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_15.VGND
flabel metal1 173619 521346 173653 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_15.VPWR
flabel nwell 173619 521346 173653 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_15.VPB
flabel pwell 173619 521890 173653 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_15.VNB
rlabel comment 173590 521907 173590 521907 2 dpga_flat_0.sr_0.FILLER_0_16_15.decap_12
flabel metal1 172239 521346 172273 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_16_Left_44.VPWR
flabel metal1 172239 521890 172273 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_16_Left_44.VGND
flabel nwell 172239 521346 172273 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_16_Left_44.VPB
flabel pwell 172239 521890 172273 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_16_Left_44.VNB
rlabel comment 172210 521907 172210 521907 2 dpga_flat_0.sr_0.PHY_EDGE_ROW_16_Left_44.decap_3
rlabel metal1 172210 521859 172486 521955 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_16_Left_44.VGND
rlabel metal1 172210 521315 172486 521411 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_16_Left_44.VPWR
flabel metal1 174716 521350 174752 521380 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_27.VPWR
flabel metal1 174716 521891 174752 521920 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_27.VGND
flabel nwell 174725 521356 174745 521373 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_27.VPB
flabel pwell 174722 521896 174746 521918 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_27.VNB
rlabel comment 174694 521907 174694 521907 2 dpga_flat_0.sr_0.FILLER_0_16_27.fill_1
rlabel metal1 174694 521859 174786 521955 5 dpga_flat_0.sr_0.FILLER_0_16_27.VGND
rlabel metal1 174694 521315 174786 521411 5 dpga_flat_0.sr_0.FILLER_0_16_27.VPWR
flabel metal1 174907 521890 174941 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_29.VGND
flabel metal1 174907 521346 174941 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_29.VPWR
flabel nwell 174907 521346 174941 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_29.VPB
flabel pwell 174907 521890 174941 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_29.VNB
rlabel comment 174878 521907 174878 521907 2 dpga_flat_0.sr_0.FILLER_0_16_29.decap_12
flabel metal1 176011 521890 176045 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_41.VGND
flabel metal1 176011 521346 176045 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_41.VPWR
flabel nwell 176011 521346 176045 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_41.VPB
flabel pwell 176011 521890 176045 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_41.VNB
rlabel comment 175982 521907 175982 521907 2 dpga_flat_0.sr_0.FILLER_0_16_41.decap_12
flabel metal1 174808 521354 174861 521383 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_16_98.VPWR
flabel metal1 174807 521887 174858 521925 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_16_98.VGND
rlabel comment 174786 521907 174786 521907 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_16_98.tapvpwrvgnd_1
rlabel metal1 174786 521859 174878 521955 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_16_98.VGND
rlabel metal1 174786 521315 174878 521411 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_16_98.VPWR
flabel metal1 177115 521890 177149 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_53.VGND
flabel metal1 177115 521346 177149 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_53.VPWR
flabel nwell 177115 521346 177149 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_53.VPB
flabel pwell 177115 521890 177149 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_53.VNB
rlabel comment 177086 521907 177086 521907 2 dpga_flat_0.sr_0.FILLER_0_16_53.decap_12
flabel metal1 178219 521890 178253 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_65.VGND
flabel metal1 178219 521346 178253 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_65.VPWR
flabel nwell 178219 521346 178253 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_65.VPB
flabel pwell 178219 521890 178253 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_65.VNB
rlabel comment 178190 521907 178190 521907 2 dpga_flat_0.sr_0.FILLER_0_16_65.decap_12
flabel metal1 179323 521346 179357 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_77.VPWR
flabel metal1 179323 521890 179357 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_77.VGND
flabel nwell 179323 521346 179357 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_77.VPB
flabel pwell 179323 521890 179357 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_77.VNB
rlabel comment 179294 521907 179294 521907 2 dpga_flat_0.sr_0.FILLER_0_16_77.decap_6
rlabel metal1 179294 521859 179846 521955 5 dpga_flat_0.sr_0.FILLER_0_16_77.VGND
rlabel metal1 179294 521315 179846 521411 5 dpga_flat_0.sr_0.FILLER_0_16_77.VPWR
flabel metal1 179868 521350 179904 521380 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_83.VPWR
flabel metal1 179868 521891 179904 521920 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_83.VGND
flabel nwell 179877 521356 179897 521373 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_83.VPB
flabel pwell 179874 521896 179898 521918 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_83.VNB
rlabel comment 179846 521907 179846 521907 2 dpga_flat_0.sr_0.FILLER_0_16_83.fill_1
rlabel metal1 179846 521859 179938 521955 5 dpga_flat_0.sr_0.FILLER_0_16_83.VGND
rlabel metal1 179846 521315 179938 521411 5 dpga_flat_0.sr_0.FILLER_0_16_83.VPWR
flabel metal1 180059 521890 180093 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_85.VGND
flabel metal1 180059 521346 180093 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_85.VPWR
flabel nwell 180059 521346 180093 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_85.VPB
flabel pwell 180059 521890 180093 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_85.VNB
rlabel comment 180030 521907 180030 521907 2 dpga_flat_0.sr_0.FILLER_0_16_85.decap_12
flabel metal1 181163 521890 181197 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_97.VGND
flabel metal1 181163 521346 181197 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_97.VPWR
flabel nwell 181163 521346 181197 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_97.VPB
flabel pwell 181163 521890 181197 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_97.VNB
rlabel comment 181134 521907 181134 521907 2 dpga_flat_0.sr_0.FILLER_0_16_97.decap_12
flabel metal1 179960 521354 180013 521383 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_16_99.VPWR
flabel metal1 179959 521887 180010 521925 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_16_99.VGND
rlabel comment 179938 521907 179938 521907 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_16_99.tapvpwrvgnd_1
rlabel metal1 179938 521859 180030 521955 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_16_99.VGND
rlabel metal1 179938 521315 180030 521411 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_16_99.VPWR
flabel metal1 182267 521890 182301 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_109.VGND
flabel metal1 182267 521346 182301 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_109.VPWR
flabel nwell 182267 521346 182301 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_109.VPB
flabel pwell 182267 521890 182301 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_109.VNB
rlabel comment 182238 521907 182238 521907 2 dpga_flat_0.sr_0.FILLER_0_16_109.decap_12
flabel metal1 183371 521890 183405 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_121.VGND
flabel metal1 183371 521346 183405 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_121.VPWR
flabel nwell 183371 521346 183405 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_121.VPB
flabel pwell 183371 521890 183405 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_121.VNB
rlabel comment 183342 521907 183342 521907 2 dpga_flat_0.sr_0.FILLER_0_16_121.decap_12
flabel metal1 184475 521346 184509 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_133.VPWR
flabel metal1 184475 521890 184509 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_133.VGND
flabel nwell 184475 521346 184509 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_133.VPB
flabel pwell 184475 521890 184509 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_133.VNB
rlabel comment 184446 521907 184446 521907 2 dpga_flat_0.sr_0.FILLER_0_16_133.decap_6
rlabel metal1 184446 521859 184998 521955 5 dpga_flat_0.sr_0.FILLER_0_16_133.VGND
rlabel metal1 184446 521315 184998 521411 5 dpga_flat_0.sr_0.FILLER_0_16_133.VPWR
flabel metal1 185020 521350 185056 521380 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_139.VPWR
flabel metal1 185020 521891 185056 521920 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_139.VGND
flabel nwell 185029 521356 185049 521373 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_139.VPB
flabel pwell 185026 521896 185050 521918 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_139.VNB
rlabel comment 184998 521907 184998 521907 2 dpga_flat_0.sr_0.FILLER_0_16_139.fill_1
rlabel metal1 184998 521859 185090 521955 5 dpga_flat_0.sr_0.FILLER_0_16_139.VGND
rlabel metal1 184998 521315 185090 521411 5 dpga_flat_0.sr_0.FILLER_0_16_139.VPWR
flabel metal1 185211 521890 185245 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_141.VGND
flabel metal1 185211 521346 185245 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_141.VPWR
flabel nwell 185211 521346 185245 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_141.VPB
flabel pwell 185211 521890 185245 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_141.VNB
rlabel comment 185182 521907 185182 521907 2 dpga_flat_0.sr_0.FILLER_0_16_141.decap_12
flabel metal1 185112 521354 185165 521383 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_16_100.VPWR
flabel metal1 185111 521887 185162 521925 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_16_100.VGND
rlabel comment 185090 521907 185090 521907 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_16_100.tapvpwrvgnd_1
rlabel metal1 185090 521859 185182 521955 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_16_100.VGND
rlabel metal1 185090 521315 185182 521411 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_16_100.VPWR
flabel metal1 186315 521346 186349 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_153.VPWR
flabel metal1 186315 521890 186349 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_153.VGND
flabel nwell 186315 521346 186349 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_153.VPB
flabel pwell 186315 521890 186349 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_153.VNB
rlabel comment 186286 521907 186286 521907 2 dpga_flat_0.sr_0.FILLER_0_16_153.decap_8
rlabel metal1 186286 521859 187022 521955 5 dpga_flat_0.sr_0.FILLER_0_16_153.VGND
rlabel metal1 186286 521315 187022 521411 5 dpga_flat_0.sr_0.FILLER_0_16_153.VPWR
flabel metal1 187042 521889 187095 521921 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_161.VGND
flabel metal1 187043 521346 187095 521377 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_161.VPWR
flabel nwell 187050 521354 187084 521372 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_161.VPB
flabel pwell 187053 521895 187085 521917 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_16_161.VNB
rlabel comment 187022 521907 187022 521907 2 dpga_flat_0.sr_0.FILLER_0_16_161.fill_2
rlabel metal1 187022 521859 187206 521955 5 dpga_flat_0.sr_0.FILLER_0_16_161.VGND
rlabel metal1 187022 521315 187206 521411 5 dpga_flat_0.sr_0.FILLER_0_16_161.VPWR
flabel metal1 187419 521346 187453 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_16_Right_16.VPWR
flabel metal1 187419 521890 187453 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_16_Right_16.VGND
flabel nwell 187419 521346 187453 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_16_Right_16.VPB
flabel pwell 187419 521890 187453 521924 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_16_Right_16.VNB
rlabel comment 187482 521907 187482 521907 8 dpga_flat_0.sr_0.PHY_EDGE_ROW_16_Right_16.decap_3
rlabel metal1 187206 521859 187482 521955 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_16_Right_16.VGND
rlabel metal1 187206 521315 187482 521411 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_16_Right_16.VPWR
flabel metal1 172515 520802 172549 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_3.VGND
flabel metal1 172515 521346 172549 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_3.VPWR
flabel nwell 172515 521346 172549 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_3.VPB
flabel pwell 172515 520802 172549 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_3.VNB
rlabel comment 172486 520819 172486 520819 4 dpga_flat_0.sr_0.FILLER_0_17_3.decap_12
flabel metal1 173619 520802 173653 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_15.VGND
flabel metal1 173619 521346 173653 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_15.VPWR
flabel nwell 173619 521346 173653 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_15.VPB
flabel pwell 173619 520802 173653 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_15.VNB
rlabel comment 173590 520819 173590 520819 4 dpga_flat_0.sr_0.FILLER_0_17_15.decap_12
flabel metal1 172239 521346 172273 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_17_Left_45.VPWR
flabel metal1 172239 520802 172273 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_17_Left_45.VGND
flabel nwell 172239 521346 172273 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_17_Left_45.VPB
flabel pwell 172239 520802 172273 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_17_Left_45.VNB
rlabel comment 172210 520819 172210 520819 4 dpga_flat_0.sr_0.PHY_EDGE_ROW_17_Left_45.decap_3
rlabel metal1 172210 520771 172486 520867 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_17_Left_45.VGND
rlabel metal1 172210 521315 172486 521411 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_17_Left_45.VPWR
flabel metal1 174723 520802 174757 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_27.VGND
flabel metal1 174723 521346 174757 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_27.VPWR
flabel nwell 174723 521346 174757 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_27.VPB
flabel pwell 174723 520802 174757 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_27.VNB
rlabel comment 174694 520819 174694 520819 4 dpga_flat_0.sr_0.FILLER_0_17_27.decap_12
flabel metal1 175827 520802 175861 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_39.VGND
flabel metal1 175827 521346 175861 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_39.VPWR
flabel nwell 175827 521346 175861 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_39.VPB
flabel pwell 175827 520802 175861 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_39.VNB
rlabel comment 175798 520819 175798 520819 4 dpga_flat_0.sr_0.FILLER_0_17_39.decap_12
flabel metal1 176931 520802 176965 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_51.VGND
flabel metal1 176931 521346 176965 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_51.VPWR
flabel nwell 176931 521346 176965 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_51.VPB
flabel pwell 176931 520802 176965 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_51.VNB
rlabel comment 176902 520819 176902 520819 4 dpga_flat_0.sr_0.FILLER_0_17_51.decap_4
rlabel metal1 176902 520771 177270 520867 1 dpga_flat_0.sr_0.FILLER_0_17_51.VGND
rlabel metal1 176902 521315 177270 521411 1 dpga_flat_0.sr_0.FILLER_0_17_51.VPWR
flabel metal1 177292 521346 177328 521376 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_55.VPWR
flabel metal1 177292 520806 177328 520835 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_55.VGND
flabel nwell 177301 521353 177321 521370 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_55.VPB
flabel pwell 177298 520808 177322 520830 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_55.VNB
rlabel comment 177270 520819 177270 520819 4 dpga_flat_0.sr_0.FILLER_0_17_55.fill_1
rlabel metal1 177270 520771 177362 520867 1 dpga_flat_0.sr_0.FILLER_0_17_55.VGND
rlabel metal1 177270 521315 177362 521411 1 dpga_flat_0.sr_0.FILLER_0_17_55.VPWR
flabel metal1 177483 520802 177517 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_57.VGND
flabel metal1 177483 521346 177517 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_57.VPWR
flabel nwell 177483 521346 177517 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_57.VPB
flabel pwell 177483 520802 177517 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_57.VNB
rlabel comment 177454 520819 177454 520819 4 dpga_flat_0.sr_0.FILLER_0_17_57.decap_12
flabel metal1 177384 521343 177437 521372 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_17_101.VPWR
flabel metal1 177383 520801 177434 520839 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_17_101.VGND
rlabel comment 177362 520819 177362 520819 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_17_101.tapvpwrvgnd_1
rlabel metal1 177362 520771 177454 520867 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_17_101.VGND
rlabel metal1 177362 521315 177454 521411 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_17_101.VPWR
flabel metal1 178587 520802 178621 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_69.VGND
flabel metal1 178587 521346 178621 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_69.VPWR
flabel nwell 178587 521346 178621 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_69.VPB
flabel pwell 178587 520802 178621 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_69.VNB
rlabel comment 178558 520819 178558 520819 4 dpga_flat_0.sr_0.FILLER_0_17_69.decap_12
flabel metal1 179691 520802 179725 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_81.VGND
flabel metal1 179691 521346 179725 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_81.VPWR
flabel nwell 179691 521346 179725 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_81.VPB
flabel pwell 179691 520802 179725 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_81.VNB
rlabel comment 179662 520819 179662 520819 4 dpga_flat_0.sr_0.FILLER_0_17_81.decap_12
flabel metal1 180795 520802 180829 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_93.VGND
flabel metal1 180795 521346 180829 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_93.VPWR
flabel nwell 180795 521346 180829 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_93.VPB
flabel pwell 180795 520802 180829 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_93.VNB
rlabel comment 180766 520819 180766 520819 4 dpga_flat_0.sr_0.FILLER_0_17_93.decap_12
flabel metal1 181899 521346 181933 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_105.VPWR
flabel metal1 181899 520802 181933 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_105.VGND
flabel nwell 181899 521346 181933 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_105.VPB
flabel pwell 181899 520802 181933 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_105.VNB
rlabel comment 181870 520819 181870 520819 4 dpga_flat_0.sr_0.FILLER_0_17_105.decap_6
rlabel metal1 181870 520771 182422 520867 1 dpga_flat_0.sr_0.FILLER_0_17_105.VGND
rlabel metal1 181870 521315 182422 521411 1 dpga_flat_0.sr_0.FILLER_0_17_105.VPWR
flabel metal1 182444 521346 182480 521376 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_111.VPWR
flabel metal1 182444 520806 182480 520835 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_111.VGND
flabel nwell 182453 521353 182473 521370 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_111.VPB
flabel pwell 182450 520808 182474 520830 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_111.VNB
rlabel comment 182422 520819 182422 520819 4 dpga_flat_0.sr_0.FILLER_0_17_111.fill_1
rlabel metal1 182422 520771 182514 520867 1 dpga_flat_0.sr_0.FILLER_0_17_111.VGND
rlabel metal1 182422 521315 182514 521411 1 dpga_flat_0.sr_0.FILLER_0_17_111.VPWR
flabel metal1 182635 520802 182669 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_113.VGND
flabel metal1 182635 521346 182669 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_113.VPWR
flabel nwell 182635 521346 182669 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_113.VPB
flabel pwell 182635 520802 182669 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_113.VNB
rlabel comment 182606 520819 182606 520819 4 dpga_flat_0.sr_0.FILLER_0_17_113.decap_12
flabel metal1 183739 520802 183773 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_125.VGND
flabel metal1 183739 521346 183773 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_125.VPWR
flabel nwell 183739 521346 183773 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_125.VPB
flabel pwell 183739 520802 183773 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_125.VNB
rlabel comment 183710 520819 183710 520819 4 dpga_flat_0.sr_0.FILLER_0_17_125.decap_12
flabel metal1 182536 521343 182589 521372 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_17_102.VPWR
flabel metal1 182535 520801 182586 520839 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_17_102.VGND
rlabel comment 182514 520819 182514 520819 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_17_102.tapvpwrvgnd_1
rlabel metal1 182514 520771 182606 520867 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_17_102.VGND
rlabel metal1 182514 521315 182606 521411 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_17_102.VPWR
flabel metal1 184843 520802 184877 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_137.VGND
flabel metal1 184843 521346 184877 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_137.VPWR
flabel nwell 184843 521346 184877 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_137.VPB
flabel pwell 184843 520802 184877 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_137.VNB
rlabel comment 184814 520819 184814 520819 4 dpga_flat_0.sr_0.FILLER_0_17_137.decap_12
flabel metal1 185947 520802 185981 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_149.VGND
flabel metal1 185947 521346 185981 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_149.VPWR
flabel nwell 185947 521346 185981 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_149.VPB
flabel pwell 185947 520802 185981 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_149.VNB
rlabel comment 185918 520819 185918 520819 4 dpga_flat_0.sr_0.FILLER_0_17_149.decap_12
flabel metal1 187042 520805 187095 520837 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_161.VGND
flabel metal1 187043 521349 187095 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_161.VPWR
flabel nwell 187050 521354 187084 521372 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_161.VPB
flabel pwell 187053 520809 187085 520831 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_17_161.VNB
rlabel comment 187022 520819 187022 520819 4 dpga_flat_0.sr_0.FILLER_0_17_161.fill_2
rlabel metal1 187022 520771 187206 520867 1 dpga_flat_0.sr_0.FILLER_0_17_161.VGND
rlabel metal1 187022 521315 187206 521411 1 dpga_flat_0.sr_0.FILLER_0_17_161.VPWR
flabel metal1 187419 521346 187453 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_17_Right_17.VPWR
flabel metal1 187419 520802 187453 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_17_Right_17.VGND
flabel nwell 187419 521346 187453 521380 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_17_Right_17.VPB
flabel pwell 187419 520802 187453 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_17_Right_17.VNB
rlabel comment 187482 520819 187482 520819 6 dpga_flat_0.sr_0.PHY_EDGE_ROW_17_Right_17.decap_3
rlabel metal1 187206 520771 187482 520867 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_17_Right_17.VGND
rlabel metal1 187206 521315 187482 521411 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_17_Right_17.VPWR
flabel metal1 172515 520802 172549 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_3.VGND
flabel metal1 172515 520258 172549 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_3.VPWR
flabel nwell 172515 520258 172549 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_3.VPB
flabel pwell 172515 520802 172549 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_3.VNB
rlabel comment 172486 520819 172486 520819 2 dpga_flat_0.sr_0.FILLER_0_18_3.decap_12
flabel metal1 173619 520802 173653 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_15.VGND
flabel metal1 173619 520258 173653 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_15.VPWR
flabel nwell 173619 520258 173653 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_15.VPB
flabel pwell 173619 520802 173653 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_15.VNB
rlabel comment 173590 520819 173590 520819 2 dpga_flat_0.sr_0.FILLER_0_18_15.decap_12
flabel metal1 172239 520258 172273 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_18_Left_46.VPWR
flabel metal1 172239 520802 172273 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_18_Left_46.VGND
flabel nwell 172239 520258 172273 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_18_Left_46.VPB
flabel pwell 172239 520802 172273 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_18_Left_46.VNB
rlabel comment 172210 520819 172210 520819 2 dpga_flat_0.sr_0.PHY_EDGE_ROW_18_Left_46.decap_3
rlabel metal1 172210 520771 172486 520867 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_18_Left_46.VGND
rlabel metal1 172210 520227 172486 520323 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_18_Left_46.VPWR
flabel metal1 174716 520262 174752 520292 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_27.VPWR
flabel metal1 174716 520803 174752 520832 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_27.VGND
flabel nwell 174725 520268 174745 520285 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_27.VPB
flabel pwell 174722 520808 174746 520830 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_27.VNB
rlabel comment 174694 520819 174694 520819 2 dpga_flat_0.sr_0.FILLER_0_18_27.fill_1
rlabel metal1 174694 520771 174786 520867 5 dpga_flat_0.sr_0.FILLER_0_18_27.VGND
rlabel metal1 174694 520227 174786 520323 5 dpga_flat_0.sr_0.FILLER_0_18_27.VPWR
flabel metal1 174907 520802 174941 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_29.VGND
flabel metal1 174907 520258 174941 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_29.VPWR
flabel nwell 174907 520258 174941 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_29.VPB
flabel pwell 174907 520802 174941 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_29.VNB
rlabel comment 174878 520819 174878 520819 2 dpga_flat_0.sr_0.FILLER_0_18_29.decap_12
flabel metal1 176011 520802 176045 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_41.VGND
flabel metal1 176011 520258 176045 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_41.VPWR
flabel nwell 176011 520258 176045 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_41.VPB
flabel pwell 176011 520802 176045 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_41.VNB
rlabel comment 175982 520819 175982 520819 2 dpga_flat_0.sr_0.FILLER_0_18_41.decap_12
flabel metal1 174808 520266 174861 520295 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_18_103.VPWR
flabel metal1 174807 520799 174858 520837 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_18_103.VGND
rlabel comment 174786 520819 174786 520819 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_18_103.tapvpwrvgnd_1
rlabel metal1 174786 520771 174878 520867 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_18_103.VGND
rlabel metal1 174786 520227 174878 520323 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_18_103.VPWR
flabel metal1 177115 520802 177149 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_53.VGND
flabel metal1 177115 520258 177149 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_53.VPWR
flabel nwell 177115 520258 177149 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_53.VPB
flabel pwell 177115 520802 177149 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_53.VNB
rlabel comment 177086 520819 177086 520819 2 dpga_flat_0.sr_0.FILLER_0_18_53.decap_12
flabel metal1 178219 520802 178253 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_65.VGND
flabel metal1 178219 520258 178253 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_65.VPWR
flabel nwell 178219 520258 178253 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_65.VPB
flabel pwell 178219 520802 178253 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_65.VNB
rlabel comment 178190 520819 178190 520819 2 dpga_flat_0.sr_0.FILLER_0_18_65.decap_12
flabel metal1 179323 520258 179357 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_77.VPWR
flabel metal1 179323 520802 179357 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_77.VGND
flabel nwell 179323 520258 179357 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_77.VPB
flabel pwell 179323 520802 179357 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_77.VNB
rlabel comment 179294 520819 179294 520819 2 dpga_flat_0.sr_0.FILLER_0_18_77.decap_6
rlabel metal1 179294 520771 179846 520867 5 dpga_flat_0.sr_0.FILLER_0_18_77.VGND
rlabel metal1 179294 520227 179846 520323 5 dpga_flat_0.sr_0.FILLER_0_18_77.VPWR
flabel metal1 179868 520262 179904 520292 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_83.VPWR
flabel metal1 179868 520803 179904 520832 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_83.VGND
flabel nwell 179877 520268 179897 520285 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_83.VPB
flabel pwell 179874 520808 179898 520830 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_83.VNB
rlabel comment 179846 520819 179846 520819 2 dpga_flat_0.sr_0.FILLER_0_18_83.fill_1
rlabel metal1 179846 520771 179938 520867 5 dpga_flat_0.sr_0.FILLER_0_18_83.VGND
rlabel metal1 179846 520227 179938 520323 5 dpga_flat_0.sr_0.FILLER_0_18_83.VPWR
flabel metal1 180059 520802 180093 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_85.VGND
flabel metal1 180059 520258 180093 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_85.VPWR
flabel nwell 180059 520258 180093 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_85.VPB
flabel pwell 180059 520802 180093 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_85.VNB
rlabel comment 180030 520819 180030 520819 2 dpga_flat_0.sr_0.FILLER_0_18_85.decap_12
flabel metal1 181163 520802 181197 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_97.VGND
flabel metal1 181163 520258 181197 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_97.VPWR
flabel nwell 181163 520258 181197 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_97.VPB
flabel pwell 181163 520802 181197 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_97.VNB
rlabel comment 181134 520819 181134 520819 2 dpga_flat_0.sr_0.FILLER_0_18_97.decap_12
flabel metal1 179960 520266 180013 520295 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_18_104.VPWR
flabel metal1 179959 520799 180010 520837 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_18_104.VGND
rlabel comment 179938 520819 179938 520819 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_18_104.tapvpwrvgnd_1
rlabel metal1 179938 520771 180030 520867 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_18_104.VGND
rlabel metal1 179938 520227 180030 520323 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_18_104.VPWR
flabel metal1 182267 520802 182301 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_109.VGND
flabel metal1 182267 520258 182301 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_109.VPWR
flabel nwell 182267 520258 182301 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_109.VPB
flabel pwell 182267 520802 182301 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_109.VNB
rlabel comment 182238 520819 182238 520819 2 dpga_flat_0.sr_0.FILLER_0_18_109.decap_12
flabel metal1 183371 520802 183405 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_121.VGND
flabel metal1 183371 520258 183405 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_121.VPWR
flabel nwell 183371 520258 183405 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_121.VPB
flabel pwell 183371 520802 183405 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_121.VNB
rlabel comment 183342 520819 183342 520819 2 dpga_flat_0.sr_0.FILLER_0_18_121.decap_12
flabel metal1 184475 520258 184509 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_133.VPWR
flabel metal1 184475 520802 184509 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_133.VGND
flabel nwell 184475 520258 184509 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_133.VPB
flabel pwell 184475 520802 184509 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_133.VNB
rlabel comment 184446 520819 184446 520819 2 dpga_flat_0.sr_0.FILLER_0_18_133.decap_6
rlabel metal1 184446 520771 184998 520867 5 dpga_flat_0.sr_0.FILLER_0_18_133.VGND
rlabel metal1 184446 520227 184998 520323 5 dpga_flat_0.sr_0.FILLER_0_18_133.VPWR
flabel metal1 185020 520262 185056 520292 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_139.VPWR
flabel metal1 185020 520803 185056 520832 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_139.VGND
flabel nwell 185029 520268 185049 520285 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_139.VPB
flabel pwell 185026 520808 185050 520830 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_139.VNB
rlabel comment 184998 520819 184998 520819 2 dpga_flat_0.sr_0.FILLER_0_18_139.fill_1
rlabel metal1 184998 520771 185090 520867 5 dpga_flat_0.sr_0.FILLER_0_18_139.VGND
rlabel metal1 184998 520227 185090 520323 5 dpga_flat_0.sr_0.FILLER_0_18_139.VPWR
flabel metal1 185211 520802 185245 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_141.VGND
flabel metal1 185211 520258 185245 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_141.VPWR
flabel nwell 185211 520258 185245 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_141.VPB
flabel pwell 185211 520802 185245 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_141.VNB
rlabel comment 185182 520819 185182 520819 2 dpga_flat_0.sr_0.FILLER_0_18_141.decap_12
flabel metal1 185112 520266 185165 520295 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_18_105.VPWR
flabel metal1 185111 520799 185162 520837 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_18_105.VGND
rlabel comment 185090 520819 185090 520819 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_18_105.tapvpwrvgnd_1
rlabel metal1 185090 520771 185182 520867 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_18_105.VGND
rlabel metal1 185090 520227 185182 520323 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_18_105.VPWR
flabel metal1 186315 520258 186349 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_153.VPWR
flabel metal1 186315 520802 186349 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_153.VGND
flabel nwell 186315 520258 186349 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_153.VPB
flabel pwell 186315 520802 186349 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_153.VNB
rlabel comment 186286 520819 186286 520819 2 dpga_flat_0.sr_0.FILLER_0_18_153.decap_8
rlabel metal1 186286 520771 187022 520867 5 dpga_flat_0.sr_0.FILLER_0_18_153.VGND
rlabel metal1 186286 520227 187022 520323 5 dpga_flat_0.sr_0.FILLER_0_18_153.VPWR
flabel metal1 187042 520801 187095 520833 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_161.VGND
flabel metal1 187043 520258 187095 520289 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_161.VPWR
flabel nwell 187050 520266 187084 520284 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_161.VPB
flabel pwell 187053 520807 187085 520829 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_18_161.VNB
rlabel comment 187022 520819 187022 520819 2 dpga_flat_0.sr_0.FILLER_0_18_161.fill_2
rlabel metal1 187022 520771 187206 520867 5 dpga_flat_0.sr_0.FILLER_0_18_161.VGND
rlabel metal1 187022 520227 187206 520323 5 dpga_flat_0.sr_0.FILLER_0_18_161.VPWR
flabel metal1 187419 520258 187453 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_18_Right_18.VPWR
flabel metal1 187419 520802 187453 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_18_Right_18.VGND
flabel nwell 187419 520258 187453 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_18_Right_18.VPB
flabel pwell 187419 520802 187453 520836 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_18_Right_18.VNB
rlabel comment 187482 520819 187482 520819 8 dpga_flat_0.sr_0.PHY_EDGE_ROW_18_Right_18.decap_3
rlabel metal1 187206 520771 187482 520867 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_18_Right_18.VGND
rlabel metal1 187206 520227 187482 520323 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_18_Right_18.VPWR
flabel metal1 172515 519714 172549 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_3.VGND
flabel metal1 172515 520258 172549 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_3.VPWR
flabel nwell 172515 520258 172549 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_3.VPB
flabel pwell 172515 519714 172549 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_3.VNB
rlabel comment 172486 519731 172486 519731 4 dpga_flat_0.sr_0.FILLER_0_19_3.decap_12
flabel metal1 173619 519714 173653 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_15.VGND
flabel metal1 173619 520258 173653 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_15.VPWR
flabel nwell 173619 520258 173653 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_15.VPB
flabel pwell 173619 519714 173653 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_15.VNB
rlabel comment 173590 519731 173590 519731 4 dpga_flat_0.sr_0.FILLER_0_19_15.decap_12
flabel metal1 172515 519714 172549 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_3.VGND
flabel metal1 172515 519170 172549 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_3.VPWR
flabel nwell 172515 519170 172549 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_3.VPB
flabel pwell 172515 519714 172549 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_3.VNB
rlabel comment 172486 519731 172486 519731 2 dpga_flat_0.sr_0.FILLER_0_20_3.decap_12
flabel metal1 173619 519714 173653 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_15.VGND
flabel metal1 173619 519170 173653 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_15.VPWR
flabel nwell 173619 519170 173653 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_15.VPB
flabel pwell 173619 519714 173653 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_15.VNB
rlabel comment 173590 519731 173590 519731 2 dpga_flat_0.sr_0.FILLER_0_20_15.decap_12
flabel metal1 172239 520258 172273 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_19_Left_47.VPWR
flabel metal1 172239 519714 172273 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_19_Left_47.VGND
flabel nwell 172239 520258 172273 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_19_Left_47.VPB
flabel pwell 172239 519714 172273 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_19_Left_47.VNB
rlabel comment 172210 519731 172210 519731 4 dpga_flat_0.sr_0.PHY_EDGE_ROW_19_Left_47.decap_3
rlabel metal1 172210 519683 172486 519779 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_19_Left_47.VGND
rlabel metal1 172210 520227 172486 520323 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_19_Left_47.VPWR
flabel metal1 172239 519170 172273 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_20_Left_48.VPWR
flabel metal1 172239 519714 172273 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_20_Left_48.VGND
flabel nwell 172239 519170 172273 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_20_Left_48.VPB
flabel pwell 172239 519714 172273 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_20_Left_48.VNB
rlabel comment 172210 519731 172210 519731 2 dpga_flat_0.sr_0.PHY_EDGE_ROW_20_Left_48.decap_3
rlabel metal1 172210 519683 172486 519779 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_20_Left_48.VGND
rlabel metal1 172210 519139 172486 519235 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_20_Left_48.VPWR
flabel metal1 174723 519714 174757 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_27.VGND
flabel metal1 174723 520258 174757 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_27.VPWR
flabel nwell 174723 520258 174757 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_27.VPB
flabel pwell 174723 519714 174757 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_27.VNB
rlabel comment 174694 519731 174694 519731 4 dpga_flat_0.sr_0.FILLER_0_19_27.decap_12
flabel metal1 175827 519714 175861 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_39.VGND
flabel metal1 175827 520258 175861 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_39.VPWR
flabel nwell 175827 520258 175861 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_39.VPB
flabel pwell 175827 519714 175861 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_39.VNB
rlabel comment 175798 519731 175798 519731 4 dpga_flat_0.sr_0.FILLER_0_19_39.decap_12
flabel metal1 174716 519174 174752 519204 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_27.VPWR
flabel metal1 174716 519715 174752 519744 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_27.VGND
flabel nwell 174725 519180 174745 519197 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_27.VPB
flabel pwell 174722 519720 174746 519742 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_27.VNB
rlabel comment 174694 519731 174694 519731 2 dpga_flat_0.sr_0.FILLER_0_20_27.fill_1
rlabel metal1 174694 519683 174786 519779 5 dpga_flat_0.sr_0.FILLER_0_20_27.VGND
rlabel metal1 174694 519139 174786 519235 5 dpga_flat_0.sr_0.FILLER_0_20_27.VPWR
flabel metal1 174907 519714 174941 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_29.VGND
flabel metal1 174907 519170 174941 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_29.VPWR
flabel nwell 174907 519170 174941 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_29.VPB
flabel pwell 174907 519714 174941 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_29.VNB
rlabel comment 174878 519731 174878 519731 2 dpga_flat_0.sr_0.FILLER_0_20_29.decap_12
flabel metal1 176011 519714 176045 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_41.VGND
flabel metal1 176011 519170 176045 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_41.VPWR
flabel nwell 176011 519170 176045 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_41.VPB
flabel pwell 176011 519714 176045 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_41.VNB
rlabel comment 175982 519731 175982 519731 2 dpga_flat_0.sr_0.FILLER_0_20_41.decap_12
flabel metal1 174808 519178 174861 519207 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_20_108.VPWR
flabel metal1 174807 519711 174858 519749 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_20_108.VGND
rlabel comment 174786 519731 174786 519731 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_20_108.tapvpwrvgnd_1
rlabel metal1 174786 519683 174878 519779 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_20_108.VGND
rlabel metal1 174786 519139 174878 519235 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_20_108.VPWR
flabel metal1 176931 519714 176965 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_51.VGND
flabel metal1 176931 520258 176965 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_51.VPWR
flabel nwell 176931 520258 176965 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_51.VPB
flabel pwell 176931 519714 176965 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_51.VNB
rlabel comment 176902 519731 176902 519731 4 dpga_flat_0.sr_0.FILLER_0_19_51.decap_4
rlabel metal1 176902 519683 177270 519779 1 dpga_flat_0.sr_0.FILLER_0_19_51.VGND
rlabel metal1 176902 520227 177270 520323 1 dpga_flat_0.sr_0.FILLER_0_19_51.VPWR
flabel metal1 177292 520258 177328 520288 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_55.VPWR
flabel metal1 177292 519718 177328 519747 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_55.VGND
flabel nwell 177301 520265 177321 520282 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_55.VPB
flabel pwell 177298 519720 177322 519742 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_55.VNB
rlabel comment 177270 519731 177270 519731 4 dpga_flat_0.sr_0.FILLER_0_19_55.fill_1
rlabel metal1 177270 519683 177362 519779 1 dpga_flat_0.sr_0.FILLER_0_19_55.VGND
rlabel metal1 177270 520227 177362 520323 1 dpga_flat_0.sr_0.FILLER_0_19_55.VPWR
flabel metal1 177483 519714 177517 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_57.VGND
flabel metal1 177483 520258 177517 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_57.VPWR
flabel nwell 177483 520258 177517 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_57.VPB
flabel pwell 177483 519714 177517 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_57.VNB
rlabel comment 177454 519731 177454 519731 4 dpga_flat_0.sr_0.FILLER_0_19_57.decap_12
flabel metal1 177115 519714 177149 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_53.VGND
flabel metal1 177115 519170 177149 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_53.VPWR
flabel nwell 177115 519170 177149 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_53.VPB
flabel pwell 177115 519714 177149 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_53.VNB
rlabel comment 177086 519731 177086 519731 2 dpga_flat_0.sr_0.FILLER_0_20_53.decap_12
flabel metal1 177384 520255 177437 520284 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_19_106.VPWR
flabel metal1 177383 519713 177434 519751 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_19_106.VGND
rlabel comment 177362 519731 177362 519731 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_19_106.tapvpwrvgnd_1
rlabel metal1 177362 519683 177454 519779 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_19_106.VGND
rlabel metal1 177362 520227 177454 520323 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_19_106.VPWR
flabel metal1 178587 519714 178621 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_69.VGND
flabel metal1 178587 520258 178621 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_69.VPWR
flabel nwell 178587 520258 178621 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_69.VPB
flabel pwell 178587 519714 178621 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_69.VNB
rlabel comment 178558 519731 178558 519731 4 dpga_flat_0.sr_0.FILLER_0_19_69.decap_12
flabel metal1 179691 519714 179725 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_81.VGND
flabel metal1 179691 520258 179725 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_81.VPWR
flabel nwell 179691 520258 179725 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_81.VPB
flabel pwell 179691 519714 179725 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_81.VNB
rlabel comment 179662 519731 179662 519731 4 dpga_flat_0.sr_0.FILLER_0_19_81.decap_12
flabel metal1 178219 519714 178253 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_65.VGND
flabel metal1 178219 519170 178253 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_65.VPWR
flabel nwell 178219 519170 178253 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_65.VPB
flabel pwell 178219 519714 178253 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_65.VNB
rlabel comment 178190 519731 178190 519731 2 dpga_flat_0.sr_0.FILLER_0_20_65.decap_12
flabel metal1 179323 519170 179357 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_77.VPWR
flabel metal1 179323 519714 179357 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_77.VGND
flabel nwell 179323 519170 179357 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_77.VPB
flabel pwell 179323 519714 179357 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_77.VNB
rlabel comment 179294 519731 179294 519731 2 dpga_flat_0.sr_0.FILLER_0_20_77.decap_6
rlabel metal1 179294 519683 179846 519779 5 dpga_flat_0.sr_0.FILLER_0_20_77.VGND
rlabel metal1 179294 519139 179846 519235 5 dpga_flat_0.sr_0.FILLER_0_20_77.VPWR
flabel metal1 179868 519174 179904 519204 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_83.VPWR
flabel metal1 179868 519715 179904 519744 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_83.VGND
flabel nwell 179877 519180 179897 519197 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_83.VPB
flabel pwell 179874 519720 179898 519742 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_83.VNB
rlabel comment 179846 519731 179846 519731 2 dpga_flat_0.sr_0.FILLER_0_20_83.fill_1
rlabel metal1 179846 519683 179938 519779 5 dpga_flat_0.sr_0.FILLER_0_20_83.VGND
rlabel metal1 179846 519139 179938 519235 5 dpga_flat_0.sr_0.FILLER_0_20_83.VPWR
flabel metal1 180795 519714 180829 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_93.VGND
flabel metal1 180795 520258 180829 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_93.VPWR
flabel nwell 180795 520258 180829 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_93.VPB
flabel pwell 180795 519714 180829 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_93.VNB
rlabel comment 180766 519731 180766 519731 4 dpga_flat_0.sr_0.FILLER_0_19_93.decap_12
flabel metal1 180059 519714 180093 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_85.VGND
flabel metal1 180059 519170 180093 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_85.VPWR
flabel nwell 180059 519170 180093 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_85.VPB
flabel pwell 180059 519714 180093 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_85.VNB
rlabel comment 180030 519731 180030 519731 2 dpga_flat_0.sr_0.FILLER_0_20_85.decap_12
flabel metal1 181163 519714 181197 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_97.VGND
flabel metal1 181163 519170 181197 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_97.VPWR
flabel nwell 181163 519170 181197 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_97.VPB
flabel pwell 181163 519714 181197 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_97.VNB
rlabel comment 181134 519731 181134 519731 2 dpga_flat_0.sr_0.FILLER_0_20_97.decap_12
flabel metal1 179960 519178 180013 519207 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_20_109.VPWR
flabel metal1 179959 519711 180010 519749 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_20_109.VGND
rlabel comment 179938 519731 179938 519731 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_20_109.tapvpwrvgnd_1
rlabel metal1 179938 519683 180030 519779 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_20_109.VGND
rlabel metal1 179938 519139 180030 519235 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_20_109.VPWR
flabel metal1 181899 520258 181933 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_105.VPWR
flabel metal1 181899 519714 181933 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_105.VGND
flabel nwell 181899 520258 181933 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_105.VPB
flabel pwell 181899 519714 181933 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_105.VNB
rlabel comment 181870 519731 181870 519731 4 dpga_flat_0.sr_0.FILLER_0_19_105.decap_6
rlabel metal1 181870 519683 182422 519779 1 dpga_flat_0.sr_0.FILLER_0_19_105.VGND
rlabel metal1 181870 520227 182422 520323 1 dpga_flat_0.sr_0.FILLER_0_19_105.VPWR
flabel metal1 182444 520258 182480 520288 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_111.VPWR
flabel metal1 182444 519718 182480 519747 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_111.VGND
flabel nwell 182453 520265 182473 520282 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_111.VPB
flabel pwell 182450 519720 182474 519742 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_111.VNB
rlabel comment 182422 519731 182422 519731 4 dpga_flat_0.sr_0.FILLER_0_19_111.fill_1
rlabel metal1 182422 519683 182514 519779 1 dpga_flat_0.sr_0.FILLER_0_19_111.VGND
rlabel metal1 182422 520227 182514 520323 1 dpga_flat_0.sr_0.FILLER_0_19_111.VPWR
flabel metal1 182635 519714 182669 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_113.VGND
flabel metal1 182635 520258 182669 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_113.VPWR
flabel nwell 182635 520258 182669 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_113.VPB
flabel pwell 182635 519714 182669 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_113.VNB
rlabel comment 182606 519731 182606 519731 4 dpga_flat_0.sr_0.FILLER_0_19_113.decap_12
flabel metal1 183739 519714 183773 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_125.VGND
flabel metal1 183739 520258 183773 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_125.VPWR
flabel nwell 183739 520258 183773 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_125.VPB
flabel pwell 183739 519714 183773 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_125.VNB
rlabel comment 183710 519731 183710 519731 4 dpga_flat_0.sr_0.FILLER_0_19_125.decap_12
flabel metal1 182267 519714 182301 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_109.VGND
flabel metal1 182267 519170 182301 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_109.VPWR
flabel nwell 182267 519170 182301 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_109.VPB
flabel pwell 182267 519714 182301 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_109.VNB
rlabel comment 182238 519731 182238 519731 2 dpga_flat_0.sr_0.FILLER_0_20_109.decap_12
flabel metal1 183371 519714 183405 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_121.VGND
flabel metal1 183371 519170 183405 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_121.VPWR
flabel nwell 183371 519170 183405 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_121.VPB
flabel pwell 183371 519714 183405 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_121.VNB
rlabel comment 183342 519731 183342 519731 2 dpga_flat_0.sr_0.FILLER_0_20_121.decap_12
flabel metal1 182536 520255 182589 520284 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_19_107.VPWR
flabel metal1 182535 519713 182586 519751 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_19_107.VGND
rlabel comment 182514 519731 182514 519731 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_19_107.tapvpwrvgnd_1
rlabel metal1 182514 519683 182606 519779 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_19_107.VGND
rlabel metal1 182514 520227 182606 520323 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_19_107.VPWR
flabel metal1 184843 519714 184877 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_137.VGND
flabel metal1 184843 520258 184877 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_137.VPWR
flabel nwell 184843 520258 184877 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_137.VPB
flabel pwell 184843 519714 184877 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_137.VNB
rlabel comment 184814 519731 184814 519731 4 dpga_flat_0.sr_0.FILLER_0_19_137.decap_12
flabel metal1 184475 519170 184509 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_133.VPWR
flabel metal1 184475 519714 184509 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_133.VGND
flabel nwell 184475 519170 184509 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_133.VPB
flabel pwell 184475 519714 184509 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_133.VNB
rlabel comment 184446 519731 184446 519731 2 dpga_flat_0.sr_0.FILLER_0_20_133.decap_6
rlabel metal1 184446 519683 184998 519779 5 dpga_flat_0.sr_0.FILLER_0_20_133.VGND
rlabel metal1 184446 519139 184998 519235 5 dpga_flat_0.sr_0.FILLER_0_20_133.VPWR
flabel metal1 185020 519174 185056 519204 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_139.VPWR
flabel metal1 185020 519715 185056 519744 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_139.VGND
flabel nwell 185029 519180 185049 519197 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_139.VPB
flabel pwell 185026 519720 185050 519742 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_139.VNB
rlabel comment 184998 519731 184998 519731 2 dpga_flat_0.sr_0.FILLER_0_20_139.fill_1
rlabel metal1 184998 519683 185090 519779 5 dpga_flat_0.sr_0.FILLER_0_20_139.VGND
rlabel metal1 184998 519139 185090 519235 5 dpga_flat_0.sr_0.FILLER_0_20_139.VPWR
flabel metal1 185211 519714 185245 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_141.VGND
flabel metal1 185211 519170 185245 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_141.VPWR
flabel nwell 185211 519170 185245 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_141.VPB
flabel pwell 185211 519714 185245 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_141.VNB
rlabel comment 185182 519731 185182 519731 2 dpga_flat_0.sr_0.FILLER_0_20_141.decap_12
flabel metal1 185112 519178 185165 519207 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_20_110.VPWR
flabel metal1 185111 519711 185162 519749 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_20_110.VGND
rlabel comment 185090 519731 185090 519731 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_20_110.tapvpwrvgnd_1
rlabel metal1 185090 519683 185182 519779 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_20_110.VGND
rlabel metal1 185090 519139 185182 519235 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_20_110.VPWR
flabel metal1 185947 519714 185981 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_149.VGND
flabel metal1 185947 520258 185981 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_149.VPWR
flabel nwell 185947 520258 185981 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_149.VPB
flabel pwell 185947 519714 185981 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_149.VNB
rlabel comment 185918 519731 185918 519731 4 dpga_flat_0.sr_0.FILLER_0_19_149.decap_12
flabel metal1 187042 519717 187095 519749 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_161.VGND
flabel metal1 187043 520261 187095 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_161.VPWR
flabel nwell 187050 520266 187084 520284 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_161.VPB
flabel pwell 187053 519721 187085 519743 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_19_161.VNB
rlabel comment 187022 519731 187022 519731 4 dpga_flat_0.sr_0.FILLER_0_19_161.fill_2
rlabel metal1 187022 519683 187206 519779 1 dpga_flat_0.sr_0.FILLER_0_19_161.VGND
rlabel metal1 187022 520227 187206 520323 1 dpga_flat_0.sr_0.FILLER_0_19_161.VPWR
flabel metal1 186315 519170 186349 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_153.VPWR
flabel metal1 186315 519714 186349 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_153.VGND
flabel nwell 186315 519170 186349 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_153.VPB
flabel pwell 186315 519714 186349 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_153.VNB
rlabel comment 186286 519731 186286 519731 2 dpga_flat_0.sr_0.FILLER_0_20_153.decap_8
rlabel metal1 186286 519683 187022 519779 5 dpga_flat_0.sr_0.FILLER_0_20_153.VGND
rlabel metal1 186286 519139 187022 519235 5 dpga_flat_0.sr_0.FILLER_0_20_153.VPWR
flabel metal1 187042 519713 187095 519745 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_161.VGND
flabel metal1 187043 519170 187095 519201 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_161.VPWR
flabel nwell 187050 519178 187084 519196 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_161.VPB
flabel pwell 187053 519719 187085 519741 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_20_161.VNB
rlabel comment 187022 519731 187022 519731 2 dpga_flat_0.sr_0.FILLER_0_20_161.fill_2
rlabel metal1 187022 519683 187206 519779 5 dpga_flat_0.sr_0.FILLER_0_20_161.VGND
rlabel metal1 187022 519139 187206 519235 5 dpga_flat_0.sr_0.FILLER_0_20_161.VPWR
flabel metal1 187419 520258 187453 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_19_Right_19.VPWR
flabel metal1 187419 519714 187453 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_19_Right_19.VGND
flabel nwell 187419 520258 187453 520292 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_19_Right_19.VPB
flabel pwell 187419 519714 187453 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_19_Right_19.VNB
rlabel comment 187482 519731 187482 519731 6 dpga_flat_0.sr_0.PHY_EDGE_ROW_19_Right_19.decap_3
rlabel metal1 187206 519683 187482 519779 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_19_Right_19.VGND
rlabel metal1 187206 520227 187482 520323 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_19_Right_19.VPWR
flabel metal1 187419 519170 187453 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_20_Right_20.VPWR
flabel metal1 187419 519714 187453 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_20_Right_20.VGND
flabel nwell 187419 519170 187453 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_20_Right_20.VPB
flabel pwell 187419 519714 187453 519748 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_20_Right_20.VNB
rlabel comment 187482 519731 187482 519731 8 dpga_flat_0.sr_0.PHY_EDGE_ROW_20_Right_20.decap_3
rlabel metal1 187206 519683 187482 519779 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_20_Right_20.VGND
rlabel metal1 187206 519139 187482 519235 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_20_Right_20.VPWR
flabel metal1 172515 518626 172549 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_3.VGND
flabel metal1 172515 519170 172549 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_3.VPWR
flabel nwell 172515 519170 172549 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_3.VPB
flabel pwell 172515 518626 172549 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_3.VNB
rlabel comment 172486 518643 172486 518643 4 dpga_flat_0.sr_0.FILLER_0_21_3.decap_12
flabel metal1 173619 518626 173653 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_15.VGND
flabel metal1 173619 519170 173653 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_15.VPWR
flabel nwell 173619 519170 173653 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_15.VPB
flabel pwell 173619 518626 173653 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_15.VNB
rlabel comment 173590 518643 173590 518643 4 dpga_flat_0.sr_0.FILLER_0_21_15.decap_12
flabel metal1 172239 519170 172273 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_21_Left_49.VPWR
flabel metal1 172239 518626 172273 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_21_Left_49.VGND
flabel nwell 172239 519170 172273 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_21_Left_49.VPB
flabel pwell 172239 518626 172273 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_21_Left_49.VNB
rlabel comment 172210 518643 172210 518643 4 dpga_flat_0.sr_0.PHY_EDGE_ROW_21_Left_49.decap_3
rlabel metal1 172210 518595 172486 518691 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_21_Left_49.VGND
rlabel metal1 172210 519139 172486 519235 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_21_Left_49.VPWR
flabel metal1 174723 518626 174757 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_27.VGND
flabel metal1 174723 519170 174757 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_27.VPWR
flabel nwell 174723 519170 174757 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_27.VPB
flabel pwell 174723 518626 174757 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_27.VNB
rlabel comment 174694 518643 174694 518643 4 dpga_flat_0.sr_0.FILLER_0_21_27.decap_12
flabel metal1 175827 518626 175861 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_39.VGND
flabel metal1 175827 519170 175861 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_39.VPWR
flabel nwell 175827 519170 175861 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_39.VPB
flabel pwell 175827 518626 175861 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_39.VNB
rlabel comment 175798 518643 175798 518643 4 dpga_flat_0.sr_0.FILLER_0_21_39.decap_12
flabel metal1 176931 518626 176965 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_51.VGND
flabel metal1 176931 519170 176965 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_51.VPWR
flabel nwell 176931 519170 176965 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_51.VPB
flabel pwell 176931 518626 176965 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_51.VNB
rlabel comment 176902 518643 176902 518643 4 dpga_flat_0.sr_0.FILLER_0_21_51.decap_4
rlabel metal1 176902 518595 177270 518691 1 dpga_flat_0.sr_0.FILLER_0_21_51.VGND
rlabel metal1 176902 519139 177270 519235 1 dpga_flat_0.sr_0.FILLER_0_21_51.VPWR
flabel metal1 177292 519170 177328 519200 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_55.VPWR
flabel metal1 177292 518630 177328 518659 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_55.VGND
flabel nwell 177301 519177 177321 519194 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_55.VPB
flabel pwell 177298 518632 177322 518654 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_55.VNB
rlabel comment 177270 518643 177270 518643 4 dpga_flat_0.sr_0.FILLER_0_21_55.fill_1
rlabel metal1 177270 518595 177362 518691 1 dpga_flat_0.sr_0.FILLER_0_21_55.VGND
rlabel metal1 177270 519139 177362 519235 1 dpga_flat_0.sr_0.FILLER_0_21_55.VPWR
flabel metal1 177483 518626 177517 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_57.VGND
flabel metal1 177483 519170 177517 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_57.VPWR
flabel nwell 177483 519170 177517 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_57.VPB
flabel pwell 177483 518626 177517 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_57.VNB
rlabel comment 177454 518643 177454 518643 4 dpga_flat_0.sr_0.FILLER_0_21_57.decap_12
flabel metal1 177384 519167 177437 519196 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_21_111.VPWR
flabel metal1 177383 518625 177434 518663 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_21_111.VGND
rlabel comment 177362 518643 177362 518643 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_21_111.tapvpwrvgnd_1
rlabel metal1 177362 518595 177454 518691 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_21_111.VGND
rlabel metal1 177362 519139 177454 519235 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_21_111.VPWR
flabel metal1 178587 518626 178621 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_69.VGND
flabel metal1 178587 519170 178621 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_69.VPWR
flabel nwell 178587 519170 178621 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_69.VPB
flabel pwell 178587 518626 178621 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_69.VNB
rlabel comment 178558 518643 178558 518643 4 dpga_flat_0.sr_0.FILLER_0_21_69.decap_12
flabel metal1 179691 518626 179725 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_81.VGND
flabel metal1 179691 519170 179725 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_81.VPWR
flabel nwell 179691 519170 179725 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_81.VPB
flabel pwell 179691 518626 179725 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_81.VNB
rlabel comment 179662 518643 179662 518643 4 dpga_flat_0.sr_0.FILLER_0_21_81.decap_12
flabel metal1 180795 518626 180829 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_93.VGND
flabel metal1 180795 519170 180829 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_93.VPWR
flabel nwell 180795 519170 180829 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_93.VPB
flabel pwell 180795 518626 180829 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_93.VNB
rlabel comment 180766 518643 180766 518643 4 dpga_flat_0.sr_0.FILLER_0_21_93.decap_12
flabel metal1 181899 519170 181933 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_105.VPWR
flabel metal1 181899 518626 181933 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_105.VGND
flabel nwell 181899 519170 181933 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_105.VPB
flabel pwell 181899 518626 181933 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_105.VNB
rlabel comment 181870 518643 181870 518643 4 dpga_flat_0.sr_0.FILLER_0_21_105.decap_6
rlabel metal1 181870 518595 182422 518691 1 dpga_flat_0.sr_0.FILLER_0_21_105.VGND
rlabel metal1 181870 519139 182422 519235 1 dpga_flat_0.sr_0.FILLER_0_21_105.VPWR
flabel metal1 182444 519170 182480 519200 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_111.VPWR
flabel metal1 182444 518630 182480 518659 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_111.VGND
flabel nwell 182453 519177 182473 519194 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_111.VPB
flabel pwell 182450 518632 182474 518654 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_111.VNB
rlabel comment 182422 518643 182422 518643 4 dpga_flat_0.sr_0.FILLER_0_21_111.fill_1
rlabel metal1 182422 518595 182514 518691 1 dpga_flat_0.sr_0.FILLER_0_21_111.VGND
rlabel metal1 182422 519139 182514 519235 1 dpga_flat_0.sr_0.FILLER_0_21_111.VPWR
flabel metal1 182635 518626 182669 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_113.VGND
flabel metal1 182635 519170 182669 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_113.VPWR
flabel nwell 182635 519170 182669 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_113.VPB
flabel pwell 182635 518626 182669 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_113.VNB
rlabel comment 182606 518643 182606 518643 4 dpga_flat_0.sr_0.FILLER_0_21_113.decap_12
flabel metal1 183739 518626 183773 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_125.VGND
flabel metal1 183739 519170 183773 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_125.VPWR
flabel nwell 183739 519170 183773 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_125.VPB
flabel pwell 183739 518626 183773 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_125.VNB
rlabel comment 183710 518643 183710 518643 4 dpga_flat_0.sr_0.FILLER_0_21_125.decap_12
flabel metal1 182536 519167 182589 519196 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_21_112.VPWR
flabel metal1 182535 518625 182586 518663 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_21_112.VGND
rlabel comment 182514 518643 182514 518643 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_21_112.tapvpwrvgnd_1
rlabel metal1 182514 518595 182606 518691 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_21_112.VGND
rlabel metal1 182514 519139 182606 519235 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_21_112.VPWR
flabel metal1 184843 518626 184877 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_137.VGND
flabel metal1 184843 519170 184877 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_137.VPWR
flabel nwell 184843 519170 184877 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_137.VPB
flabel pwell 184843 518626 184877 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_137.VNB
rlabel comment 184814 518643 184814 518643 4 dpga_flat_0.sr_0.FILLER_0_21_137.decap_12
flabel metal1 185947 518626 185981 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_149.VGND
flabel metal1 185947 519170 185981 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_149.VPWR
flabel nwell 185947 519170 185981 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_149.VPB
flabel pwell 185947 518626 185981 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_149.VNB
rlabel comment 185918 518643 185918 518643 4 dpga_flat_0.sr_0.FILLER_0_21_149.decap_12
flabel metal1 187042 518629 187095 518661 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_161.VGND
flabel metal1 187043 519173 187095 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_161.VPWR
flabel nwell 187050 519178 187084 519196 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_161.VPB
flabel pwell 187053 518633 187085 518655 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_21_161.VNB
rlabel comment 187022 518643 187022 518643 4 dpga_flat_0.sr_0.FILLER_0_21_161.fill_2
rlabel metal1 187022 518595 187206 518691 1 dpga_flat_0.sr_0.FILLER_0_21_161.VGND
rlabel metal1 187022 519139 187206 519235 1 dpga_flat_0.sr_0.FILLER_0_21_161.VPWR
flabel metal1 187419 519170 187453 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_21_Right_21.VPWR
flabel metal1 187419 518626 187453 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_21_Right_21.VGND
flabel nwell 187419 519170 187453 519204 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_21_Right_21.VPB
flabel pwell 187419 518626 187453 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_21_Right_21.VNB
rlabel comment 187482 518643 187482 518643 6 dpga_flat_0.sr_0.PHY_EDGE_ROW_21_Right_21.decap_3
rlabel metal1 187206 518595 187482 518691 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_21_Right_21.VGND
rlabel metal1 187206 519139 187482 519235 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_21_Right_21.VPWR
flabel metal1 172515 518626 172549 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_3.VGND
flabel metal1 172515 518082 172549 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_3.VPWR
flabel nwell 172515 518082 172549 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_3.VPB
flabel pwell 172515 518626 172549 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_3.VNB
rlabel comment 172486 518643 172486 518643 2 dpga_flat_0.sr_0.FILLER_0_22_3.decap_12
flabel metal1 173619 518626 173653 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_15.VGND
flabel metal1 173619 518082 173653 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_15.VPWR
flabel nwell 173619 518082 173653 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_15.VPB
flabel pwell 173619 518626 173653 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_15.VNB
rlabel comment 173590 518643 173590 518643 2 dpga_flat_0.sr_0.FILLER_0_22_15.decap_12
flabel metal1 172239 518082 172273 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_22_Left_50.VPWR
flabel metal1 172239 518626 172273 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_22_Left_50.VGND
flabel nwell 172239 518082 172273 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_22_Left_50.VPB
flabel pwell 172239 518626 172273 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_22_Left_50.VNB
rlabel comment 172210 518643 172210 518643 2 dpga_flat_0.sr_0.PHY_EDGE_ROW_22_Left_50.decap_3
rlabel metal1 172210 518595 172486 518691 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_22_Left_50.VGND
rlabel metal1 172210 518051 172486 518147 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_22_Left_50.VPWR
flabel metal1 174716 518086 174752 518116 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_27.VPWR
flabel metal1 174716 518627 174752 518656 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_27.VGND
flabel nwell 174725 518092 174745 518109 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_27.VPB
flabel pwell 174722 518632 174746 518654 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_27.VNB
rlabel comment 174694 518643 174694 518643 2 dpga_flat_0.sr_0.FILLER_0_22_27.fill_1
rlabel metal1 174694 518595 174786 518691 5 dpga_flat_0.sr_0.FILLER_0_22_27.VGND
rlabel metal1 174694 518051 174786 518147 5 dpga_flat_0.sr_0.FILLER_0_22_27.VPWR
flabel metal1 174907 518626 174941 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_29.VGND
flabel metal1 174907 518082 174941 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_29.VPWR
flabel nwell 174907 518082 174941 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_29.VPB
flabel pwell 174907 518626 174941 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_29.VNB
rlabel comment 174878 518643 174878 518643 2 dpga_flat_0.sr_0.FILLER_0_22_29.decap_12
flabel metal1 176011 518626 176045 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_41.VGND
flabel metal1 176011 518082 176045 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_41.VPWR
flabel nwell 176011 518082 176045 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_41.VPB
flabel pwell 176011 518626 176045 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_41.VNB
rlabel comment 175982 518643 175982 518643 2 dpga_flat_0.sr_0.FILLER_0_22_41.decap_12
flabel metal1 174808 518090 174861 518119 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_22_113.VPWR
flabel metal1 174807 518623 174858 518661 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_22_113.VGND
rlabel comment 174786 518643 174786 518643 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_22_113.tapvpwrvgnd_1
rlabel metal1 174786 518595 174878 518691 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_22_113.VGND
rlabel metal1 174786 518051 174878 518147 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_22_113.VPWR
flabel metal1 177115 518626 177149 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_53.VGND
flabel metal1 177115 518082 177149 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_53.VPWR
flabel nwell 177115 518082 177149 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_53.VPB
flabel pwell 177115 518626 177149 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_53.VNB
rlabel comment 177086 518643 177086 518643 2 dpga_flat_0.sr_0.FILLER_0_22_53.decap_12
flabel metal1 178219 518626 178253 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_65.VGND
flabel metal1 178219 518082 178253 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_65.VPWR
flabel nwell 178219 518082 178253 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_65.VPB
flabel pwell 178219 518626 178253 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_65.VNB
rlabel comment 178190 518643 178190 518643 2 dpga_flat_0.sr_0.FILLER_0_22_65.decap_12
flabel metal1 179323 518082 179357 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_77.VPWR
flabel metal1 179323 518626 179357 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_77.VGND
flabel nwell 179323 518082 179357 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_77.VPB
flabel pwell 179323 518626 179357 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_77.VNB
rlabel comment 179294 518643 179294 518643 2 dpga_flat_0.sr_0.FILLER_0_22_77.decap_6
rlabel metal1 179294 518595 179846 518691 5 dpga_flat_0.sr_0.FILLER_0_22_77.VGND
rlabel metal1 179294 518051 179846 518147 5 dpga_flat_0.sr_0.FILLER_0_22_77.VPWR
flabel metal1 179868 518086 179904 518116 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_83.VPWR
flabel metal1 179868 518627 179904 518656 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_83.VGND
flabel nwell 179877 518092 179897 518109 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_83.VPB
flabel pwell 179874 518632 179898 518654 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_83.VNB
rlabel comment 179846 518643 179846 518643 2 dpga_flat_0.sr_0.FILLER_0_22_83.fill_1
rlabel metal1 179846 518595 179938 518691 5 dpga_flat_0.sr_0.FILLER_0_22_83.VGND
rlabel metal1 179846 518051 179938 518147 5 dpga_flat_0.sr_0.FILLER_0_22_83.VPWR
flabel metal1 180059 518626 180093 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_85.VGND
flabel metal1 180059 518082 180093 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_85.VPWR
flabel nwell 180059 518082 180093 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_85.VPB
flabel pwell 180059 518626 180093 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_85.VNB
rlabel comment 180030 518643 180030 518643 2 dpga_flat_0.sr_0.FILLER_0_22_85.decap_12
flabel metal1 181163 518626 181197 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_97.VGND
flabel metal1 181163 518082 181197 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_97.VPWR
flabel nwell 181163 518082 181197 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_97.VPB
flabel pwell 181163 518626 181197 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_97.VNB
rlabel comment 181134 518643 181134 518643 2 dpga_flat_0.sr_0.FILLER_0_22_97.decap_12
flabel metal1 179960 518090 180013 518119 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_22_114.VPWR
flabel metal1 179959 518623 180010 518661 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_22_114.VGND
rlabel comment 179938 518643 179938 518643 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_22_114.tapvpwrvgnd_1
rlabel metal1 179938 518595 180030 518691 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_22_114.VGND
rlabel metal1 179938 518051 180030 518147 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_22_114.VPWR
flabel metal1 182267 518626 182301 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_109.VGND
flabel metal1 182267 518082 182301 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_109.VPWR
flabel nwell 182267 518082 182301 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_109.VPB
flabel pwell 182267 518626 182301 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_109.VNB
rlabel comment 182238 518643 182238 518643 2 dpga_flat_0.sr_0.FILLER_0_22_109.decap_12
flabel metal1 183371 518626 183405 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_121.VGND
flabel metal1 183371 518082 183405 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_121.VPWR
flabel nwell 183371 518082 183405 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_121.VPB
flabel pwell 183371 518626 183405 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_121.VNB
rlabel comment 183342 518643 183342 518643 2 dpga_flat_0.sr_0.FILLER_0_22_121.decap_12
flabel metal1 184475 518082 184509 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_133.VPWR
flabel metal1 184475 518626 184509 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_133.VGND
flabel nwell 184475 518082 184509 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_133.VPB
flabel pwell 184475 518626 184509 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_133.VNB
rlabel comment 184446 518643 184446 518643 2 dpga_flat_0.sr_0.FILLER_0_22_133.decap_6
rlabel metal1 184446 518595 184998 518691 5 dpga_flat_0.sr_0.FILLER_0_22_133.VGND
rlabel metal1 184446 518051 184998 518147 5 dpga_flat_0.sr_0.FILLER_0_22_133.VPWR
flabel metal1 185020 518086 185056 518116 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_139.VPWR
flabel metal1 185020 518627 185056 518656 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_139.VGND
flabel nwell 185029 518092 185049 518109 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_139.VPB
flabel pwell 185026 518632 185050 518654 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_139.VNB
rlabel comment 184998 518643 184998 518643 2 dpga_flat_0.sr_0.FILLER_0_22_139.fill_1
rlabel metal1 184998 518595 185090 518691 5 dpga_flat_0.sr_0.FILLER_0_22_139.VGND
rlabel metal1 184998 518051 185090 518147 5 dpga_flat_0.sr_0.FILLER_0_22_139.VPWR
flabel metal1 185211 518626 185245 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_141.VGND
flabel metal1 185211 518082 185245 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_141.VPWR
flabel nwell 185211 518082 185245 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_141.VPB
flabel pwell 185211 518626 185245 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_141.VNB
rlabel comment 185182 518643 185182 518643 2 dpga_flat_0.sr_0.FILLER_0_22_141.decap_12
flabel metal1 185112 518090 185165 518119 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_22_115.VPWR
flabel metal1 185111 518623 185162 518661 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_22_115.VGND
rlabel comment 185090 518643 185090 518643 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_22_115.tapvpwrvgnd_1
rlabel metal1 185090 518595 185182 518691 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_22_115.VGND
rlabel metal1 185090 518051 185182 518147 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_22_115.VPWR
flabel metal1 186315 518082 186349 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_153.VPWR
flabel metal1 186315 518626 186349 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_153.VGND
flabel nwell 186315 518082 186349 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_153.VPB
flabel pwell 186315 518626 186349 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_153.VNB
rlabel comment 186286 518643 186286 518643 2 dpga_flat_0.sr_0.FILLER_0_22_153.decap_8
rlabel metal1 186286 518595 187022 518691 5 dpga_flat_0.sr_0.FILLER_0_22_153.VGND
rlabel metal1 186286 518051 187022 518147 5 dpga_flat_0.sr_0.FILLER_0_22_153.VPWR
flabel metal1 187042 518625 187095 518657 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_161.VGND
flabel metal1 187043 518082 187095 518113 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_161.VPWR
flabel nwell 187050 518090 187084 518108 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_161.VPB
flabel pwell 187053 518631 187085 518653 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_22_161.VNB
rlabel comment 187022 518643 187022 518643 2 dpga_flat_0.sr_0.FILLER_0_22_161.fill_2
rlabel metal1 187022 518595 187206 518691 5 dpga_flat_0.sr_0.FILLER_0_22_161.VGND
rlabel metal1 187022 518051 187206 518147 5 dpga_flat_0.sr_0.FILLER_0_22_161.VPWR
flabel metal1 187419 518082 187453 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_22_Right_22.VPWR
flabel metal1 187419 518626 187453 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_22_Right_22.VGND
flabel nwell 187419 518082 187453 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_22_Right_22.VPB
flabel pwell 187419 518626 187453 518660 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_22_Right_22.VNB
rlabel comment 187482 518643 187482 518643 8 dpga_flat_0.sr_0.PHY_EDGE_ROW_22_Right_22.decap_3
rlabel metal1 187206 518595 187482 518691 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_22_Right_22.VGND
rlabel metal1 187206 518051 187482 518147 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_22_Right_22.VPWR
flabel metal1 172515 517538 172549 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_3.VGND
flabel metal1 172515 518082 172549 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_3.VPWR
flabel nwell 172515 518082 172549 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_3.VPB
flabel pwell 172515 517538 172549 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_3.VNB
rlabel comment 172486 517555 172486 517555 4 dpga_flat_0.sr_0.FILLER_0_23_3.decap_12
flabel metal1 173619 517538 173653 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_15.VGND
flabel metal1 173619 518082 173653 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_15.VPWR
flabel nwell 173619 518082 173653 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_15.VPB
flabel pwell 173619 517538 173653 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_15.VNB
rlabel comment 173590 517555 173590 517555 4 dpga_flat_0.sr_0.FILLER_0_23_15.decap_12
flabel metal1 172239 518082 172273 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_23_Left_51.VPWR
flabel metal1 172239 517538 172273 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_23_Left_51.VGND
flabel nwell 172239 518082 172273 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_23_Left_51.VPB
flabel pwell 172239 517538 172273 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_23_Left_51.VNB
rlabel comment 172210 517555 172210 517555 4 dpga_flat_0.sr_0.PHY_EDGE_ROW_23_Left_51.decap_3
rlabel metal1 172210 517507 172486 517603 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_23_Left_51.VGND
rlabel metal1 172210 518051 172486 518147 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_23_Left_51.VPWR
flabel metal1 174723 517538 174757 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_27.VGND
flabel metal1 174723 518082 174757 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_27.VPWR
flabel nwell 174723 518082 174757 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_27.VPB
flabel pwell 174723 517538 174757 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_27.VNB
rlabel comment 174694 517555 174694 517555 4 dpga_flat_0.sr_0.FILLER_0_23_27.decap_12
flabel metal1 175827 517538 175861 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_39.VGND
flabel metal1 175827 518082 175861 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_39.VPWR
flabel nwell 175827 518082 175861 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_39.VPB
flabel pwell 175827 517538 175861 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_39.VNB
rlabel comment 175798 517555 175798 517555 4 dpga_flat_0.sr_0.FILLER_0_23_39.decap_12
flabel metal1 176931 517538 176965 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_51.VGND
flabel metal1 176931 518082 176965 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_51.VPWR
flabel nwell 176931 518082 176965 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_51.VPB
flabel pwell 176931 517538 176965 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_51.VNB
rlabel comment 176902 517555 176902 517555 4 dpga_flat_0.sr_0.FILLER_0_23_51.decap_4
rlabel metal1 176902 517507 177270 517603 1 dpga_flat_0.sr_0.FILLER_0_23_51.VGND
rlabel metal1 176902 518051 177270 518147 1 dpga_flat_0.sr_0.FILLER_0_23_51.VPWR
flabel metal1 177292 518082 177328 518112 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_55.VPWR
flabel metal1 177292 517542 177328 517571 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_55.VGND
flabel nwell 177301 518089 177321 518106 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_55.VPB
flabel pwell 177298 517544 177322 517566 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_55.VNB
rlabel comment 177270 517555 177270 517555 4 dpga_flat_0.sr_0.FILLER_0_23_55.fill_1
rlabel metal1 177270 517507 177362 517603 1 dpga_flat_0.sr_0.FILLER_0_23_55.VGND
rlabel metal1 177270 518051 177362 518147 1 dpga_flat_0.sr_0.FILLER_0_23_55.VPWR
flabel metal1 177483 517538 177517 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_57.VGND
flabel metal1 177483 518082 177517 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_57.VPWR
flabel nwell 177483 518082 177517 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_57.VPB
flabel pwell 177483 517538 177517 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_57.VNB
rlabel comment 177454 517555 177454 517555 4 dpga_flat_0.sr_0.FILLER_0_23_57.decap_12
flabel metal1 177384 518079 177437 518108 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_23_116.VPWR
flabel metal1 177383 517537 177434 517575 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_23_116.VGND
rlabel comment 177362 517555 177362 517555 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_23_116.tapvpwrvgnd_1
rlabel metal1 177362 517507 177454 517603 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_23_116.VGND
rlabel metal1 177362 518051 177454 518147 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_23_116.VPWR
flabel metal1 178587 517538 178621 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_69.VGND
flabel metal1 178587 518082 178621 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_69.VPWR
flabel nwell 178587 518082 178621 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_69.VPB
flabel pwell 178587 517538 178621 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_69.VNB
rlabel comment 178558 517555 178558 517555 4 dpga_flat_0.sr_0.FILLER_0_23_69.decap_12
flabel metal1 179691 517538 179725 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_81.VGND
flabel metal1 179691 518082 179725 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_81.VPWR
flabel nwell 179691 518082 179725 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_81.VPB
flabel pwell 179691 517538 179725 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_81.VNB
rlabel comment 179662 517555 179662 517555 4 dpga_flat_0.sr_0.FILLER_0_23_81.decap_12
flabel metal1 180795 517538 180829 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_93.VGND
flabel metal1 180795 518082 180829 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_93.VPWR
flabel nwell 180795 518082 180829 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_93.VPB
flabel pwell 180795 517538 180829 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_93.VNB
rlabel comment 180766 517555 180766 517555 4 dpga_flat_0.sr_0.FILLER_0_23_93.decap_12
flabel metal1 181899 518082 181933 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_105.VPWR
flabel metal1 181899 517538 181933 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_105.VGND
flabel nwell 181899 518082 181933 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_105.VPB
flabel pwell 181899 517538 181933 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_105.VNB
rlabel comment 181870 517555 181870 517555 4 dpga_flat_0.sr_0.FILLER_0_23_105.decap_6
rlabel metal1 181870 517507 182422 517603 1 dpga_flat_0.sr_0.FILLER_0_23_105.VGND
rlabel metal1 181870 518051 182422 518147 1 dpga_flat_0.sr_0.FILLER_0_23_105.VPWR
flabel metal1 182444 518082 182480 518112 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_111.VPWR
flabel metal1 182444 517542 182480 517571 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_111.VGND
flabel nwell 182453 518089 182473 518106 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_111.VPB
flabel pwell 182450 517544 182474 517566 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_111.VNB
rlabel comment 182422 517555 182422 517555 4 dpga_flat_0.sr_0.FILLER_0_23_111.fill_1
rlabel metal1 182422 517507 182514 517603 1 dpga_flat_0.sr_0.FILLER_0_23_111.VGND
rlabel metal1 182422 518051 182514 518147 1 dpga_flat_0.sr_0.FILLER_0_23_111.VPWR
flabel metal1 182635 517538 182669 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_113.VGND
flabel metal1 182635 518082 182669 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_113.VPWR
flabel nwell 182635 518082 182669 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_113.VPB
flabel pwell 182635 517538 182669 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_113.VNB
rlabel comment 182606 517555 182606 517555 4 dpga_flat_0.sr_0.FILLER_0_23_113.decap_12
flabel metal1 183739 517538 183773 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_125.VGND
flabel metal1 183739 518082 183773 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_125.VPWR
flabel nwell 183739 518082 183773 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_125.VPB
flabel pwell 183739 517538 183773 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_125.VNB
rlabel comment 183710 517555 183710 517555 4 dpga_flat_0.sr_0.FILLER_0_23_125.decap_12
flabel metal1 182536 518079 182589 518108 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_23_117.VPWR
flabel metal1 182535 517537 182586 517575 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_23_117.VGND
rlabel comment 182514 517555 182514 517555 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_23_117.tapvpwrvgnd_1
rlabel metal1 182514 517507 182606 517603 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_23_117.VGND
rlabel metal1 182514 518051 182606 518147 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_23_117.VPWR
flabel metal1 184843 517538 184877 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_137.VGND
flabel metal1 184843 518082 184877 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_137.VPWR
flabel nwell 184843 518082 184877 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_137.VPB
flabel pwell 184843 517538 184877 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_137.VNB
rlabel comment 184814 517555 184814 517555 4 dpga_flat_0.sr_0.FILLER_0_23_137.decap_12
flabel metal1 185947 517538 185981 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_149.VGND
flabel metal1 185947 518082 185981 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_149.VPWR
flabel nwell 185947 518082 185981 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_149.VPB
flabel pwell 185947 517538 185981 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_149.VNB
rlabel comment 185918 517555 185918 517555 4 dpga_flat_0.sr_0.FILLER_0_23_149.decap_12
flabel metal1 187042 517541 187095 517573 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_161.VGND
flabel metal1 187043 518085 187095 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_161.VPWR
flabel nwell 187050 518090 187084 518108 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_161.VPB
flabel pwell 187053 517545 187085 517567 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_23_161.VNB
rlabel comment 187022 517555 187022 517555 4 dpga_flat_0.sr_0.FILLER_0_23_161.fill_2
rlabel metal1 187022 517507 187206 517603 1 dpga_flat_0.sr_0.FILLER_0_23_161.VGND
rlabel metal1 187022 518051 187206 518147 1 dpga_flat_0.sr_0.FILLER_0_23_161.VPWR
flabel metal1 187419 518082 187453 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_23_Right_23.VPWR
flabel metal1 187419 517538 187453 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_23_Right_23.VGND
flabel nwell 187419 518082 187453 518116 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_23_Right_23.VPB
flabel pwell 187419 517538 187453 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_23_Right_23.VNB
rlabel comment 187482 517555 187482 517555 6 dpga_flat_0.sr_0.PHY_EDGE_ROW_23_Right_23.decap_3
rlabel metal1 187206 517507 187482 517603 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_23_Right_23.VGND
rlabel metal1 187206 518051 187482 518147 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_23_Right_23.VPWR
flabel metal1 172515 517538 172549 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_3.VGND
flabel metal1 172515 516994 172549 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_3.VPWR
flabel nwell 172515 516994 172549 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_3.VPB
flabel pwell 172515 517538 172549 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_3.VNB
rlabel comment 172486 517555 172486 517555 2 dpga_flat_0.sr_0.FILLER_0_24_3.decap_12
flabel metal1 173619 517538 173653 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_15.VGND
flabel metal1 173619 516994 173653 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_15.VPWR
flabel nwell 173619 516994 173653 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_15.VPB
flabel pwell 173619 517538 173653 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_15.VNB
rlabel comment 173590 517555 173590 517555 2 dpga_flat_0.sr_0.FILLER_0_24_15.decap_12
flabel metal1 172239 516994 172273 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_24_Left_52.VPWR
flabel metal1 172239 517538 172273 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_24_Left_52.VGND
flabel nwell 172239 516994 172273 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_24_Left_52.VPB
flabel pwell 172239 517538 172273 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_24_Left_52.VNB
rlabel comment 172210 517555 172210 517555 2 dpga_flat_0.sr_0.PHY_EDGE_ROW_24_Left_52.decap_3
rlabel metal1 172210 517507 172486 517603 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_24_Left_52.VGND
rlabel metal1 172210 516963 172486 517059 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_24_Left_52.VPWR
flabel metal1 174716 516998 174752 517028 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_27.VPWR
flabel metal1 174716 517539 174752 517568 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_27.VGND
flabel nwell 174725 517004 174745 517021 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_27.VPB
flabel pwell 174722 517544 174746 517566 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_27.VNB
rlabel comment 174694 517555 174694 517555 2 dpga_flat_0.sr_0.FILLER_0_24_27.fill_1
rlabel metal1 174694 517507 174786 517603 5 dpga_flat_0.sr_0.FILLER_0_24_27.VGND
rlabel metal1 174694 516963 174786 517059 5 dpga_flat_0.sr_0.FILLER_0_24_27.VPWR
flabel metal1 174907 517538 174941 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_29.VGND
flabel metal1 174907 516994 174941 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_29.VPWR
flabel nwell 174907 516994 174941 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_29.VPB
flabel pwell 174907 517538 174941 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_29.VNB
rlabel comment 174878 517555 174878 517555 2 dpga_flat_0.sr_0.FILLER_0_24_29.decap_12
flabel metal1 176011 517538 176045 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_41.VGND
flabel metal1 176011 516994 176045 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_41.VPWR
flabel nwell 176011 516994 176045 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_41.VPB
flabel pwell 176011 517538 176045 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_41.VNB
rlabel comment 175982 517555 175982 517555 2 dpga_flat_0.sr_0.FILLER_0_24_41.decap_12
flabel metal1 174808 517002 174861 517031 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_24_118.VPWR
flabel metal1 174807 517535 174858 517573 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_24_118.VGND
rlabel comment 174786 517555 174786 517555 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_24_118.tapvpwrvgnd_1
rlabel metal1 174786 517507 174878 517603 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_24_118.VGND
rlabel metal1 174786 516963 174878 517059 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_24_118.VPWR
flabel metal1 177115 517538 177149 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_53.VGND
flabel metal1 177115 516994 177149 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_53.VPWR
flabel nwell 177115 516994 177149 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_53.VPB
flabel pwell 177115 517538 177149 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_53.VNB
rlabel comment 177086 517555 177086 517555 2 dpga_flat_0.sr_0.FILLER_0_24_53.decap_12
flabel metal1 178219 517538 178253 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_65.VGND
flabel metal1 178219 516994 178253 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_65.VPWR
flabel nwell 178219 516994 178253 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_65.VPB
flabel pwell 178219 517538 178253 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_65.VNB
rlabel comment 178190 517555 178190 517555 2 dpga_flat_0.sr_0.FILLER_0_24_65.decap_12
flabel metal1 179323 516994 179357 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_77.VPWR
flabel metal1 179323 517538 179357 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_77.VGND
flabel nwell 179323 516994 179357 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_77.VPB
flabel pwell 179323 517538 179357 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_77.VNB
rlabel comment 179294 517555 179294 517555 2 dpga_flat_0.sr_0.FILLER_0_24_77.decap_6
rlabel metal1 179294 517507 179846 517603 5 dpga_flat_0.sr_0.FILLER_0_24_77.VGND
rlabel metal1 179294 516963 179846 517059 5 dpga_flat_0.sr_0.FILLER_0_24_77.VPWR
flabel metal1 179868 516998 179904 517028 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_83.VPWR
flabel metal1 179868 517539 179904 517568 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_83.VGND
flabel nwell 179877 517004 179897 517021 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_83.VPB
flabel pwell 179874 517544 179898 517566 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_83.VNB
rlabel comment 179846 517555 179846 517555 2 dpga_flat_0.sr_0.FILLER_0_24_83.fill_1
rlabel metal1 179846 517507 179938 517603 5 dpga_flat_0.sr_0.FILLER_0_24_83.VGND
rlabel metal1 179846 516963 179938 517059 5 dpga_flat_0.sr_0.FILLER_0_24_83.VPWR
flabel metal1 180059 517538 180093 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_85.VGND
flabel metal1 180059 516994 180093 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_85.VPWR
flabel nwell 180059 516994 180093 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_85.VPB
flabel pwell 180059 517538 180093 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_85.VNB
rlabel comment 180030 517555 180030 517555 2 dpga_flat_0.sr_0.FILLER_0_24_85.decap_12
flabel metal1 181163 517538 181197 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_97.VGND
flabel metal1 181163 516994 181197 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_97.VPWR
flabel nwell 181163 516994 181197 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_97.VPB
flabel pwell 181163 517538 181197 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_97.VNB
rlabel comment 181134 517555 181134 517555 2 dpga_flat_0.sr_0.FILLER_0_24_97.decap_12
flabel metal1 179960 517002 180013 517031 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_24_119.VPWR
flabel metal1 179959 517535 180010 517573 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_24_119.VGND
rlabel comment 179938 517555 179938 517555 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_24_119.tapvpwrvgnd_1
rlabel metal1 179938 517507 180030 517603 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_24_119.VGND
rlabel metal1 179938 516963 180030 517059 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_24_119.VPWR
flabel metal1 182267 517538 182301 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_109.VGND
flabel metal1 182267 516994 182301 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_109.VPWR
flabel nwell 182267 516994 182301 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_109.VPB
flabel pwell 182267 517538 182301 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_109.VNB
rlabel comment 182238 517555 182238 517555 2 dpga_flat_0.sr_0.FILLER_0_24_109.decap_12
flabel metal1 183371 517538 183405 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_121.VGND
flabel metal1 183371 516994 183405 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_121.VPWR
flabel nwell 183371 516994 183405 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_121.VPB
flabel pwell 183371 517538 183405 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_121.VNB
rlabel comment 183342 517555 183342 517555 2 dpga_flat_0.sr_0.FILLER_0_24_121.decap_12
flabel metal1 184475 516994 184509 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_133.VPWR
flabel metal1 184475 517538 184509 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_133.VGND
flabel nwell 184475 516994 184509 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_133.VPB
flabel pwell 184475 517538 184509 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_133.VNB
rlabel comment 184446 517555 184446 517555 2 dpga_flat_0.sr_0.FILLER_0_24_133.decap_6
rlabel metal1 184446 517507 184998 517603 5 dpga_flat_0.sr_0.FILLER_0_24_133.VGND
rlabel metal1 184446 516963 184998 517059 5 dpga_flat_0.sr_0.FILLER_0_24_133.VPWR
flabel metal1 185020 516998 185056 517028 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_139.VPWR
flabel metal1 185020 517539 185056 517568 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_139.VGND
flabel nwell 185029 517004 185049 517021 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_139.VPB
flabel pwell 185026 517544 185050 517566 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_139.VNB
rlabel comment 184998 517555 184998 517555 2 dpga_flat_0.sr_0.FILLER_0_24_139.fill_1
rlabel metal1 184998 517507 185090 517603 5 dpga_flat_0.sr_0.FILLER_0_24_139.VGND
rlabel metal1 184998 516963 185090 517059 5 dpga_flat_0.sr_0.FILLER_0_24_139.VPWR
flabel metal1 185211 517538 185245 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_141.VGND
flabel metal1 185211 516994 185245 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_141.VPWR
flabel nwell 185211 516994 185245 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_141.VPB
flabel pwell 185211 517538 185245 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_141.VNB
rlabel comment 185182 517555 185182 517555 2 dpga_flat_0.sr_0.FILLER_0_24_141.decap_12
flabel metal1 185112 517002 185165 517031 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_24_120.VPWR
flabel metal1 185111 517535 185162 517573 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_24_120.VGND
rlabel comment 185090 517555 185090 517555 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_24_120.tapvpwrvgnd_1
rlabel metal1 185090 517507 185182 517603 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_24_120.VGND
rlabel metal1 185090 516963 185182 517059 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_24_120.VPWR
flabel metal1 186315 516994 186349 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_153.VPWR
flabel metal1 186315 517538 186349 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_153.VGND
flabel nwell 186315 516994 186349 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_153.VPB
flabel pwell 186315 517538 186349 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_153.VNB
rlabel comment 186286 517555 186286 517555 2 dpga_flat_0.sr_0.FILLER_0_24_153.decap_8
rlabel metal1 186286 517507 187022 517603 5 dpga_flat_0.sr_0.FILLER_0_24_153.VGND
rlabel metal1 186286 516963 187022 517059 5 dpga_flat_0.sr_0.FILLER_0_24_153.VPWR
flabel metal1 187042 517537 187095 517569 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_161.VGND
flabel metal1 187043 516994 187095 517025 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_161.VPWR
flabel nwell 187050 517002 187084 517020 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_161.VPB
flabel pwell 187053 517543 187085 517565 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_24_161.VNB
rlabel comment 187022 517555 187022 517555 2 dpga_flat_0.sr_0.FILLER_0_24_161.fill_2
rlabel metal1 187022 517507 187206 517603 5 dpga_flat_0.sr_0.FILLER_0_24_161.VGND
rlabel metal1 187022 516963 187206 517059 5 dpga_flat_0.sr_0.FILLER_0_24_161.VPWR
flabel metal1 187419 516994 187453 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_24_Right_24.VPWR
flabel metal1 187419 517538 187453 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_24_Right_24.VGND
flabel nwell 187419 516994 187453 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_24_Right_24.VPB
flabel pwell 187419 517538 187453 517572 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_24_Right_24.VNB
rlabel comment 187482 517555 187482 517555 8 dpga_flat_0.sr_0.PHY_EDGE_ROW_24_Right_24.decap_3
rlabel metal1 187206 517507 187482 517603 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_24_Right_24.VGND
rlabel metal1 187206 516963 187482 517059 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_24_Right_24.VPWR
flabel metal1 172515 516450 172549 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_3.VGND
flabel metal1 172515 516994 172549 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_3.VPWR
flabel nwell 172515 516994 172549 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_3.VPB
flabel pwell 172515 516450 172549 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_3.VNB
rlabel comment 172486 516467 172486 516467 4 dpga_flat_0.sr_0.FILLER_0_25_3.decap_12
flabel metal1 173619 516450 173653 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_15.VGND
flabel metal1 173619 516994 173653 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_15.VPWR
flabel nwell 173619 516994 173653 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_15.VPB
flabel pwell 173619 516450 173653 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_15.VNB
rlabel comment 173590 516467 173590 516467 4 dpga_flat_0.sr_0.FILLER_0_25_15.decap_12
flabel metal1 172239 516994 172273 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_25_Left_53.VPWR
flabel metal1 172239 516450 172273 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_25_Left_53.VGND
flabel nwell 172239 516994 172273 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_25_Left_53.VPB
flabel pwell 172239 516450 172273 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_25_Left_53.VNB
rlabel comment 172210 516467 172210 516467 4 dpga_flat_0.sr_0.PHY_EDGE_ROW_25_Left_53.decap_3
rlabel metal1 172210 516419 172486 516515 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_25_Left_53.VGND
rlabel metal1 172210 516963 172486 517059 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_25_Left_53.VPWR
flabel metal1 174723 516450 174757 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_27.VGND
flabel metal1 174723 516994 174757 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_27.VPWR
flabel nwell 174723 516994 174757 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_27.VPB
flabel pwell 174723 516450 174757 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_27.VNB
rlabel comment 174694 516467 174694 516467 4 dpga_flat_0.sr_0.FILLER_0_25_27.decap_12
flabel metal1 175827 516450 175861 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_39.VGND
flabel metal1 175827 516994 175861 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_39.VPWR
flabel nwell 175827 516994 175861 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_39.VPB
flabel pwell 175827 516450 175861 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_39.VNB
rlabel comment 175798 516467 175798 516467 4 dpga_flat_0.sr_0.FILLER_0_25_39.decap_12
flabel metal1 176931 516450 176965 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_51.VGND
flabel metal1 176931 516994 176965 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_51.VPWR
flabel nwell 176931 516994 176965 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_51.VPB
flabel pwell 176931 516450 176965 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_51.VNB
rlabel comment 176902 516467 176902 516467 4 dpga_flat_0.sr_0.FILLER_0_25_51.decap_4
rlabel metal1 176902 516419 177270 516515 1 dpga_flat_0.sr_0.FILLER_0_25_51.VGND
rlabel metal1 176902 516963 177270 517059 1 dpga_flat_0.sr_0.FILLER_0_25_51.VPWR
flabel metal1 177292 516994 177328 517024 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_55.VPWR
flabel metal1 177292 516454 177328 516483 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_55.VGND
flabel nwell 177301 517001 177321 517018 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_55.VPB
flabel pwell 177298 516456 177322 516478 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_55.VNB
rlabel comment 177270 516467 177270 516467 4 dpga_flat_0.sr_0.FILLER_0_25_55.fill_1
rlabel metal1 177270 516419 177362 516515 1 dpga_flat_0.sr_0.FILLER_0_25_55.VGND
rlabel metal1 177270 516963 177362 517059 1 dpga_flat_0.sr_0.FILLER_0_25_55.VPWR
flabel metal1 177483 516450 177517 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_57.VGND
flabel metal1 177483 516994 177517 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_57.VPWR
flabel nwell 177483 516994 177517 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_57.VPB
flabel pwell 177483 516450 177517 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_57.VNB
rlabel comment 177454 516467 177454 516467 4 dpga_flat_0.sr_0.FILLER_0_25_57.decap_12
flabel metal1 177384 516991 177437 517020 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_25_121.VPWR
flabel metal1 177383 516449 177434 516487 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_25_121.VGND
rlabel comment 177362 516467 177362 516467 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_25_121.tapvpwrvgnd_1
rlabel metal1 177362 516419 177454 516515 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_25_121.VGND
rlabel metal1 177362 516963 177454 517059 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_25_121.VPWR
flabel metal1 178587 516450 178621 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_69.VGND
flabel metal1 178587 516994 178621 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_69.VPWR
flabel nwell 178587 516994 178621 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_69.VPB
flabel pwell 178587 516450 178621 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_69.VNB
rlabel comment 178558 516467 178558 516467 4 dpga_flat_0.sr_0.FILLER_0_25_69.decap_12
flabel metal1 179691 516450 179725 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_81.VGND
flabel metal1 179691 516994 179725 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_81.VPWR
flabel nwell 179691 516994 179725 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_81.VPB
flabel pwell 179691 516450 179725 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_81.VNB
rlabel comment 179662 516467 179662 516467 4 dpga_flat_0.sr_0.FILLER_0_25_81.decap_12
flabel metal1 180795 516450 180829 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_93.VGND
flabel metal1 180795 516994 180829 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_93.VPWR
flabel nwell 180795 516994 180829 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_93.VPB
flabel pwell 180795 516450 180829 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_93.VNB
rlabel comment 180766 516467 180766 516467 4 dpga_flat_0.sr_0.FILLER_0_25_93.decap_12
flabel metal1 181899 516994 181933 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_105.VPWR
flabel metal1 181899 516450 181933 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_105.VGND
flabel nwell 181899 516994 181933 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_105.VPB
flabel pwell 181899 516450 181933 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_105.VNB
rlabel comment 181870 516467 181870 516467 4 dpga_flat_0.sr_0.FILLER_0_25_105.decap_6
rlabel metal1 181870 516419 182422 516515 1 dpga_flat_0.sr_0.FILLER_0_25_105.VGND
rlabel metal1 181870 516963 182422 517059 1 dpga_flat_0.sr_0.FILLER_0_25_105.VPWR
flabel metal1 182444 516994 182480 517024 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_111.VPWR
flabel metal1 182444 516454 182480 516483 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_111.VGND
flabel nwell 182453 517001 182473 517018 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_111.VPB
flabel pwell 182450 516456 182474 516478 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_111.VNB
rlabel comment 182422 516467 182422 516467 4 dpga_flat_0.sr_0.FILLER_0_25_111.fill_1
rlabel metal1 182422 516419 182514 516515 1 dpga_flat_0.sr_0.FILLER_0_25_111.VGND
rlabel metal1 182422 516963 182514 517059 1 dpga_flat_0.sr_0.FILLER_0_25_111.VPWR
flabel metal1 182635 516450 182669 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_113.VGND
flabel metal1 182635 516994 182669 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_113.VPWR
flabel nwell 182635 516994 182669 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_113.VPB
flabel pwell 182635 516450 182669 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_113.VNB
rlabel comment 182606 516467 182606 516467 4 dpga_flat_0.sr_0.FILLER_0_25_113.decap_12
flabel metal1 183739 516450 183773 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_125.VGND
flabel metal1 183739 516994 183773 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_125.VPWR
flabel nwell 183739 516994 183773 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_125.VPB
flabel pwell 183739 516450 183773 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_125.VNB
rlabel comment 183710 516467 183710 516467 4 dpga_flat_0.sr_0.FILLER_0_25_125.decap_12
flabel metal1 182536 516991 182589 517020 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_25_122.VPWR
flabel metal1 182535 516449 182586 516487 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_25_122.VGND
rlabel comment 182514 516467 182514 516467 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_25_122.tapvpwrvgnd_1
rlabel metal1 182514 516419 182606 516515 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_25_122.VGND
rlabel metal1 182514 516963 182606 517059 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_25_122.VPWR
flabel metal1 184843 516450 184877 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_137.VGND
flabel metal1 184843 516994 184877 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_137.VPWR
flabel nwell 184843 516994 184877 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_137.VPB
flabel pwell 184843 516450 184877 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_137.VNB
rlabel comment 184814 516467 184814 516467 4 dpga_flat_0.sr_0.FILLER_0_25_137.decap_12
flabel metal1 185947 516450 185981 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_149.VGND
flabel metal1 185947 516994 185981 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_149.VPWR
flabel nwell 185947 516994 185981 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_149.VPB
flabel pwell 185947 516450 185981 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_149.VNB
rlabel comment 185918 516467 185918 516467 4 dpga_flat_0.sr_0.FILLER_0_25_149.decap_12
flabel metal1 187042 516453 187095 516485 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_161.VGND
flabel metal1 187043 516997 187095 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_161.VPWR
flabel nwell 187050 517002 187084 517020 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_161.VPB
flabel pwell 187053 516457 187085 516479 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_25_161.VNB
rlabel comment 187022 516467 187022 516467 4 dpga_flat_0.sr_0.FILLER_0_25_161.fill_2
rlabel metal1 187022 516419 187206 516515 1 dpga_flat_0.sr_0.FILLER_0_25_161.VGND
rlabel metal1 187022 516963 187206 517059 1 dpga_flat_0.sr_0.FILLER_0_25_161.VPWR
flabel metal1 187419 516994 187453 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_25_Right_25.VPWR
flabel metal1 187419 516450 187453 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_25_Right_25.VGND
flabel nwell 187419 516994 187453 517028 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_25_Right_25.VPB
flabel pwell 187419 516450 187453 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_25_Right_25.VNB
rlabel comment 187482 516467 187482 516467 6 dpga_flat_0.sr_0.PHY_EDGE_ROW_25_Right_25.decap_3
rlabel metal1 187206 516419 187482 516515 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_25_Right_25.VGND
rlabel metal1 187206 516963 187482 517059 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_25_Right_25.VPWR
flabel metal1 172515 516450 172549 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_3.VGND
flabel metal1 172515 515906 172549 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_3.VPWR
flabel nwell 172515 515906 172549 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_3.VPB
flabel pwell 172515 516450 172549 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_3.VNB
rlabel comment 172486 516467 172486 516467 2 dpga_flat_0.sr_0.FILLER_0_26_3.decap_12
flabel metal1 173619 516450 173653 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_15.VGND
flabel metal1 173619 515906 173653 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_15.VPWR
flabel nwell 173619 515906 173653 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_15.VPB
flabel pwell 173619 516450 173653 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_15.VNB
rlabel comment 173590 516467 173590 516467 2 dpga_flat_0.sr_0.FILLER_0_26_15.decap_12
flabel metal1 172515 515906 172549 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_3.VPWR
flabel metal1 172515 515362 172549 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_3.VGND
flabel nwell 172515 515906 172549 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_3.VPB
flabel pwell 172515 515362 172549 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_3.VNB
rlabel comment 172486 515379 172486 515379 4 dpga_flat_0.sr_0.FILLER_0_27_3.decap_8
rlabel metal1 172486 515331 173222 515427 1 dpga_flat_0.sr_0.FILLER_0_27_3.VGND
rlabel metal1 172486 515875 173222 515971 1 dpga_flat_0.sr_0.FILLER_0_27_3.VPWR
flabel metal1 173242 515365 173295 515397 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_11.VGND
flabel metal1 173243 515909 173295 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_11.VPWR
flabel nwell 173250 515914 173284 515932 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_11.VPB
flabel pwell 173253 515369 173285 515391 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_11.VNB
rlabel comment 173222 515379 173222 515379 4 dpga_flat_0.sr_0.FILLER_0_27_11.fill_2
rlabel metal1 173222 515331 173406 515427 1 dpga_flat_0.sr_0.FILLER_0_27_11.VGND
rlabel metal1 173222 515875 173406 515971 1 dpga_flat_0.sr_0.FILLER_0_27_11.VPWR
flabel metal1 173987 515906 174021 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_19.VPWR
flabel metal1 173987 515362 174021 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_19.VGND
flabel nwell 173987 515906 174021 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_19.VPB
flabel pwell 173987 515362 174021 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_19.VNB
rlabel comment 173958 515379 173958 515379 4 dpga_flat_0.sr_0.FILLER_0_27_19.decap_8
rlabel metal1 173958 515331 174694 515427 1 dpga_flat_0.sr_0.FILLER_0_27_19.VGND
rlabel metal1 173958 515875 174694 515971 1 dpga_flat_0.sr_0.FILLER_0_27_19.VPWR
flabel metal1 172239 515906 172273 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_26_Left_54.VPWR
flabel metal1 172239 516450 172273 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_26_Left_54.VGND
flabel nwell 172239 515906 172273 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_26_Left_54.VPB
flabel pwell 172239 516450 172273 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_26_Left_54.VNB
rlabel comment 172210 516467 172210 516467 2 dpga_flat_0.sr_0.PHY_EDGE_ROW_26_Left_54.decap_3
rlabel metal1 172210 516419 172486 516515 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_26_Left_54.VGND
rlabel metal1 172210 515875 172486 515971 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_26_Left_54.VPWR
flabel metal1 172239 515906 172273 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_27_Left_55.VPWR
flabel metal1 172239 515362 172273 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_27_Left_55.VGND
flabel nwell 172239 515906 172273 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_27_Left_55.VPB
flabel pwell 172239 515362 172273 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_27_Left_55.VNB
rlabel comment 172210 515379 172210 515379 4 dpga_flat_0.sr_0.PHY_EDGE_ROW_27_Left_55.decap_3
rlabel metal1 172210 515331 172486 515427 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_27_Left_55.VGND
rlabel metal1 172210 515875 172486 515971 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_27_Left_55.VPWR
flabel locali 173803 515668 173837 515702 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input3.X
flabel locali 173527 515532 173561 515566 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input3.A
flabel locali 173895 515532 173929 515566 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input3.X
flabel locali 173527 515600 173561 515634 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input3.A
flabel locali 173895 515600 173929 515634 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input3.X
flabel metal1 173435 515362 173469 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input3.VGND
flabel metal1 173435 515906 173469 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input3.VPWR
flabel nwell 173435 515906 173469 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input3.VPB
flabel pwell 173435 515362 173469 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input3.VNB
rlabel comment 173406 515379 173406 515379 4 dpga_flat_0.sr_0.input3.clkbuf_4
rlabel metal1 173406 515331 173958 515427 1 dpga_flat_0.sr_0.input3.VGND
rlabel metal1 173406 515875 173958 515971 1 dpga_flat_0.sr_0.input3.VPWR
flabel metal1 174716 515910 174752 515940 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_27.VPWR
flabel metal1 174716 516451 174752 516480 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_27.VGND
flabel nwell 174725 515916 174745 515933 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_27.VPB
flabel pwell 174722 516456 174746 516478 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_27.VNB
rlabel comment 174694 516467 174694 516467 2 dpga_flat_0.sr_0.FILLER_0_26_27.fill_1
rlabel metal1 174694 516419 174786 516515 5 dpga_flat_0.sr_0.FILLER_0_26_27.VGND
rlabel metal1 174694 515875 174786 515971 5 dpga_flat_0.sr_0.FILLER_0_26_27.VPWR
flabel metal1 174907 516450 174941 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_29.VGND
flabel metal1 174907 515906 174941 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_29.VPWR
flabel nwell 174907 515906 174941 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_29.VPB
flabel pwell 174907 516450 174941 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_29.VNB
rlabel comment 174878 516467 174878 516467 2 dpga_flat_0.sr_0.FILLER_0_26_29.decap_12
flabel metal1 176011 516450 176045 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_41.VGND
flabel metal1 176011 515906 176045 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_41.VPWR
flabel nwell 176011 515906 176045 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_41.VPB
flabel pwell 176011 516450 176045 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_41.VNB
rlabel comment 175982 516467 175982 516467 2 dpga_flat_0.sr_0.FILLER_0_26_41.decap_12
flabel metal1 174716 515906 174752 515936 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_27.VPWR
flabel metal1 174716 515366 174752 515395 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_27.VGND
flabel nwell 174725 515913 174745 515930 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_27.VPB
flabel pwell 174722 515368 174746 515390 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_27.VNB
rlabel comment 174694 515379 174694 515379 4 dpga_flat_0.sr_0.FILLER_0_27_27.fill_1
rlabel metal1 174694 515331 174786 515427 1 dpga_flat_0.sr_0.FILLER_0_27_27.VGND
rlabel metal1 174694 515875 174786 515971 1 dpga_flat_0.sr_0.FILLER_0_27_27.VPWR
flabel metal1 174907 515362 174941 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_29.VGND
flabel metal1 174907 515906 174941 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_29.VPWR
flabel nwell 174907 515906 174941 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_29.VPB
flabel pwell 174907 515362 174941 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_29.VNB
rlabel comment 174878 515379 174878 515379 4 dpga_flat_0.sr_0.FILLER_0_27_29.decap_12
flabel metal1 176011 515362 176045 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_41.VGND
flabel metal1 176011 515906 176045 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_41.VPWR
flabel nwell 176011 515906 176045 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_41.VPB
flabel pwell 176011 515362 176045 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_41.VNB
rlabel comment 175982 515379 175982 515379 4 dpga_flat_0.sr_0.FILLER_0_27_41.decap_12
flabel metal1 174808 515914 174861 515943 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_26_123.VPWR
flabel metal1 174807 516447 174858 516485 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_26_123.VGND
rlabel comment 174786 516467 174786 516467 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_26_123.tapvpwrvgnd_1
rlabel metal1 174786 516419 174878 516515 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_26_123.VGND
rlabel metal1 174786 515875 174878 515971 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_26_123.VPWR
flabel metal1 174808 515903 174861 515932 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_126.VPWR
flabel metal1 174807 515361 174858 515399 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_126.VGND
rlabel comment 174786 515379 174786 515379 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_126.tapvpwrvgnd_1
rlabel metal1 174786 515331 174878 515427 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_126.VGND
rlabel metal1 174786 515875 174878 515971 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_126.VPWR
flabel metal1 177115 516450 177149 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_53.VGND
flabel metal1 177115 515906 177149 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_53.VPWR
flabel nwell 177115 515906 177149 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_53.VPB
flabel pwell 177115 516450 177149 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_53.VNB
rlabel comment 177086 516467 177086 516467 2 dpga_flat_0.sr_0.FILLER_0_26_53.decap_12
flabel metal1 177115 515906 177149 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_53.VPWR
flabel metal1 177115 515362 177149 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_53.VGND
flabel nwell 177115 515906 177149 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_53.VPB
flabel pwell 177115 515362 177149 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_53.VNB
rlabel comment 177086 515379 177086 515379 4 dpga_flat_0.sr_0.FILLER_0_27_53.decap_3
rlabel metal1 177086 515331 177362 515427 1 dpga_flat_0.sr_0.FILLER_0_27_53.VGND
rlabel metal1 177086 515875 177362 515971 1 dpga_flat_0.sr_0.FILLER_0_27_53.VPWR
flabel metal1 177483 515362 177517 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_57.VGND
flabel metal1 177483 515906 177517 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_57.VPWR
flabel nwell 177483 515906 177517 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_57.VPB
flabel pwell 177483 515362 177517 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_57.VNB
rlabel comment 177454 515379 177454 515379 4 dpga_flat_0.sr_0.FILLER_0_27_57.decap_12
flabel metal1 177384 515903 177437 515932 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_127.VPWR
flabel metal1 177383 515361 177434 515399 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_127.VGND
rlabel comment 177362 515379 177362 515379 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_127.tapvpwrvgnd_1
rlabel metal1 177362 515331 177454 515427 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_127.VGND
rlabel metal1 177362 515875 177454 515971 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_127.VPWR
flabel metal1 178219 516450 178253 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_65.VGND
flabel metal1 178219 515906 178253 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_65.VPWR
flabel nwell 178219 515906 178253 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_65.VPB
flabel pwell 178219 516450 178253 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_65.VNB
rlabel comment 178190 516467 178190 516467 2 dpga_flat_0.sr_0.FILLER_0_26_65.decap_12
flabel metal1 179323 515906 179357 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_77.VPWR
flabel metal1 179323 516450 179357 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_77.VGND
flabel nwell 179323 515906 179357 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_77.VPB
flabel pwell 179323 516450 179357 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_77.VNB
rlabel comment 179294 516467 179294 516467 2 dpga_flat_0.sr_0.FILLER_0_26_77.decap_6
rlabel metal1 179294 516419 179846 516515 5 dpga_flat_0.sr_0.FILLER_0_26_77.VGND
rlabel metal1 179294 515875 179846 515971 5 dpga_flat_0.sr_0.FILLER_0_26_77.VPWR
flabel metal1 179868 515910 179904 515940 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_83.VPWR
flabel metal1 179868 516451 179904 516480 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_83.VGND
flabel nwell 179877 515916 179897 515933 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_83.VPB
flabel pwell 179874 516456 179898 516478 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_83.VNB
rlabel comment 179846 516467 179846 516467 2 dpga_flat_0.sr_0.FILLER_0_26_83.fill_1
rlabel metal1 179846 516419 179938 516515 5 dpga_flat_0.sr_0.FILLER_0_26_83.VGND
rlabel metal1 179846 515875 179938 515971 5 dpga_flat_0.sr_0.FILLER_0_26_83.VPWR
flabel metal1 178587 515362 178621 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_69.VGND
flabel metal1 178587 515906 178621 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_69.VPWR
flabel nwell 178587 515906 178621 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_69.VPB
flabel pwell 178587 515362 178621 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_69.VNB
rlabel comment 178558 515379 178558 515379 4 dpga_flat_0.sr_0.FILLER_0_27_69.decap_12
flabel metal1 179691 515906 179725 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_81.VPWR
flabel metal1 179691 515362 179725 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_81.VGND
flabel nwell 179691 515906 179725 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_81.VPB
flabel pwell 179691 515362 179725 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_81.VNB
rlabel comment 179662 515379 179662 515379 4 dpga_flat_0.sr_0.FILLER_0_27_81.decap_3
rlabel metal1 179662 515331 179938 515427 1 dpga_flat_0.sr_0.FILLER_0_27_81.VGND
rlabel metal1 179662 515875 179938 515971 1 dpga_flat_0.sr_0.FILLER_0_27_81.VPWR
flabel metal1 180059 516450 180093 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_85.VGND
flabel metal1 180059 515906 180093 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_85.VPWR
flabel nwell 180059 515906 180093 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_85.VPB
flabel pwell 180059 516450 180093 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_85.VNB
rlabel comment 180030 516467 180030 516467 2 dpga_flat_0.sr_0.FILLER_0_26_85.decap_12
flabel metal1 181163 516450 181197 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_97.VGND
flabel metal1 181163 515906 181197 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_97.VPWR
flabel nwell 181163 515906 181197 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_97.VPB
flabel pwell 181163 516450 181197 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_97.VNB
rlabel comment 181134 516467 181134 516467 2 dpga_flat_0.sr_0.FILLER_0_26_97.decap_12
flabel metal1 180059 515362 180093 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_85.VGND
flabel metal1 180059 515906 180093 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_85.VPWR
flabel nwell 180059 515906 180093 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_85.VPB
flabel pwell 180059 515362 180093 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_85.VNB
rlabel comment 180030 515379 180030 515379 4 dpga_flat_0.sr_0.FILLER_0_27_85.decap_12
flabel metal1 181163 515906 181197 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_97.VPWR
flabel metal1 181163 515362 181197 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_97.VGND
flabel nwell 181163 515906 181197 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_97.VPB
flabel pwell 181163 515362 181197 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_97.VNB
rlabel comment 181134 515379 181134 515379 4 dpga_flat_0.sr_0.FILLER_0_27_97.decap_8
rlabel metal1 181134 515331 181870 515427 1 dpga_flat_0.sr_0.FILLER_0_27_97.VGND
rlabel metal1 181134 515875 181870 515971 1 dpga_flat_0.sr_0.FILLER_0_27_97.VPWR
flabel metal1 179960 515914 180013 515943 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_26_124.VPWR
flabel metal1 179959 516447 180010 516485 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_26_124.VGND
rlabel comment 179938 516467 179938 516467 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_26_124.tapvpwrvgnd_1
rlabel metal1 179938 516419 180030 516515 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_26_124.VGND
rlabel metal1 179938 515875 180030 515971 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_26_124.VPWR
flabel metal1 179960 515903 180013 515932 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_128.VPWR
flabel metal1 179959 515361 180010 515399 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_128.VGND
rlabel comment 179938 515379 179938 515379 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_128.tapvpwrvgnd_1
rlabel metal1 179938 515331 180030 515427 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_128.VGND
rlabel metal1 179938 515875 180030 515971 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_128.VPWR
flabel metal1 182267 516450 182301 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_109.VGND
flabel metal1 182267 515906 182301 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_109.VPWR
flabel nwell 182267 515906 182301 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_109.VPB
flabel pwell 182267 516450 182301 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_109.VNB
rlabel comment 182238 516467 182238 516467 2 dpga_flat_0.sr_0.FILLER_0_26_109.decap_12
flabel metal1 183371 516450 183405 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_121.VGND
flabel metal1 183371 515906 183405 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_121.VPWR
flabel nwell 183371 515906 183405 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_121.VPB
flabel pwell 183371 516450 183405 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_121.VNB
rlabel comment 183342 516467 183342 516467 2 dpga_flat_0.sr_0.FILLER_0_26_121.decap_12
flabel metal1 181890 515365 181943 515397 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_105.VGND
flabel metal1 181891 515909 181943 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_105.VPWR
flabel nwell 181898 515914 181932 515932 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_105.VPB
flabel pwell 181901 515369 181933 515391 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_105.VNB
rlabel comment 181870 515379 181870 515379 4 dpga_flat_0.sr_0.FILLER_0_27_105.fill_2
rlabel metal1 181870 515331 182054 515427 1 dpga_flat_0.sr_0.FILLER_0_27_105.VGND
rlabel metal1 181870 515875 182054 515971 1 dpga_flat_0.sr_0.FILLER_0_27_105.VPWR
flabel metal1 182350 515365 182403 515397 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_110.VGND
flabel metal1 182351 515909 182403 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_110.VPWR
flabel nwell 182358 515914 182392 515932 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_110.VPB
flabel pwell 182361 515369 182393 515391 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_110.VNB
rlabel comment 182330 515379 182330 515379 4 dpga_flat_0.sr_0.FILLER_0_27_110.fill_2
rlabel metal1 182330 515331 182514 515427 1 dpga_flat_0.sr_0.FILLER_0_27_110.VGND
rlabel metal1 182330 515875 182514 515971 1 dpga_flat_0.sr_0.FILLER_0_27_110.VPWR
flabel metal1 182635 515362 182669 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_113.VGND
flabel metal1 182635 515906 182669 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_113.VPWR
flabel nwell 182635 515906 182669 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_113.VPB
flabel pwell 182635 515362 182669 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_113.VNB
rlabel comment 182606 515379 182606 515379 4 dpga_flat_0.sr_0.FILLER_0_27_113.decap_12
flabel metal1 183739 515362 183773 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_125.VGND
flabel metal1 183739 515906 183773 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_125.VPWR
flabel nwell 183739 515906 183773 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_125.VPB
flabel pwell 183739 515362 183773 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_125.VNB
rlabel comment 183710 515379 183710 515379 4 dpga_flat_0.sr_0.FILLER_0_27_125.decap_12
flabel metal1 182536 515903 182589 515932 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_129.VPWR
flabel metal1 182535 515361 182586 515399 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_129.VGND
rlabel comment 182514 515379 182514 515379 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_129.tapvpwrvgnd_1
rlabel metal1 182514 515331 182606 515427 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_129.VGND
rlabel metal1 182514 515875 182606 515971 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_129.VPWR
flabel metal1 182265 515362 182299 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input2.VGND
flabel metal1 182267 515906 182301 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input2.VPWR
flabel locali 182267 515906 182301 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input2.VPWR
flabel locali 182265 515362 182299 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input2.VGND
flabel locali 182085 515464 182119 515498 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input2.X
flabel locali 182085 515736 182119 515770 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input2.X
flabel locali 182085 515804 182119 515838 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input2.X
flabel locali 182267 515600 182301 515634 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input2.A
flabel nwell 182267 515906 182301 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input2.VPB
flabel pwell 182265 515362 182299 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input2.VNB
rlabel comment 182330 515379 182330 515379 6 dpga_flat_0.sr_0.input2.buf_1
rlabel metal1 182054 515331 182330 515427 1 dpga_flat_0.sr_0.input2.VGND
rlabel metal1 182054 515875 182330 515971 1 dpga_flat_0.sr_0.input2.VPWR
flabel metal1 184475 515906 184509 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_133.VPWR
flabel metal1 184475 516450 184509 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_133.VGND
flabel nwell 184475 515906 184509 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_133.VPB
flabel pwell 184475 516450 184509 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_133.VNB
rlabel comment 184446 516467 184446 516467 2 dpga_flat_0.sr_0.FILLER_0_26_133.decap_6
rlabel metal1 184446 516419 184998 516515 5 dpga_flat_0.sr_0.FILLER_0_26_133.VGND
rlabel metal1 184446 515875 184998 515971 5 dpga_flat_0.sr_0.FILLER_0_26_133.VPWR
flabel metal1 185020 515910 185056 515940 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_139.VPWR
flabel metal1 185020 516451 185056 516480 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_139.VGND
flabel nwell 185029 515916 185049 515933 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_139.VPB
flabel pwell 185026 516456 185050 516478 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_139.VNB
rlabel comment 184998 516467 184998 516467 2 dpga_flat_0.sr_0.FILLER_0_26_139.fill_1
rlabel metal1 184998 516419 185090 516515 5 dpga_flat_0.sr_0.FILLER_0_26_139.VGND
rlabel metal1 184998 515875 185090 515971 5 dpga_flat_0.sr_0.FILLER_0_26_139.VPWR
flabel metal1 185211 516450 185245 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_141.VGND
flabel metal1 185211 515906 185245 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_141.VPWR
flabel nwell 185211 515906 185245 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_141.VPB
flabel pwell 185211 516450 185245 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_141.VNB
rlabel comment 185182 516467 185182 516467 2 dpga_flat_0.sr_0.FILLER_0_26_141.decap_12
flabel metal1 184843 515906 184877 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_137.VPWR
flabel metal1 184843 515362 184877 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_137.VGND
flabel nwell 184843 515906 184877 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_137.VPB
flabel pwell 184843 515362 184877 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_137.VNB
rlabel comment 184814 515379 184814 515379 4 dpga_flat_0.sr_0.FILLER_0_27_137.decap_3
rlabel metal1 184814 515331 185090 515427 1 dpga_flat_0.sr_0.FILLER_0_27_137.VGND
rlabel metal1 184814 515875 185090 515971 1 dpga_flat_0.sr_0.FILLER_0_27_137.VPWR
flabel metal1 185211 515362 185245 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_141.VGND
flabel metal1 185211 515906 185245 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_141.VPWR
flabel nwell 185211 515906 185245 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_141.VPB
flabel pwell 185211 515362 185245 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_141.VNB
rlabel comment 185182 515379 185182 515379 4 dpga_flat_0.sr_0.FILLER_0_27_141.decap_12
flabel metal1 185112 515914 185165 515943 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_26_125.VPWR
flabel metal1 185111 516447 185162 516485 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_26_125.VGND
rlabel comment 185090 516467 185090 516467 2 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_26_125.tapvpwrvgnd_1
rlabel metal1 185090 516419 185182 516515 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_26_125.VGND
rlabel metal1 185090 515875 185182 515971 5 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_26_125.VPWR
flabel metal1 185112 515903 185165 515932 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_130.VPWR
flabel metal1 185111 515361 185162 515399 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_130.VGND
rlabel comment 185090 515379 185090 515379 4 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_130.tapvpwrvgnd_1
rlabel metal1 185090 515331 185182 515427 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_130.VGND
rlabel metal1 185090 515875 185182 515971 1 dpga_flat_0.sr_0.TAP_TAPCELL_ROW_27_130.VPWR
flabel metal1 186315 515906 186349 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_153.VPWR
flabel metal1 186315 516450 186349 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_153.VGND
flabel nwell 186315 515906 186349 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_153.VPB
flabel pwell 186315 516450 186349 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_153.VNB
rlabel comment 186286 516467 186286 516467 2 dpga_flat_0.sr_0.FILLER_0_26_153.decap_8
rlabel metal1 186286 516419 187022 516515 5 dpga_flat_0.sr_0.FILLER_0_26_153.VGND
rlabel metal1 186286 515875 187022 515971 5 dpga_flat_0.sr_0.FILLER_0_26_153.VPWR
flabel metal1 187042 516449 187095 516481 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_161.VGND
flabel metal1 187043 515906 187095 515937 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_161.VPWR
flabel nwell 187050 515914 187084 515932 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_161.VPB
flabel pwell 187053 516455 187085 516477 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_26_161.VNB
rlabel comment 187022 516467 187022 516467 2 dpga_flat_0.sr_0.FILLER_0_26_161.fill_2
rlabel metal1 187022 516419 187206 516515 5 dpga_flat_0.sr_0.FILLER_0_26_161.VGND
rlabel metal1 187022 515875 187206 515971 5 dpga_flat_0.sr_0.FILLER_0_26_161.VPWR
flabel metal1 186308 515906 186344 515936 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_153.VPWR
flabel metal1 186308 515366 186344 515395 0 FreeSans 250 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_153.VGND
flabel nwell 186317 515913 186337 515930 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_153.VPB
flabel pwell 186314 515368 186338 515390 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_153.VNB
rlabel comment 186286 515379 186286 515379 4 dpga_flat_0.sr_0.FILLER_0_27_153.fill_1
rlabel metal1 186286 515331 186378 515427 1 dpga_flat_0.sr_0.FILLER_0_27_153.VGND
rlabel metal1 186286 515875 186378 515971 1 dpga_flat_0.sr_0.FILLER_0_27_153.VPWR
flabel metal1 186959 515906 186993 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_160.VPWR
flabel metal1 186959 515362 186993 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_160.VGND
flabel nwell 186959 515906 186993 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_160.VPB
flabel pwell 186959 515362 186993 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.FILLER_0_27_160.VNB
rlabel comment 186930 515379 186930 515379 4 dpga_flat_0.sr_0.FILLER_0_27_160.decap_3
rlabel metal1 186930 515331 187206 515427 1 dpga_flat_0.sr_0.FILLER_0_27_160.VGND
rlabel metal1 186930 515875 187206 515971 1 dpga_flat_0.sr_0.FILLER_0_27_160.VPWR
flabel metal1 187419 515906 187453 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_26_Right_26.VPWR
flabel metal1 187419 516450 187453 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_26_Right_26.VGND
flabel nwell 187419 515906 187453 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_26_Right_26.VPB
flabel pwell 187419 516450 187453 516484 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_26_Right_26.VNB
rlabel comment 187482 516467 187482 516467 8 dpga_flat_0.sr_0.PHY_EDGE_ROW_26_Right_26.decap_3
rlabel metal1 187206 516419 187482 516515 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_26_Right_26.VGND
rlabel metal1 187206 515875 187482 515971 5 dpga_flat_0.sr_0.PHY_EDGE_ROW_26_Right_26.VPWR
flabel metal1 187419 515906 187453 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_27_Right_27.VPWR
flabel metal1 187419 515362 187453 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_27_Right_27.VGND
flabel nwell 187419 515906 187453 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_27_Right_27.VPB
flabel pwell 187419 515362 187453 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.PHY_EDGE_ROW_27_Right_27.VNB
rlabel comment 187482 515379 187482 515379 6 dpga_flat_0.sr_0.PHY_EDGE_ROW_27_Right_27.decap_3
rlabel metal1 187206 515331 187482 515427 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_27_Right_27.VGND
rlabel metal1 187206 515875 187482 515971 1 dpga_flat_0.sr_0.PHY_EDGE_ROW_27_Right_27.VPWR
flabel locali 186775 515668 186809 515702 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input1.X
flabel locali 186499 515532 186533 515566 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input1.A
flabel locali 186867 515532 186901 515566 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input1.X
flabel locali 186499 515600 186533 515634 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input1.A
flabel locali 186867 515600 186901 515634 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input1.X
flabel metal1 186407 515362 186441 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input1.VGND
flabel metal1 186407 515906 186441 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input1.VPWR
flabel nwell 186407 515906 186441 515940 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input1.VPB
flabel pwell 186407 515362 186441 515396 0 FreeSans 200 0 0 0 dpga_flat_0.sr_0.input1.VNB
rlabel comment 186378 515379 186378 515379 4 dpga_flat_0.sr_0.input1.clkbuf_4
rlabel metal1 186378 515331 186930 515427 1 dpga_flat_0.sr_0.input1.VGND
rlabel metal1 186378 515875 186930 515971 1 dpga_flat_0.sr_0.input1.VPWR
flabel metal1 157000 536797 157200 536987 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.out
flabel metal1 192230 540097 192430 540287 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.gnd
flabel metal1 192230 539147 192430 539347 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.vd
flabel metal1 163530 542597 163730 542787 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.inp
flabel metal1 178180 542557 178380 542747 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.inn
flabel metal1 163030 533347 163230 533537 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.ib
flabel metal1 167520 533337 167720 533537 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.c0
flabel metal1 171050 533337 171250 533537 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.c1
flabel metal1 174680 533337 174880 533537 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.c2
flabel metal1 178220 533337 178420 533537 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.c3
flabel metal1 181730 533337 181930 533537 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.c4
flabel metal1 184970 533337 185170 533537 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.c5
flabel metal1 188200 533337 188400 533537 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.c6
flabel metal1 191480 533337 191680 533537 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.c7
flabel metal1 163030 538707 163230 538907 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.ota_0.vs
flabel metal1 163020 537027 163220 537227 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.ota_0.inn
flabel metal1 163020 537867 163220 538067 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.ota_0.inp
flabel metal1 163030 536597 163230 536797 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.ota_0.ib
flabel metal1 160180 535417 160380 535617 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.ota_0.vd
flabel metal1 157200 536787 157400 536987 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.ota_0.out
flabel metal1 161450 538077 161490 538097 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.ota_0.d
flabel metal1 162190 538077 162190 538097 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.ota_0.c
flabel metal2 161650 536857 161670 536877 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.ota_0.b
flabel metal1 167520 535247 167720 535447 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.c0
flabel metal1 171050 535247 171250 535447 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.c1
flabel metal1 174680 535247 174880 535447 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.c2
flabel metal1 178220 535247 178420 535447 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.c3
flabel metal1 181730 535247 181930 535447 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.c4
flabel metal1 184970 535247 185170 535447 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.c5
flabel metal1 188200 535247 188400 535447 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.c6
flabel metal1 191480 535247 191680 535447 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.c7
flabel metal1 178180 542097 178380 542297 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.n0
flabel metal1 163530 536037 163730 536237 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.n8
flabel metal1 192030 540087 192230 540287 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.gnd
flabel metal1 192030 539147 192230 539347 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.vd
flabel metal1 170480 539147 170680 539347 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_7.vd
flabel metal1 168080 539587 168280 539787 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_7.b
flabel metal1 170480 540087 170680 540287 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_7.vgnd
flabel metal1 170480 540727 170680 540927 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_7.ctrl
flabel metal1 168080 540867 168280 541067 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_7.a
flabel metal1 169940 538517 169960 538527 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_7.nctrl
flabel metal1 174180 539147 174380 539347 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_6.vd
flabel metal1 171780 539587 171980 539787 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_6.b
flabel metal1 174180 540087 174380 540287 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_6.vgnd
flabel metal1 174180 540727 174380 540927 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_6.ctrl
flabel metal1 171780 540867 171980 541067 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_6.a
flabel metal1 173640 538517 173660 538527 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_6.nctrl
flabel metal1 177680 539147 177880 539347 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_5.vd
flabel metal1 175280 539587 175480 539787 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_5.b
flabel metal1 177680 540087 177880 540287 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_5.vgnd
flabel metal1 177680 540727 177880 540927 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_5.ctrl
flabel metal1 175280 540867 175480 541067 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_5.a
flabel metal1 177140 538517 177160 538527 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_5.nctrl
flabel metal1 166680 539147 166880 539347 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_4.vd
flabel metal1 164280 539587 164480 539787 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_4.b
flabel metal1 166680 540087 166880 540287 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_4.vgnd
flabel metal1 166680 540727 166880 540927 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_4.ctrl
flabel metal1 164280 540867 164480 541067 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_4.a
flabel metal1 166140 538517 166160 538527 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_4.nctrl
flabel metal1 181280 539147 181480 539347 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_3.vd
flabel metal1 178880 539587 179080 539787 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_3.b
flabel metal1 181280 540087 181480 540287 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_3.vgnd
flabel metal1 181280 540727 181480 540927 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_3.ctrl
flabel metal1 178880 540867 179080 541067 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_3.a
flabel metal1 180740 538517 180760 538527 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_3.nctrl
flabel metal1 184580 539147 184780 539347 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_2.vd
flabel metal1 182180 539587 182380 539787 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_2.b
flabel metal1 184580 540087 184780 540287 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_2.vgnd
flabel metal1 184580 540727 184780 540927 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_2.ctrl
flabel metal1 182180 540867 182380 541067 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_2.a
flabel metal1 184040 538517 184060 538527 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_2.nctrl
flabel metal1 191180 539147 191380 539347 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_1.vd
flabel metal1 188780 539587 188980 539787 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_1.b
flabel metal1 191180 540087 191380 540287 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_1.vgnd
flabel metal1 191180 540727 191380 540927 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_1.ctrl
flabel metal1 188780 540867 188980 541067 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_1.a
flabel metal1 190640 538517 190660 538527 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_1.nctrl
flabel metal1 187880 539147 188080 539347 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_0.vd
flabel metal1 185480 539587 185680 539787 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_0.b
flabel metal1 187880 540087 188080 540287 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_0.vgnd
flabel metal1 187880 540727 188080 540927 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_0.ctrl
flabel metal1 185480 540867 185680 541067 0 FreeSans 256 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_0.a
flabel metal1 187340 538517 187360 538527 0 FreeSans 1600 0 0 0 dpga_flat_0.ota_digpot_0.digpotp_0.tg_0.nctrl
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1699065138
use cafeina_top_level  cafeina_top_level_0
timestamp 1699054617
transform 1 0 0 0 1 9
box 217294 450753 583581 703284
use dpga_wires_flat  dpga_wires_flat_0
timestamp 1699064461
transform 1 0 -2 0 1 2
box 600 377990 195000 703400
use gme_cefet_top_level  gme_cefet_top_level_0
timestamp 1699054617
transform 1 0 78 0 1 -9
box 326 15091 583606 406686
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
